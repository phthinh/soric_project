VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO flexbex_ibex_core
  CLASS BLOCK ;
  FOREIGN flexbex_ibex_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN boot_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 74.160 1200.000 74.760 ;
    END
  END boot_addr_i[0]
  PIN boot_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END boot_addr_i[10]
  PIN boot_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 1196.000 426.330 1200.000 ;
    END
  END boot_addr_i[11]
  PIN boot_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END boot_addr_i[12]
  PIN boot_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END boot_addr_i[13]
  PIN boot_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 1196.000 546.390 1200.000 ;
    END
  END boot_addr_i[14]
  PIN boot_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 605.240 1200.000 605.840 ;
    END
  END boot_addr_i[15]
  PIN boot_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 1196.000 678.410 1200.000 ;
    END
  END boot_addr_i[16]
  PIN boot_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 674.600 1200.000 675.200 ;
    END
  END boot_addr_i[17]
  PIN boot_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 1196.000 714.290 1200.000 ;
    END
  END boot_addr_i[18]
  PIN boot_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 723.560 4.000 724.160 ;
    END
  END boot_addr_i[19]
  PIN boot_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 131.960 1200.000 132.560 ;
    END
  END boot_addr_i[1]
  PIN boot_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END boot_addr_i[20]
  PIN boot_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 1196.000 822.390 1200.000 ;
    END
  END boot_addr_i[21]
  PIN boot_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END boot_addr_i[22]
  PIN boot_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.830 1196.000 906.110 1200.000 ;
    END
  END boot_addr_i[23]
  PIN boot_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 0.000 942.910 4.000 ;
    END
  END boot_addr_i[24]
  PIN boot_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 1196.000 966.370 1200.000 ;
    END
  END boot_addr_i[25]
  PIN boot_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 0.000 999.950 4.000 ;
    END
  END boot_addr_i[26]
  PIN boot_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1043.840 1200.000 1044.440 ;
    END
  END boot_addr_i[27]
  PIN boot_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.720 4.000 1089.320 ;
    END
  END boot_addr_i[28]
  PIN boot_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.080 4.000 1141.680 ;
    END
  END boot_addr_i[29]
  PIN boot_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END boot_addr_i[2]
  PIN boot_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.250 0.000 1148.530 4.000 ;
    END
  END boot_addr_i[30]
  PIN boot_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.990 1196.000 1134.270 1200.000 ;
    END
  END boot_addr_i[31]
  PIN boot_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 178.200 1200.000 178.800 ;
    END
  END boot_addr_i[3]
  PIN boot_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 247.560 1200.000 248.160 ;
    END
  END boot_addr_i[4]
  PIN boot_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 1196.000 246.010 1200.000 ;
    END
  END boot_addr_i[5]
  PIN boot_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 340.040 1200.000 340.640 ;
    END
  END boot_addr_i[6]
  PIN boot_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 397.840 1200.000 398.440 ;
    END
  END boot_addr_i[7]
  PIN boot_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 1196.000 401.950 1200.000 ;
    END
  END boot_addr_i[8]
  PIN boot_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END boot_addr_i[9]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 5.480 1200.000 6.080 ;
    END
  END clk_i
  PIN cluster_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END cluster_id_i[0]
  PIN cluster_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END cluster_id_i[1]
  PIN cluster_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END cluster_id_i[2]
  PIN cluster_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END cluster_id_i[3]
  PIN cluster_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END cluster_id_i[4]
  PIN cluster_id_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 1196.000 257.970 1200.000 ;
    END
  END cluster_id_i[5]
  PIN core_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END core_id_i[0]
  PIN core_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END core_id_i[1]
  PIN core_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END core_id_i[2]
  PIN core_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 1196.000 186.210 1200.000 ;
    END
  END core_id_i[3]
  PIN data_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END data_addr_o[0]
  PIN data_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 1196.000 414.370 1200.000 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 1196.000 462.210 1200.000 ;
    END
  END data_addr_o[12]
  PIN data_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 1196.000 498.090 1200.000 ;
    END
  END data_addr_o[13]
  PIN data_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 582.120 1200.000 582.720 ;
    END
  END data_addr_o[14]
  PIN data_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 1196.000 618.150 1200.000 ;
    END
  END data_addr_o[15]
  PIN data_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 0.000 771.330 4.000 ;
    END
  END data_addr_o[16]
  PIN data_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END data_addr_o[17]
  PIN data_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 1196.000 726.250 1200.000 ;
    END
  END data_addr_o[18]
  PIN data_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 736.480 4.000 737.080 ;
    END
  END data_addr_o[19]
  PIN data_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 1196.000 78.110 1200.000 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 1196.000 786.050 1200.000 ;
    END
  END data_addr_o[20]
  PIN data_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 812.640 1200.000 813.240 ;
    END
  END data_addr_o[21]
  PIN data_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 1196.000 858.270 1200.000 ;
    END
  END data_addr_o[22]
  PIN data_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END data_addr_o[23]
  PIN data_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 1196.000 954.410 1200.000 ;
    END
  END data_addr_o[24]
  PIN data_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 986.040 1200.000 986.640 ;
    END
  END data_addr_o[25]
  PIN data_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1010.520 4.000 1011.120 ;
    END
  END data_addr_o[26]
  PIN data_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1055.400 1200.000 1056.000 ;
    END
  END data_addr_o[27]
  PIN data_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END data_addr_o[28]
  PIN data_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 4.000 ;
    END
  END data_addr_o[29]
  PIN data_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1154.000 4.000 1154.600 ;
    END
  END data_addr_o[30]
  PIN data_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1171.000 1200.000 1171.600 ;
    END
  END data_addr_o[31]
  PIN data_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 189.760 1200.000 190.360 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 259.120 1200.000 259.720 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 1196.000 318.230 1200.000 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 408.720 1200.000 409.320 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END data_addr_o[9]
  PIN data_be_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 1196.000 42.230 1200.000 ;
    END
  END data_be_o[0]
  PIN data_be_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 1196.000 90.070 1200.000 ;
    END
  END data_be_o[1]
  PIN data_be_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 1196.000 137.910 1200.000 ;
    END
  END data_be_o[2]
  PIN data_be_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 201.320 1200.000 201.920 ;
    END
  END data_be_o[3]
  PIN data_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END data_err_i
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END data_gnt_i
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END data_rdata_i[0]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 512.760 1200.000 513.360 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 535.880 1200.000 536.480 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 1196.000 558.350 1200.000 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 1196.000 630.110 1200.000 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 686.160 1200.000 686.760 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 1196.000 102.030 1200.000 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 1196.000 834.350 1200.000 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 893.560 1200.000 894.160 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.960 4.000 880.560 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 932.320 4.000 932.920 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 997.600 1200.000 998.200 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.800 4.000 1076.400 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1090.080 1200.000 1090.680 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.770 1196.000 1062.050 1200.000 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 1196.000 150.330 1200.000 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 1196.000 1098.390 1200.000 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1182.560 1200.000 1183.160 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 212.880 1200.000 213.480 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 270.680 1200.000 271.280 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 1196.000 269.930 1200.000 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 466.520 1200.000 467.120 ;
    END
  END data_rdata_i[9]
  PIN data_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 16.360 1200.000 16.960 ;
    END
  END data_req_o
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 27.920 1200.000 28.520 ;
    END
  END data_rvalid_i
  PIN data_wdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END data_wdata_o[0]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 1196.000 510.050 1200.000 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 1196.000 570.310 1200.000 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 1196.000 642.070 1200.000 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 628.360 1200.000 628.960 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 697.720 1200.000 698.320 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 0.000 862.870 4.000 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 1196.000 798.010 1200.000 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 824.200 1200.000 824.800 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.950 1196.000 870.230 1200.000 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 1196.000 918.070 1200.000 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.630 0.000 965.910 4.000 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.670 0.000 1045.950 4.000 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1114.560 4.000 1115.160 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.710 0.000 1102.990 4.000 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 1196.000 162.290 1200.000 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.750 0.000 1160.030 4.000 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 1196.000 1146.230 1200.000 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 1196.000 282.350 1200.000 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 0.000 565.710 4.000 ;
    END
  END data_wdata_o[9]
  PIN data_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 1196.000 6.350 1200.000 ;
    END
  END data_we_o
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END debug_req_i
  PIN eFPGA_delay_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 1196.000 54.190 1200.000 ;
    END
  END eFPGA_delay_o[0]
  PIN eFPGA_delay_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 1196.000 113.990 1200.000 ;
    END
  END eFPGA_delay_o[1]
  PIN eFPGA_delay_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END eFPGA_delay_o[2]
  PIN eFPGA_delay_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 1196.000 198.170 1200.000 ;
    END
  END eFPGA_delay_o[3]
  PIN eFPGA_en_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END eFPGA_en_o
  PIN eFPGA_fpga_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END eFPGA_fpga_done_i
  PIN eFPGA_operand_a_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 85.720 1200.000 86.320 ;
    END
  END eFPGA_operand_a_o[0]
  PIN eFPGA_operand_a_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 0.000 645.750 4.000 ;
    END
  END eFPGA_operand_a_o[10]
  PIN eFPGA_operand_a_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 547.440 1200.000 548.040 ;
    END
  END eFPGA_operand_a_o[11]
  PIN eFPGA_operand_a_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END eFPGA_operand_a_o[12]
  PIN eFPGA_operand_a_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END eFPGA_operand_a_o[13]
  PIN eFPGA_operand_a_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END eFPGA_operand_a_o[14]
  PIN eFPGA_operand_a_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END eFPGA_operand_a_o[15]
  PIN eFPGA_operand_a_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 1196.000 690.370 1200.000 ;
    END
  END eFPGA_operand_a_o[16]
  PIN eFPGA_operand_a_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 709.280 1200.000 709.880 ;
    END
  END eFPGA_operand_a_o[17]
  PIN eFPGA_operand_a_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END eFPGA_operand_a_o[18]
  PIN eFPGA_operand_a_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 767.080 1200.000 767.680 ;
    END
  END eFPGA_operand_a_o[19]
  PIN eFPGA_operand_a_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END eFPGA_operand_a_o[1]
  PIN eFPGA_operand_a_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 0.000 897.370 4.000 ;
    END
  END eFPGA_operand_a_o[20]
  PIN eFPGA_operand_a_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 835.760 1200.000 836.360 ;
    END
  END eFPGA_operand_a_o[21]
  PIN eFPGA_operand_a_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 827.600 4.000 828.200 ;
    END
  END eFPGA_operand_a_o[22]
  PIN eFPGA_operand_a_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 928.240 1200.000 928.840 ;
    END
  END eFPGA_operand_a_o[23]
  PIN eFPGA_operand_a_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 939.800 1200.000 940.400 ;
    END
  END eFPGA_operand_a_o[24]
  PIN eFPGA_operand_a_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 4.000 ;
    END
  END eFPGA_operand_a_o[25]
  PIN eFPGA_operand_a_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.280 4.000 1049.880 ;
    END
  END eFPGA_operand_a_o[26]
  PIN eFPGA_operand_a_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1066.960 1200.000 1067.560 ;
    END
  END eFPGA_operand_a_o[27]
  PIN eFPGA_operand_a_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 1196.000 1038.130 1200.000 ;
    END
  END eFPGA_operand_a_o[28]
  PIN eFPGA_operand_a_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.190 1196.000 1074.470 1200.000 ;
    END
  END eFPGA_operand_a_o[29]
  PIN eFPGA_operand_a_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END eFPGA_operand_a_o[2]
  PIN eFPGA_operand_a_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.250 0.000 1171.530 4.000 ;
    END
  END eFPGA_operand_a_o[30]
  PIN eFPGA_operand_a_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.840 4.000 1180.440 ;
    END
  END eFPGA_operand_a_o[31]
  PIN eFPGA_operand_a_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END eFPGA_operand_a_o[3]
  PIN eFPGA_operand_a_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 282.240 1200.000 282.840 ;
    END
  END eFPGA_operand_a_o[4]
  PIN eFPGA_operand_a_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 328.480 1200.000 329.080 ;
    END
  END eFPGA_operand_a_o[5]
  PIN eFPGA_operand_a_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 1196.000 330.190 1200.000 ;
    END
  END eFPGA_operand_a_o[6]
  PIN eFPGA_operand_a_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END eFPGA_operand_a_o[7]
  PIN eFPGA_operand_a_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 443.400 1200.000 444.000 ;
    END
  END eFPGA_operand_a_o[8]
  PIN eFPGA_operand_a_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END eFPGA_operand_a_o[9]
  PIN eFPGA_operand_b_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END eFPGA_operand_b_o[0]
  PIN eFPGA_operand_b_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 524.320 1200.000 524.920 ;
    END
  END eFPGA_operand_b_o[10]
  PIN eFPGA_operand_b_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 1196.000 438.290 1200.000 ;
    END
  END eFPGA_operand_b_o[11]
  PIN eFPGA_operand_b_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 570.560 1200.000 571.160 ;
    END
  END eFPGA_operand_b_o[12]
  PIN eFPGA_operand_b_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END eFPGA_operand_b_o[13]
  PIN eFPGA_operand_b_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 593.680 1200.000 594.280 ;
    END
  END eFPGA_operand_b_o[14]
  PIN eFPGA_operand_b_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 616.800 1200.000 617.400 ;
    END
  END eFPGA_operand_b_o[15]
  PIN eFPGA_operand_b_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 1196.000 702.330 1200.000 ;
    END
  END eFPGA_operand_b_o[16]
  PIN eFPGA_operand_b_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END eFPGA_operand_b_o[17]
  PIN eFPGA_operand_b_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 743.960 1200.000 744.560 ;
    END
  END eFPGA_operand_b_o[18]
  PIN eFPGA_operand_b_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 1196.000 762.130 1200.000 ;
    END
  END eFPGA_operand_b_o[19]
  PIN eFPGA_operand_b_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 1196.000 125.950 1200.000 ;
    END
  END eFPGA_operand_b_o[1]
  PIN eFPGA_operand_b_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 790.200 1200.000 790.800 ;
    END
  END eFPGA_operand_b_o[20]
  PIN eFPGA_operand_b_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 847.320 1200.000 847.920 ;
    END
  END eFPGA_operand_b_o[21]
  PIN eFPGA_operand_b_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END eFPGA_operand_b_o[22]
  PIN eFPGA_operand_b_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 1196.000 930.030 1200.000 ;
    END
  END eFPGA_operand_b_o[23]
  PIN eFPGA_operand_b_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.160 4.000 958.760 ;
    END
  END eFPGA_operand_b_o[24]
  PIN eFPGA_operand_b_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 984.000 4.000 984.600 ;
    END
  END eFPGA_operand_b_o[25]
  PIN eFPGA_operand_b_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.200 4.000 1062.800 ;
    END
  END eFPGA_operand_b_o[26]
  PIN eFPGA_operand_b_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 1196.000 1002.250 1200.000 ;
    END
  END eFPGA_operand_b_o[27]
  PIN eFPGA_operand_b_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1101.640 1200.000 1102.240 ;
    END
  END eFPGA_operand_b_o[28]
  PIN eFPGA_operand_b_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END eFPGA_operand_b_o[29]
  PIN eFPGA_operand_b_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 166.640 1200.000 167.240 ;
    END
  END eFPGA_operand_b_o[2]
  PIN eFPGA_operand_b_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.750 0.000 1183.030 4.000 ;
    END
  END eFPGA_operand_b_o[30]
  PIN eFPGA_operand_b_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1194.120 1200.000 1194.720 ;
    END
  END eFPGA_operand_b_o[31]
  PIN eFPGA_operand_b_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 224.440 1200.000 225.040 ;
    END
  END eFPGA_operand_b_o[3]
  PIN eFPGA_operand_b_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 1196.000 222.090 1200.000 ;
    END
  END eFPGA_operand_b_o[4]
  PIN eFPGA_operand_b_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END eFPGA_operand_b_o[5]
  PIN eFPGA_operand_b_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 351.600 1200.000 352.200 ;
    END
  END eFPGA_operand_b_o[6]
  PIN eFPGA_operand_b_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END eFPGA_operand_b_o[7]
  PIN eFPGA_operand_b_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END eFPGA_operand_b_o[8]
  PIN eFPGA_operand_b_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END eFPGA_operand_b_o[9]
  PIN eFPGA_operator_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END eFPGA_operator_o[0]
  PIN eFPGA_operator_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END eFPGA_operator_o[1]
  PIN eFPGA_result_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 97.280 1200.000 97.880 ;
    END
  END eFPGA_result_a_i[0]
  PIN eFPGA_result_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END eFPGA_result_a_i[10]
  PIN eFPGA_result_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 1196.000 450.250 1200.000 ;
    END
  END eFPGA_result_a_i[11]
  PIN eFPGA_result_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END eFPGA_result_a_i[12]
  PIN eFPGA_result_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END eFPGA_result_a_i[13]
  PIN eFPGA_result_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 1196.000 582.270 1200.000 ;
    END
  END eFPGA_result_a_i[14]
  PIN eFPGA_result_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 0.000 759.830 4.000 ;
    END
  END eFPGA_result_a_i[15]
  PIN eFPGA_result_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 639.920 1200.000 640.520 ;
    END
  END eFPGA_result_a_i[16]
  PIN eFPGA_result_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.200 4.000 671.800 ;
    END
  END eFPGA_result_a_i[17]
  PIN eFPGA_result_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 4.000 ;
    END
  END eFPGA_result_a_i[18]
  PIN eFPGA_result_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END eFPGA_result_a_i[19]
  PIN eFPGA_result_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 143.520 1200.000 144.120 ;
    END
  END eFPGA_result_a_i[1]
  PIN eFPGA_result_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END eFPGA_result_a_i[20]
  PIN eFPGA_result_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 858.880 1200.000 859.480 ;
    END
  END eFPGA_result_a_i[21]
  PIN eFPGA_result_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 905.120 1200.000 905.720 ;
    END
  END eFPGA_result_a_i[22]
  PIN eFPGA_result_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 1196.000 942.450 1200.000 ;
    END
  END eFPGA_result_a_i[23]
  PIN eFPGA_result_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 951.360 1200.000 951.960 ;
    END
  END eFPGA_result_a_i[24]
  PIN eFPGA_result_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1009.160 1200.000 1009.760 ;
    END
  END eFPGA_result_a_i[25]
  PIN eFPGA_result_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1032.280 1200.000 1032.880 ;
    END
  END eFPGA_result_a_i[26]
  PIN eFPGA_result_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 0.000 1056.990 4.000 ;
    END
  END eFPGA_result_a_i[27]
  PIN eFPGA_result_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1127.480 4.000 1128.080 ;
    END
  END eFPGA_result_a_i[28]
  PIN eFPGA_result_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1136.320 1200.000 1136.920 ;
    END
  END eFPGA_result_a_i[29]
  PIN eFPGA_result_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END eFPGA_result_a_i[2]
  PIN eFPGA_result_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 1196.000 1110.350 1200.000 ;
    END
  END eFPGA_result_a_i[30]
  PIN eFPGA_result_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.910 1196.000 1158.190 1200.000 ;
    END
  END eFPGA_result_a_i[31]
  PIN eFPGA_result_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 236.000 1200.000 236.600 ;
    END
  END eFPGA_result_a_i[3]
  PIN eFPGA_result_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 293.800 1200.000 294.400 ;
    END
  END eFPGA_result_a_i[4]
  PIN eFPGA_result_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END eFPGA_result_a_i[5]
  PIN eFPGA_result_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 1196.000 342.150 1200.000 ;
    END
  END eFPGA_result_a_i[6]
  PIN eFPGA_result_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 420.280 1200.000 420.880 ;
    END
  END eFPGA_result_a_i[7]
  PIN eFPGA_result_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END eFPGA_result_a_i[8]
  PIN eFPGA_result_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 478.080 1200.000 478.680 ;
    END
  END eFPGA_result_a_i[9]
  PIN eFPGA_result_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 1196.000 66.150 1200.000 ;
    END
  END eFPGA_result_b_i[0]
  PIN eFPGA_result_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END eFPGA_result_b_i[10]
  PIN eFPGA_result_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 559.000 1200.000 559.600 ;
    END
  END eFPGA_result_b_i[11]
  PIN eFPGA_result_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 475.360 4.000 475.960 ;
    END
  END eFPGA_result_b_i[12]
  PIN eFPGA_result_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END eFPGA_result_b_i[13]
  PIN eFPGA_result_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 1196.000 594.230 1200.000 ;
    END
  END eFPGA_result_b_i[14]
  PIN eFPGA_result_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1196.000 654.030 1200.000 ;
    END
  END eFPGA_result_b_i[15]
  PIN eFPGA_result_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 651.480 1200.000 652.080 ;
    END
  END eFPGA_result_b_i[16]
  PIN eFPGA_result_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 720.840 1200.000 721.440 ;
    END
  END eFPGA_result_b_i[17]
  PIN eFPGA_result_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 1196.000 738.210 1200.000 ;
    END
  END eFPGA_result_b_i[18]
  PIN eFPGA_result_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 1196.000 774.090 1200.000 ;
    END
  END eFPGA_result_b_i[19]
  PIN eFPGA_result_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END eFPGA_result_b_i[1]
  PIN eFPGA_result_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 801.760 1200.000 802.360 ;
    END
  END eFPGA_result_b_i[20]
  PIN eFPGA_result_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.760 4.000 802.360 ;
    END
  END eFPGA_result_b_i[21]
  PIN eFPGA_result_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.120 4.000 854.720 ;
    END
  END eFPGA_result_b_i[22]
  PIN eFPGA_result_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.880 4.000 893.480 ;
    END
  END eFPGA_result_b_i[23]
  PIN eFPGA_result_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 962.920 1200.000 963.520 ;
    END
  END eFPGA_result_b_i[24]
  PIN eFPGA_result_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 0.000 988.450 4.000 ;
    END
  END eFPGA_result_b_i[25]
  PIN eFPGA_result_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 1196.000 990.290 1200.000 ;
    END
  END eFPGA_result_b_i[26]
  PIN eFPGA_result_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1078.520 1200.000 1079.120 ;
    END
  END eFPGA_result_b_i[27]
  PIN eFPGA_result_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1113.200 1200.000 1113.800 ;
    END
  END eFPGA_result_b_i[28]
  PIN eFPGA_result_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1147.880 1200.000 1148.480 ;
    END
  END eFPGA_result_b_i[29]
  PIN eFPGA_result_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1196.000 174.250 1200.000 ;
    END
  END eFPGA_result_b_i[2]
  PIN eFPGA_result_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.030 1196.000 1122.310 1200.000 ;
    END
  END eFPGA_result_b_i[30]
  PIN eFPGA_result_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1192.760 4.000 1193.360 ;
    END
  END eFPGA_result_b_i[31]
  PIN eFPGA_result_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END eFPGA_result_b_i[3]
  PIN eFPGA_result_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 4.000 ;
    END
  END eFPGA_result_b_i[4]
  PIN eFPGA_result_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END eFPGA_result_b_i[5]
  PIN eFPGA_result_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 1196.000 354.110 1200.000 ;
    END
  END eFPGA_result_b_i[6]
  PIN eFPGA_result_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 1196.000 366.070 1200.000 ;
    END
  END eFPGA_result_b_i[7]
  PIN eFPGA_result_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 4.000 ;
    END
  END eFPGA_result_b_i[8]
  PIN eFPGA_result_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 489.640 1200.000 490.240 ;
    END
  END eFPGA_result_b_i[9]
  PIN eFPGA_result_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 108.840 1200.000 109.440 ;
    END
  END eFPGA_result_c_i[0]
  PIN eFPGA_result_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END eFPGA_result_c_i[10]
  PIN eFPGA_result_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END eFPGA_result_c_i[11]
  PIN eFPGA_result_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 0.000 725.790 4.000 ;
    END
  END eFPGA_result_c_i[12]
  PIN eFPGA_result_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 1196.000 522.010 1200.000 ;
    END
  END eFPGA_result_c_i[13]
  PIN eFPGA_result_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.080 4.000 580.680 ;
    END
  END eFPGA_result_c_i[14]
  PIN eFPGA_result_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 4.000 606.520 ;
    END
  END eFPGA_result_c_i[15]
  PIN eFPGA_result_c_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END eFPGA_result_c_i[16]
  PIN eFPGA_result_c_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 4.000 ;
    END
  END eFPGA_result_c_i[17]
  PIN eFPGA_result_c_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 0.000 839.870 4.000 ;
    END
  END eFPGA_result_c_i[18]
  PIN eFPGA_result_c_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 0.000 874.370 4.000 ;
    END
  END eFPGA_result_c_i[19]
  PIN eFPGA_result_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 155.080 1200.000 155.680 ;
    END
  END eFPGA_result_c_i[1]
  PIN eFPGA_result_c_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 1196.000 810.430 1200.000 ;
    END
  END eFPGA_result_c_i[20]
  PIN eFPGA_result_c_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 870.440 1200.000 871.040 ;
    END
  END eFPGA_result_c_i[21]
  PIN eFPGA_result_c_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.910 1196.000 882.190 1200.000 ;
    END
  END eFPGA_result_c_i[22]
  PIN eFPGA_result_c_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 0.000 931.410 4.000 ;
    END
  END eFPGA_result_c_i[23]
  PIN eFPGA_result_c_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 0.000 954.410 4.000 ;
    END
  END eFPGA_result_c_i[24]
  PIN eFPGA_result_c_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 997.600 4.000 998.200 ;
    END
  END eFPGA_result_c_i[25]
  PIN eFPGA_result_c_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END eFPGA_result_c_i[26]
  PIN eFPGA_result_c_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 1196.000 1014.210 1200.000 ;
    END
  END eFPGA_result_c_i[27]
  PIN eFPGA_result_c_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 0.000 1079.990 4.000 ;
    END
  END eFPGA_result_c_i[28]
  PIN eFPGA_result_c_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END eFPGA_result_c_i[29]
  PIN eFPGA_result_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END eFPGA_result_c_i[2]
  PIN eFPGA_result_c_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1159.440 1200.000 1160.040 ;
    END
  END eFPGA_result_c_i[30]
  PIN eFPGA_result_c_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 1196.000 1170.150 1200.000 ;
    END
  END eFPGA_result_c_i[31]
  PIN eFPGA_result_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 1196.000 210.130 1200.000 ;
    END
  END eFPGA_result_c_i[3]
  PIN eFPGA_result_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 305.360 1200.000 305.960 ;
    END
  END eFPGA_result_c_i[4]
  PIN eFPGA_result_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END eFPGA_result_c_i[5]
  PIN eFPGA_result_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 363.160 1200.000 363.760 ;
    END
  END eFPGA_result_c_i[6]
  PIN eFPGA_result_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 1196.000 378.030 1200.000 ;
    END
  END eFPGA_result_c_i[7]
  PIN eFPGA_result_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END eFPGA_result_c_i[8]
  PIN eFPGA_result_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 501.200 1200.000 501.800 ;
    END
  END eFPGA_result_c_i[9]
  PIN eFPGA_write_strobe_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END eFPGA_write_strobe_o
  PIN ext_perf_counters_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END ext_perf_counters_i
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 39.480 1200.000 40.080 ;
    END
  END fetch_enable_i
  PIN instr_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 120.400 1200.000 121.000 ;
    END
  END instr_addr_o[0]
  PIN instr_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 0.000 668.750 4.000 ;
    END
  END instr_addr_o[10]
  PIN instr_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END instr_addr_o[11]
  PIN instr_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 1196.000 474.170 1200.000 ;
    END
  END instr_addr_o[12]
  PIN instr_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 1196.000 533.970 1200.000 ;
    END
  END instr_addr_o[13]
  PIN instr_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END instr_addr_o[14]
  PIN instr_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 1196.000 665.990 1200.000 ;
    END
  END instr_addr_o[15]
  PIN instr_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 645.360 4.000 645.960 ;
    END
  END instr_addr_o[16]
  PIN instr_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 732.400 1200.000 733.000 ;
    END
  END instr_addr_o[17]
  PIN instr_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 1196.000 750.170 1200.000 ;
    END
  END instr_addr_o[18]
  PIN instr_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 762.320 4.000 762.920 ;
    END
  END instr_addr_o[19]
  PIN instr_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END instr_addr_o[1]
  PIN instr_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END instr_addr_o[20]
  PIN instr_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 882.000 1200.000 882.600 ;
    END
  END instr_addr_o[21]
  PIN instr_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 1196.000 894.150 1200.000 ;
    END
  END instr_addr_o[22]
  PIN instr_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END instr_addr_o[23]
  PIN instr_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 974.480 1200.000 975.080 ;
    END
  END instr_addr_o[24]
  PIN instr_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.050 1196.000 978.330 1200.000 ;
    END
  END instr_addr_o[25]
  PIN instr_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.670 0.000 1022.950 4.000 ;
    END
  END instr_addr_o[26]
  PIN instr_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.210 0.000 1068.490 4.000 ;
    END
  END instr_addr_o[27]
  PIN instr_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 1196.000 1050.090 1200.000 ;
    END
  END instr_addr_o[28]
  PIN instr_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 1196.000 1086.430 1200.000 ;
    END
  END instr_addr_o[29]
  PIN instr_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END instr_addr_o[2]
  PIN instr_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.920 4.000 1167.520 ;
    END
  END instr_addr_o[30]
  PIN instr_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 1196.000 1182.110 1200.000 ;
    END
  END instr_addr_o[31]
  PIN instr_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END instr_addr_o[3]
  PIN instr_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 1196.000 234.050 1200.000 ;
    END
  END instr_addr_o[4]
  PIN instr_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 1196.000 294.310 1200.000 ;
    END
  END instr_addr_o[5]
  PIN instr_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 374.720 1200.000 375.320 ;
    END
  END instr_addr_o[6]
  PIN instr_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 1196.000 389.990 1200.000 ;
    END
  END instr_addr_o[7]
  PIN instr_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 0.000 531.210 4.000 ;
    END
  END instr_addr_o[8]
  PIN instr_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END instr_addr_o[9]
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 51.040 1200.000 51.640 ;
    END
  END instr_gnt_i
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END instr_rdata_i[0]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 1196.000 486.130 1200.000 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 4.000 567.080 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 1196.000 606.190 1200.000 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 663.040 1200.000 663.640 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 755.520 1200.000 756.120 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 778.640 1200.000 779.240 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.630 0.000 919.910 4.000 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 1196.000 846.310 1200.000 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 916.680 1200.000 917.280 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.720 4.000 919.320 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1020.720 1200.000 1021.320 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 0.000 1034.450 4.000 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.890 1196.000 1026.170 1200.000 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1124.760 1200.000 1125.360 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 4.000 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.790 1196.000 1194.070 1200.000 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 316.920 1200.000 317.520 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 1196.000 306.270 1200.000 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 386.280 1200.000 386.880 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 431.840 1200.000 432.440 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 454.960 1200.000 455.560 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 0.000 611.250 4.000 ;
    END
  END instr_rdata_i[9]
  PIN instr_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 62.600 1200.000 63.200 ;
    END
  END instr_req_o
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 1196.000 18.310 1200.000 ;
    END
  END instr_rvalid_i
  PIN irq_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END irq_ack_o
  PIN irq_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END irq_i
  PIN irq_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END irq_id_i[0]
  PIN irq_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END irq_id_i[1]
  PIN irq_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END irq_id_i[2]
  PIN irq_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END irq_id_i[3]
  PIN irq_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END irq_id_i[4]
  PIN irq_id_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END irq_id_o[0]
  PIN irq_id_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END irq_id_o[1]
  PIN irq_id_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END irq_id_o[2]
  PIN irq_id_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END irq_id_o[3]
  PIN irq_id_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END irq_id_o[4]
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 1196.000 30.270 1200.000 ;
    END
  END test_en_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 1188.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.040 10.640 147.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 10.640 247.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.040 10.640 297.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.040 10.640 347.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 10.640 397.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.040 10.640 447.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.040 10.640 497.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 10.640 547.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.040 10.640 597.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.040 10.640 647.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 10.640 697.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.040 10.640 747.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.040 10.640 797.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 10.640 847.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 896.040 10.640 897.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.040 10.640 947.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.040 10.640 997.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1046.040 10.640 1047.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.040 10.640 1097.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.040 10.640 1147.640 1188.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 8.585 1194.935 1188.725 ;
      LAYER met1 ;
        RECT 0.070 6.500 1194.995 1188.880 ;
      LAYER met2 ;
        RECT 0.100 1195.720 5.790 1196.530 ;
        RECT 6.630 1195.720 17.750 1196.530 ;
        RECT 18.590 1195.720 29.710 1196.530 ;
        RECT 30.550 1195.720 41.670 1196.530 ;
        RECT 42.510 1195.720 53.630 1196.530 ;
        RECT 54.470 1195.720 65.590 1196.530 ;
        RECT 66.430 1195.720 77.550 1196.530 ;
        RECT 78.390 1195.720 89.510 1196.530 ;
        RECT 90.350 1195.720 101.470 1196.530 ;
        RECT 102.310 1195.720 113.430 1196.530 ;
        RECT 114.270 1195.720 125.390 1196.530 ;
        RECT 126.230 1195.720 137.350 1196.530 ;
        RECT 138.190 1195.720 149.770 1196.530 ;
        RECT 150.610 1195.720 161.730 1196.530 ;
        RECT 162.570 1195.720 173.690 1196.530 ;
        RECT 174.530 1195.720 185.650 1196.530 ;
        RECT 186.490 1195.720 197.610 1196.530 ;
        RECT 198.450 1195.720 209.570 1196.530 ;
        RECT 210.410 1195.720 221.530 1196.530 ;
        RECT 222.370 1195.720 233.490 1196.530 ;
        RECT 234.330 1195.720 245.450 1196.530 ;
        RECT 246.290 1195.720 257.410 1196.530 ;
        RECT 258.250 1195.720 269.370 1196.530 ;
        RECT 270.210 1195.720 281.790 1196.530 ;
        RECT 282.630 1195.720 293.750 1196.530 ;
        RECT 294.590 1195.720 305.710 1196.530 ;
        RECT 306.550 1195.720 317.670 1196.530 ;
        RECT 318.510 1195.720 329.630 1196.530 ;
        RECT 330.470 1195.720 341.590 1196.530 ;
        RECT 342.430 1195.720 353.550 1196.530 ;
        RECT 354.390 1195.720 365.510 1196.530 ;
        RECT 366.350 1195.720 377.470 1196.530 ;
        RECT 378.310 1195.720 389.430 1196.530 ;
        RECT 390.270 1195.720 401.390 1196.530 ;
        RECT 402.230 1195.720 413.810 1196.530 ;
        RECT 414.650 1195.720 425.770 1196.530 ;
        RECT 426.610 1195.720 437.730 1196.530 ;
        RECT 438.570 1195.720 449.690 1196.530 ;
        RECT 450.530 1195.720 461.650 1196.530 ;
        RECT 462.490 1195.720 473.610 1196.530 ;
        RECT 474.450 1195.720 485.570 1196.530 ;
        RECT 486.410 1195.720 497.530 1196.530 ;
        RECT 498.370 1195.720 509.490 1196.530 ;
        RECT 510.330 1195.720 521.450 1196.530 ;
        RECT 522.290 1195.720 533.410 1196.530 ;
        RECT 534.250 1195.720 545.830 1196.530 ;
        RECT 546.670 1195.720 557.790 1196.530 ;
        RECT 558.630 1195.720 569.750 1196.530 ;
        RECT 570.590 1195.720 581.710 1196.530 ;
        RECT 582.550 1195.720 593.670 1196.530 ;
        RECT 594.510 1195.720 605.630 1196.530 ;
        RECT 606.470 1195.720 617.590 1196.530 ;
        RECT 618.430 1195.720 629.550 1196.530 ;
        RECT 630.390 1195.720 641.510 1196.530 ;
        RECT 642.350 1195.720 653.470 1196.530 ;
        RECT 654.310 1195.720 665.430 1196.530 ;
        RECT 666.270 1195.720 677.850 1196.530 ;
        RECT 678.690 1195.720 689.810 1196.530 ;
        RECT 690.650 1195.720 701.770 1196.530 ;
        RECT 702.610 1195.720 713.730 1196.530 ;
        RECT 714.570 1195.720 725.690 1196.530 ;
        RECT 726.530 1195.720 737.650 1196.530 ;
        RECT 738.490 1195.720 749.610 1196.530 ;
        RECT 750.450 1195.720 761.570 1196.530 ;
        RECT 762.410 1195.720 773.530 1196.530 ;
        RECT 774.370 1195.720 785.490 1196.530 ;
        RECT 786.330 1195.720 797.450 1196.530 ;
        RECT 798.290 1195.720 809.870 1196.530 ;
        RECT 810.710 1195.720 821.830 1196.530 ;
        RECT 822.670 1195.720 833.790 1196.530 ;
        RECT 834.630 1195.720 845.750 1196.530 ;
        RECT 846.590 1195.720 857.710 1196.530 ;
        RECT 858.550 1195.720 869.670 1196.530 ;
        RECT 870.510 1195.720 881.630 1196.530 ;
        RECT 882.470 1195.720 893.590 1196.530 ;
        RECT 894.430 1195.720 905.550 1196.530 ;
        RECT 906.390 1195.720 917.510 1196.530 ;
        RECT 918.350 1195.720 929.470 1196.530 ;
        RECT 930.310 1195.720 941.890 1196.530 ;
        RECT 942.730 1195.720 953.850 1196.530 ;
        RECT 954.690 1195.720 965.810 1196.530 ;
        RECT 966.650 1195.720 977.770 1196.530 ;
        RECT 978.610 1195.720 989.730 1196.530 ;
        RECT 990.570 1195.720 1001.690 1196.530 ;
        RECT 1002.530 1195.720 1013.650 1196.530 ;
        RECT 1014.490 1195.720 1025.610 1196.530 ;
        RECT 1026.450 1195.720 1037.570 1196.530 ;
        RECT 1038.410 1195.720 1049.530 1196.530 ;
        RECT 1050.370 1195.720 1061.490 1196.530 ;
        RECT 1062.330 1195.720 1073.910 1196.530 ;
        RECT 1074.750 1195.720 1085.870 1196.530 ;
        RECT 1086.710 1195.720 1097.830 1196.530 ;
        RECT 1098.670 1195.720 1109.790 1196.530 ;
        RECT 1110.630 1195.720 1121.750 1196.530 ;
        RECT 1122.590 1195.720 1133.710 1196.530 ;
        RECT 1134.550 1195.720 1145.670 1196.530 ;
        RECT 1146.510 1195.720 1157.630 1196.530 ;
        RECT 1158.470 1195.720 1169.590 1196.530 ;
        RECT 1170.430 1195.720 1181.550 1196.530 ;
        RECT 1182.390 1195.720 1193.510 1196.530 ;
        RECT 1194.350 1195.720 1194.520 1196.530 ;
        RECT 0.100 4.280 1194.520 1195.720 ;
        RECT 0.100 3.670 5.330 4.280 ;
        RECT 6.170 3.670 16.370 4.280 ;
        RECT 17.210 3.670 27.870 4.280 ;
        RECT 28.710 3.670 39.370 4.280 ;
        RECT 40.210 3.670 50.870 4.280 ;
        RECT 51.710 3.670 62.370 4.280 ;
        RECT 63.210 3.670 73.870 4.280 ;
        RECT 74.710 3.670 84.910 4.280 ;
        RECT 85.750 3.670 96.410 4.280 ;
        RECT 97.250 3.670 107.910 4.280 ;
        RECT 108.750 3.670 119.410 4.280 ;
        RECT 120.250 3.670 130.910 4.280 ;
        RECT 131.750 3.670 142.410 4.280 ;
        RECT 143.250 3.670 153.910 4.280 ;
        RECT 154.750 3.670 164.950 4.280 ;
        RECT 165.790 3.670 176.450 4.280 ;
        RECT 177.290 3.670 187.950 4.280 ;
        RECT 188.790 3.670 199.450 4.280 ;
        RECT 200.290 3.670 210.950 4.280 ;
        RECT 211.790 3.670 222.450 4.280 ;
        RECT 223.290 3.670 233.490 4.280 ;
        RECT 234.330 3.670 244.990 4.280 ;
        RECT 245.830 3.670 256.490 4.280 ;
        RECT 257.330 3.670 267.990 4.280 ;
        RECT 268.830 3.670 279.490 4.280 ;
        RECT 280.330 3.670 290.990 4.280 ;
        RECT 291.830 3.670 302.490 4.280 ;
        RECT 303.330 3.670 313.530 4.280 ;
        RECT 314.370 3.670 325.030 4.280 ;
        RECT 325.870 3.670 336.530 4.280 ;
        RECT 337.370 3.670 348.030 4.280 ;
        RECT 348.870 3.670 359.530 4.280 ;
        RECT 360.370 3.670 371.030 4.280 ;
        RECT 371.870 3.670 382.070 4.280 ;
        RECT 382.910 3.670 393.570 4.280 ;
        RECT 394.410 3.670 405.070 4.280 ;
        RECT 405.910 3.670 416.570 4.280 ;
        RECT 417.410 3.670 428.070 4.280 ;
        RECT 428.910 3.670 439.570 4.280 ;
        RECT 440.410 3.670 451.070 4.280 ;
        RECT 451.910 3.670 462.110 4.280 ;
        RECT 462.950 3.670 473.610 4.280 ;
        RECT 474.450 3.670 485.110 4.280 ;
        RECT 485.950 3.670 496.610 4.280 ;
        RECT 497.450 3.670 508.110 4.280 ;
        RECT 508.950 3.670 519.610 4.280 ;
        RECT 520.450 3.670 530.650 4.280 ;
        RECT 531.490 3.670 542.150 4.280 ;
        RECT 542.990 3.670 553.650 4.280 ;
        RECT 554.490 3.670 565.150 4.280 ;
        RECT 565.990 3.670 576.650 4.280 ;
        RECT 577.490 3.670 588.150 4.280 ;
        RECT 588.990 3.670 599.650 4.280 ;
        RECT 600.490 3.670 610.690 4.280 ;
        RECT 611.530 3.670 622.190 4.280 ;
        RECT 623.030 3.670 633.690 4.280 ;
        RECT 634.530 3.670 645.190 4.280 ;
        RECT 646.030 3.670 656.690 4.280 ;
        RECT 657.530 3.670 668.190 4.280 ;
        RECT 669.030 3.670 679.690 4.280 ;
        RECT 680.530 3.670 690.730 4.280 ;
        RECT 691.570 3.670 702.230 4.280 ;
        RECT 703.070 3.670 713.730 4.280 ;
        RECT 714.570 3.670 725.230 4.280 ;
        RECT 726.070 3.670 736.730 4.280 ;
        RECT 737.570 3.670 748.230 4.280 ;
        RECT 749.070 3.670 759.270 4.280 ;
        RECT 760.110 3.670 770.770 4.280 ;
        RECT 771.610 3.670 782.270 4.280 ;
        RECT 783.110 3.670 793.770 4.280 ;
        RECT 794.610 3.670 805.270 4.280 ;
        RECT 806.110 3.670 816.770 4.280 ;
        RECT 817.610 3.670 828.270 4.280 ;
        RECT 829.110 3.670 839.310 4.280 ;
        RECT 840.150 3.670 850.810 4.280 ;
        RECT 851.650 3.670 862.310 4.280 ;
        RECT 863.150 3.670 873.810 4.280 ;
        RECT 874.650 3.670 885.310 4.280 ;
        RECT 886.150 3.670 896.810 4.280 ;
        RECT 897.650 3.670 907.850 4.280 ;
        RECT 908.690 3.670 919.350 4.280 ;
        RECT 920.190 3.670 930.850 4.280 ;
        RECT 931.690 3.670 942.350 4.280 ;
        RECT 943.190 3.670 953.850 4.280 ;
        RECT 954.690 3.670 965.350 4.280 ;
        RECT 966.190 3.670 976.850 4.280 ;
        RECT 977.690 3.670 987.890 4.280 ;
        RECT 988.730 3.670 999.390 4.280 ;
        RECT 1000.230 3.670 1010.890 4.280 ;
        RECT 1011.730 3.670 1022.390 4.280 ;
        RECT 1023.230 3.670 1033.890 4.280 ;
        RECT 1034.730 3.670 1045.390 4.280 ;
        RECT 1046.230 3.670 1056.430 4.280 ;
        RECT 1057.270 3.670 1067.930 4.280 ;
        RECT 1068.770 3.670 1079.430 4.280 ;
        RECT 1080.270 3.670 1090.930 4.280 ;
        RECT 1091.770 3.670 1102.430 4.280 ;
        RECT 1103.270 3.670 1113.930 4.280 ;
        RECT 1114.770 3.670 1125.430 4.280 ;
        RECT 1126.270 3.670 1136.470 4.280 ;
        RECT 1137.310 3.670 1147.970 4.280 ;
        RECT 1148.810 3.670 1159.470 4.280 ;
        RECT 1160.310 3.670 1170.970 4.280 ;
        RECT 1171.810 3.670 1182.470 4.280 ;
        RECT 1183.310 3.670 1193.970 4.280 ;
      LAYER met3 ;
        RECT 4.000 1193.760 1195.600 1194.585 ;
        RECT 4.400 1193.720 1195.600 1193.760 ;
        RECT 4.400 1192.360 1196.610 1193.720 ;
        RECT 4.000 1183.560 1196.610 1192.360 ;
        RECT 4.000 1182.160 1195.600 1183.560 ;
        RECT 4.000 1180.840 1196.610 1182.160 ;
        RECT 4.400 1179.440 1196.610 1180.840 ;
        RECT 4.000 1172.000 1196.610 1179.440 ;
        RECT 4.000 1170.600 1195.600 1172.000 ;
        RECT 4.000 1167.920 1196.610 1170.600 ;
        RECT 4.400 1166.520 1196.610 1167.920 ;
        RECT 4.000 1160.440 1196.610 1166.520 ;
        RECT 4.000 1159.040 1195.600 1160.440 ;
        RECT 4.000 1155.000 1196.610 1159.040 ;
        RECT 4.400 1153.600 1196.610 1155.000 ;
        RECT 4.000 1148.880 1196.610 1153.600 ;
        RECT 4.000 1147.480 1195.600 1148.880 ;
        RECT 4.000 1142.080 1196.610 1147.480 ;
        RECT 4.400 1140.680 1196.610 1142.080 ;
        RECT 4.000 1137.320 1196.610 1140.680 ;
        RECT 4.000 1135.920 1195.600 1137.320 ;
        RECT 4.000 1128.480 1196.610 1135.920 ;
        RECT 4.400 1127.080 1196.610 1128.480 ;
        RECT 4.000 1125.760 1196.610 1127.080 ;
        RECT 4.000 1124.360 1195.600 1125.760 ;
        RECT 4.000 1115.560 1196.610 1124.360 ;
        RECT 4.400 1114.200 1196.610 1115.560 ;
        RECT 4.400 1114.160 1195.600 1114.200 ;
        RECT 4.000 1112.800 1195.600 1114.160 ;
        RECT 4.000 1102.640 1196.610 1112.800 ;
        RECT 4.400 1101.240 1195.600 1102.640 ;
        RECT 4.000 1091.080 1196.610 1101.240 ;
        RECT 4.000 1089.720 1195.600 1091.080 ;
        RECT 4.400 1089.680 1195.600 1089.720 ;
        RECT 4.400 1088.320 1196.610 1089.680 ;
        RECT 4.000 1079.520 1196.610 1088.320 ;
        RECT 4.000 1078.120 1195.600 1079.520 ;
        RECT 4.000 1076.800 1196.610 1078.120 ;
        RECT 4.400 1075.400 1196.610 1076.800 ;
        RECT 4.000 1067.960 1196.610 1075.400 ;
        RECT 4.000 1066.560 1195.600 1067.960 ;
        RECT 4.000 1063.200 1196.610 1066.560 ;
        RECT 4.400 1061.800 1196.610 1063.200 ;
        RECT 4.000 1056.400 1196.610 1061.800 ;
        RECT 4.000 1055.000 1195.600 1056.400 ;
        RECT 4.000 1050.280 1196.610 1055.000 ;
        RECT 4.400 1048.880 1196.610 1050.280 ;
        RECT 4.000 1044.840 1196.610 1048.880 ;
        RECT 4.000 1043.440 1195.600 1044.840 ;
        RECT 4.000 1037.360 1196.610 1043.440 ;
        RECT 4.400 1035.960 1196.610 1037.360 ;
        RECT 4.000 1033.280 1196.610 1035.960 ;
        RECT 4.000 1031.880 1195.600 1033.280 ;
        RECT 4.000 1024.440 1196.610 1031.880 ;
        RECT 4.400 1023.040 1196.610 1024.440 ;
        RECT 4.000 1021.720 1196.610 1023.040 ;
        RECT 4.000 1020.320 1195.600 1021.720 ;
        RECT 4.000 1011.520 1196.610 1020.320 ;
        RECT 4.400 1010.160 1196.610 1011.520 ;
        RECT 4.400 1010.120 1195.600 1010.160 ;
        RECT 4.000 1008.760 1195.600 1010.120 ;
        RECT 4.000 998.600 1196.610 1008.760 ;
        RECT 4.400 997.200 1195.600 998.600 ;
        RECT 4.000 987.040 1196.610 997.200 ;
        RECT 4.000 985.640 1195.600 987.040 ;
        RECT 4.000 985.000 1196.610 985.640 ;
        RECT 4.400 983.600 1196.610 985.000 ;
        RECT 4.000 975.480 1196.610 983.600 ;
        RECT 4.000 974.080 1195.600 975.480 ;
        RECT 4.000 972.080 1196.610 974.080 ;
        RECT 4.400 970.680 1196.610 972.080 ;
        RECT 4.000 963.920 1196.610 970.680 ;
        RECT 4.000 962.520 1195.600 963.920 ;
        RECT 4.000 959.160 1196.610 962.520 ;
        RECT 4.400 957.760 1196.610 959.160 ;
        RECT 4.000 952.360 1196.610 957.760 ;
        RECT 4.000 950.960 1195.600 952.360 ;
        RECT 4.000 946.240 1196.610 950.960 ;
        RECT 4.400 944.840 1196.610 946.240 ;
        RECT 4.000 940.800 1196.610 944.840 ;
        RECT 4.000 939.400 1195.600 940.800 ;
        RECT 4.000 933.320 1196.610 939.400 ;
        RECT 4.400 931.920 1196.610 933.320 ;
        RECT 4.000 929.240 1196.610 931.920 ;
        RECT 4.000 927.840 1195.600 929.240 ;
        RECT 4.000 919.720 1196.610 927.840 ;
        RECT 4.400 918.320 1196.610 919.720 ;
        RECT 4.000 917.680 1196.610 918.320 ;
        RECT 4.000 916.280 1195.600 917.680 ;
        RECT 4.000 906.800 1196.610 916.280 ;
        RECT 4.400 906.120 1196.610 906.800 ;
        RECT 4.400 905.400 1195.600 906.120 ;
        RECT 4.000 904.720 1195.600 905.400 ;
        RECT 4.000 894.560 1196.610 904.720 ;
        RECT 4.000 893.880 1195.600 894.560 ;
        RECT 4.400 893.160 1195.600 893.880 ;
        RECT 4.400 892.480 1196.610 893.160 ;
        RECT 4.000 883.000 1196.610 892.480 ;
        RECT 4.000 881.600 1195.600 883.000 ;
        RECT 4.000 880.960 1196.610 881.600 ;
        RECT 4.400 879.560 1196.610 880.960 ;
        RECT 4.000 871.440 1196.610 879.560 ;
        RECT 4.000 870.040 1195.600 871.440 ;
        RECT 4.000 868.040 1196.610 870.040 ;
        RECT 4.400 866.640 1196.610 868.040 ;
        RECT 4.000 859.880 1196.610 866.640 ;
        RECT 4.000 858.480 1195.600 859.880 ;
        RECT 4.000 855.120 1196.610 858.480 ;
        RECT 4.400 853.720 1196.610 855.120 ;
        RECT 4.000 848.320 1196.610 853.720 ;
        RECT 4.000 846.920 1195.600 848.320 ;
        RECT 4.000 841.520 1196.610 846.920 ;
        RECT 4.400 840.120 1196.610 841.520 ;
        RECT 4.000 836.760 1196.610 840.120 ;
        RECT 4.000 835.360 1195.600 836.760 ;
        RECT 4.000 828.600 1196.610 835.360 ;
        RECT 4.400 827.200 1196.610 828.600 ;
        RECT 4.000 825.200 1196.610 827.200 ;
        RECT 4.000 823.800 1195.600 825.200 ;
        RECT 4.000 815.680 1196.610 823.800 ;
        RECT 4.400 814.280 1196.610 815.680 ;
        RECT 4.000 813.640 1196.610 814.280 ;
        RECT 4.000 812.240 1195.600 813.640 ;
        RECT 4.000 802.760 1196.610 812.240 ;
        RECT 4.400 801.360 1195.600 802.760 ;
        RECT 4.000 791.200 1196.610 801.360 ;
        RECT 4.000 789.840 1195.600 791.200 ;
        RECT 4.400 789.800 1195.600 789.840 ;
        RECT 4.400 788.440 1196.610 789.800 ;
        RECT 4.000 779.640 1196.610 788.440 ;
        RECT 4.000 778.240 1195.600 779.640 ;
        RECT 4.000 776.240 1196.610 778.240 ;
        RECT 4.400 774.840 1196.610 776.240 ;
        RECT 4.000 768.080 1196.610 774.840 ;
        RECT 4.000 766.680 1195.600 768.080 ;
        RECT 4.000 763.320 1196.610 766.680 ;
        RECT 4.400 761.920 1196.610 763.320 ;
        RECT 4.000 756.520 1196.610 761.920 ;
        RECT 4.000 755.120 1195.600 756.520 ;
        RECT 4.000 750.400 1196.610 755.120 ;
        RECT 4.400 749.000 1196.610 750.400 ;
        RECT 4.000 744.960 1196.610 749.000 ;
        RECT 4.000 743.560 1195.600 744.960 ;
        RECT 4.000 737.480 1196.610 743.560 ;
        RECT 4.400 736.080 1196.610 737.480 ;
        RECT 4.000 733.400 1196.610 736.080 ;
        RECT 4.000 732.000 1195.600 733.400 ;
        RECT 4.000 724.560 1196.610 732.000 ;
        RECT 4.400 723.160 1196.610 724.560 ;
        RECT 4.000 721.840 1196.610 723.160 ;
        RECT 4.000 720.440 1195.600 721.840 ;
        RECT 4.000 710.960 1196.610 720.440 ;
        RECT 4.400 710.280 1196.610 710.960 ;
        RECT 4.400 709.560 1195.600 710.280 ;
        RECT 4.000 708.880 1195.600 709.560 ;
        RECT 4.000 698.720 1196.610 708.880 ;
        RECT 4.000 698.040 1195.600 698.720 ;
        RECT 4.400 697.320 1195.600 698.040 ;
        RECT 4.400 696.640 1196.610 697.320 ;
        RECT 4.000 687.160 1196.610 696.640 ;
        RECT 4.000 685.760 1195.600 687.160 ;
        RECT 4.000 685.120 1196.610 685.760 ;
        RECT 4.400 683.720 1196.610 685.120 ;
        RECT 4.000 675.600 1196.610 683.720 ;
        RECT 4.000 674.200 1195.600 675.600 ;
        RECT 4.000 672.200 1196.610 674.200 ;
        RECT 4.400 670.800 1196.610 672.200 ;
        RECT 4.000 664.040 1196.610 670.800 ;
        RECT 4.000 662.640 1195.600 664.040 ;
        RECT 4.000 659.280 1196.610 662.640 ;
        RECT 4.400 657.880 1196.610 659.280 ;
        RECT 4.000 652.480 1196.610 657.880 ;
        RECT 4.000 651.080 1195.600 652.480 ;
        RECT 4.000 646.360 1196.610 651.080 ;
        RECT 4.400 644.960 1196.610 646.360 ;
        RECT 4.000 640.920 1196.610 644.960 ;
        RECT 4.000 639.520 1195.600 640.920 ;
        RECT 4.000 632.760 1196.610 639.520 ;
        RECT 4.400 631.360 1196.610 632.760 ;
        RECT 4.000 629.360 1196.610 631.360 ;
        RECT 4.000 627.960 1195.600 629.360 ;
        RECT 4.000 619.840 1196.610 627.960 ;
        RECT 4.400 618.440 1196.610 619.840 ;
        RECT 4.000 617.800 1196.610 618.440 ;
        RECT 4.000 616.400 1195.600 617.800 ;
        RECT 4.000 606.920 1196.610 616.400 ;
        RECT 4.400 606.240 1196.610 606.920 ;
        RECT 4.400 605.520 1195.600 606.240 ;
        RECT 4.000 604.840 1195.600 605.520 ;
        RECT 4.000 594.680 1196.610 604.840 ;
        RECT 4.000 594.000 1195.600 594.680 ;
        RECT 4.400 593.280 1195.600 594.000 ;
        RECT 4.400 592.600 1196.610 593.280 ;
        RECT 4.000 583.120 1196.610 592.600 ;
        RECT 4.000 581.720 1195.600 583.120 ;
        RECT 4.000 581.080 1196.610 581.720 ;
        RECT 4.400 579.680 1196.610 581.080 ;
        RECT 4.000 571.560 1196.610 579.680 ;
        RECT 4.000 570.160 1195.600 571.560 ;
        RECT 4.000 567.480 1196.610 570.160 ;
        RECT 4.400 566.080 1196.610 567.480 ;
        RECT 4.000 560.000 1196.610 566.080 ;
        RECT 4.000 558.600 1195.600 560.000 ;
        RECT 4.000 554.560 1196.610 558.600 ;
        RECT 4.400 553.160 1196.610 554.560 ;
        RECT 4.000 548.440 1196.610 553.160 ;
        RECT 4.000 547.040 1195.600 548.440 ;
        RECT 4.000 541.640 1196.610 547.040 ;
        RECT 4.400 540.240 1196.610 541.640 ;
        RECT 4.000 536.880 1196.610 540.240 ;
        RECT 4.000 535.480 1195.600 536.880 ;
        RECT 4.000 528.720 1196.610 535.480 ;
        RECT 4.400 527.320 1196.610 528.720 ;
        RECT 4.000 525.320 1196.610 527.320 ;
        RECT 4.000 523.920 1195.600 525.320 ;
        RECT 4.000 515.800 1196.610 523.920 ;
        RECT 4.400 514.400 1196.610 515.800 ;
        RECT 4.000 513.760 1196.610 514.400 ;
        RECT 4.000 512.360 1195.600 513.760 ;
        RECT 4.000 502.880 1196.610 512.360 ;
        RECT 4.400 502.200 1196.610 502.880 ;
        RECT 4.400 501.480 1195.600 502.200 ;
        RECT 4.000 500.800 1195.600 501.480 ;
        RECT 4.000 490.640 1196.610 500.800 ;
        RECT 4.000 489.280 1195.600 490.640 ;
        RECT 4.400 489.240 1195.600 489.280 ;
        RECT 4.400 487.880 1196.610 489.240 ;
        RECT 4.000 479.080 1196.610 487.880 ;
        RECT 4.000 477.680 1195.600 479.080 ;
        RECT 4.000 476.360 1196.610 477.680 ;
        RECT 4.400 474.960 1196.610 476.360 ;
        RECT 4.000 467.520 1196.610 474.960 ;
        RECT 4.000 466.120 1195.600 467.520 ;
        RECT 4.000 463.440 1196.610 466.120 ;
        RECT 4.400 462.040 1196.610 463.440 ;
        RECT 4.000 455.960 1196.610 462.040 ;
        RECT 4.000 454.560 1195.600 455.960 ;
        RECT 4.000 450.520 1196.610 454.560 ;
        RECT 4.400 449.120 1196.610 450.520 ;
        RECT 4.000 444.400 1196.610 449.120 ;
        RECT 4.000 443.000 1195.600 444.400 ;
        RECT 4.000 437.600 1196.610 443.000 ;
        RECT 4.400 436.200 1196.610 437.600 ;
        RECT 4.000 432.840 1196.610 436.200 ;
        RECT 4.000 431.440 1195.600 432.840 ;
        RECT 4.000 424.000 1196.610 431.440 ;
        RECT 4.400 422.600 1196.610 424.000 ;
        RECT 4.000 421.280 1196.610 422.600 ;
        RECT 4.000 419.880 1195.600 421.280 ;
        RECT 4.000 411.080 1196.610 419.880 ;
        RECT 4.400 409.720 1196.610 411.080 ;
        RECT 4.400 409.680 1195.600 409.720 ;
        RECT 4.000 408.320 1195.600 409.680 ;
        RECT 4.000 398.840 1196.610 408.320 ;
        RECT 4.000 398.160 1195.600 398.840 ;
        RECT 4.400 397.440 1195.600 398.160 ;
        RECT 4.400 396.760 1196.610 397.440 ;
        RECT 4.000 387.280 1196.610 396.760 ;
        RECT 4.000 385.880 1195.600 387.280 ;
        RECT 4.000 385.240 1196.610 385.880 ;
        RECT 4.400 383.840 1196.610 385.240 ;
        RECT 4.000 375.720 1196.610 383.840 ;
        RECT 4.000 374.320 1195.600 375.720 ;
        RECT 4.000 372.320 1196.610 374.320 ;
        RECT 4.400 370.920 1196.610 372.320 ;
        RECT 4.000 364.160 1196.610 370.920 ;
        RECT 4.000 362.760 1195.600 364.160 ;
        RECT 4.000 358.720 1196.610 362.760 ;
        RECT 4.400 357.320 1196.610 358.720 ;
        RECT 4.000 352.600 1196.610 357.320 ;
        RECT 4.000 351.200 1195.600 352.600 ;
        RECT 4.000 345.800 1196.610 351.200 ;
        RECT 4.400 344.400 1196.610 345.800 ;
        RECT 4.000 341.040 1196.610 344.400 ;
        RECT 4.000 339.640 1195.600 341.040 ;
        RECT 4.000 332.880 1196.610 339.640 ;
        RECT 4.400 331.480 1196.610 332.880 ;
        RECT 4.000 329.480 1196.610 331.480 ;
        RECT 4.000 328.080 1195.600 329.480 ;
        RECT 4.000 319.960 1196.610 328.080 ;
        RECT 4.400 318.560 1196.610 319.960 ;
        RECT 4.000 317.920 1196.610 318.560 ;
        RECT 4.000 316.520 1195.600 317.920 ;
        RECT 4.000 307.040 1196.610 316.520 ;
        RECT 4.400 306.360 1196.610 307.040 ;
        RECT 4.400 305.640 1195.600 306.360 ;
        RECT 4.000 304.960 1195.600 305.640 ;
        RECT 4.000 294.800 1196.610 304.960 ;
        RECT 4.000 294.120 1195.600 294.800 ;
        RECT 4.400 293.400 1195.600 294.120 ;
        RECT 4.400 292.720 1196.610 293.400 ;
        RECT 4.000 283.240 1196.610 292.720 ;
        RECT 4.000 281.840 1195.600 283.240 ;
        RECT 4.000 280.520 1196.610 281.840 ;
        RECT 4.400 279.120 1196.610 280.520 ;
        RECT 4.000 271.680 1196.610 279.120 ;
        RECT 4.000 270.280 1195.600 271.680 ;
        RECT 4.000 267.600 1196.610 270.280 ;
        RECT 4.400 266.200 1196.610 267.600 ;
        RECT 4.000 260.120 1196.610 266.200 ;
        RECT 4.000 258.720 1195.600 260.120 ;
        RECT 4.000 254.680 1196.610 258.720 ;
        RECT 4.400 253.280 1196.610 254.680 ;
        RECT 4.000 248.560 1196.610 253.280 ;
        RECT 4.000 247.160 1195.600 248.560 ;
        RECT 4.000 241.760 1196.610 247.160 ;
        RECT 4.400 240.360 1196.610 241.760 ;
        RECT 4.000 237.000 1196.610 240.360 ;
        RECT 4.000 235.600 1195.600 237.000 ;
        RECT 4.000 228.840 1196.610 235.600 ;
        RECT 4.400 227.440 1196.610 228.840 ;
        RECT 4.000 225.440 1196.610 227.440 ;
        RECT 4.000 224.040 1195.600 225.440 ;
        RECT 4.000 215.240 1196.610 224.040 ;
        RECT 4.400 213.880 1196.610 215.240 ;
        RECT 4.400 213.840 1195.600 213.880 ;
        RECT 4.000 212.480 1195.600 213.840 ;
        RECT 4.000 202.320 1196.610 212.480 ;
        RECT 4.400 200.920 1195.600 202.320 ;
        RECT 4.000 190.760 1196.610 200.920 ;
        RECT 4.000 189.400 1195.600 190.760 ;
        RECT 4.400 189.360 1195.600 189.400 ;
        RECT 4.400 188.000 1196.610 189.360 ;
        RECT 4.000 179.200 1196.610 188.000 ;
        RECT 4.000 177.800 1195.600 179.200 ;
        RECT 4.000 176.480 1196.610 177.800 ;
        RECT 4.400 175.080 1196.610 176.480 ;
        RECT 4.000 167.640 1196.610 175.080 ;
        RECT 4.000 166.240 1195.600 167.640 ;
        RECT 4.000 163.560 1196.610 166.240 ;
        RECT 4.400 162.160 1196.610 163.560 ;
        RECT 4.000 156.080 1196.610 162.160 ;
        RECT 4.000 154.680 1195.600 156.080 ;
        RECT 4.000 150.640 1196.610 154.680 ;
        RECT 4.400 149.240 1196.610 150.640 ;
        RECT 4.000 144.520 1196.610 149.240 ;
        RECT 4.000 143.120 1195.600 144.520 ;
        RECT 4.000 137.040 1196.610 143.120 ;
        RECT 4.400 135.640 1196.610 137.040 ;
        RECT 4.000 132.960 1196.610 135.640 ;
        RECT 4.000 131.560 1195.600 132.960 ;
        RECT 4.000 124.120 1196.610 131.560 ;
        RECT 4.400 122.720 1196.610 124.120 ;
        RECT 4.000 121.400 1196.610 122.720 ;
        RECT 4.000 120.000 1195.600 121.400 ;
        RECT 4.000 111.200 1196.610 120.000 ;
        RECT 4.400 109.840 1196.610 111.200 ;
        RECT 4.400 109.800 1195.600 109.840 ;
        RECT 4.000 108.440 1195.600 109.800 ;
        RECT 4.000 98.280 1196.610 108.440 ;
        RECT 4.400 96.880 1195.600 98.280 ;
        RECT 4.000 86.720 1196.610 96.880 ;
        RECT 4.000 85.360 1195.600 86.720 ;
        RECT 4.400 85.320 1195.600 85.360 ;
        RECT 4.400 83.960 1196.610 85.320 ;
        RECT 4.000 75.160 1196.610 83.960 ;
        RECT 4.000 73.760 1195.600 75.160 ;
        RECT 4.000 71.760 1196.610 73.760 ;
        RECT 4.400 70.360 1196.610 71.760 ;
        RECT 4.000 63.600 1196.610 70.360 ;
        RECT 4.000 62.200 1195.600 63.600 ;
        RECT 4.000 58.840 1196.610 62.200 ;
        RECT 4.400 57.440 1196.610 58.840 ;
        RECT 4.000 52.040 1196.610 57.440 ;
        RECT 4.000 50.640 1195.600 52.040 ;
        RECT 4.000 45.920 1196.610 50.640 ;
        RECT 4.400 44.520 1196.610 45.920 ;
        RECT 4.000 40.480 1196.610 44.520 ;
        RECT 4.000 39.080 1195.600 40.480 ;
        RECT 4.000 33.000 1196.610 39.080 ;
        RECT 4.400 31.600 1196.610 33.000 ;
        RECT 4.000 28.920 1196.610 31.600 ;
        RECT 4.000 27.520 1195.600 28.920 ;
        RECT 4.000 20.080 1196.610 27.520 ;
        RECT 4.400 18.680 1196.610 20.080 ;
        RECT 4.000 17.360 1196.610 18.680 ;
        RECT 4.000 15.960 1195.600 17.360 ;
        RECT 4.000 7.160 1196.610 15.960 ;
        RECT 4.400 6.480 1196.610 7.160 ;
        RECT 4.400 5.760 1195.600 6.480 ;
        RECT 4.000 5.615 1195.600 5.760 ;
      LAYER met4 ;
        RECT 177.855 127.335 195.640 1034.785 ;
        RECT 198.040 127.335 220.640 1034.785 ;
        RECT 223.040 127.335 245.640 1034.785 ;
        RECT 248.040 127.335 270.640 1034.785 ;
        RECT 273.040 127.335 295.640 1034.785 ;
        RECT 298.040 127.335 320.640 1034.785 ;
        RECT 323.040 127.335 345.640 1034.785 ;
        RECT 348.040 127.335 370.640 1034.785 ;
        RECT 373.040 127.335 395.640 1034.785 ;
        RECT 398.040 127.335 420.640 1034.785 ;
        RECT 423.040 127.335 445.640 1034.785 ;
        RECT 448.040 127.335 470.640 1034.785 ;
        RECT 473.040 127.335 495.640 1034.785 ;
        RECT 498.040 127.335 520.640 1034.785 ;
        RECT 523.040 127.335 545.640 1034.785 ;
        RECT 548.040 127.335 570.640 1034.785 ;
        RECT 573.040 127.335 595.640 1034.785 ;
        RECT 598.040 127.335 620.640 1034.785 ;
        RECT 623.040 127.335 645.640 1034.785 ;
        RECT 648.040 127.335 670.640 1034.785 ;
        RECT 673.040 127.335 695.640 1034.785 ;
        RECT 698.040 127.335 720.640 1034.785 ;
        RECT 723.040 127.335 745.640 1034.785 ;
        RECT 748.040 127.335 770.640 1034.785 ;
        RECT 773.040 127.335 795.640 1034.785 ;
        RECT 798.040 127.335 819.425 1034.785 ;
  END
END flexbex_ibex_core
END LIBRARY

