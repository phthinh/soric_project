VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ibex_top
  CLASS BLOCK ;
  FOREIGN ibex_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN alert_major_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 9.560 1200.000 10.160 ;
    END
  END alert_major_o
  PIN alert_minor_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 4.000 ;
    END
  END alert_minor_o
  PIN boot_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 29.280 1200.000 29.880 ;
    END
  END boot_addr_i[0]
  PIN boot_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END boot_addr_i[10]
  PIN boot_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END boot_addr_i[11]
  PIN boot_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.630 1196.000 1011.910 1200.000 ;
    END
  END boot_addr_i[12]
  PIN boot_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.110 0.000 1052.390 4.000 ;
    END
  END boot_addr_i[13]
  PIN boot_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 209.480 1200.000 210.080 ;
    END
  END boot_addr_i[14]
  PIN boot_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.230 0.000 1062.510 4.000 ;
    END
  END boot_addr_i[15]
  PIN boot_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 269.320 1200.000 269.920 ;
    END
  END boot_addr_i[16]
  PIN boot_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 1196.000 1026.630 1200.000 ;
    END
  END boot_addr_i[17]
  PIN boot_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.410 1196.000 1031.690 1200.000 ;
    END
  END boot_addr_i[18]
  PIN boot_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END boot_addr_i[19]
  PIN boot_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 69.400 1200.000 70.000 ;
    END
  END boot_addr_i[1]
  PIN boot_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 1196.000 1046.870 1200.000 ;
    END
  END boot_addr_i[20]
  PIN boot_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 1196.000 1051.930 1200.000 ;
    END
  END boot_addr_i[21]
  PIN boot_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 409.400 1200.000 410.000 ;
    END
  END boot_addr_i[22]
  PIN boot_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 449.520 1200.000 450.120 ;
    END
  END boot_addr_i[23]
  PIN boot_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 469.240 1200.000 469.840 ;
    END
  END boot_addr_i[24]
  PIN boot_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 1196.000 1072.170 1200.000 ;
    END
  END boot_addr_i[25]
  PIN boot_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 489.640 1200.000 490.240 ;
    END
  END boot_addr_i[26]
  PIN boot_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.730 1196.000 1097.010 1200.000 ;
    END
  END boot_addr_i[27]
  PIN boot_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END boot_addr_i[28]
  PIN boot_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.070 0.000 1087.350 4.000 ;
    END
  END boot_addr_i[29]
  PIN boot_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END boot_addr_i[2]
  PIN boot_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.130 0.000 1092.410 4.000 ;
    END
  END boot_addr_i[30]
  PIN boot_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END boot_addr_i[31]
  PIN boot_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END boot_addr_i[3]
  PIN boot_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END boot_addr_i[4]
  PIN boot_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 1196.000 966.370 1200.000 ;
    END
  END boot_addr_i[5]
  PIN boot_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 1196.000 976.490 1200.000 ;
    END
  END boot_addr_i[6]
  PIN boot_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 0.000 1032.610 4.000 ;
    END
  END boot_addr_i[7]
  PIN boot_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 129.240 1200.000 129.840 ;
    END
  END boot_addr_i[8]
  PIN boot_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 1196.000 996.730 1200.000 ;
    END
  END boot_addr_i[9]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 4.000 ;
    END
  END clk_i
  PIN core_sleep_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END core_sleep_o
  PIN crash_dump_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.370 0.000 997.650 4.000 ;
    END
  END crash_dump_o[0]
  PIN crash_dump_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1049.280 1200.000 1049.880 ;
    END
  END crash_dump_o[100]
  PIN crash_dump_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 1196.000 1172.450 1200.000 ;
    END
  END crash_dump_o[101]
  PIN crash_dump_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END crash_dump_o[102]
  PIN crash_dump_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 1196.000 1177.510 1200.000 ;
    END
  END crash_dump_o[103]
  PIN crash_dump_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.110 0.000 1167.390 4.000 ;
    END
  END crash_dump_o[104]
  PIN crash_dump_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1069.680 1200.000 1070.280 ;
    END
  END crash_dump_o[105]
  PIN crash_dump_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1052.680 4.000 1053.280 ;
    END
  END crash_dump_o[106]
  PIN crash_dump_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1079.200 4.000 1079.800 ;
    END
  END crash_dump_o[107]
  PIN crash_dump_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 0.000 1172.450 4.000 ;
    END
  END crash_dump_o[108]
  PIN crash_dump_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1106.400 4.000 1107.000 ;
    END
  END crash_dump_o[109]
  PIN crash_dump_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.570 1196.000 1006.850 1200.000 ;
    END
  END crash_dump_o[10]
  PIN crash_dump_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.290 1196.000 1182.570 1200.000 ;
    END
  END crash_dump_o[110]
  PIN crash_dump_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.350 1196.000 1187.630 1200.000 ;
    END
  END crash_dump_o[111]
  PIN crash_dump_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1089.400 1200.000 1090.000 ;
    END
  END crash_dump_o[112]
  PIN crash_dump_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.920 4.000 1133.520 ;
    END
  END crash_dump_o[113]
  PIN crash_dump_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 0.000 1177.510 4.000 ;
    END
  END crash_dump_o[114]
  PIN crash_dump_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1109.120 1200.000 1109.720 ;
    END
  END crash_dump_o[115]
  PIN crash_dump_o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1129.520 1200.000 1130.120 ;
    END
  END crash_dump_o[116]
  PIN crash_dump_o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1149.240 1200.000 1149.840 ;
    END
  END crash_dump_o[117]
  PIN crash_dump_o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.290 0.000 1182.570 4.000 ;
    END
  END crash_dump_o[118]
  PIN crash_dump_o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1169.640 1200.000 1170.240 ;
    END
  END crash_dump_o[119]
  PIN crash_dump_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 169.360 1200.000 169.960 ;
    END
  END crash_dump_o[11]
  PIN crash_dump_o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.410 1196.000 1192.690 1200.000 ;
    END
  END crash_dump_o[120]
  PIN crash_dump_o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.350 0.000 1187.630 4.000 ;
    END
  END crash_dump_o[121]
  PIN crash_dump_o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.410 0.000 1192.690 4.000 ;
    END
  END crash_dump_o[122]
  PIN crash_dump_o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.470 0.000 1197.750 4.000 ;
    END
  END crash_dump_o[123]
  PIN crash_dump_o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1189.360 1200.000 1189.960 ;
    END
  END crash_dump_o[124]
  PIN crash_dump_o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END crash_dump_o[125]
  PIN crash_dump_o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1185.960 4.000 1186.560 ;
    END
  END crash_dump_o[126]
  PIN crash_dump_o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.470 1196.000 1197.750 1200.000 ;
    END
  END crash_dump_o[127]
  PIN crash_dump_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 1196.000 1016.970 1200.000 ;
    END
  END crash_dump_o[12]
  PIN crash_dump_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 189.080 1200.000 189.680 ;
    END
  END crash_dump_o[13]
  PIN crash_dump_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END crash_dump_o[14]
  PIN crash_dump_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 229.200 1200.000 229.800 ;
    END
  END crash_dump_o[15]
  PIN crash_dump_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 289.040 1200.000 289.640 ;
    END
  END crash_dump_o[16]
  PIN crash_dump_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 329.160 1200.000 329.760 ;
    END
  END crash_dump_o[17]
  PIN crash_dump_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.470 1196.000 1036.750 1200.000 ;
    END
  END crash_dump_o[18]
  PIN crash_dump_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 369.280 1200.000 369.880 ;
    END
  END crash_dump_o[19]
  PIN crash_dump_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 0.000 1002.710 4.000 ;
    END
  END crash_dump_o[1]
  PIN crash_dump_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END crash_dump_o[20]
  PIN crash_dump_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END crash_dump_o[21]
  PIN crash_dump_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 429.120 1200.000 429.720 ;
    END
  END crash_dump_o[22]
  PIN crash_dump_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 1196.000 1056.990 1200.000 ;
    END
  END crash_dump_o[23]
  PIN crash_dump_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.770 1196.000 1062.050 1200.000 ;
    END
  END crash_dump_o[24]
  PIN crash_dump_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 1196.000 1077.230 1200.000 ;
    END
  END crash_dump_o[25]
  PIN crash_dump_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.610 1196.000 1086.890 1200.000 ;
    END
  END crash_dump_o[26]
  PIN crash_dump_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.470 0.000 1082.750 4.000 ;
    END
  END crash_dump_o[27]
  PIN crash_dump_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 509.360 1200.000 509.960 ;
    END
  END crash_dump_o[28]
  PIN crash_dump_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 529.080 1200.000 529.680 ;
    END
  END crash_dump_o[29]
  PIN crash_dump_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 89.120 1200.000 89.720 ;
    END
  END crash_dump_o[2]
  PIN crash_dump_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 1196.000 1102.070 1200.000 ;
    END
  END crash_dump_o[30]
  PIN crash_dump_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 549.480 1200.000 550.080 ;
    END
  END crash_dump_o[31]
  PIN crash_dump_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 1196.000 1112.190 1200.000 ;
    END
  END crash_dump_o[32]
  PIN crash_dump_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 569.200 1200.000 569.800 ;
    END
  END crash_dump_o[33]
  PIN crash_dump_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.080 4.000 546.680 ;
    END
  END crash_dump_o[34]
  PIN crash_dump_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.190 0.000 1097.470 4.000 ;
    END
  END crash_dump_o[35]
  PIN crash_dump_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 589.600 1200.000 590.200 ;
    END
  END crash_dump_o[36]
  PIN crash_dump_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.970 1196.000 1117.250 1200.000 ;
    END
  END crash_dump_o[37]
  PIN crash_dump_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 0.000 1102.530 4.000 ;
    END
  END crash_dump_o[38]
  PIN crash_dump_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 609.320 1200.000 609.920 ;
    END
  END crash_dump_o[39]
  PIN crash_dump_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 0.000 1007.770 4.000 ;
    END
  END crash_dump_o[3]
  PIN crash_dump_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.030 1196.000 1122.310 1200.000 ;
    END
  END crash_dump_o[40]
  PIN crash_dump_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END crash_dump_o[41]
  PIN crash_dump_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END crash_dump_o[42]
  PIN crash_dump_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 626.320 4.000 626.920 ;
    END
  END crash_dump_o[43]
  PIN crash_dump_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END crash_dump_o[44]
  PIN crash_dump_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 679.360 4.000 679.960 ;
    END
  END crash_dump_o[45]
  PIN crash_dump_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 629.040 1200.000 629.640 ;
    END
  END crash_dump_o[46]
  PIN crash_dump_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.310 0.000 1107.590 4.000 ;
    END
  END crash_dump_o[47]
  PIN crash_dump_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.370 0.000 1112.650 4.000 ;
    END
  END crash_dump_o[48]
  PIN crash_dump_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 1196.000 1127.370 1200.000 ;
    END
  END crash_dump_o[49]
  PIN crash_dump_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.090 0.000 1012.370 4.000 ;
    END
  END crash_dump_o[4]
  PIN crash_dump_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 649.440 1200.000 650.040 ;
    END
  END crash_dump_o[50]
  PIN crash_dump_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 669.160 1200.000 669.760 ;
    END
  END crash_dump_o[51]
  PIN crash_dump_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END crash_dump_o[52]
  PIN crash_dump_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END crash_dump_o[53]
  PIN crash_dump_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 689.560 1200.000 690.160 ;
    END
  END crash_dump_o[54]
  PIN crash_dump_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 709.280 1200.000 709.880 ;
    END
  END crash_dump_o[55]
  PIN crash_dump_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.150 1196.000 1132.430 1200.000 ;
    END
  END crash_dump_o[56]
  PIN crash_dump_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 4.000 ;
    END
  END crash_dump_o[57]
  PIN crash_dump_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 729.680 1200.000 730.280 ;
    END
  END crash_dump_o[58]
  PIN crash_dump_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 749.400 1200.000 750.000 ;
    END
  END crash_dump_o[59]
  PIN crash_dump_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.150 1196.000 971.430 1200.000 ;
    END
  END crash_dump_o[5]
  PIN crash_dump_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.490 0.000 1122.770 4.000 ;
    END
  END crash_dump_o[60]
  PIN crash_dump_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 769.120 1200.000 769.720 ;
    END
  END crash_dump_o[61]
  PIN crash_dump_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 759.600 4.000 760.200 ;
    END
  END crash_dump_o[62]
  PIN crash_dump_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END crash_dump_o[63]
  PIN crash_dump_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 1196.000 1137.490 1200.000 ;
    END
  END crash_dump_o[64]
  PIN crash_dump_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 789.520 1200.000 790.120 ;
    END
  END crash_dump_o[65]
  PIN crash_dump_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.270 1196.000 1142.550 1200.000 ;
    END
  END crash_dump_o[66]
  PIN crash_dump_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END crash_dump_o[67]
  PIN crash_dump_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 809.240 1200.000 809.840 ;
    END
  END crash_dump_o[68]
  PIN crash_dump_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 829.640 1200.000 830.240 ;
    END
  END crash_dump_o[69]
  PIN crash_dump_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 0.000 1022.490 4.000 ;
    END
  END crash_dump_o[6]
  PIN crash_dump_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 849.360 1200.000 849.960 ;
    END
  END crash_dump_o[70]
  PIN crash_dump_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.150 0.000 1132.430 4.000 ;
    END
  END crash_dump_o[71]
  PIN crash_dump_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 869.080 1200.000 869.680 ;
    END
  END crash_dump_o[72]
  PIN crash_dump_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 889.480 1200.000 890.080 ;
    END
  END crash_dump_o[73]
  PIN crash_dump_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 0.000 1137.490 4.000 ;
    END
  END crash_dump_o[74]
  PIN crash_dump_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.870 1196.000 1147.150 1200.000 ;
    END
  END crash_dump_o[75]
  PIN crash_dump_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END crash_dump_o[76]
  PIN crash_dump_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END crash_dump_o[77]
  PIN crash_dump_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 909.200 1200.000 909.800 ;
    END
  END crash_dump_o[78]
  PIN crash_dump_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.930 1196.000 1152.210 1200.000 ;
    END
  END crash_dump_o[79]
  PIN crash_dump_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 1196.000 981.550 1200.000 ;
    END
  END crash_dump_o[7]
  PIN crash_dump_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 929.600 1200.000 930.200 ;
    END
  END crash_dump_o[80]
  PIN crash_dump_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END crash_dump_o[81]
  PIN crash_dump_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.270 0.000 1142.550 4.000 ;
    END
  END crash_dump_o[82]
  PIN crash_dump_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.330 0.000 1147.610 4.000 ;
    END
  END crash_dump_o[83]
  PIN crash_dump_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 949.320 1200.000 949.920 ;
    END
  END crash_dump_o[84]
  PIN crash_dump_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.880 4.000 893.480 ;
    END
  END crash_dump_o[85]
  PIN crash_dump_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 919.400 4.000 920.000 ;
    END
  END crash_dump_o[86]
  PIN crash_dump_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 969.720 1200.000 970.320 ;
    END
  END crash_dump_o[87]
  PIN crash_dump_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.990 1196.000 1157.270 1200.000 ;
    END
  END crash_dump_o[88]
  PIN crash_dump_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.050 1196.000 1162.330 1200.000 ;
    END
  END crash_dump_o[89]
  PIN crash_dump_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END crash_dump_o[8]
  PIN crash_dump_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.920 4.000 946.520 ;
    END
  END crash_dump_o[90]
  PIN crash_dump_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.390 0.000 1152.670 4.000 ;
    END
  END crash_dump_o[91]
  PIN crash_dump_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.110 1196.000 1167.390 1200.000 ;
    END
  END crash_dump_o[92]
  PIN crash_dump_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 989.440 1200.000 990.040 ;
    END
  END crash_dump_o[93]
  PIN crash_dump_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.120 4.000 973.720 ;
    END
  END crash_dump_o[94]
  PIN crash_dump_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1009.160 1200.000 1009.760 ;
    END
  END crash_dump_o[95]
  PIN crash_dump_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END crash_dump_o[96]
  PIN crash_dump_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1029.560 1200.000 1030.160 ;
    END
  END crash_dump_o[97]
  PIN crash_dump_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.160 4.000 1026.760 ;
    END
  END crash_dump_o[98]
  PIN crash_dump_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 0.000 1157.730 4.000 ;
    END
  END crash_dump_o[99]
  PIN crash_dump_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END crash_dump_o[9]
  PIN data_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END data_addr_o[0]
  PIN data_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 0.000 642.530 4.000 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 0.000 672.430 4.000 ;
    END
  END data_addr_o[12]
  PIN data_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END data_addr_o[13]
  PIN data_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END data_addr_o[14]
  PIN data_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 0.000 717.510 4.000 ;
    END
  END data_addr_o[15]
  PIN data_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 4.000 ;
    END
  END data_addr_o[16]
  PIN data_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END data_addr_o[17]
  PIN data_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 0.000 762.590 4.000 ;
    END
  END data_addr_o[18]
  PIN data_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END data_addr_o[19]
  PIN data_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END data_addr_o[20]
  PIN data_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 0.000 807.670 4.000 ;
    END
  END data_addr_o[21]
  PIN data_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END data_addr_o[22]
  PIN data_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END data_addr_o[23]
  PIN data_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 0.000 852.750 4.000 ;
    END
  END data_addr_o[24]
  PIN data_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.190 0.000 867.470 4.000 ;
    END
  END data_addr_o[25]
  PIN data_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END data_addr_o[26]
  PIN data_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 0.000 897.370 4.000 ;
    END
  END data_addr_o[27]
  PIN data_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 0.000 912.550 4.000 ;
    END
  END data_addr_o[28]
  PIN data_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END data_addr_o[29]
  PIN data_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END data_addr_o[30]
  PIN data_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 0.000 957.630 4.000 ;
    END
  END data_addr_o[31]
  PIN data_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 0.000 597.450 4.000 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 0.000 627.350 4.000 ;
    END
  END data_addr_o[9]
  PIN data_be_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END data_be_o[0]
  PIN data_be_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END data_be_o[1]
  PIN data_be_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END data_be_o[2]
  PIN data_be_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END data_be_o[3]
  PIN data_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END data_err_i
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END data_gnt_i
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END data_rdata_i[0]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 0.000 662.310 4.000 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 0.000 677.490 4.000 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 0.000 707.390 4.000 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 4.000 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 4.000 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.170 0.000 827.450 4.000 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 0.000 842.630 4.000 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070 0.000 857.350 4.000 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 0.000 887.710 4.000 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.150 0.000 902.430 4.000 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.330 0.000 917.610 4.000 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 0.000 947.510 4.000 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 0.000 962.690 4.000 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END data_rdata_i[9]
  PIN data_rdata_intg_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END data_rdata_intg_i[0]
  PIN data_rdata_intg_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END data_rdata_intg_i[1]
  PIN data_rdata_intg_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END data_rdata_intg_i[2]
  PIN data_rdata_intg_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END data_rdata_intg_i[3]
  PIN data_rdata_intg_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END data_rdata_intg_i[4]
  PIN data_rdata_intg_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END data_rdata_intg_i[5]
  PIN data_rdata_intg_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END data_rdata_intg_i[6]
  PIN data_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END data_req_o
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END data_rvalid_i
  PIN data_wdata_intg_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END data_wdata_intg_o[0]
  PIN data_wdata_intg_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END data_wdata_intg_o[1]
  PIN data_wdata_intg_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END data_wdata_intg_o[2]
  PIN data_wdata_intg_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END data_wdata_intg_o[3]
  PIN data_wdata_intg_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END data_wdata_intg_o[4]
  PIN data_wdata_intg_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END data_wdata_intg_o[5]
  PIN data_wdata_intg_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END data_wdata_intg_o[6]
  PIN data_wdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END data_wdata_o[0]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 0.000 742.350 4.000 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.430 0.000 772.710 4.000 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.230 0.000 832.510 4.000 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 0.000 847.690 4.000 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 0.000 862.410 4.000 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 0.000 877.590 4.000 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 0.000 892.770 4.000 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 0.000 922.670 4.000 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 0.000 952.570 4.000 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 4.000 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END data_wdata_o[9]
  PIN data_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END data_we_o
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END debug_req_i
  PIN eFPGA_delay_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 1196.000 17.390 1200.000 ;
    END
  END eFPGA_delay_o[0]
  PIN eFPGA_delay_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 1196.000 52.810 1200.000 ;
    END
  END eFPGA_delay_o[1]
  PIN eFPGA_delay_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 1196.000 87.770 1200.000 ;
    END
  END eFPGA_delay_o[2]
  PIN eFPGA_delay_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 1196.000 118.130 1200.000 ;
    END
  END eFPGA_delay_o[3]
  PIN eFPGA_en_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 1196.000 2.670 1200.000 ;
    END
  END eFPGA_en_o
  PIN eFPGA_fpga_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 1196.000 7.270 1200.000 ;
    END
  END eFPGA_fpga_done_i
  PIN eFPGA_operand_a_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 1196.000 22.450 1200.000 ;
    END
  END eFPGA_operand_a_o[0]
  PIN eFPGA_operand_a_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 1196.000 298.910 1200.000 ;
    END
  END eFPGA_operand_a_o[10]
  PIN eFPGA_operand_a_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 1196.000 323.750 1200.000 ;
    END
  END eFPGA_operand_a_o[11]
  PIN eFPGA_operand_a_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 1196.000 349.050 1200.000 ;
    END
  END eFPGA_operand_a_o[12]
  PIN eFPGA_operand_a_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 1196.000 373.890 1200.000 ;
    END
  END eFPGA_operand_a_o[13]
  PIN eFPGA_operand_a_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 1196.000 399.190 1200.000 ;
    END
  END eFPGA_operand_a_o[14]
  PIN eFPGA_operand_a_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 1196.000 424.030 1200.000 ;
    END
  END eFPGA_operand_a_o[15]
  PIN eFPGA_operand_a_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 1196.000 449.330 1200.000 ;
    END
  END eFPGA_operand_a_o[16]
  PIN eFPGA_operand_a_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 1196.000 474.630 1200.000 ;
    END
  END eFPGA_operand_a_o[17]
  PIN eFPGA_operand_a_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 1196.000 499.470 1200.000 ;
    END
  END eFPGA_operand_a_o[18]
  PIN eFPGA_operand_a_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 1196.000 524.770 1200.000 ;
    END
  END eFPGA_operand_a_o[19]
  PIN eFPGA_operand_a_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 1196.000 57.870 1200.000 ;
    END
  END eFPGA_operand_a_o[1]
  PIN eFPGA_operand_a_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 1196.000 549.610 1200.000 ;
    END
  END eFPGA_operand_a_o[20]
  PIN eFPGA_operand_a_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 1196.000 574.910 1200.000 ;
    END
  END eFPGA_operand_a_o[21]
  PIN eFPGA_operand_a_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 1196.000 600.210 1200.000 ;
    END
  END eFPGA_operand_a_o[22]
  PIN eFPGA_operand_a_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 1196.000 625.050 1200.000 ;
    END
  END eFPGA_operand_a_o[23]
  PIN eFPGA_operand_a_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 1196.000 650.350 1200.000 ;
    END
  END eFPGA_operand_a_o[24]
  PIN eFPGA_operand_a_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 1196.000 675.190 1200.000 ;
    END
  END eFPGA_operand_a_o[25]
  PIN eFPGA_operand_a_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 1196.000 700.490 1200.000 ;
    END
  END eFPGA_operand_a_o[26]
  PIN eFPGA_operand_a_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 1196.000 725.330 1200.000 ;
    END
  END eFPGA_operand_a_o[27]
  PIN eFPGA_operand_a_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 1196.000 750.630 1200.000 ;
    END
  END eFPGA_operand_a_o[28]
  PIN eFPGA_operand_a_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 1196.000 775.930 1200.000 ;
    END
  END eFPGA_operand_a_o[29]
  PIN eFPGA_operand_a_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 1196.000 92.830 1200.000 ;
    END
  END eFPGA_operand_a_o[2]
  PIN eFPGA_operand_a_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 1196.000 800.770 1200.000 ;
    END
  END eFPGA_operand_a_o[30]
  PIN eFPGA_operand_a_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 1196.000 826.070 1200.000 ;
    END
  END eFPGA_operand_a_o[31]
  PIN eFPGA_operand_a_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1196.000 122.730 1200.000 ;
    END
  END eFPGA_operand_a_o[3]
  PIN eFPGA_operand_a_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 1196.000 148.030 1200.000 ;
    END
  END eFPGA_operand_a_o[4]
  PIN eFPGA_operand_a_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 1196.000 173.330 1200.000 ;
    END
  END eFPGA_operand_a_o[5]
  PIN eFPGA_operand_a_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 1196.000 198.170 1200.000 ;
    END
  END eFPGA_operand_a_o[6]
  PIN eFPGA_operand_a_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 1196.000 223.470 1200.000 ;
    END
  END eFPGA_operand_a_o[7]
  PIN eFPGA_operand_a_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 1196.000 248.310 1200.000 ;
    END
  END eFPGA_operand_a_o[8]
  PIN eFPGA_operand_a_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 1196.000 273.610 1200.000 ;
    END
  END eFPGA_operand_a_o[9]
  PIN eFPGA_operand_b_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 1196.000 27.510 1200.000 ;
    END
  END eFPGA_operand_b_o[0]
  PIN eFPGA_operand_b_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 1196.000 303.510 1200.000 ;
    END
  END eFPGA_operand_b_o[10]
  PIN eFPGA_operand_b_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 1196.000 328.810 1200.000 ;
    END
  END eFPGA_operand_b_o[11]
  PIN eFPGA_operand_b_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 1196.000 354.110 1200.000 ;
    END
  END eFPGA_operand_b_o[12]
  PIN eFPGA_operand_b_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 1196.000 378.950 1200.000 ;
    END
  END eFPGA_operand_b_o[13]
  PIN eFPGA_operand_b_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 1196.000 404.250 1200.000 ;
    END
  END eFPGA_operand_b_o[14]
  PIN eFPGA_operand_b_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 1196.000 429.090 1200.000 ;
    END
  END eFPGA_operand_b_o[15]
  PIN eFPGA_operand_b_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1196.000 454.390 1200.000 ;
    END
  END eFPGA_operand_b_o[16]
  PIN eFPGA_operand_b_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 1196.000 479.690 1200.000 ;
    END
  END eFPGA_operand_b_o[17]
  PIN eFPGA_operand_b_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 1196.000 504.530 1200.000 ;
    END
  END eFPGA_operand_b_o[18]
  PIN eFPGA_operand_b_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 1196.000 529.830 1200.000 ;
    END
  END eFPGA_operand_b_o[19]
  PIN eFPGA_operand_b_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 1196.000 62.470 1200.000 ;
    END
  END eFPGA_operand_b_o[1]
  PIN eFPGA_operand_b_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 1196.000 554.670 1200.000 ;
    END
  END eFPGA_operand_b_o[20]
  PIN eFPGA_operand_b_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 1196.000 579.970 1200.000 ;
    END
  END eFPGA_operand_b_o[21]
  PIN eFPGA_operand_b_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1196.000 604.810 1200.000 ;
    END
  END eFPGA_operand_b_o[22]
  PIN eFPGA_operand_b_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 1196.000 630.110 1200.000 ;
    END
  END eFPGA_operand_b_o[23]
  PIN eFPGA_operand_b_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 1196.000 655.410 1200.000 ;
    END
  END eFPGA_operand_b_o[24]
  PIN eFPGA_operand_b_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 1196.000 680.250 1200.000 ;
    END
  END eFPGA_operand_b_o[25]
  PIN eFPGA_operand_b_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 1196.000 705.550 1200.000 ;
    END
  END eFPGA_operand_b_o[26]
  PIN eFPGA_operand_b_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 1196.000 730.390 1200.000 ;
    END
  END eFPGA_operand_b_o[27]
  PIN eFPGA_operand_b_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 1196.000 755.690 1200.000 ;
    END
  END eFPGA_operand_b_o[28]
  PIN eFPGA_operand_b_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 1196.000 780.990 1200.000 ;
    END
  END eFPGA_operand_b_o[29]
  PIN eFPGA_operand_b_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 1196.000 97.890 1200.000 ;
    END
  END eFPGA_operand_b_o[2]
  PIN eFPGA_operand_b_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 1196.000 805.830 1200.000 ;
    END
  END eFPGA_operand_b_o[30]
  PIN eFPGA_operand_b_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 1196.000 831.130 1200.000 ;
    END
  END eFPGA_operand_b_o[31]
  PIN eFPGA_operand_b_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 1196.000 127.790 1200.000 ;
    END
  END eFPGA_operand_b_o[3]
  PIN eFPGA_operand_b_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 1196.000 153.090 1200.000 ;
    END
  END eFPGA_operand_b_o[4]
  PIN eFPGA_operand_b_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 1196.000 178.390 1200.000 ;
    END
  END eFPGA_operand_b_o[5]
  PIN eFPGA_operand_b_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 1196.000 203.230 1200.000 ;
    END
  END eFPGA_operand_b_o[6]
  PIN eFPGA_operand_b_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 1196.000 228.530 1200.000 ;
    END
  END eFPGA_operand_b_o[7]
  PIN eFPGA_operand_b_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 1196.000 253.370 1200.000 ;
    END
  END eFPGA_operand_b_o[8]
  PIN eFPGA_operand_b_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 1196.000 278.670 1200.000 ;
    END
  END eFPGA_operand_b_o[9]
  PIN eFPGA_operator_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 1196.000 32.570 1200.000 ;
    END
  END eFPGA_operator_o[0]
  PIN eFPGA_operator_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 1196.000 67.530 1200.000 ;
    END
  END eFPGA_operator_o[1]
  PIN eFPGA_result_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 1196.000 37.630 1200.000 ;
    END
  END eFPGA_result_a_i[0]
  PIN eFPGA_result_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 1196.000 308.570 1200.000 ;
    END
  END eFPGA_result_a_i[10]
  PIN eFPGA_result_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 1196.000 333.870 1200.000 ;
    END
  END eFPGA_result_a_i[11]
  PIN eFPGA_result_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 1196.000 359.170 1200.000 ;
    END
  END eFPGA_result_a_i[12]
  PIN eFPGA_result_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 1196.000 384.010 1200.000 ;
    END
  END eFPGA_result_a_i[13]
  PIN eFPGA_result_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 1196.000 409.310 1200.000 ;
    END
  END eFPGA_result_a_i[14]
  PIN eFPGA_result_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 1196.000 434.150 1200.000 ;
    END
  END eFPGA_result_a_i[15]
  PIN eFPGA_result_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 1196.000 459.450 1200.000 ;
    END
  END eFPGA_result_a_i[16]
  PIN eFPGA_result_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 1196.000 484.290 1200.000 ;
    END
  END eFPGA_result_a_i[17]
  PIN eFPGA_result_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 1196.000 509.590 1200.000 ;
    END
  END eFPGA_result_a_i[18]
  PIN eFPGA_result_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 1196.000 534.890 1200.000 ;
    END
  END eFPGA_result_a_i[19]
  PIN eFPGA_result_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 1196.000 72.590 1200.000 ;
    END
  END eFPGA_result_a_i[1]
  PIN eFPGA_result_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 1196.000 559.730 1200.000 ;
    END
  END eFPGA_result_a_i[20]
  PIN eFPGA_result_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 1196.000 585.030 1200.000 ;
    END
  END eFPGA_result_a_i[21]
  PIN eFPGA_result_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 1196.000 609.870 1200.000 ;
    END
  END eFPGA_result_a_i[22]
  PIN eFPGA_result_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 1196.000 635.170 1200.000 ;
    END
  END eFPGA_result_a_i[23]
  PIN eFPGA_result_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 1196.000 660.470 1200.000 ;
    END
  END eFPGA_result_a_i[24]
  PIN eFPGA_result_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 1196.000 685.310 1200.000 ;
    END
  END eFPGA_result_a_i[25]
  PIN eFPGA_result_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 1196.000 710.610 1200.000 ;
    END
  END eFPGA_result_a_i[26]
  PIN eFPGA_result_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 1196.000 735.450 1200.000 ;
    END
  END eFPGA_result_a_i[27]
  PIN eFPGA_result_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 1196.000 760.750 1200.000 ;
    END
  END eFPGA_result_a_i[28]
  PIN eFPGA_result_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 1196.000 785.590 1200.000 ;
    END
  END eFPGA_result_a_i[29]
  PIN eFPGA_result_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 1196.000 102.950 1200.000 ;
    END
  END eFPGA_result_a_i[2]
  PIN eFPGA_result_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 1196.000 810.890 1200.000 ;
    END
  END eFPGA_result_a_i[30]
  PIN eFPGA_result_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.910 1196.000 836.190 1200.000 ;
    END
  END eFPGA_result_a_i[31]
  PIN eFPGA_result_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 1196.000 132.850 1200.000 ;
    END
  END eFPGA_result_a_i[3]
  PIN eFPGA_result_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 1196.000 158.150 1200.000 ;
    END
  END eFPGA_result_a_i[4]
  PIN eFPGA_result_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 1196.000 182.990 1200.000 ;
    END
  END eFPGA_result_a_i[5]
  PIN eFPGA_result_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 1196.000 208.290 1200.000 ;
    END
  END eFPGA_result_a_i[6]
  PIN eFPGA_result_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 1196.000 233.590 1200.000 ;
    END
  END eFPGA_result_a_i[7]
  PIN eFPGA_result_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 1196.000 258.430 1200.000 ;
    END
  END eFPGA_result_a_i[8]
  PIN eFPGA_result_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1196.000 283.730 1200.000 ;
    END
  END eFPGA_result_a_i[9]
  PIN eFPGA_result_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 1196.000 42.690 1200.000 ;
    END
  END eFPGA_result_b_i[0]
  PIN eFPGA_result_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 1196.000 313.630 1200.000 ;
    END
  END eFPGA_result_b_i[10]
  PIN eFPGA_result_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 1196.000 338.930 1200.000 ;
    END
  END eFPGA_result_b_i[11]
  PIN eFPGA_result_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 1196.000 363.770 1200.000 ;
    END
  END eFPGA_result_b_i[12]
  PIN eFPGA_result_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 1196.000 389.070 1200.000 ;
    END
  END eFPGA_result_b_i[13]
  PIN eFPGA_result_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 1196.000 414.370 1200.000 ;
    END
  END eFPGA_result_b_i[14]
  PIN eFPGA_result_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 1196.000 439.210 1200.000 ;
    END
  END eFPGA_result_b_i[15]
  PIN eFPGA_result_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 1196.000 464.510 1200.000 ;
    END
  END eFPGA_result_b_i[16]
  PIN eFPGA_result_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 1196.000 489.350 1200.000 ;
    END
  END eFPGA_result_b_i[17]
  PIN eFPGA_result_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 1196.000 514.650 1200.000 ;
    END
  END eFPGA_result_b_i[18]
  PIN eFPGA_result_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 1196.000 539.950 1200.000 ;
    END
  END eFPGA_result_b_i[19]
  PIN eFPGA_result_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1196.000 77.650 1200.000 ;
    END
  END eFPGA_result_b_i[1]
  PIN eFPGA_result_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 1196.000 564.790 1200.000 ;
    END
  END eFPGA_result_b_i[20]
  PIN eFPGA_result_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 1196.000 590.090 1200.000 ;
    END
  END eFPGA_result_b_i[21]
  PIN eFPGA_result_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 1196.000 614.930 1200.000 ;
    END
  END eFPGA_result_b_i[22]
  PIN eFPGA_result_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 1196.000 640.230 1200.000 ;
    END
  END eFPGA_result_b_i[23]
  PIN eFPGA_result_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 1196.000 665.070 1200.000 ;
    END
  END eFPGA_result_b_i[24]
  PIN eFPGA_result_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 1196.000 690.370 1200.000 ;
    END
  END eFPGA_result_b_i[25]
  PIN eFPGA_result_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 1196.000 715.670 1200.000 ;
    END
  END eFPGA_result_b_i[26]
  PIN eFPGA_result_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 1196.000 740.510 1200.000 ;
    END
  END eFPGA_result_b_i[27]
  PIN eFPGA_result_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 1196.000 765.810 1200.000 ;
    END
  END eFPGA_result_b_i[28]
  PIN eFPGA_result_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 1196.000 790.650 1200.000 ;
    END
  END eFPGA_result_b_i[29]
  PIN eFPGA_result_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 1196.000 108.010 1200.000 ;
    END
  END eFPGA_result_b_i[2]
  PIN eFPGA_result_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 1196.000 815.950 1200.000 ;
    END
  END eFPGA_result_b_i[30]
  PIN eFPGA_result_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.970 1196.000 841.250 1200.000 ;
    END
  END eFPGA_result_b_i[31]
  PIN eFPGA_result_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 1196.000 137.910 1200.000 ;
    END
  END eFPGA_result_b_i[3]
  PIN eFPGA_result_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 1196.000 163.210 1200.000 ;
    END
  END eFPGA_result_b_i[4]
  PIN eFPGA_result_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 1196.000 188.050 1200.000 ;
    END
  END eFPGA_result_b_i[5]
  PIN eFPGA_result_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 1196.000 213.350 1200.000 ;
    END
  END eFPGA_result_b_i[6]
  PIN eFPGA_result_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 1196.000 238.650 1200.000 ;
    END
  END eFPGA_result_b_i[7]
  PIN eFPGA_result_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 1196.000 263.490 1200.000 ;
    END
  END eFPGA_result_b_i[8]
  PIN eFPGA_result_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 1196.000 288.790 1200.000 ;
    END
  END eFPGA_result_b_i[9]
  PIN eFPGA_result_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 1196.000 47.750 1200.000 ;
    END
  END eFPGA_result_c_i[0]
  PIN eFPGA_result_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 1196.000 318.690 1200.000 ;
    END
  END eFPGA_result_c_i[10]
  PIN eFPGA_result_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 1196.000 343.990 1200.000 ;
    END
  END eFPGA_result_c_i[11]
  PIN eFPGA_result_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 1196.000 368.830 1200.000 ;
    END
  END eFPGA_result_c_i[12]
  PIN eFPGA_result_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 1196.000 394.130 1200.000 ;
    END
  END eFPGA_result_c_i[13]
  PIN eFPGA_result_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 1196.000 419.430 1200.000 ;
    END
  END eFPGA_result_c_i[14]
  PIN eFPGA_result_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 1196.000 444.270 1200.000 ;
    END
  END eFPGA_result_c_i[15]
  PIN eFPGA_result_c_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 1196.000 469.570 1200.000 ;
    END
  END eFPGA_result_c_i[16]
  PIN eFPGA_result_c_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 1196.000 494.410 1200.000 ;
    END
  END eFPGA_result_c_i[17]
  PIN eFPGA_result_c_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 1196.000 519.710 1200.000 ;
    END
  END eFPGA_result_c_i[18]
  PIN eFPGA_result_c_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 1196.000 544.550 1200.000 ;
    END
  END eFPGA_result_c_i[19]
  PIN eFPGA_result_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 1196.000 82.710 1200.000 ;
    END
  END eFPGA_result_c_i[1]
  PIN eFPGA_result_c_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 1196.000 569.850 1200.000 ;
    END
  END eFPGA_result_c_i[20]
  PIN eFPGA_result_c_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 1196.000 595.150 1200.000 ;
    END
  END eFPGA_result_c_i[21]
  PIN eFPGA_result_c_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 1196.000 619.990 1200.000 ;
    END
  END eFPGA_result_c_i[22]
  PIN eFPGA_result_c_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 1196.000 645.290 1200.000 ;
    END
  END eFPGA_result_c_i[23]
  PIN eFPGA_result_c_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 1196.000 670.130 1200.000 ;
    END
  END eFPGA_result_c_i[24]
  PIN eFPGA_result_c_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 1196.000 695.430 1200.000 ;
    END
  END eFPGA_result_c_i[25]
  PIN eFPGA_result_c_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 1196.000 720.730 1200.000 ;
    END
  END eFPGA_result_c_i[26]
  PIN eFPGA_result_c_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 1196.000 745.570 1200.000 ;
    END
  END eFPGA_result_c_i[27]
  PIN eFPGA_result_c_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 1196.000 770.870 1200.000 ;
    END
  END eFPGA_result_c_i[28]
  PIN eFPGA_result_c_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 1196.000 795.710 1200.000 ;
    END
  END eFPGA_result_c_i[29]
  PIN eFPGA_result_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1196.000 113.070 1200.000 ;
    END
  END eFPGA_result_c_i[2]
  PIN eFPGA_result_c_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 1196.000 821.010 1200.000 ;
    END
  END eFPGA_result_c_i[30]
  PIN eFPGA_result_c_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 1196.000 845.850 1200.000 ;
    END
  END eFPGA_result_c_i[31]
  PIN eFPGA_result_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 1196.000 142.970 1200.000 ;
    END
  END eFPGA_result_c_i[3]
  PIN eFPGA_result_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 1196.000 168.270 1200.000 ;
    END
  END eFPGA_result_c_i[4]
  PIN eFPGA_result_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 1196.000 193.110 1200.000 ;
    END
  END eFPGA_result_c_i[5]
  PIN eFPGA_result_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 1196.000 218.410 1200.000 ;
    END
  END eFPGA_result_c_i[6]
  PIN eFPGA_result_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 1196.000 243.250 1200.000 ;
    END
  END eFPGA_result_c_i[7]
  PIN eFPGA_result_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 1196.000 268.550 1200.000 ;
    END
  END eFPGA_result_c_i[8]
  PIN eFPGA_result_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 1196.000 293.850 1200.000 ;
    END
  END eFPGA_result_c_i[9]
  PIN eFPGA_write_strobe_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 1196.000 12.330 1200.000 ;
    END
  END eFPGA_write_strobe_o
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 1196.000 946.590 1200.000 ;
    END
  END fetch_enable_i
  PIN hart_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 49.000 1200.000 49.600 ;
    END
  END hart_id_i[0]
  PIN hart_id_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 148.960 1200.000 149.560 ;
    END
  END hart_id_i[10]
  PIN hart_id_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.450 0.000 1042.730 4.000 ;
    END
  END hart_id_i[11]
  PIN hart_id_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 0.000 1047.790 4.000 ;
    END
  END hart_id_i[12]
  PIN hart_id_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.170 0.000 1057.450 4.000 ;
    END
  END hart_id_i[13]
  PIN hart_id_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.750 1196.000 1022.030 1200.000 ;
    END
  END hart_id_i[14]
  PIN hart_id_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 249.600 1200.000 250.200 ;
    END
  END hart_id_i[15]
  PIN hart_id_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 309.440 1200.000 310.040 ;
    END
  END hart_id_i[16]
  PIN hart_id_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 349.560 1200.000 350.160 ;
    END
  END hart_id_i[17]
  PIN hart_id_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.530 1196.000 1041.810 1200.000 ;
    END
  END hart_id_i[18]
  PIN hart_id_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.290 0.000 1067.570 4.000 ;
    END
  END hart_id_i[19]
  PIN hart_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 1196.000 961.770 1200.000 ;
    END
  END hart_id_i[1]
  PIN hart_id_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END hart_id_i[20]
  PIN hart_id_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 389.000 1200.000 389.600 ;
    END
  END hart_id_i[21]
  PIN hart_id_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END hart_id_i[22]
  PIN hart_id_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.410 0.000 1077.690 4.000 ;
    END
  END hart_id_i[23]
  PIN hart_id_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.830 1196.000 1067.110 1200.000 ;
    END
  END hart_id_i[24]
  PIN hart_id_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 1196.000 1082.290 1200.000 ;
    END
  END hart_id_i[25]
  PIN hart_id_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 1196.000 1091.950 1200.000 ;
    END
  END hart_id_i[26]
  PIN hart_id_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END hart_id_i[27]
  PIN hart_id_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END hart_id_i[28]
  PIN hart_id_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END hart_id_i[29]
  PIN hart_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END hart_id_i[2]
  PIN hart_id_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END hart_id_i[30]
  PIN hart_id_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 1196.000 1107.130 1200.000 ;
    END
  END hart_id_i[31]
  PIN hart_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 109.520 1200.000 110.120 ;
    END
  END hart_id_i[3]
  PIN hart_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 0.000 1017.430 4.000 ;
    END
  END hart_id_i[4]
  PIN hart_id_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END hart_id_i[5]
  PIN hart_id_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 0.000 1027.550 4.000 ;
    END
  END hart_id_i[6]
  PIN hart_id_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330 1196.000 986.610 1200.000 ;
    END
  END hart_id_i[7]
  PIN hart_id_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 1196.000 991.670 1200.000 ;
    END
  END hart_id_i[8]
  PIN hart_id_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 1196.000 1001.790 1200.000 ;
    END
  END hart_id_i[9]
  PIN instr_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END instr_addr_o[0]
  PIN instr_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END instr_addr_o[10]
  PIN instr_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END instr_addr_o[11]
  PIN instr_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END instr_addr_o[12]
  PIN instr_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END instr_addr_o[13]
  PIN instr_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END instr_addr_o[14]
  PIN instr_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END instr_addr_o[15]
  PIN instr_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END instr_addr_o[16]
  PIN instr_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END instr_addr_o[17]
  PIN instr_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END instr_addr_o[18]
  PIN instr_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END instr_addr_o[19]
  PIN instr_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END instr_addr_o[1]
  PIN instr_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END instr_addr_o[20]
  PIN instr_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END instr_addr_o[21]
  PIN instr_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END instr_addr_o[22]
  PIN instr_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END instr_addr_o[23]
  PIN instr_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END instr_addr_o[24]
  PIN instr_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END instr_addr_o[25]
  PIN instr_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END instr_addr_o[26]
  PIN instr_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END instr_addr_o[27]
  PIN instr_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END instr_addr_o[28]
  PIN instr_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END instr_addr_o[29]
  PIN instr_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END instr_addr_o[2]
  PIN instr_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END instr_addr_o[30]
  PIN instr_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END instr_addr_o[31]
  PIN instr_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END instr_addr_o[3]
  PIN instr_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END instr_addr_o[4]
  PIN instr_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END instr_addr_o[5]
  PIN instr_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END instr_addr_o[6]
  PIN instr_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END instr_addr_o[7]
  PIN instr_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END instr_addr_o[8]
  PIN instr_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END instr_addr_o[9]
  PIN instr_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END instr_err_i
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END instr_gnt_i
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END instr_rdata_i[0]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END instr_rdata_i[9]
  PIN instr_rdata_intg_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END instr_rdata_intg_i[0]
  PIN instr_rdata_intg_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END instr_rdata_intg_i[1]
  PIN instr_rdata_intg_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END instr_rdata_intg_i[2]
  PIN instr_rdata_intg_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END instr_rdata_intg_i[3]
  PIN instr_rdata_intg_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END instr_rdata_intg_i[4]
  PIN instr_rdata_intg_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END instr_rdata_intg_i[5]
  PIN instr_rdata_intg_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END instr_rdata_intg_i[6]
  PIN instr_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END instr_req_o
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END instr_rvalid_i
  PIN irq_external_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 1196.000 850.910 1200.000 ;
    END
  END irq_external_i
  PIN irq_fast_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 1196.000 871.150 1200.000 ;
    END
  END irq_fast_i[0]
  PIN irq_fast_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 1196.000 921.290 1200.000 ;
    END
  END irq_fast_i[10]
  PIN irq_fast_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 1196.000 926.350 1200.000 ;
    END
  END irq_fast_i[11]
  PIN irq_fast_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 1196.000 931.410 1200.000 ;
    END
  END irq_fast_i[12]
  PIN irq_fast_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.190 1196.000 936.470 1200.000 ;
    END
  END irq_fast_i[13]
  PIN irq_fast_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 1196.000 941.530 1200.000 ;
    END
  END irq_fast_i[14]
  PIN irq_fast_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 1196.000 876.210 1200.000 ;
    END
  END irq_fast_i[1]
  PIN irq_fast_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 1196.000 881.270 1200.000 ;
    END
  END irq_fast_i[2]
  PIN irq_fast_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 1196.000 886.330 1200.000 ;
    END
  END irq_fast_i[3]
  PIN irq_fast_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 1196.000 891.390 1200.000 ;
    END
  END irq_fast_i[4]
  PIN irq_fast_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 1196.000 896.450 1200.000 ;
    END
  END irq_fast_i[5]
  PIN irq_fast_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 1196.000 901.510 1200.000 ;
    END
  END irq_fast_i[6]
  PIN irq_fast_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.830 1196.000 906.110 1200.000 ;
    END
  END irq_fast_i[7]
  PIN irq_fast_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 1196.000 911.170 1200.000 ;
    END
  END irq_fast_i[8]
  PIN irq_fast_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 1196.000 916.230 1200.000 ;
    END
  END irq_fast_i[9]
  PIN irq_nm_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 1196.000 855.970 1200.000 ;
    END
  END irq_nm_i
  PIN irq_software_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 1196.000 861.030 1200.000 ;
    END
  END irq_software_i
  PIN irq_timer_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 1196.000 866.090 1200.000 ;
    END
  END irq_timer_i
  PIN ram_cfg_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 1196.000 951.650 1200.000 ;
    END
  END ram_cfg_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 1196.000 956.710 1200.000 ;
    END
  END rst_ni
  PIN scan_rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END scan_rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 0.000 992.590 4.000 ;
    END
  END test_en_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1188.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1188.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 7.905 1198.615 1189.915 ;
      LAYER met1 ;
        RECT 2.370 7.520 1198.675 1190.300 ;
      LAYER met2 ;
        RECT 2.950 1195.720 6.710 1196.530 ;
        RECT 7.550 1195.720 11.770 1196.530 ;
        RECT 12.610 1195.720 16.830 1196.530 ;
        RECT 17.670 1195.720 21.890 1196.530 ;
        RECT 22.730 1195.720 26.950 1196.530 ;
        RECT 27.790 1195.720 32.010 1196.530 ;
        RECT 32.850 1195.720 37.070 1196.530 ;
        RECT 37.910 1195.720 42.130 1196.530 ;
        RECT 42.970 1195.720 47.190 1196.530 ;
        RECT 48.030 1195.720 52.250 1196.530 ;
        RECT 53.090 1195.720 57.310 1196.530 ;
        RECT 58.150 1195.720 61.910 1196.530 ;
        RECT 62.750 1195.720 66.970 1196.530 ;
        RECT 67.810 1195.720 72.030 1196.530 ;
        RECT 72.870 1195.720 77.090 1196.530 ;
        RECT 77.930 1195.720 82.150 1196.530 ;
        RECT 82.990 1195.720 87.210 1196.530 ;
        RECT 88.050 1195.720 92.270 1196.530 ;
        RECT 93.110 1195.720 97.330 1196.530 ;
        RECT 98.170 1195.720 102.390 1196.530 ;
        RECT 103.230 1195.720 107.450 1196.530 ;
        RECT 108.290 1195.720 112.510 1196.530 ;
        RECT 113.350 1195.720 117.570 1196.530 ;
        RECT 118.410 1195.720 122.170 1196.530 ;
        RECT 123.010 1195.720 127.230 1196.530 ;
        RECT 128.070 1195.720 132.290 1196.530 ;
        RECT 133.130 1195.720 137.350 1196.530 ;
        RECT 138.190 1195.720 142.410 1196.530 ;
        RECT 143.250 1195.720 147.470 1196.530 ;
        RECT 148.310 1195.720 152.530 1196.530 ;
        RECT 153.370 1195.720 157.590 1196.530 ;
        RECT 158.430 1195.720 162.650 1196.530 ;
        RECT 163.490 1195.720 167.710 1196.530 ;
        RECT 168.550 1195.720 172.770 1196.530 ;
        RECT 173.610 1195.720 177.830 1196.530 ;
        RECT 178.670 1195.720 182.430 1196.530 ;
        RECT 183.270 1195.720 187.490 1196.530 ;
        RECT 188.330 1195.720 192.550 1196.530 ;
        RECT 193.390 1195.720 197.610 1196.530 ;
        RECT 198.450 1195.720 202.670 1196.530 ;
        RECT 203.510 1195.720 207.730 1196.530 ;
        RECT 208.570 1195.720 212.790 1196.530 ;
        RECT 213.630 1195.720 217.850 1196.530 ;
        RECT 218.690 1195.720 222.910 1196.530 ;
        RECT 223.750 1195.720 227.970 1196.530 ;
        RECT 228.810 1195.720 233.030 1196.530 ;
        RECT 233.870 1195.720 238.090 1196.530 ;
        RECT 238.930 1195.720 242.690 1196.530 ;
        RECT 243.530 1195.720 247.750 1196.530 ;
        RECT 248.590 1195.720 252.810 1196.530 ;
        RECT 253.650 1195.720 257.870 1196.530 ;
        RECT 258.710 1195.720 262.930 1196.530 ;
        RECT 263.770 1195.720 267.990 1196.530 ;
        RECT 268.830 1195.720 273.050 1196.530 ;
        RECT 273.890 1195.720 278.110 1196.530 ;
        RECT 278.950 1195.720 283.170 1196.530 ;
        RECT 284.010 1195.720 288.230 1196.530 ;
        RECT 289.070 1195.720 293.290 1196.530 ;
        RECT 294.130 1195.720 298.350 1196.530 ;
        RECT 299.190 1195.720 302.950 1196.530 ;
        RECT 303.790 1195.720 308.010 1196.530 ;
        RECT 308.850 1195.720 313.070 1196.530 ;
        RECT 313.910 1195.720 318.130 1196.530 ;
        RECT 318.970 1195.720 323.190 1196.530 ;
        RECT 324.030 1195.720 328.250 1196.530 ;
        RECT 329.090 1195.720 333.310 1196.530 ;
        RECT 334.150 1195.720 338.370 1196.530 ;
        RECT 339.210 1195.720 343.430 1196.530 ;
        RECT 344.270 1195.720 348.490 1196.530 ;
        RECT 349.330 1195.720 353.550 1196.530 ;
        RECT 354.390 1195.720 358.610 1196.530 ;
        RECT 359.450 1195.720 363.210 1196.530 ;
        RECT 364.050 1195.720 368.270 1196.530 ;
        RECT 369.110 1195.720 373.330 1196.530 ;
        RECT 374.170 1195.720 378.390 1196.530 ;
        RECT 379.230 1195.720 383.450 1196.530 ;
        RECT 384.290 1195.720 388.510 1196.530 ;
        RECT 389.350 1195.720 393.570 1196.530 ;
        RECT 394.410 1195.720 398.630 1196.530 ;
        RECT 399.470 1195.720 403.690 1196.530 ;
        RECT 404.530 1195.720 408.750 1196.530 ;
        RECT 409.590 1195.720 413.810 1196.530 ;
        RECT 414.650 1195.720 418.870 1196.530 ;
        RECT 419.710 1195.720 423.470 1196.530 ;
        RECT 424.310 1195.720 428.530 1196.530 ;
        RECT 429.370 1195.720 433.590 1196.530 ;
        RECT 434.430 1195.720 438.650 1196.530 ;
        RECT 439.490 1195.720 443.710 1196.530 ;
        RECT 444.550 1195.720 448.770 1196.530 ;
        RECT 449.610 1195.720 453.830 1196.530 ;
        RECT 454.670 1195.720 458.890 1196.530 ;
        RECT 459.730 1195.720 463.950 1196.530 ;
        RECT 464.790 1195.720 469.010 1196.530 ;
        RECT 469.850 1195.720 474.070 1196.530 ;
        RECT 474.910 1195.720 479.130 1196.530 ;
        RECT 479.970 1195.720 483.730 1196.530 ;
        RECT 484.570 1195.720 488.790 1196.530 ;
        RECT 489.630 1195.720 493.850 1196.530 ;
        RECT 494.690 1195.720 498.910 1196.530 ;
        RECT 499.750 1195.720 503.970 1196.530 ;
        RECT 504.810 1195.720 509.030 1196.530 ;
        RECT 509.870 1195.720 514.090 1196.530 ;
        RECT 514.930 1195.720 519.150 1196.530 ;
        RECT 519.990 1195.720 524.210 1196.530 ;
        RECT 525.050 1195.720 529.270 1196.530 ;
        RECT 530.110 1195.720 534.330 1196.530 ;
        RECT 535.170 1195.720 539.390 1196.530 ;
        RECT 540.230 1195.720 543.990 1196.530 ;
        RECT 544.830 1195.720 549.050 1196.530 ;
        RECT 549.890 1195.720 554.110 1196.530 ;
        RECT 554.950 1195.720 559.170 1196.530 ;
        RECT 560.010 1195.720 564.230 1196.530 ;
        RECT 565.070 1195.720 569.290 1196.530 ;
        RECT 570.130 1195.720 574.350 1196.530 ;
        RECT 575.190 1195.720 579.410 1196.530 ;
        RECT 580.250 1195.720 584.470 1196.530 ;
        RECT 585.310 1195.720 589.530 1196.530 ;
        RECT 590.370 1195.720 594.590 1196.530 ;
        RECT 595.430 1195.720 599.650 1196.530 ;
        RECT 600.490 1195.720 604.250 1196.530 ;
        RECT 605.090 1195.720 609.310 1196.530 ;
        RECT 610.150 1195.720 614.370 1196.530 ;
        RECT 615.210 1195.720 619.430 1196.530 ;
        RECT 620.270 1195.720 624.490 1196.530 ;
        RECT 625.330 1195.720 629.550 1196.530 ;
        RECT 630.390 1195.720 634.610 1196.530 ;
        RECT 635.450 1195.720 639.670 1196.530 ;
        RECT 640.510 1195.720 644.730 1196.530 ;
        RECT 645.570 1195.720 649.790 1196.530 ;
        RECT 650.630 1195.720 654.850 1196.530 ;
        RECT 655.690 1195.720 659.910 1196.530 ;
        RECT 660.750 1195.720 664.510 1196.530 ;
        RECT 665.350 1195.720 669.570 1196.530 ;
        RECT 670.410 1195.720 674.630 1196.530 ;
        RECT 675.470 1195.720 679.690 1196.530 ;
        RECT 680.530 1195.720 684.750 1196.530 ;
        RECT 685.590 1195.720 689.810 1196.530 ;
        RECT 690.650 1195.720 694.870 1196.530 ;
        RECT 695.710 1195.720 699.930 1196.530 ;
        RECT 700.770 1195.720 704.990 1196.530 ;
        RECT 705.830 1195.720 710.050 1196.530 ;
        RECT 710.890 1195.720 715.110 1196.530 ;
        RECT 715.950 1195.720 720.170 1196.530 ;
        RECT 721.010 1195.720 724.770 1196.530 ;
        RECT 725.610 1195.720 729.830 1196.530 ;
        RECT 730.670 1195.720 734.890 1196.530 ;
        RECT 735.730 1195.720 739.950 1196.530 ;
        RECT 740.790 1195.720 745.010 1196.530 ;
        RECT 745.850 1195.720 750.070 1196.530 ;
        RECT 750.910 1195.720 755.130 1196.530 ;
        RECT 755.970 1195.720 760.190 1196.530 ;
        RECT 761.030 1195.720 765.250 1196.530 ;
        RECT 766.090 1195.720 770.310 1196.530 ;
        RECT 771.150 1195.720 775.370 1196.530 ;
        RECT 776.210 1195.720 780.430 1196.530 ;
        RECT 781.270 1195.720 785.030 1196.530 ;
        RECT 785.870 1195.720 790.090 1196.530 ;
        RECT 790.930 1195.720 795.150 1196.530 ;
        RECT 795.990 1195.720 800.210 1196.530 ;
        RECT 801.050 1195.720 805.270 1196.530 ;
        RECT 806.110 1195.720 810.330 1196.530 ;
        RECT 811.170 1195.720 815.390 1196.530 ;
        RECT 816.230 1195.720 820.450 1196.530 ;
        RECT 821.290 1195.720 825.510 1196.530 ;
        RECT 826.350 1195.720 830.570 1196.530 ;
        RECT 831.410 1195.720 835.630 1196.530 ;
        RECT 836.470 1195.720 840.690 1196.530 ;
        RECT 841.530 1195.720 845.290 1196.530 ;
        RECT 846.130 1195.720 850.350 1196.530 ;
        RECT 851.190 1195.720 855.410 1196.530 ;
        RECT 856.250 1195.720 860.470 1196.530 ;
        RECT 861.310 1195.720 865.530 1196.530 ;
        RECT 866.370 1195.720 870.590 1196.530 ;
        RECT 871.430 1195.720 875.650 1196.530 ;
        RECT 876.490 1195.720 880.710 1196.530 ;
        RECT 881.550 1195.720 885.770 1196.530 ;
        RECT 886.610 1195.720 890.830 1196.530 ;
        RECT 891.670 1195.720 895.890 1196.530 ;
        RECT 896.730 1195.720 900.950 1196.530 ;
        RECT 901.790 1195.720 905.550 1196.530 ;
        RECT 906.390 1195.720 910.610 1196.530 ;
        RECT 911.450 1195.720 915.670 1196.530 ;
        RECT 916.510 1195.720 920.730 1196.530 ;
        RECT 921.570 1195.720 925.790 1196.530 ;
        RECT 926.630 1195.720 930.850 1196.530 ;
        RECT 931.690 1195.720 935.910 1196.530 ;
        RECT 936.750 1195.720 940.970 1196.530 ;
        RECT 941.810 1195.720 946.030 1196.530 ;
        RECT 946.870 1195.720 951.090 1196.530 ;
        RECT 951.930 1195.720 956.150 1196.530 ;
        RECT 956.990 1195.720 961.210 1196.530 ;
        RECT 962.050 1195.720 965.810 1196.530 ;
        RECT 966.650 1195.720 970.870 1196.530 ;
        RECT 971.710 1195.720 975.930 1196.530 ;
        RECT 976.770 1195.720 980.990 1196.530 ;
        RECT 981.830 1195.720 986.050 1196.530 ;
        RECT 986.890 1195.720 991.110 1196.530 ;
        RECT 991.950 1195.720 996.170 1196.530 ;
        RECT 997.010 1195.720 1001.230 1196.530 ;
        RECT 1002.070 1195.720 1006.290 1196.530 ;
        RECT 1007.130 1195.720 1011.350 1196.530 ;
        RECT 1012.190 1195.720 1016.410 1196.530 ;
        RECT 1017.250 1195.720 1021.470 1196.530 ;
        RECT 1022.310 1195.720 1026.070 1196.530 ;
        RECT 1026.910 1195.720 1031.130 1196.530 ;
        RECT 1031.970 1195.720 1036.190 1196.530 ;
        RECT 1037.030 1195.720 1041.250 1196.530 ;
        RECT 1042.090 1195.720 1046.310 1196.530 ;
        RECT 1047.150 1195.720 1051.370 1196.530 ;
        RECT 1052.210 1195.720 1056.430 1196.530 ;
        RECT 1057.270 1195.720 1061.490 1196.530 ;
        RECT 1062.330 1195.720 1066.550 1196.530 ;
        RECT 1067.390 1195.720 1071.610 1196.530 ;
        RECT 1072.450 1195.720 1076.670 1196.530 ;
        RECT 1077.510 1195.720 1081.730 1196.530 ;
        RECT 1082.570 1195.720 1086.330 1196.530 ;
        RECT 1087.170 1195.720 1091.390 1196.530 ;
        RECT 1092.230 1195.720 1096.450 1196.530 ;
        RECT 1097.290 1195.720 1101.510 1196.530 ;
        RECT 1102.350 1195.720 1106.570 1196.530 ;
        RECT 1107.410 1195.720 1111.630 1196.530 ;
        RECT 1112.470 1195.720 1116.690 1196.530 ;
        RECT 1117.530 1195.720 1121.750 1196.530 ;
        RECT 1122.590 1195.720 1126.810 1196.530 ;
        RECT 1127.650 1195.720 1131.870 1196.530 ;
        RECT 1132.710 1195.720 1136.930 1196.530 ;
        RECT 1137.770 1195.720 1141.990 1196.530 ;
        RECT 1142.830 1195.720 1146.590 1196.530 ;
        RECT 1147.430 1195.720 1151.650 1196.530 ;
        RECT 1152.490 1195.720 1156.710 1196.530 ;
        RECT 1157.550 1195.720 1161.770 1196.530 ;
        RECT 1162.610 1195.720 1166.830 1196.530 ;
        RECT 1167.670 1195.720 1171.890 1196.530 ;
        RECT 1172.730 1195.720 1176.950 1196.530 ;
        RECT 1177.790 1195.720 1182.010 1196.530 ;
        RECT 1182.850 1195.720 1187.070 1196.530 ;
        RECT 1187.910 1195.720 1192.130 1196.530 ;
        RECT 1192.970 1195.720 1197.190 1196.530 ;
        RECT 2.400 4.280 1197.740 1195.720 ;
        RECT 2.950 3.670 6.710 4.280 ;
        RECT 7.550 3.670 11.770 4.280 ;
        RECT 12.610 3.670 16.830 4.280 ;
        RECT 17.670 3.670 21.890 4.280 ;
        RECT 22.730 3.670 26.950 4.280 ;
        RECT 27.790 3.670 32.010 4.280 ;
        RECT 32.850 3.670 37.070 4.280 ;
        RECT 37.910 3.670 41.670 4.280 ;
        RECT 42.510 3.670 46.730 4.280 ;
        RECT 47.570 3.670 51.790 4.280 ;
        RECT 52.630 3.670 56.850 4.280 ;
        RECT 57.690 3.670 61.910 4.280 ;
        RECT 62.750 3.670 66.970 4.280 ;
        RECT 67.810 3.670 72.030 4.280 ;
        RECT 72.870 3.670 77.090 4.280 ;
        RECT 77.930 3.670 81.690 4.280 ;
        RECT 82.530 3.670 86.750 4.280 ;
        RECT 87.590 3.670 91.810 4.280 ;
        RECT 92.650 3.670 96.870 4.280 ;
        RECT 97.710 3.670 101.930 4.280 ;
        RECT 102.770 3.670 106.990 4.280 ;
        RECT 107.830 3.670 112.050 4.280 ;
        RECT 112.890 3.670 117.110 4.280 ;
        RECT 117.950 3.670 121.710 4.280 ;
        RECT 122.550 3.670 126.770 4.280 ;
        RECT 127.610 3.670 131.830 4.280 ;
        RECT 132.670 3.670 136.890 4.280 ;
        RECT 137.730 3.670 141.950 4.280 ;
        RECT 142.790 3.670 147.010 4.280 ;
        RECT 147.850 3.670 152.070 4.280 ;
        RECT 152.910 3.670 156.670 4.280 ;
        RECT 157.510 3.670 161.730 4.280 ;
        RECT 162.570 3.670 166.790 4.280 ;
        RECT 167.630 3.670 171.850 4.280 ;
        RECT 172.690 3.670 176.910 4.280 ;
        RECT 177.750 3.670 181.970 4.280 ;
        RECT 182.810 3.670 187.030 4.280 ;
        RECT 187.870 3.670 192.090 4.280 ;
        RECT 192.930 3.670 196.690 4.280 ;
        RECT 197.530 3.670 201.750 4.280 ;
        RECT 202.590 3.670 206.810 4.280 ;
        RECT 207.650 3.670 211.870 4.280 ;
        RECT 212.710 3.670 216.930 4.280 ;
        RECT 217.770 3.670 221.990 4.280 ;
        RECT 222.830 3.670 227.050 4.280 ;
        RECT 227.890 3.670 232.110 4.280 ;
        RECT 232.950 3.670 236.710 4.280 ;
        RECT 237.550 3.670 241.770 4.280 ;
        RECT 242.610 3.670 246.830 4.280 ;
        RECT 247.670 3.670 251.890 4.280 ;
        RECT 252.730 3.670 256.950 4.280 ;
        RECT 257.790 3.670 262.010 4.280 ;
        RECT 262.850 3.670 267.070 4.280 ;
        RECT 267.910 3.670 272.130 4.280 ;
        RECT 272.970 3.670 276.730 4.280 ;
        RECT 277.570 3.670 281.790 4.280 ;
        RECT 282.630 3.670 286.850 4.280 ;
        RECT 287.690 3.670 291.910 4.280 ;
        RECT 292.750 3.670 296.970 4.280 ;
        RECT 297.810 3.670 302.030 4.280 ;
        RECT 302.870 3.670 307.090 4.280 ;
        RECT 307.930 3.670 311.690 4.280 ;
        RECT 312.530 3.670 316.750 4.280 ;
        RECT 317.590 3.670 321.810 4.280 ;
        RECT 322.650 3.670 326.870 4.280 ;
        RECT 327.710 3.670 331.930 4.280 ;
        RECT 332.770 3.670 336.990 4.280 ;
        RECT 337.830 3.670 342.050 4.280 ;
        RECT 342.890 3.670 347.110 4.280 ;
        RECT 347.950 3.670 351.710 4.280 ;
        RECT 352.550 3.670 356.770 4.280 ;
        RECT 357.610 3.670 361.830 4.280 ;
        RECT 362.670 3.670 366.890 4.280 ;
        RECT 367.730 3.670 371.950 4.280 ;
        RECT 372.790 3.670 377.010 4.280 ;
        RECT 377.850 3.670 382.070 4.280 ;
        RECT 382.910 3.670 387.130 4.280 ;
        RECT 387.970 3.670 391.730 4.280 ;
        RECT 392.570 3.670 396.790 4.280 ;
        RECT 397.630 3.670 401.850 4.280 ;
        RECT 402.690 3.670 406.910 4.280 ;
        RECT 407.750 3.670 411.970 4.280 ;
        RECT 412.810 3.670 417.030 4.280 ;
        RECT 417.870 3.670 422.090 4.280 ;
        RECT 422.930 3.670 427.150 4.280 ;
        RECT 427.990 3.670 431.750 4.280 ;
        RECT 432.590 3.670 436.810 4.280 ;
        RECT 437.650 3.670 441.870 4.280 ;
        RECT 442.710 3.670 446.930 4.280 ;
        RECT 447.770 3.670 451.990 4.280 ;
        RECT 452.830 3.670 457.050 4.280 ;
        RECT 457.890 3.670 462.110 4.280 ;
        RECT 462.950 3.670 466.710 4.280 ;
        RECT 467.550 3.670 471.770 4.280 ;
        RECT 472.610 3.670 476.830 4.280 ;
        RECT 477.670 3.670 481.890 4.280 ;
        RECT 482.730 3.670 486.950 4.280 ;
        RECT 487.790 3.670 492.010 4.280 ;
        RECT 492.850 3.670 497.070 4.280 ;
        RECT 497.910 3.670 502.130 4.280 ;
        RECT 502.970 3.670 506.730 4.280 ;
        RECT 507.570 3.670 511.790 4.280 ;
        RECT 512.630 3.670 516.850 4.280 ;
        RECT 517.690 3.670 521.910 4.280 ;
        RECT 522.750 3.670 526.970 4.280 ;
        RECT 527.810 3.670 532.030 4.280 ;
        RECT 532.870 3.670 537.090 4.280 ;
        RECT 537.930 3.670 542.150 4.280 ;
        RECT 542.990 3.670 546.750 4.280 ;
        RECT 547.590 3.670 551.810 4.280 ;
        RECT 552.650 3.670 556.870 4.280 ;
        RECT 557.710 3.670 561.930 4.280 ;
        RECT 562.770 3.670 566.990 4.280 ;
        RECT 567.830 3.670 572.050 4.280 ;
        RECT 572.890 3.670 577.110 4.280 ;
        RECT 577.950 3.670 582.170 4.280 ;
        RECT 583.010 3.670 586.770 4.280 ;
        RECT 587.610 3.670 591.830 4.280 ;
        RECT 592.670 3.670 596.890 4.280 ;
        RECT 597.730 3.670 601.950 4.280 ;
        RECT 602.790 3.670 607.010 4.280 ;
        RECT 607.850 3.670 612.070 4.280 ;
        RECT 612.910 3.670 617.130 4.280 ;
        RECT 617.970 3.670 621.730 4.280 ;
        RECT 622.570 3.670 626.790 4.280 ;
        RECT 627.630 3.670 631.850 4.280 ;
        RECT 632.690 3.670 636.910 4.280 ;
        RECT 637.750 3.670 641.970 4.280 ;
        RECT 642.810 3.670 647.030 4.280 ;
        RECT 647.870 3.670 652.090 4.280 ;
        RECT 652.930 3.670 657.150 4.280 ;
        RECT 657.990 3.670 661.750 4.280 ;
        RECT 662.590 3.670 666.810 4.280 ;
        RECT 667.650 3.670 671.870 4.280 ;
        RECT 672.710 3.670 676.930 4.280 ;
        RECT 677.770 3.670 681.990 4.280 ;
        RECT 682.830 3.670 687.050 4.280 ;
        RECT 687.890 3.670 692.110 4.280 ;
        RECT 692.950 3.670 697.170 4.280 ;
        RECT 698.010 3.670 701.770 4.280 ;
        RECT 702.610 3.670 706.830 4.280 ;
        RECT 707.670 3.670 711.890 4.280 ;
        RECT 712.730 3.670 716.950 4.280 ;
        RECT 717.790 3.670 722.010 4.280 ;
        RECT 722.850 3.670 727.070 4.280 ;
        RECT 727.910 3.670 732.130 4.280 ;
        RECT 732.970 3.670 737.190 4.280 ;
        RECT 738.030 3.670 741.790 4.280 ;
        RECT 742.630 3.670 746.850 4.280 ;
        RECT 747.690 3.670 751.910 4.280 ;
        RECT 752.750 3.670 756.970 4.280 ;
        RECT 757.810 3.670 762.030 4.280 ;
        RECT 762.870 3.670 767.090 4.280 ;
        RECT 767.930 3.670 772.150 4.280 ;
        RECT 772.990 3.670 776.750 4.280 ;
        RECT 777.590 3.670 781.810 4.280 ;
        RECT 782.650 3.670 786.870 4.280 ;
        RECT 787.710 3.670 791.930 4.280 ;
        RECT 792.770 3.670 796.990 4.280 ;
        RECT 797.830 3.670 802.050 4.280 ;
        RECT 802.890 3.670 807.110 4.280 ;
        RECT 807.950 3.670 812.170 4.280 ;
        RECT 813.010 3.670 816.770 4.280 ;
        RECT 817.610 3.670 821.830 4.280 ;
        RECT 822.670 3.670 826.890 4.280 ;
        RECT 827.730 3.670 831.950 4.280 ;
        RECT 832.790 3.670 837.010 4.280 ;
        RECT 837.850 3.670 842.070 4.280 ;
        RECT 842.910 3.670 847.130 4.280 ;
        RECT 847.970 3.670 852.190 4.280 ;
        RECT 853.030 3.670 856.790 4.280 ;
        RECT 857.630 3.670 861.850 4.280 ;
        RECT 862.690 3.670 866.910 4.280 ;
        RECT 867.750 3.670 871.970 4.280 ;
        RECT 872.810 3.670 877.030 4.280 ;
        RECT 877.870 3.670 882.090 4.280 ;
        RECT 882.930 3.670 887.150 4.280 ;
        RECT 887.990 3.670 892.210 4.280 ;
        RECT 893.050 3.670 896.810 4.280 ;
        RECT 897.650 3.670 901.870 4.280 ;
        RECT 902.710 3.670 906.930 4.280 ;
        RECT 907.770 3.670 911.990 4.280 ;
        RECT 912.830 3.670 917.050 4.280 ;
        RECT 917.890 3.670 922.110 4.280 ;
        RECT 922.950 3.670 927.170 4.280 ;
        RECT 928.010 3.670 931.770 4.280 ;
        RECT 932.610 3.670 936.830 4.280 ;
        RECT 937.670 3.670 941.890 4.280 ;
        RECT 942.730 3.670 946.950 4.280 ;
        RECT 947.790 3.670 952.010 4.280 ;
        RECT 952.850 3.670 957.070 4.280 ;
        RECT 957.910 3.670 962.130 4.280 ;
        RECT 962.970 3.670 967.190 4.280 ;
        RECT 968.030 3.670 971.790 4.280 ;
        RECT 972.630 3.670 976.850 4.280 ;
        RECT 977.690 3.670 981.910 4.280 ;
        RECT 982.750 3.670 986.970 4.280 ;
        RECT 987.810 3.670 992.030 4.280 ;
        RECT 992.870 3.670 997.090 4.280 ;
        RECT 997.930 3.670 1002.150 4.280 ;
        RECT 1002.990 3.670 1007.210 4.280 ;
        RECT 1008.050 3.670 1011.810 4.280 ;
        RECT 1012.650 3.670 1016.870 4.280 ;
        RECT 1017.710 3.670 1021.930 4.280 ;
        RECT 1022.770 3.670 1026.990 4.280 ;
        RECT 1027.830 3.670 1032.050 4.280 ;
        RECT 1032.890 3.670 1037.110 4.280 ;
        RECT 1037.950 3.670 1042.170 4.280 ;
        RECT 1043.010 3.670 1047.230 4.280 ;
        RECT 1048.070 3.670 1051.830 4.280 ;
        RECT 1052.670 3.670 1056.890 4.280 ;
        RECT 1057.730 3.670 1061.950 4.280 ;
        RECT 1062.790 3.670 1067.010 4.280 ;
        RECT 1067.850 3.670 1072.070 4.280 ;
        RECT 1072.910 3.670 1077.130 4.280 ;
        RECT 1077.970 3.670 1082.190 4.280 ;
        RECT 1083.030 3.670 1086.790 4.280 ;
        RECT 1087.630 3.670 1091.850 4.280 ;
        RECT 1092.690 3.670 1096.910 4.280 ;
        RECT 1097.750 3.670 1101.970 4.280 ;
        RECT 1102.810 3.670 1107.030 4.280 ;
        RECT 1107.870 3.670 1112.090 4.280 ;
        RECT 1112.930 3.670 1117.150 4.280 ;
        RECT 1117.990 3.670 1122.210 4.280 ;
        RECT 1123.050 3.670 1126.810 4.280 ;
        RECT 1127.650 3.670 1131.870 4.280 ;
        RECT 1132.710 3.670 1136.930 4.280 ;
        RECT 1137.770 3.670 1141.990 4.280 ;
        RECT 1142.830 3.670 1147.050 4.280 ;
        RECT 1147.890 3.670 1152.110 4.280 ;
        RECT 1152.950 3.670 1157.170 4.280 ;
        RECT 1158.010 3.670 1162.230 4.280 ;
        RECT 1163.070 3.670 1166.830 4.280 ;
        RECT 1167.670 3.670 1171.890 4.280 ;
        RECT 1172.730 3.670 1176.950 4.280 ;
        RECT 1177.790 3.670 1182.010 4.280 ;
        RECT 1182.850 3.670 1187.070 4.280 ;
        RECT 1187.910 3.670 1192.130 4.280 ;
        RECT 1192.970 3.670 1197.190 4.280 ;
      LAYER met3 ;
        RECT 4.000 1188.960 1195.600 1189.825 ;
        RECT 4.000 1186.960 1196.000 1188.960 ;
        RECT 4.400 1185.560 1196.000 1186.960 ;
        RECT 4.000 1170.640 1196.000 1185.560 ;
        RECT 4.000 1169.240 1195.600 1170.640 ;
        RECT 4.000 1160.440 1196.000 1169.240 ;
        RECT 4.400 1159.040 1196.000 1160.440 ;
        RECT 4.000 1150.240 1196.000 1159.040 ;
        RECT 4.000 1148.840 1195.600 1150.240 ;
        RECT 4.000 1133.920 1196.000 1148.840 ;
        RECT 4.400 1132.520 1196.000 1133.920 ;
        RECT 4.000 1130.520 1196.000 1132.520 ;
        RECT 4.000 1129.120 1195.600 1130.520 ;
        RECT 4.000 1110.120 1196.000 1129.120 ;
        RECT 4.000 1108.720 1195.600 1110.120 ;
        RECT 4.000 1107.400 1196.000 1108.720 ;
        RECT 4.400 1106.000 1196.000 1107.400 ;
        RECT 4.000 1090.400 1196.000 1106.000 ;
        RECT 4.000 1089.000 1195.600 1090.400 ;
        RECT 4.000 1080.200 1196.000 1089.000 ;
        RECT 4.400 1078.800 1196.000 1080.200 ;
        RECT 4.000 1070.680 1196.000 1078.800 ;
        RECT 4.000 1069.280 1195.600 1070.680 ;
        RECT 4.000 1053.680 1196.000 1069.280 ;
        RECT 4.400 1052.280 1196.000 1053.680 ;
        RECT 4.000 1050.280 1196.000 1052.280 ;
        RECT 4.000 1048.880 1195.600 1050.280 ;
        RECT 4.000 1030.560 1196.000 1048.880 ;
        RECT 4.000 1029.160 1195.600 1030.560 ;
        RECT 4.000 1027.160 1196.000 1029.160 ;
        RECT 4.400 1025.760 1196.000 1027.160 ;
        RECT 4.000 1010.160 1196.000 1025.760 ;
        RECT 4.000 1008.760 1195.600 1010.160 ;
        RECT 4.000 1000.640 1196.000 1008.760 ;
        RECT 4.400 999.240 1196.000 1000.640 ;
        RECT 4.000 990.440 1196.000 999.240 ;
        RECT 4.000 989.040 1195.600 990.440 ;
        RECT 4.000 974.120 1196.000 989.040 ;
        RECT 4.400 972.720 1196.000 974.120 ;
        RECT 4.000 970.720 1196.000 972.720 ;
        RECT 4.000 969.320 1195.600 970.720 ;
        RECT 4.000 950.320 1196.000 969.320 ;
        RECT 4.000 948.920 1195.600 950.320 ;
        RECT 4.000 946.920 1196.000 948.920 ;
        RECT 4.400 945.520 1196.000 946.920 ;
        RECT 4.000 930.600 1196.000 945.520 ;
        RECT 4.000 929.200 1195.600 930.600 ;
        RECT 4.000 920.400 1196.000 929.200 ;
        RECT 4.400 919.000 1196.000 920.400 ;
        RECT 4.000 910.200 1196.000 919.000 ;
        RECT 4.000 908.800 1195.600 910.200 ;
        RECT 4.000 893.880 1196.000 908.800 ;
        RECT 4.400 892.480 1196.000 893.880 ;
        RECT 4.000 890.480 1196.000 892.480 ;
        RECT 4.000 889.080 1195.600 890.480 ;
        RECT 4.000 870.080 1196.000 889.080 ;
        RECT 4.000 868.680 1195.600 870.080 ;
        RECT 4.000 867.360 1196.000 868.680 ;
        RECT 4.400 865.960 1196.000 867.360 ;
        RECT 4.000 850.360 1196.000 865.960 ;
        RECT 4.000 848.960 1195.600 850.360 ;
        RECT 4.000 840.160 1196.000 848.960 ;
        RECT 4.400 838.760 1196.000 840.160 ;
        RECT 4.000 830.640 1196.000 838.760 ;
        RECT 4.000 829.240 1195.600 830.640 ;
        RECT 4.000 813.640 1196.000 829.240 ;
        RECT 4.400 812.240 1196.000 813.640 ;
        RECT 4.000 810.240 1196.000 812.240 ;
        RECT 4.000 808.840 1195.600 810.240 ;
        RECT 4.000 790.520 1196.000 808.840 ;
        RECT 4.000 789.120 1195.600 790.520 ;
        RECT 4.000 787.120 1196.000 789.120 ;
        RECT 4.400 785.720 1196.000 787.120 ;
        RECT 4.000 770.120 1196.000 785.720 ;
        RECT 4.000 768.720 1195.600 770.120 ;
        RECT 4.000 760.600 1196.000 768.720 ;
        RECT 4.400 759.200 1196.000 760.600 ;
        RECT 4.000 750.400 1196.000 759.200 ;
        RECT 4.000 749.000 1195.600 750.400 ;
        RECT 4.000 734.080 1196.000 749.000 ;
        RECT 4.400 732.680 1196.000 734.080 ;
        RECT 4.000 730.680 1196.000 732.680 ;
        RECT 4.000 729.280 1195.600 730.680 ;
        RECT 4.000 710.280 1196.000 729.280 ;
        RECT 4.000 708.880 1195.600 710.280 ;
        RECT 4.000 706.880 1196.000 708.880 ;
        RECT 4.400 705.480 1196.000 706.880 ;
        RECT 4.000 690.560 1196.000 705.480 ;
        RECT 4.000 689.160 1195.600 690.560 ;
        RECT 4.000 680.360 1196.000 689.160 ;
        RECT 4.400 678.960 1196.000 680.360 ;
        RECT 4.000 670.160 1196.000 678.960 ;
        RECT 4.000 668.760 1195.600 670.160 ;
        RECT 4.000 653.840 1196.000 668.760 ;
        RECT 4.400 652.440 1196.000 653.840 ;
        RECT 4.000 650.440 1196.000 652.440 ;
        RECT 4.000 649.040 1195.600 650.440 ;
        RECT 4.000 630.040 1196.000 649.040 ;
        RECT 4.000 628.640 1195.600 630.040 ;
        RECT 4.000 627.320 1196.000 628.640 ;
        RECT 4.400 625.920 1196.000 627.320 ;
        RECT 4.000 610.320 1196.000 625.920 ;
        RECT 4.000 608.920 1195.600 610.320 ;
        RECT 4.000 600.120 1196.000 608.920 ;
        RECT 4.400 598.720 1196.000 600.120 ;
        RECT 4.000 590.600 1196.000 598.720 ;
        RECT 4.000 589.200 1195.600 590.600 ;
        RECT 4.000 573.600 1196.000 589.200 ;
        RECT 4.400 572.200 1196.000 573.600 ;
        RECT 4.000 570.200 1196.000 572.200 ;
        RECT 4.000 568.800 1195.600 570.200 ;
        RECT 4.000 550.480 1196.000 568.800 ;
        RECT 4.000 549.080 1195.600 550.480 ;
        RECT 4.000 547.080 1196.000 549.080 ;
        RECT 4.400 545.680 1196.000 547.080 ;
        RECT 4.000 530.080 1196.000 545.680 ;
        RECT 4.000 528.680 1195.600 530.080 ;
        RECT 4.000 520.560 1196.000 528.680 ;
        RECT 4.400 519.160 1196.000 520.560 ;
        RECT 4.000 510.360 1196.000 519.160 ;
        RECT 4.000 508.960 1195.600 510.360 ;
        RECT 4.000 494.040 1196.000 508.960 ;
        RECT 4.400 492.640 1196.000 494.040 ;
        RECT 4.000 490.640 1196.000 492.640 ;
        RECT 4.000 489.240 1195.600 490.640 ;
        RECT 4.000 470.240 1196.000 489.240 ;
        RECT 4.000 468.840 1195.600 470.240 ;
        RECT 4.000 466.840 1196.000 468.840 ;
        RECT 4.400 465.440 1196.000 466.840 ;
        RECT 4.000 450.520 1196.000 465.440 ;
        RECT 4.000 449.120 1195.600 450.520 ;
        RECT 4.000 440.320 1196.000 449.120 ;
        RECT 4.400 438.920 1196.000 440.320 ;
        RECT 4.000 430.120 1196.000 438.920 ;
        RECT 4.000 428.720 1195.600 430.120 ;
        RECT 4.000 413.800 1196.000 428.720 ;
        RECT 4.400 412.400 1196.000 413.800 ;
        RECT 4.000 410.400 1196.000 412.400 ;
        RECT 4.000 409.000 1195.600 410.400 ;
        RECT 4.000 390.000 1196.000 409.000 ;
        RECT 4.000 388.600 1195.600 390.000 ;
        RECT 4.000 387.280 1196.000 388.600 ;
        RECT 4.400 385.880 1196.000 387.280 ;
        RECT 4.000 370.280 1196.000 385.880 ;
        RECT 4.000 368.880 1195.600 370.280 ;
        RECT 4.000 360.080 1196.000 368.880 ;
        RECT 4.400 358.680 1196.000 360.080 ;
        RECT 4.000 350.560 1196.000 358.680 ;
        RECT 4.000 349.160 1195.600 350.560 ;
        RECT 4.000 333.560 1196.000 349.160 ;
        RECT 4.400 332.160 1196.000 333.560 ;
        RECT 4.000 330.160 1196.000 332.160 ;
        RECT 4.000 328.760 1195.600 330.160 ;
        RECT 4.000 310.440 1196.000 328.760 ;
        RECT 4.000 309.040 1195.600 310.440 ;
        RECT 4.000 307.040 1196.000 309.040 ;
        RECT 4.400 305.640 1196.000 307.040 ;
        RECT 4.000 290.040 1196.000 305.640 ;
        RECT 4.000 288.640 1195.600 290.040 ;
        RECT 4.000 280.520 1196.000 288.640 ;
        RECT 4.400 279.120 1196.000 280.520 ;
        RECT 4.000 270.320 1196.000 279.120 ;
        RECT 4.000 268.920 1195.600 270.320 ;
        RECT 4.000 254.000 1196.000 268.920 ;
        RECT 4.400 252.600 1196.000 254.000 ;
        RECT 4.000 250.600 1196.000 252.600 ;
        RECT 4.000 249.200 1195.600 250.600 ;
        RECT 4.000 230.200 1196.000 249.200 ;
        RECT 4.000 228.800 1195.600 230.200 ;
        RECT 4.000 226.800 1196.000 228.800 ;
        RECT 4.400 225.400 1196.000 226.800 ;
        RECT 4.000 210.480 1196.000 225.400 ;
        RECT 4.000 209.080 1195.600 210.480 ;
        RECT 4.000 200.280 1196.000 209.080 ;
        RECT 4.400 198.880 1196.000 200.280 ;
        RECT 4.000 190.080 1196.000 198.880 ;
        RECT 4.000 188.680 1195.600 190.080 ;
        RECT 4.000 173.760 1196.000 188.680 ;
        RECT 4.400 172.360 1196.000 173.760 ;
        RECT 4.000 170.360 1196.000 172.360 ;
        RECT 4.000 168.960 1195.600 170.360 ;
        RECT 4.000 149.960 1196.000 168.960 ;
        RECT 4.000 148.560 1195.600 149.960 ;
        RECT 4.000 147.240 1196.000 148.560 ;
        RECT 4.400 145.840 1196.000 147.240 ;
        RECT 4.000 130.240 1196.000 145.840 ;
        RECT 4.000 128.840 1195.600 130.240 ;
        RECT 4.000 120.040 1196.000 128.840 ;
        RECT 4.400 118.640 1196.000 120.040 ;
        RECT 4.000 110.520 1196.000 118.640 ;
        RECT 4.000 109.120 1195.600 110.520 ;
        RECT 4.000 93.520 1196.000 109.120 ;
        RECT 4.400 92.120 1196.000 93.520 ;
        RECT 4.000 90.120 1196.000 92.120 ;
        RECT 4.000 88.720 1195.600 90.120 ;
        RECT 4.000 70.400 1196.000 88.720 ;
        RECT 4.000 69.000 1195.600 70.400 ;
        RECT 4.000 67.000 1196.000 69.000 ;
        RECT 4.400 65.600 1196.000 67.000 ;
        RECT 4.000 50.000 1196.000 65.600 ;
        RECT 4.000 48.600 1195.600 50.000 ;
        RECT 4.000 40.480 1196.000 48.600 ;
        RECT 4.400 39.080 1196.000 40.480 ;
        RECT 4.000 30.280 1196.000 39.080 ;
        RECT 4.000 28.880 1195.600 30.280 ;
        RECT 4.000 13.960 1196.000 28.880 ;
        RECT 4.400 12.560 1196.000 13.960 ;
        RECT 4.000 10.560 1196.000 12.560 ;
        RECT 4.000 9.695 1195.600 10.560 ;
      LAYER met4 ;
        RECT 517.335 219.135 558.240 1187.785 ;
        RECT 560.640 219.135 635.040 1187.785 ;
        RECT 637.440 219.135 711.840 1187.785 ;
        RECT 714.240 219.135 788.640 1187.785 ;
        RECT 791.040 219.135 865.440 1187.785 ;
        RECT 867.840 219.135 942.240 1187.785 ;
        RECT 944.640 219.135 1019.040 1187.785 ;
        RECT 1021.440 219.135 1067.825 1187.785 ;
  END
END ibex_top
END LIBRARY

