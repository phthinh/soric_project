magic
tech sky130A
magscale 1 2
timestamp 1640739197
<< obsli1 >>
rect 1104 1241 259135 258179
<< obsm1 >>
rect 1104 1235 259242 258188
<< metal2 >>
rect 1766 259200 1822 260000
rect 5354 259200 5410 260000
rect 9034 259200 9090 260000
rect 12714 259200 12770 260000
rect 16394 259200 16450 260000
rect 20074 259200 20130 260000
rect 23662 259200 23718 260000
rect 27342 259200 27398 260000
rect 31022 259200 31078 260000
rect 34702 259200 34758 260000
rect 38382 259200 38438 260000
rect 41970 259200 42026 260000
rect 45650 259200 45706 260000
rect 49330 259200 49386 260000
rect 53010 259200 53066 260000
rect 56690 259200 56746 260000
rect 60278 259200 60334 260000
rect 63958 259200 64014 260000
rect 67638 259200 67694 260000
rect 71318 259200 71374 260000
rect 74998 259200 75054 260000
rect 78586 259200 78642 260000
rect 82266 259200 82322 260000
rect 85946 259200 86002 260000
rect 89626 259200 89682 260000
rect 93306 259200 93362 260000
rect 96894 259200 96950 260000
rect 100574 259200 100630 260000
rect 104254 259200 104310 260000
rect 107934 259200 107990 260000
rect 111614 259200 111670 260000
rect 115202 259200 115258 260000
rect 118882 259200 118938 260000
rect 122562 259200 122618 260000
rect 126242 259200 126298 260000
rect 129922 259200 129978 260000
rect 133510 259200 133566 260000
rect 137190 259200 137246 260000
rect 140870 259200 140926 260000
rect 144550 259200 144606 260000
rect 148230 259200 148286 260000
rect 151818 259200 151874 260000
rect 155498 259200 155554 260000
rect 159178 259200 159234 260000
rect 162858 259200 162914 260000
rect 166538 259200 166594 260000
rect 170126 259200 170182 260000
rect 173806 259200 173862 260000
rect 177486 259200 177542 260000
rect 181166 259200 181222 260000
rect 184846 259200 184902 260000
rect 188434 259200 188490 260000
rect 192114 259200 192170 260000
rect 195794 259200 195850 260000
rect 199474 259200 199530 260000
rect 203154 259200 203210 260000
rect 206742 259200 206798 260000
rect 210422 259200 210478 260000
rect 214102 259200 214158 260000
rect 217782 259200 217838 260000
rect 221462 259200 221518 260000
rect 225050 259200 225106 260000
rect 228730 259200 228786 260000
rect 232410 259200 232466 260000
rect 236090 259200 236146 260000
rect 239770 259200 239826 260000
rect 243358 259200 243414 260000
rect 247038 259200 247094 260000
rect 250718 259200 250774 260000
rect 254398 259200 254454 260000
rect 258078 259200 258134 260000
rect 662 0 718 800
rect 2042 0 2098 800
rect 3422 0 3478 800
rect 4894 0 4950 800
rect 6274 0 6330 800
rect 7746 0 7802 800
rect 9126 0 9182 800
rect 10598 0 10654 800
rect 11978 0 12034 800
rect 13358 0 13414 800
rect 14830 0 14886 800
rect 16210 0 16266 800
rect 17682 0 17738 800
rect 19062 0 19118 800
rect 20534 0 20590 800
rect 21914 0 21970 800
rect 23386 0 23442 800
rect 24766 0 24822 800
rect 26146 0 26202 800
rect 27618 0 27674 800
rect 28998 0 29054 800
rect 30470 0 30526 800
rect 31850 0 31906 800
rect 33322 0 33378 800
rect 34702 0 34758 800
rect 36174 0 36230 800
rect 37554 0 37610 800
rect 38934 0 38990 800
rect 40406 0 40462 800
rect 41786 0 41842 800
rect 43258 0 43314 800
rect 44638 0 44694 800
rect 46110 0 46166 800
rect 47490 0 47546 800
rect 48962 0 49018 800
rect 50342 0 50398 800
rect 51722 0 51778 800
rect 53194 0 53250 800
rect 54574 0 54630 800
rect 56046 0 56102 800
rect 57426 0 57482 800
rect 58898 0 58954 800
rect 60278 0 60334 800
rect 61750 0 61806 800
rect 63130 0 63186 800
rect 64510 0 64566 800
rect 65982 0 66038 800
rect 67362 0 67418 800
rect 68834 0 68890 800
rect 70214 0 70270 800
rect 71686 0 71742 800
rect 73066 0 73122 800
rect 74538 0 74594 800
rect 75918 0 75974 800
rect 77298 0 77354 800
rect 78770 0 78826 800
rect 80150 0 80206 800
rect 81622 0 81678 800
rect 83002 0 83058 800
rect 84474 0 84530 800
rect 85854 0 85910 800
rect 87326 0 87382 800
rect 88706 0 88762 800
rect 90086 0 90142 800
rect 91558 0 91614 800
rect 92938 0 92994 800
rect 94410 0 94466 800
rect 95790 0 95846 800
rect 97262 0 97318 800
rect 98642 0 98698 800
rect 100022 0 100078 800
rect 101494 0 101550 800
rect 102874 0 102930 800
rect 104346 0 104402 800
rect 105726 0 105782 800
rect 107198 0 107254 800
rect 108578 0 108634 800
rect 110050 0 110106 800
rect 111430 0 111486 800
rect 112810 0 112866 800
rect 114282 0 114338 800
rect 115662 0 115718 800
rect 117134 0 117190 800
rect 118514 0 118570 800
rect 119986 0 120042 800
rect 121366 0 121422 800
rect 122838 0 122894 800
rect 124218 0 124274 800
rect 125598 0 125654 800
rect 127070 0 127126 800
rect 128450 0 128506 800
rect 129922 0 129978 800
rect 131302 0 131358 800
rect 132774 0 132830 800
rect 134154 0 134210 800
rect 135626 0 135682 800
rect 137006 0 137062 800
rect 138386 0 138442 800
rect 139858 0 139914 800
rect 141238 0 141294 800
rect 142710 0 142766 800
rect 144090 0 144146 800
rect 145562 0 145618 800
rect 146942 0 146998 800
rect 148414 0 148470 800
rect 149794 0 149850 800
rect 151174 0 151230 800
rect 152646 0 152702 800
rect 154026 0 154082 800
rect 155498 0 155554 800
rect 156878 0 156934 800
rect 158350 0 158406 800
rect 159730 0 159786 800
rect 161202 0 161258 800
rect 162582 0 162638 800
rect 163962 0 164018 800
rect 165434 0 165490 800
rect 166814 0 166870 800
rect 168286 0 168342 800
rect 169666 0 169722 800
rect 171138 0 171194 800
rect 172518 0 172574 800
rect 173990 0 174046 800
rect 175370 0 175426 800
rect 176750 0 176806 800
rect 178222 0 178278 800
rect 179602 0 179658 800
rect 181074 0 181130 800
rect 182454 0 182510 800
rect 183926 0 183982 800
rect 185306 0 185362 800
rect 186686 0 186742 800
rect 188158 0 188214 800
rect 189538 0 189594 800
rect 191010 0 191066 800
rect 192390 0 192446 800
rect 193862 0 193918 800
rect 195242 0 195298 800
rect 196714 0 196770 800
rect 198094 0 198150 800
rect 199474 0 199530 800
rect 200946 0 201002 800
rect 202326 0 202382 800
rect 203798 0 203854 800
rect 205178 0 205234 800
rect 206650 0 206706 800
rect 208030 0 208086 800
rect 209502 0 209558 800
rect 210882 0 210938 800
rect 212262 0 212318 800
rect 213734 0 213790 800
rect 215114 0 215170 800
rect 216586 0 216642 800
rect 217966 0 218022 800
rect 219438 0 219494 800
rect 220818 0 220874 800
rect 222290 0 222346 800
rect 223670 0 223726 800
rect 225050 0 225106 800
rect 226522 0 226578 800
rect 227902 0 227958 800
rect 229374 0 229430 800
rect 230754 0 230810 800
rect 232226 0 232282 800
rect 233606 0 233662 800
rect 235078 0 235134 800
rect 236458 0 236514 800
rect 237838 0 237894 800
rect 239310 0 239366 800
rect 240690 0 240746 800
rect 242162 0 242218 800
rect 243542 0 243598 800
rect 245014 0 245070 800
rect 246394 0 246450 800
rect 247866 0 247922 800
rect 249246 0 249302 800
rect 250626 0 250682 800
rect 252098 0 252154 800
rect 253478 0 253534 800
rect 254950 0 255006 800
rect 256330 0 256386 800
rect 257802 0 257858 800
rect 259182 0 259238 800
<< obsm2 >>
rect 1398 259144 1710 259298
rect 1878 259144 5298 259298
rect 5466 259144 8978 259298
rect 9146 259144 12658 259298
rect 12826 259144 16338 259298
rect 16506 259144 20018 259298
rect 20186 259144 23606 259298
rect 23774 259144 27286 259298
rect 27454 259144 30966 259298
rect 31134 259144 34646 259298
rect 34814 259144 38326 259298
rect 38494 259144 41914 259298
rect 42082 259144 45594 259298
rect 45762 259144 49274 259298
rect 49442 259144 52954 259298
rect 53122 259144 56634 259298
rect 56802 259144 60222 259298
rect 60390 259144 63902 259298
rect 64070 259144 67582 259298
rect 67750 259144 71262 259298
rect 71430 259144 74942 259298
rect 75110 259144 78530 259298
rect 78698 259144 82210 259298
rect 82378 259144 85890 259298
rect 86058 259144 89570 259298
rect 89738 259144 93250 259298
rect 93418 259144 96838 259298
rect 97006 259144 100518 259298
rect 100686 259144 104198 259298
rect 104366 259144 107878 259298
rect 108046 259144 111558 259298
rect 111726 259144 115146 259298
rect 115314 259144 118826 259298
rect 118994 259144 122506 259298
rect 122674 259144 126186 259298
rect 126354 259144 129866 259298
rect 130034 259144 133454 259298
rect 133622 259144 137134 259298
rect 137302 259144 140814 259298
rect 140982 259144 144494 259298
rect 144662 259144 148174 259298
rect 148342 259144 151762 259298
rect 151930 259144 155442 259298
rect 155610 259144 159122 259298
rect 159290 259144 162802 259298
rect 162970 259144 166482 259298
rect 166650 259144 170070 259298
rect 170238 259144 173750 259298
rect 173918 259144 177430 259298
rect 177598 259144 181110 259298
rect 181278 259144 184790 259298
rect 184958 259144 188378 259298
rect 188546 259144 192058 259298
rect 192226 259144 195738 259298
rect 195906 259144 199418 259298
rect 199586 259144 203098 259298
rect 203266 259144 206686 259298
rect 206854 259144 210366 259298
rect 210534 259144 214046 259298
rect 214214 259144 217726 259298
rect 217894 259144 221406 259298
rect 221574 259144 224994 259298
rect 225162 259144 228674 259298
rect 228842 259144 232354 259298
rect 232522 259144 236034 259298
rect 236202 259144 239714 259298
rect 239882 259144 243302 259298
rect 243470 259144 246982 259298
rect 247150 259144 250662 259298
rect 250830 259144 254342 259298
rect 254510 259144 258022 259298
rect 258190 259144 259236 259298
rect 1398 856 259236 259144
rect 1398 734 1986 856
rect 2154 734 3366 856
rect 3534 734 4838 856
rect 5006 734 6218 856
rect 6386 734 7690 856
rect 7858 734 9070 856
rect 9238 734 10542 856
rect 10710 734 11922 856
rect 12090 734 13302 856
rect 13470 734 14774 856
rect 14942 734 16154 856
rect 16322 734 17626 856
rect 17794 734 19006 856
rect 19174 734 20478 856
rect 20646 734 21858 856
rect 22026 734 23330 856
rect 23498 734 24710 856
rect 24878 734 26090 856
rect 26258 734 27562 856
rect 27730 734 28942 856
rect 29110 734 30414 856
rect 30582 734 31794 856
rect 31962 734 33266 856
rect 33434 734 34646 856
rect 34814 734 36118 856
rect 36286 734 37498 856
rect 37666 734 38878 856
rect 39046 734 40350 856
rect 40518 734 41730 856
rect 41898 734 43202 856
rect 43370 734 44582 856
rect 44750 734 46054 856
rect 46222 734 47434 856
rect 47602 734 48906 856
rect 49074 734 50286 856
rect 50454 734 51666 856
rect 51834 734 53138 856
rect 53306 734 54518 856
rect 54686 734 55990 856
rect 56158 734 57370 856
rect 57538 734 58842 856
rect 59010 734 60222 856
rect 60390 734 61694 856
rect 61862 734 63074 856
rect 63242 734 64454 856
rect 64622 734 65926 856
rect 66094 734 67306 856
rect 67474 734 68778 856
rect 68946 734 70158 856
rect 70326 734 71630 856
rect 71798 734 73010 856
rect 73178 734 74482 856
rect 74650 734 75862 856
rect 76030 734 77242 856
rect 77410 734 78714 856
rect 78882 734 80094 856
rect 80262 734 81566 856
rect 81734 734 82946 856
rect 83114 734 84418 856
rect 84586 734 85798 856
rect 85966 734 87270 856
rect 87438 734 88650 856
rect 88818 734 90030 856
rect 90198 734 91502 856
rect 91670 734 92882 856
rect 93050 734 94354 856
rect 94522 734 95734 856
rect 95902 734 97206 856
rect 97374 734 98586 856
rect 98754 734 99966 856
rect 100134 734 101438 856
rect 101606 734 102818 856
rect 102986 734 104290 856
rect 104458 734 105670 856
rect 105838 734 107142 856
rect 107310 734 108522 856
rect 108690 734 109994 856
rect 110162 734 111374 856
rect 111542 734 112754 856
rect 112922 734 114226 856
rect 114394 734 115606 856
rect 115774 734 117078 856
rect 117246 734 118458 856
rect 118626 734 119930 856
rect 120098 734 121310 856
rect 121478 734 122782 856
rect 122950 734 124162 856
rect 124330 734 125542 856
rect 125710 734 127014 856
rect 127182 734 128394 856
rect 128562 734 129866 856
rect 130034 734 131246 856
rect 131414 734 132718 856
rect 132886 734 134098 856
rect 134266 734 135570 856
rect 135738 734 136950 856
rect 137118 734 138330 856
rect 138498 734 139802 856
rect 139970 734 141182 856
rect 141350 734 142654 856
rect 142822 734 144034 856
rect 144202 734 145506 856
rect 145674 734 146886 856
rect 147054 734 148358 856
rect 148526 734 149738 856
rect 149906 734 151118 856
rect 151286 734 152590 856
rect 152758 734 153970 856
rect 154138 734 155442 856
rect 155610 734 156822 856
rect 156990 734 158294 856
rect 158462 734 159674 856
rect 159842 734 161146 856
rect 161314 734 162526 856
rect 162694 734 163906 856
rect 164074 734 165378 856
rect 165546 734 166758 856
rect 166926 734 168230 856
rect 168398 734 169610 856
rect 169778 734 171082 856
rect 171250 734 172462 856
rect 172630 734 173934 856
rect 174102 734 175314 856
rect 175482 734 176694 856
rect 176862 734 178166 856
rect 178334 734 179546 856
rect 179714 734 181018 856
rect 181186 734 182398 856
rect 182566 734 183870 856
rect 184038 734 185250 856
rect 185418 734 186630 856
rect 186798 734 188102 856
rect 188270 734 189482 856
rect 189650 734 190954 856
rect 191122 734 192334 856
rect 192502 734 193806 856
rect 193974 734 195186 856
rect 195354 734 196658 856
rect 196826 734 198038 856
rect 198206 734 199418 856
rect 199586 734 200890 856
rect 201058 734 202270 856
rect 202438 734 203742 856
rect 203910 734 205122 856
rect 205290 734 206594 856
rect 206762 734 207974 856
rect 208142 734 209446 856
rect 209614 734 210826 856
rect 210994 734 212206 856
rect 212374 734 213678 856
rect 213846 734 215058 856
rect 215226 734 216530 856
rect 216698 734 217910 856
rect 218078 734 219382 856
rect 219550 734 220762 856
rect 220930 734 222234 856
rect 222402 734 223614 856
rect 223782 734 224994 856
rect 225162 734 226466 856
rect 226634 734 227846 856
rect 228014 734 229318 856
rect 229486 734 230698 856
rect 230866 734 232170 856
rect 232338 734 233550 856
rect 233718 734 235022 856
rect 235190 734 236402 856
rect 236570 734 237782 856
rect 237950 734 239254 856
rect 239422 734 240634 856
rect 240802 734 242106 856
rect 242274 734 243486 856
rect 243654 734 244958 856
rect 245126 734 246338 856
rect 246506 734 247810 856
rect 247978 734 249190 856
rect 249358 734 250570 856
rect 250738 734 252042 856
rect 252210 734 253422 856
rect 253590 734 254894 856
rect 255062 734 256274 856
rect 256442 734 257746 856
rect 257914 734 259126 856
<< metal3 >>
rect 0 258136 800 258256
rect 259200 258136 260000 258256
rect 259200 254736 260000 254856
rect 0 254464 800 254584
rect 259200 251336 260000 251456
rect 0 250792 800 250912
rect 259200 247936 260000 248056
rect 0 247120 800 247240
rect 259200 244536 260000 244656
rect 0 243448 800 243568
rect 259200 241136 260000 241256
rect 0 239776 800 239896
rect 259200 237600 260000 237720
rect 0 236104 800 236224
rect 259200 234200 260000 234320
rect 0 232432 800 232552
rect 259200 230800 260000 230920
rect 0 228760 800 228880
rect 259200 227400 260000 227520
rect 0 225088 800 225208
rect 259200 224000 260000 224120
rect 0 221416 800 221536
rect 259200 220600 260000 220720
rect 0 217744 800 217864
rect 259200 217064 260000 217184
rect 0 214072 800 214192
rect 259200 213664 260000 213784
rect 0 210400 800 210520
rect 259200 210264 260000 210384
rect 0 206864 800 206984
rect 259200 206864 260000 206984
rect 259200 203464 260000 203584
rect 0 203192 800 203312
rect 259200 200064 260000 200184
rect 0 199520 800 199640
rect 259200 196664 260000 196784
rect 0 195848 800 195968
rect 259200 193128 260000 193248
rect 0 192176 800 192296
rect 259200 189728 260000 189848
rect 0 188504 800 188624
rect 259200 186328 260000 186448
rect 0 184832 800 184952
rect 259200 182928 260000 183048
rect 0 181160 800 181280
rect 259200 179528 260000 179648
rect 0 177488 800 177608
rect 259200 176128 260000 176248
rect 0 173816 800 173936
rect 259200 172592 260000 172712
rect 0 170144 800 170264
rect 259200 169192 260000 169312
rect 0 166472 800 166592
rect 259200 165792 260000 165912
rect 0 162800 800 162920
rect 259200 162392 260000 162512
rect 0 159128 800 159248
rect 259200 158992 260000 159112
rect 0 155592 800 155712
rect 259200 155592 260000 155712
rect 0 151920 800 152040
rect 259200 152056 260000 152176
rect 259200 148656 260000 148776
rect 0 148248 800 148368
rect 259200 145256 260000 145376
rect 0 144576 800 144696
rect 259200 141856 260000 141976
rect 0 140904 800 141024
rect 259200 138456 260000 138576
rect 0 137232 800 137352
rect 259200 135056 260000 135176
rect 0 133560 800 133680
rect 259200 131656 260000 131776
rect 0 129888 800 130008
rect 259200 128120 260000 128240
rect 0 126216 800 126336
rect 259200 124720 260000 124840
rect 0 122544 800 122664
rect 259200 121320 260000 121440
rect 0 118872 800 118992
rect 259200 117920 260000 118040
rect 0 115200 800 115320
rect 259200 114520 260000 114640
rect 0 111528 800 111648
rect 259200 111120 260000 111240
rect 0 107856 800 107976
rect 259200 107584 260000 107704
rect 0 104320 800 104440
rect 259200 104184 260000 104304
rect 0 100648 800 100768
rect 259200 100784 260000 100904
rect 259200 97384 260000 97504
rect 0 96976 800 97096
rect 259200 93984 260000 94104
rect 0 93304 800 93424
rect 259200 90584 260000 90704
rect 0 89632 800 89752
rect 259200 87048 260000 87168
rect 0 85960 800 86080
rect 259200 83648 260000 83768
rect 0 82288 800 82408
rect 259200 80248 260000 80368
rect 0 78616 800 78736
rect 259200 76848 260000 76968
rect 0 74944 800 75064
rect 259200 73448 260000 73568
rect 0 71272 800 71392
rect 259200 70048 260000 70168
rect 0 67600 800 67720
rect 259200 66648 260000 66768
rect 0 63928 800 64048
rect 259200 63112 260000 63232
rect 0 60256 800 60376
rect 259200 59712 260000 59832
rect 0 56584 800 56704
rect 259200 56312 260000 56432
rect 0 53048 800 53168
rect 259200 52912 260000 53032
rect 0 49376 800 49496
rect 259200 49512 260000 49632
rect 259200 46112 260000 46232
rect 0 45704 800 45824
rect 259200 42576 260000 42696
rect 0 42032 800 42152
rect 259200 39176 260000 39296
rect 0 38360 800 38480
rect 259200 35776 260000 35896
rect 0 34688 800 34808
rect 259200 32376 260000 32496
rect 0 31016 800 31136
rect 259200 28976 260000 29096
rect 0 27344 800 27464
rect 259200 25576 260000 25696
rect 0 23672 800 23792
rect 259200 22040 260000 22160
rect 0 20000 800 20120
rect 259200 18640 260000 18760
rect 0 16328 800 16448
rect 259200 15240 260000 15360
rect 0 12656 800 12776
rect 259200 11840 260000 11960
rect 0 8984 800 9104
rect 259200 8440 260000 8560
rect 0 5312 800 5432
rect 259200 5040 260000 5160
rect 0 1776 800 1896
rect 259200 1640 260000 1760
<< obsm3 >>
rect 880 258056 259120 258229
rect 800 254936 259200 258056
rect 800 254664 259120 254936
rect 880 254656 259120 254664
rect 880 254384 259200 254656
rect 800 251536 259200 254384
rect 800 251256 259120 251536
rect 800 250992 259200 251256
rect 880 250712 259200 250992
rect 800 248136 259200 250712
rect 800 247856 259120 248136
rect 800 247320 259200 247856
rect 880 247040 259200 247320
rect 800 244736 259200 247040
rect 800 244456 259120 244736
rect 800 243648 259200 244456
rect 880 243368 259200 243648
rect 800 241336 259200 243368
rect 800 241056 259120 241336
rect 800 239976 259200 241056
rect 880 239696 259200 239976
rect 800 237800 259200 239696
rect 800 237520 259120 237800
rect 800 236304 259200 237520
rect 880 236024 259200 236304
rect 800 234400 259200 236024
rect 800 234120 259120 234400
rect 800 232632 259200 234120
rect 880 232352 259200 232632
rect 800 231000 259200 232352
rect 800 230720 259120 231000
rect 800 228960 259200 230720
rect 880 228680 259200 228960
rect 800 227600 259200 228680
rect 800 227320 259120 227600
rect 800 225288 259200 227320
rect 880 225008 259200 225288
rect 800 224200 259200 225008
rect 800 223920 259120 224200
rect 800 221616 259200 223920
rect 880 221336 259200 221616
rect 800 220800 259200 221336
rect 800 220520 259120 220800
rect 800 217944 259200 220520
rect 880 217664 259200 217944
rect 800 217264 259200 217664
rect 800 216984 259120 217264
rect 800 214272 259200 216984
rect 880 213992 259200 214272
rect 800 213864 259200 213992
rect 800 213584 259120 213864
rect 800 210600 259200 213584
rect 880 210464 259200 210600
rect 880 210320 259120 210464
rect 800 210184 259120 210320
rect 800 207064 259200 210184
rect 880 206784 259120 207064
rect 800 203664 259200 206784
rect 800 203392 259120 203664
rect 880 203384 259120 203392
rect 880 203112 259200 203384
rect 800 200264 259200 203112
rect 800 199984 259120 200264
rect 800 199720 259200 199984
rect 880 199440 259200 199720
rect 800 196864 259200 199440
rect 800 196584 259120 196864
rect 800 196048 259200 196584
rect 880 195768 259200 196048
rect 800 193328 259200 195768
rect 800 193048 259120 193328
rect 800 192376 259200 193048
rect 880 192096 259200 192376
rect 800 189928 259200 192096
rect 800 189648 259120 189928
rect 800 188704 259200 189648
rect 880 188424 259200 188704
rect 800 186528 259200 188424
rect 800 186248 259120 186528
rect 800 185032 259200 186248
rect 880 184752 259200 185032
rect 800 183128 259200 184752
rect 800 182848 259120 183128
rect 800 181360 259200 182848
rect 880 181080 259200 181360
rect 800 179728 259200 181080
rect 800 179448 259120 179728
rect 800 177688 259200 179448
rect 880 177408 259200 177688
rect 800 176328 259200 177408
rect 800 176048 259120 176328
rect 800 174016 259200 176048
rect 880 173736 259200 174016
rect 800 172792 259200 173736
rect 800 172512 259120 172792
rect 800 170344 259200 172512
rect 880 170064 259200 170344
rect 800 169392 259200 170064
rect 800 169112 259120 169392
rect 800 166672 259200 169112
rect 880 166392 259200 166672
rect 800 165992 259200 166392
rect 800 165712 259120 165992
rect 800 163000 259200 165712
rect 880 162720 259200 163000
rect 800 162592 259200 162720
rect 800 162312 259120 162592
rect 800 159328 259200 162312
rect 880 159192 259200 159328
rect 880 159048 259120 159192
rect 800 158912 259120 159048
rect 800 155792 259200 158912
rect 880 155512 259120 155792
rect 800 152256 259200 155512
rect 800 152120 259120 152256
rect 880 151976 259120 152120
rect 880 151840 259200 151976
rect 800 148856 259200 151840
rect 800 148576 259120 148856
rect 800 148448 259200 148576
rect 880 148168 259200 148448
rect 800 145456 259200 148168
rect 800 145176 259120 145456
rect 800 144776 259200 145176
rect 880 144496 259200 144776
rect 800 142056 259200 144496
rect 800 141776 259120 142056
rect 800 141104 259200 141776
rect 880 140824 259200 141104
rect 800 138656 259200 140824
rect 800 138376 259120 138656
rect 800 137432 259200 138376
rect 880 137152 259200 137432
rect 800 135256 259200 137152
rect 800 134976 259120 135256
rect 800 133760 259200 134976
rect 880 133480 259200 133760
rect 800 131856 259200 133480
rect 800 131576 259120 131856
rect 800 130088 259200 131576
rect 880 129808 259200 130088
rect 800 128320 259200 129808
rect 800 128040 259120 128320
rect 800 126416 259200 128040
rect 880 126136 259200 126416
rect 800 124920 259200 126136
rect 800 124640 259120 124920
rect 800 122744 259200 124640
rect 880 122464 259200 122744
rect 800 121520 259200 122464
rect 800 121240 259120 121520
rect 800 119072 259200 121240
rect 880 118792 259200 119072
rect 800 118120 259200 118792
rect 800 117840 259120 118120
rect 800 115400 259200 117840
rect 880 115120 259200 115400
rect 800 114720 259200 115120
rect 800 114440 259120 114720
rect 800 111728 259200 114440
rect 880 111448 259200 111728
rect 800 111320 259200 111448
rect 800 111040 259120 111320
rect 800 108056 259200 111040
rect 880 107784 259200 108056
rect 880 107776 259120 107784
rect 800 107504 259120 107776
rect 800 104520 259200 107504
rect 880 104384 259200 104520
rect 880 104240 259120 104384
rect 800 104104 259120 104240
rect 800 100984 259200 104104
rect 800 100848 259120 100984
rect 880 100704 259120 100848
rect 880 100568 259200 100704
rect 800 97584 259200 100568
rect 800 97304 259120 97584
rect 800 97176 259200 97304
rect 880 96896 259200 97176
rect 800 94184 259200 96896
rect 800 93904 259120 94184
rect 800 93504 259200 93904
rect 880 93224 259200 93504
rect 800 90784 259200 93224
rect 800 90504 259120 90784
rect 800 89832 259200 90504
rect 880 89552 259200 89832
rect 800 87248 259200 89552
rect 800 86968 259120 87248
rect 800 86160 259200 86968
rect 880 85880 259200 86160
rect 800 83848 259200 85880
rect 800 83568 259120 83848
rect 800 82488 259200 83568
rect 880 82208 259200 82488
rect 800 80448 259200 82208
rect 800 80168 259120 80448
rect 800 78816 259200 80168
rect 880 78536 259200 78816
rect 800 77048 259200 78536
rect 800 76768 259120 77048
rect 800 75144 259200 76768
rect 880 74864 259200 75144
rect 800 73648 259200 74864
rect 800 73368 259120 73648
rect 800 71472 259200 73368
rect 880 71192 259200 71472
rect 800 70248 259200 71192
rect 800 69968 259120 70248
rect 800 67800 259200 69968
rect 880 67520 259200 67800
rect 800 66848 259200 67520
rect 800 66568 259120 66848
rect 800 64128 259200 66568
rect 880 63848 259200 64128
rect 800 63312 259200 63848
rect 800 63032 259120 63312
rect 800 60456 259200 63032
rect 880 60176 259200 60456
rect 800 59912 259200 60176
rect 800 59632 259120 59912
rect 800 56784 259200 59632
rect 880 56512 259200 56784
rect 880 56504 259120 56512
rect 800 56232 259120 56504
rect 800 53248 259200 56232
rect 880 53112 259200 53248
rect 880 52968 259120 53112
rect 800 52832 259120 52968
rect 800 49712 259200 52832
rect 800 49576 259120 49712
rect 880 49432 259120 49576
rect 880 49296 259200 49432
rect 800 46312 259200 49296
rect 800 46032 259120 46312
rect 800 45904 259200 46032
rect 880 45624 259200 45904
rect 800 42776 259200 45624
rect 800 42496 259120 42776
rect 800 42232 259200 42496
rect 880 41952 259200 42232
rect 800 39376 259200 41952
rect 800 39096 259120 39376
rect 800 38560 259200 39096
rect 880 38280 259200 38560
rect 800 35976 259200 38280
rect 800 35696 259120 35976
rect 800 34888 259200 35696
rect 880 34608 259200 34888
rect 800 32576 259200 34608
rect 800 32296 259120 32576
rect 800 31216 259200 32296
rect 880 30936 259200 31216
rect 800 29176 259200 30936
rect 800 28896 259120 29176
rect 800 27544 259200 28896
rect 880 27264 259200 27544
rect 800 25776 259200 27264
rect 800 25496 259120 25776
rect 800 23872 259200 25496
rect 880 23592 259200 23872
rect 800 22240 259200 23592
rect 800 21960 259120 22240
rect 800 20200 259200 21960
rect 880 19920 259200 20200
rect 800 18840 259200 19920
rect 800 18560 259120 18840
rect 800 16528 259200 18560
rect 880 16248 259200 16528
rect 800 15440 259200 16248
rect 800 15160 259120 15440
rect 800 12856 259200 15160
rect 880 12576 259200 12856
rect 800 12040 259200 12576
rect 800 11760 259120 12040
rect 800 9184 259200 11760
rect 880 8904 259200 9184
rect 800 8640 259200 8904
rect 800 8360 259120 8640
rect 800 5512 259200 8360
rect 880 5240 259200 5512
rect 880 5232 259120 5240
rect 800 4960 259120 5232
rect 800 1976 259200 4960
rect 880 1840 259200 1976
rect 880 1696 259120 1840
rect 800 1560 259120 1696
rect 800 1395 259200 1560
<< metal4 >>
rect 4208 2128 4528 257360
rect 9208 2128 9528 257360
rect 14208 2128 14528 257360
rect 19208 2128 19528 257360
rect 24208 2128 24528 257360
rect 29208 2128 29528 257360
rect 34208 2128 34528 257360
rect 39208 2128 39528 257360
rect 44208 2128 44528 257360
rect 49208 2128 49528 257360
rect 54208 2128 54528 257360
rect 59208 2128 59528 257360
rect 64208 2128 64528 257360
rect 69208 2128 69528 257360
rect 74208 2128 74528 257360
rect 79208 2128 79528 257360
rect 84208 2128 84528 257360
rect 89208 2128 89528 257360
rect 94208 2128 94528 257360
rect 99208 2128 99528 257360
rect 104208 2128 104528 257360
rect 109208 2128 109528 257360
rect 114208 2128 114528 257360
rect 119208 2128 119528 257360
rect 124208 2128 124528 257360
rect 129208 2128 129528 257360
rect 134208 2128 134528 257360
rect 139208 2128 139528 257360
rect 144208 2128 144528 257360
rect 149208 2128 149528 257360
rect 154208 2128 154528 257360
rect 159208 2128 159528 257360
rect 164208 2128 164528 257360
rect 169208 2128 169528 257360
rect 174208 2128 174528 257360
rect 179208 2128 179528 257360
rect 184208 2128 184528 257360
rect 189208 2128 189528 257360
rect 194208 2128 194528 257360
rect 199208 2128 199528 257360
rect 204208 2128 204528 257360
rect 209208 2128 209528 257360
rect 214208 2128 214528 257360
rect 219208 2128 219528 257360
rect 224208 2128 224528 257360
rect 229208 2128 229528 257360
rect 234208 2128 234528 257360
rect 239208 2128 239528 257360
rect 244208 2128 244528 257360
rect 249208 2128 249528 257360
rect 254208 2128 254528 257360
<< obsm4 >>
rect 82123 13907 84128 183701
rect 84608 13907 89128 183701
rect 89608 13907 94128 183701
rect 94608 13907 99128 183701
rect 99608 13907 104128 183701
rect 104608 13907 109128 183701
rect 109608 13907 114128 183701
rect 114608 13907 119128 183701
rect 119608 13907 124128 183701
rect 124608 13907 129128 183701
rect 129608 13907 134128 183701
rect 134608 13907 139128 183701
rect 139608 13907 144128 183701
rect 144608 13907 149128 183701
rect 149608 13907 154128 183701
rect 154608 13907 159128 183701
rect 159608 13907 164128 183701
rect 164608 13907 169128 183701
rect 169608 13907 174128 183701
rect 174608 13907 179128 183701
rect 179608 13907 184128 183701
rect 184608 13907 189128 183701
rect 189608 13907 194128 183701
rect 194608 13907 199128 183701
rect 199608 13907 204128 183701
rect 204608 13907 208781 183701
<< labels >>
rlabel metal2 s 12714 259200 12770 260000 6 boot_addr_i[0]
port 1 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 boot_addr_i[10]
port 2 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 boot_addr_i[11]
port 3 nsew signal input
rlabel metal3 s 259200 114520 260000 114640 6 boot_addr_i[12]
port 4 nsew signal input
rlabel metal2 s 196714 0 196770 800 6 boot_addr_i[13]
port 5 nsew signal input
rlabel metal2 s 148230 259200 148286 260000 6 boot_addr_i[14]
port 6 nsew signal input
rlabel metal3 s 259200 152056 260000 152176 6 boot_addr_i[15]
port 7 nsew signal input
rlabel metal3 s 259200 165792 260000 165912 6 boot_addr_i[16]
port 8 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 boot_addr_i[17]
port 9 nsew signal input
rlabel metal2 s 173806 259200 173862 260000 6 boot_addr_i[18]
port 10 nsew signal input
rlabel metal3 s 0 162800 800 162920 6 boot_addr_i[19]
port 11 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 boot_addr_i[1]
port 12 nsew signal input
rlabel metal3 s 0 173816 800 173936 6 boot_addr_i[20]
port 13 nsew signal input
rlabel metal3 s 0 184832 800 184952 6 boot_addr_i[21]
port 14 nsew signal input
rlabel metal2 s 220818 0 220874 800 6 boot_addr_i[22]
port 15 nsew signal input
rlabel metal2 s 206742 259200 206798 260000 6 boot_addr_i[23]
port 16 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 boot_addr_i[24]
port 17 nsew signal input
rlabel metal3 s 259200 220600 260000 220720 6 boot_addr_i[25]
port 18 nsew signal input
rlabel metal3 s 259200 230800 260000 230920 6 boot_addr_i[26]
port 19 nsew signal input
rlabel metal3 s 259200 237600 260000 237720 6 boot_addr_i[27]
port 20 nsew signal input
rlabel metal3 s 259200 244536 260000 244656 6 boot_addr_i[28]
port 21 nsew signal input
rlabel metal2 s 245014 0 245070 800 6 boot_addr_i[29]
port 22 nsew signal input
rlabel metal3 s 0 27344 800 27464 6 boot_addr_i[2]
port 23 nsew signal input
rlabel metal2 s 249246 0 249302 800 6 boot_addr_i[30]
port 24 nsew signal input
rlabel metal2 s 254950 0 255006 800 6 boot_addr_i[31]
port 25 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 boot_addr_i[3]
port 26 nsew signal input
rlabel metal3 s 259200 70048 260000 70168 6 boot_addr_i[4]
port 27 nsew signal input
rlabel metal2 s 89626 259200 89682 260000 6 boot_addr_i[5]
port 28 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 boot_addr_i[6]
port 29 nsew signal input
rlabel metal3 s 259200 83648 260000 83768 6 boot_addr_i[7]
port 30 nsew signal input
rlabel metal2 s 182454 0 182510 800 6 boot_addr_i[8]
port 31 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 boot_addr_i[9]
port 32 nsew signal input
rlabel metal3 s 259200 1640 260000 1760 6 clk_i
port 33 nsew signal input
rlabel metal2 s 16394 259200 16450 260000 6 cluster_id_i[0]
port 34 nsew signal input
rlabel metal3 s 259200 39176 260000 39296 6 cluster_id_i[1]
port 35 nsew signal input
rlabel metal3 s 259200 49512 260000 49632 6 cluster_id_i[2]
port 36 nsew signal input
rlabel metal2 s 67638 259200 67694 260000 6 cluster_id_i[3]
port 37 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 cluster_id_i[4]
port 38 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 cluster_id_i[5]
port 39 nsew signal input
rlabel metal2 s 20074 259200 20130 260000 6 core_id_i[0]
port 40 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 core_id_i[1]
port 41 nsew signal input
rlabel metal2 s 49330 259200 49386 260000 6 core_id_i[2]
port 42 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 core_id_i[3]
port 43 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 data_addr_o[0]
port 44 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 data_addr_o[10]
port 45 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 data_addr_o[11]
port 46 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 data_addr_o[12]
port 47 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 data_addr_o[13]
port 48 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 data_addr_o[14]
port 49 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 data_addr_o[15]
port 50 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 data_addr_o[16]
port 51 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 data_addr_o[17]
port 52 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 data_addr_o[18]
port 53 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 data_addr_o[19]
port 54 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 data_addr_o[1]
port 55 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 data_addr_o[20]
port 56 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 data_addr_o[21]
port 57 nsew signal output
rlabel metal2 s 107198 0 107254 800 6 data_addr_o[22]
port 58 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 data_addr_o[23]
port 59 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 data_addr_o[24]
port 60 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 data_addr_o[25]
port 61 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 data_addr_o[26]
port 62 nsew signal output
rlabel metal2 s 128450 0 128506 800 6 data_addr_o[27]
port 63 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 data_addr_o[28]
port 64 nsew signal output
rlabel metal2 s 137006 0 137062 800 6 data_addr_o[29]
port 65 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 data_addr_o[2]
port 66 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 data_addr_o[30]
port 67 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 data_addr_o[31]
port 68 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 data_addr_o[3]
port 69 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 data_addr_o[4]
port 70 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 data_addr_o[5]
port 71 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 data_addr_o[6]
port 72 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 data_addr_o[7]
port 73 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 data_addr_o[8]
port 74 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 data_addr_o[9]
port 75 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 data_be_o[0]
port 76 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 data_be_o[1]
port 77 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 data_be_o[2]
port 78 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 data_be_o[3]
port 79 nsew signal output
rlabel metal2 s 662 0 718 800 6 data_err_i
port 80 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 data_gnt_i
port 81 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 data_rdata_i[0]
port 82 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 data_rdata_i[10]
port 83 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 data_rdata_i[11]
port 84 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 data_rdata_i[12]
port 85 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 data_rdata_i[13]
port 86 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 data_rdata_i[14]
port 87 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 data_rdata_i[15]
port 88 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 data_rdata_i[16]
port 89 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 data_rdata_i[17]
port 90 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 data_rdata_i[18]
port 91 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 data_rdata_i[19]
port 92 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 data_rdata_i[1]
port 93 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 data_rdata_i[20]
port 94 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 data_rdata_i[21]
port 95 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 data_rdata_i[22]
port 96 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 data_rdata_i[23]
port 97 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 data_rdata_i[24]
port 98 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 data_rdata_i[25]
port 99 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 data_rdata_i[26]
port 100 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 data_rdata_i[27]
port 101 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 data_rdata_i[28]
port 102 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 data_rdata_i[29]
port 103 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 data_rdata_i[2]
port 104 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 data_rdata_i[30]
port 105 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 data_rdata_i[31]
port 106 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 data_rdata_i[3]
port 107 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 data_rdata_i[4]
port 108 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 data_rdata_i[5]
port 109 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 data_rdata_i[6]
port 110 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 data_rdata_i[7]
port 111 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 data_rdata_i[8]
port 112 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 data_rdata_i[9]
port 113 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 data_req_o
port 114 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 data_rvalid_i
port 115 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 data_wdata_o[0]
port 116 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 data_wdata_o[10]
port 117 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 data_wdata_o[11]
port 118 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 data_wdata_o[12]
port 119 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 data_wdata_o[13]
port 120 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 data_wdata_o[14]
port 121 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 data_wdata_o[15]
port 122 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 data_wdata_o[16]
port 123 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 data_wdata_o[17]
port 124 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 data_wdata_o[18]
port 125 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 data_wdata_o[19]
port 126 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 data_wdata_o[1]
port 127 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 data_wdata_o[20]
port 128 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 data_wdata_o[21]
port 129 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 data_wdata_o[22]
port 130 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 data_wdata_o[23]
port 131 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 data_wdata_o[24]
port 132 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 data_wdata_o[25]
port 133 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 data_wdata_o[26]
port 134 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 data_wdata_o[27]
port 135 nsew signal output
rlabel metal2 s 135626 0 135682 800 6 data_wdata_o[28]
port 136 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 data_wdata_o[29]
port 137 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 data_wdata_o[2]
port 138 nsew signal output
rlabel metal2 s 144090 0 144146 800 6 data_wdata_o[30]
port 139 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 data_wdata_o[31]
port 140 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 data_wdata_o[3]
port 141 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 data_wdata_o[4]
port 142 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 data_wdata_o[5]
port 143 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 data_wdata_o[6]
port 144 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 data_wdata_o[7]
port 145 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 data_wdata_o[8]
port 146 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 data_wdata_o[9]
port 147 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 data_we_o
port 148 nsew signal output
rlabel metal3 s 259200 5040 260000 5160 6 debug_req_i
port 149 nsew signal input
rlabel metal2 s 23662 259200 23718 260000 6 eFPGA_delay_o[0]
port 150 nsew signal output
rlabel metal3 s 259200 42576 260000 42696 6 eFPGA_delay_o[1]
port 151 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 eFPGA_delay_o[2]
port 152 nsew signal output
rlabel metal3 s 259200 52912 260000 53032 6 eFPGA_delay_o[3]
port 153 nsew signal output
rlabel metal2 s 1766 259200 1822 260000 6 eFPGA_en_o
port 154 nsew signal output
rlabel metal2 s 149794 0 149850 800 6 eFPGA_fpga_done_i
port 155 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 eFPGA_operand_a_o[0]
port 156 nsew signal output
rlabel metal3 s 259200 100784 260000 100904 6 eFPGA_operand_a_o[10]
port 157 nsew signal output
rlabel metal3 s 0 107856 800 107976 6 eFPGA_operand_a_o[11]
port 158 nsew signal output
rlabel metal2 s 192390 0 192446 800 6 eFPGA_operand_a_o[12]
port 159 nsew signal output
rlabel metal3 s 259200 128120 260000 128240 6 eFPGA_operand_a_o[13]
port 160 nsew signal output
rlabel metal2 s 151818 259200 151874 260000 6 eFPGA_operand_a_o[14]
port 161 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 eFPGA_operand_a_o[15]
port 162 nsew signal output
rlabel metal2 s 162858 259200 162914 260000 6 eFPGA_operand_a_o[16]
port 163 nsew signal output
rlabel metal3 s 259200 176128 260000 176248 6 eFPGA_operand_a_o[17]
port 164 nsew signal output
rlabel metal3 s 0 151920 800 152040 6 eFPGA_operand_a_o[18]
port 165 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 eFPGA_operand_a_o[19]
port 166 nsew signal output
rlabel metal3 s 259200 46112 260000 46232 6 eFPGA_operand_a_o[1]
port 167 nsew signal output
rlabel metal3 s 259200 196664 260000 196784 6 eFPGA_operand_a_o[20]
port 168 nsew signal output
rlabel metal3 s 0 188504 800 188624 6 eFPGA_operand_a_o[21]
port 169 nsew signal output
rlabel metal3 s 0 203192 800 203312 6 eFPGA_operand_a_o[22]
port 170 nsew signal output
rlabel metal2 s 210422 259200 210478 260000 6 eFPGA_operand_a_o[23]
port 171 nsew signal output
rlabel metal3 s 259200 213664 260000 213784 6 eFPGA_operand_a_o[24]
port 172 nsew signal output
rlabel metal2 s 228730 259200 228786 260000 6 eFPGA_operand_a_o[25]
port 173 nsew signal output
rlabel metal2 s 236090 259200 236146 260000 6 eFPGA_operand_a_o[26]
port 174 nsew signal output
rlabel metal2 s 236458 0 236514 800 6 eFPGA_operand_a_o[27]
port 175 nsew signal output
rlabel metal3 s 0 225088 800 225208 6 eFPGA_operand_a_o[28]
port 176 nsew signal output
rlabel metal3 s 0 232432 800 232552 6 eFPGA_operand_a_o[29]
port 177 nsew signal output
rlabel metal2 s 162582 0 162638 800 6 eFPGA_operand_a_o[2]
port 178 nsew signal output
rlabel metal2 s 250626 0 250682 800 6 eFPGA_operand_a_o[30]
port 179 nsew signal output
rlabel metal2 s 256330 0 256386 800 6 eFPGA_operand_a_o[31]
port 180 nsew signal output
rlabel metal2 s 71318 259200 71374 260000 6 eFPGA_operand_a_o[3]
port 181 nsew signal output
rlabel metal3 s 0 49376 800 49496 6 eFPGA_operand_a_o[4]
port 182 nsew signal output
rlabel metal2 s 175370 0 175426 800 6 eFPGA_operand_a_o[5]
port 183 nsew signal output
rlabel metal2 s 104254 259200 104310 260000 6 eFPGA_operand_a_o[6]
port 184 nsew signal output
rlabel metal2 s 179602 0 179658 800 6 eFPGA_operand_a_o[7]
port 185 nsew signal output
rlabel metal2 s 122562 259200 122618 260000 6 eFPGA_operand_a_o[8]
port 186 nsew signal output
rlabel metal3 s 259200 93984 260000 94104 6 eFPGA_operand_a_o[9]
port 187 nsew signal output
rlabel metal2 s 27342 259200 27398 260000 6 eFPGA_operand_b_o[0]
port 188 nsew signal output
rlabel metal3 s 259200 104184 260000 104304 6 eFPGA_operand_b_o[10]
port 189 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 eFPGA_operand_b_o[11]
port 190 nsew signal output
rlabel metal3 s 259200 117920 260000 118040 6 eFPGA_operand_b_o[12]
port 191 nsew signal output
rlabel metal3 s 259200 131656 260000 131776 6 eFPGA_operand_b_o[13]
port 192 nsew signal output
rlabel metal2 s 155498 259200 155554 260000 6 eFPGA_operand_b_o[14]
port 193 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 eFPGA_operand_b_o[15]
port 194 nsew signal output
rlabel metal2 s 202326 0 202382 800 6 eFPGA_operand_b_o[16]
port 195 nsew signal output
rlabel metal2 s 205178 0 205234 800 6 eFPGA_operand_b_o[17]
port 196 nsew signal output
rlabel metal3 s 259200 186328 260000 186448 6 eFPGA_operand_b_o[18]
port 197 nsew signal output
rlabel metal2 s 212262 0 212318 800 6 eFPGA_operand_b_o[19]
port 198 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 eFPGA_operand_b_o[1]
port 199 nsew signal output
rlabel metal2 s 215114 0 215170 800 6 eFPGA_operand_b_o[20]
port 200 nsew signal output
rlabel metal2 s 184846 259200 184902 260000 6 eFPGA_operand_b_o[21]
port 201 nsew signal output
rlabel metal2 s 192114 259200 192170 260000 6 eFPGA_operand_b_o[22]
port 202 nsew signal output
rlabel metal3 s 259200 206864 260000 206984 6 eFPGA_operand_b_o[23]
port 203 nsew signal output
rlabel metal2 s 226522 0 226578 800 6 eFPGA_operand_b_o[24]
port 204 nsew signal output
rlabel metal3 s 259200 224000 260000 224120 6 eFPGA_operand_b_o[25]
port 205 nsew signal output
rlabel metal3 s 259200 234200 260000 234320 6 eFPGA_operand_b_o[26]
port 206 nsew signal output
rlabel metal2 s 237838 0 237894 800 6 eFPGA_operand_b_o[27]
port 207 nsew signal output
rlabel metal2 s 242162 0 242218 800 6 eFPGA_operand_b_o[28]
port 208 nsew signal output
rlabel metal2 s 246394 0 246450 800 6 eFPGA_operand_b_o[29]
port 209 nsew signal output
rlabel metal2 s 53010 259200 53066 260000 6 eFPGA_operand_b_o[2]
port 210 nsew signal output
rlabel metal3 s 0 247120 800 247240 6 eFPGA_operand_b_o[30]
port 211 nsew signal output
rlabel metal3 s 259200 258136 260000 258256 6 eFPGA_operand_b_o[31]
port 212 nsew signal output
rlabel metal3 s 259200 56312 260000 56432 6 eFPGA_operand_b_o[3]
port 213 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 eFPGA_operand_b_o[4]
port 214 nsew signal output
rlabel metal2 s 93306 259200 93362 260000 6 eFPGA_operand_b_o[5]
port 215 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 eFPGA_operand_b_o[6]
port 216 nsew signal output
rlabel metal2 s 115202 259200 115258 260000 6 eFPGA_operand_b_o[7]
port 217 nsew signal output
rlabel metal2 s 183926 0 183982 800 6 eFPGA_operand_b_o[8]
port 218 nsew signal output
rlabel metal3 s 259200 97384 260000 97504 6 eFPGA_operand_b_o[9]
port 219 nsew signal output
rlabel metal3 s 259200 22040 260000 22160 6 eFPGA_operator_o[0]
port 220 nsew signal output
rlabel metal2 s 31022 259200 31078 260000 6 eFPGA_operator_o[1]
port 221 nsew signal output
rlabel metal3 s 259200 25576 260000 25696 6 eFPGA_result_a_i[0]
port 222 nsew signal input
rlabel metal3 s 259200 107584 260000 107704 6 eFPGA_result_a_i[10]
port 223 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 eFPGA_result_a_i[11]
port 224 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 eFPGA_result_a_i[12]
port 225 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 eFPGA_result_a_i[13]
port 226 nsew signal input
rlabel metal3 s 259200 141856 260000 141976 6 eFPGA_result_a_i[14]
port 227 nsew signal input
rlabel metal3 s 259200 155592 260000 155712 6 eFPGA_result_a_i[15]
port 228 nsew signal input
rlabel metal3 s 0 144576 800 144696 6 eFPGA_result_a_i[16]
port 229 nsew signal input
rlabel metal2 s 206650 0 206706 800 6 eFPGA_result_a_i[17]
port 230 nsew signal input
rlabel metal3 s 0 155592 800 155712 6 eFPGA_result_a_i[18]
port 231 nsew signal input
rlabel metal2 s 181166 259200 181222 260000 6 eFPGA_result_a_i[19]
port 232 nsew signal input
rlabel metal2 s 34702 259200 34758 260000 6 eFPGA_result_a_i[1]
port 233 nsew signal input
rlabel metal3 s 0 177488 800 177608 6 eFPGA_result_a_i[20]
port 234 nsew signal input
rlabel metal3 s 0 192176 800 192296 6 eFPGA_result_a_i[21]
port 235 nsew signal input
rlabel metal2 s 222290 0 222346 800 6 eFPGA_result_a_i[22]
port 236 nsew signal input
rlabel metal2 s 214102 259200 214158 260000 6 eFPGA_result_a_i[23]
port 237 nsew signal input
rlabel metal2 s 227902 0 227958 800 6 eFPGA_result_a_i[24]
port 238 nsew signal input
rlabel metal2 s 230754 0 230810 800 6 eFPGA_result_a_i[25]
port 239 nsew signal input
rlabel metal2 s 233606 0 233662 800 6 eFPGA_result_a_i[26]
port 240 nsew signal input
rlabel metal3 s 0 217744 800 217864 6 eFPGA_result_a_i[27]
port 241 nsew signal input
rlabel metal3 s 259200 247936 260000 248056 6 eFPGA_result_a_i[28]
port 242 nsew signal input
rlabel metal3 s 0 236104 800 236224 6 eFPGA_result_a_i[29]
port 243 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 eFPGA_result_a_i[2]
port 244 nsew signal input
rlabel metal3 s 0 250792 800 250912 6 eFPGA_result_a_i[30]
port 245 nsew signal input
rlabel metal2 s 257802 0 257858 800 6 eFPGA_result_a_i[31]
port 246 nsew signal input
rlabel metal3 s 259200 59712 260000 59832 6 eFPGA_result_a_i[3]
port 247 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 eFPGA_result_a_i[4]
port 248 nsew signal input
rlabel metal2 s 96894 259200 96950 260000 6 eFPGA_result_a_i[5]
port 249 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 eFPGA_result_a_i[6]
port 250 nsew signal input
rlabel metal2 s 118882 259200 118938 260000 6 eFPGA_result_a_i[7]
port 251 nsew signal input
rlabel metal2 s 126242 259200 126298 260000 6 eFPGA_result_a_i[8]
port 252 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 eFPGA_result_a_i[9]
port 253 nsew signal input
rlabel metal3 s 259200 28976 260000 29096 6 eFPGA_result_b_i[0]
port 254 nsew signal input
rlabel metal2 s 133510 259200 133566 260000 6 eFPGA_result_b_i[10]
port 255 nsew signal input
rlabel metal3 s 0 115200 800 115320 6 eFPGA_result_b_i[11]
port 256 nsew signal input
rlabel metal3 s 0 126216 800 126336 6 eFPGA_result_b_i[12]
port 257 nsew signal input
rlabel metal2 s 199474 0 199530 800 6 eFPGA_result_b_i[13]
port 258 nsew signal input
rlabel metal3 s 259200 145256 260000 145376 6 eFPGA_result_b_i[14]
port 259 nsew signal input
rlabel metal3 s 0 137232 800 137352 6 eFPGA_result_b_i[15]
port 260 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 eFPGA_result_b_i[16]
port 261 nsew signal input
rlabel metal3 s 259200 179528 260000 179648 6 eFPGA_result_b_i[17]
port 262 nsew signal input
rlabel metal3 s 259200 189728 260000 189848 6 eFPGA_result_b_i[18]
port 263 nsew signal input
rlabel metal2 s 213734 0 213790 800 6 eFPGA_result_b_i[19]
port 264 nsew signal input
rlabel metal2 s 38382 259200 38438 260000 6 eFPGA_result_b_i[1]
port 265 nsew signal input
rlabel metal3 s 259200 200064 260000 200184 6 eFPGA_result_b_i[20]
port 266 nsew signal input
rlabel metal2 s 188434 259200 188490 260000 6 eFPGA_result_b_i[21]
port 267 nsew signal input
rlabel metal2 s 195794 259200 195850 260000 6 eFPGA_result_b_i[22]
port 268 nsew signal input
rlabel metal3 s 259200 210264 260000 210384 6 eFPGA_result_b_i[23]
port 269 nsew signal input
rlabel metal2 s 225050 259200 225106 260000 6 eFPGA_result_b_i[24]
port 270 nsew signal input
rlabel metal3 s 259200 227400 260000 227520 6 eFPGA_result_b_i[25]
port 271 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 eFPGA_result_b_i[26]
port 272 nsew signal input
rlabel metal2 s 239310 0 239366 800 6 eFPGA_result_b_i[27]
port 273 nsew signal input
rlabel metal3 s 259200 251336 260000 251456 6 eFPGA_result_b_i[28]
port 274 nsew signal input
rlabel metal2 s 247866 0 247922 800 6 eFPGA_result_b_i[29]
port 275 nsew signal input
rlabel metal2 s 56690 259200 56746 260000 6 eFPGA_result_b_i[2]
port 276 nsew signal input
rlabel metal2 s 252098 0 252154 800 6 eFPGA_result_b_i[30]
port 277 nsew signal input
rlabel metal2 s 258078 259200 258134 260000 6 eFPGA_result_b_i[31]
port 278 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 eFPGA_result_b_i[3]
port 279 nsew signal input
rlabel metal2 s 82266 259200 82322 260000 6 eFPGA_result_b_i[4]
port 280 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 eFPGA_result_b_i[5]
port 281 nsew signal input
rlabel metal2 s 107934 259200 107990 260000 6 eFPGA_result_b_i[6]
port 282 nsew signal input
rlabel metal2 s 181074 0 181130 800 6 eFPGA_result_b_i[7]
port 283 nsew signal input
rlabel metal2 s 185306 0 185362 800 6 eFPGA_result_b_i[8]
port 284 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 eFPGA_result_b_i[9]
port 285 nsew signal input
rlabel metal3 s 259200 32376 260000 32496 6 eFPGA_result_c_i[0]
port 286 nsew signal input
rlabel metal3 s 0 104320 800 104440 6 eFPGA_result_c_i[10]
port 287 nsew signal input
rlabel metal2 s 140870 259200 140926 260000 6 eFPGA_result_c_i[11]
port 288 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 eFPGA_result_c_i[12]
port 289 nsew signal input
rlabel metal3 s 259200 135056 260000 135176 6 eFPGA_result_c_i[13]
port 290 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 eFPGA_result_c_i[14]
port 291 nsew signal input
rlabel metal3 s 259200 158992 260000 159112 6 eFPGA_result_c_i[15]
port 292 nsew signal input
rlabel metal3 s 259200 169192 260000 169312 6 eFPGA_result_c_i[16]
port 293 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 eFPGA_result_c_i[17]
port 294 nsew signal input
rlabel metal2 s 209502 0 209558 800 6 eFPGA_result_c_i[18]
port 295 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 eFPGA_result_c_i[19]
port 296 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 eFPGA_result_c_i[1]
port 297 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 eFPGA_result_c_i[20]
port 298 nsew signal input
rlabel metal2 s 219438 0 219494 800 6 eFPGA_result_c_i[21]
port 299 nsew signal input
rlabel metal3 s 259200 203464 260000 203584 6 eFPGA_result_c_i[22]
port 300 nsew signal input
rlabel metal2 s 217782 259200 217838 260000 6 eFPGA_result_c_i[23]
port 301 nsew signal input
rlabel metal2 s 229374 0 229430 800 6 eFPGA_result_c_i[24]
port 302 nsew signal input
rlabel metal2 s 232226 0 232282 800 6 eFPGA_result_c_i[25]
port 303 nsew signal input
rlabel metal2 s 239770 259200 239826 260000 6 eFPGA_result_c_i[26]
port 304 nsew signal input
rlabel metal3 s 259200 241136 260000 241256 6 eFPGA_result_c_i[27]
port 305 nsew signal input
rlabel metal3 s 0 228760 800 228880 6 eFPGA_result_c_i[28]
port 306 nsew signal input
rlabel metal2 s 250718 259200 250774 260000 6 eFPGA_result_c_i[29]
port 307 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 eFPGA_result_c_i[2]
port 308 nsew signal input
rlabel metal2 s 253478 0 253534 800 6 eFPGA_result_c_i[30]
port 309 nsew signal input
rlabel metal2 s 259182 0 259238 800 6 eFPGA_result_c_i[31]
port 310 nsew signal input
rlabel metal2 s 74998 259200 75054 260000 6 eFPGA_result_c_i[3]
port 311 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 eFPGA_result_c_i[4]
port 312 nsew signal input
rlabel metal3 s 0 60256 800 60376 6 eFPGA_result_c_i[5]
port 313 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 eFPGA_result_c_i[6]
port 314 nsew signal input
rlabel metal3 s 259200 87048 260000 87168 6 eFPGA_result_c_i[7]
port 315 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 eFPGA_result_c_i[8]
port 316 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 eFPGA_result_c_i[9]
port 317 nsew signal input
rlabel metal2 s 5354 259200 5410 260000 6 eFPGA_write_strobe_o
port 318 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 ext_perf_counters_i
port 319 nsew signal input
rlabel metal3 s 259200 8440 260000 8560 6 fetch_enable_i
port 320 nsew signal input
rlabel metal3 s 259200 35776 260000 35896 6 instr_addr_o[0]
port 321 nsew signal output
rlabel metal3 s 259200 111120 260000 111240 6 instr_addr_o[10]
port 322 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 instr_addr_o[11]
port 323 nsew signal output
rlabel metal3 s 259200 121320 260000 121440 6 instr_addr_o[12]
port 324 nsew signal output
rlabel metal3 s 259200 138456 260000 138576 6 instr_addr_o[13]
port 325 nsew signal output
rlabel metal3 s 259200 148656 260000 148776 6 instr_addr_o[14]
port 326 nsew signal output
rlabel metal3 s 259200 162392 260000 162512 6 instr_addr_o[15]
port 327 nsew signal output
rlabel metal2 s 166538 259200 166594 260000 6 instr_addr_o[16]
port 328 nsew signal output
rlabel metal2 s 170126 259200 170182 260000 6 instr_addr_o[17]
port 329 nsew signal output
rlabel metal3 s 0 159128 800 159248 6 instr_addr_o[18]
port 330 nsew signal output
rlabel metal3 s 259200 193128 260000 193248 6 instr_addr_o[19]
port 331 nsew signal output
rlabel metal2 s 41970 259200 42026 260000 6 instr_addr_o[1]
port 332 nsew signal output
rlabel metal2 s 216586 0 216642 800 6 instr_addr_o[20]
port 333 nsew signal output
rlabel metal3 s 0 195848 800 195968 6 instr_addr_o[21]
port 334 nsew signal output
rlabel metal2 s 199474 259200 199530 260000 6 instr_addr_o[22]
port 335 nsew signal output
rlabel metal2 s 223670 0 223726 800 6 instr_addr_o[23]
port 336 nsew signal output
rlabel metal3 s 259200 217064 260000 217184 6 instr_addr_o[24]
port 337 nsew signal output
rlabel metal3 s 0 210400 800 210520 6 instr_addr_o[25]
port 338 nsew signal output
rlabel metal2 s 243358 259200 243414 260000 6 instr_addr_o[26]
port 339 nsew signal output
rlabel metal3 s 0 221416 800 221536 6 instr_addr_o[27]
port 340 nsew signal output
rlabel metal2 s 243542 0 243598 800 6 instr_addr_o[28]
port 341 nsew signal output
rlabel metal3 s 0 239776 800 239896 6 instr_addr_o[29]
port 342 nsew signal output
rlabel metal2 s 60278 259200 60334 260000 6 instr_addr_o[2]
port 343 nsew signal output
rlabel metal3 s 259200 254736 260000 254856 6 instr_addr_o[30]
port 344 nsew signal output
rlabel metal3 s 0 254464 800 254584 6 instr_addr_o[31]
port 345 nsew signal output
rlabel metal3 s 259200 63112 260000 63232 6 instr_addr_o[3]
port 346 nsew signal output
rlabel metal2 s 85946 259200 86002 260000 6 instr_addr_o[4]
port 347 nsew signal output
rlabel metal2 s 100574 259200 100630 260000 6 instr_addr_o[5]
port 348 nsew signal output
rlabel metal2 s 111614 259200 111670 260000 6 instr_addr_o[6]
port 349 nsew signal output
rlabel metal3 s 0 74944 800 75064 6 instr_addr_o[7]
port 350 nsew signal output
rlabel metal3 s 0 85960 800 86080 6 instr_addr_o[8]
port 351 nsew signal output
rlabel metal2 s 129922 259200 129978 260000 6 instr_addr_o[9]
port 352 nsew signal output
rlabel metal2 s 9034 259200 9090 260000 6 instr_gnt_i
port 353 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 instr_rdata_i[0]
port 354 nsew signal input
rlabel metal2 s 137190 259200 137246 260000 6 instr_rdata_i[10]
port 355 nsew signal input
rlabel metal3 s 0 122544 800 122664 6 instr_rdata_i[11]
port 356 nsew signal input
rlabel metal3 s 259200 124720 260000 124840 6 instr_rdata_i[12]
port 357 nsew signal input
rlabel metal2 s 144550 259200 144606 260000 6 instr_rdata_i[13]
port 358 nsew signal input
rlabel metal2 s 159178 259200 159234 260000 6 instr_rdata_i[14]
port 359 nsew signal input
rlabel metal3 s 0 140904 800 141024 6 instr_rdata_i[15]
port 360 nsew signal input
rlabel metal3 s 259200 172592 260000 172712 6 instr_rdata_i[16]
port 361 nsew signal input
rlabel metal3 s 259200 182928 260000 183048 6 instr_rdata_i[17]
port 362 nsew signal input
rlabel metal2 s 177486 259200 177542 260000 6 instr_rdata_i[18]
port 363 nsew signal input
rlabel metal3 s 0 170144 800 170264 6 instr_rdata_i[19]
port 364 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 instr_rdata_i[1]
port 365 nsew signal input
rlabel metal2 s 217966 0 218022 800 6 instr_rdata_i[20]
port 366 nsew signal input
rlabel metal3 s 0 199520 800 199640 6 instr_rdata_i[21]
port 367 nsew signal input
rlabel metal2 s 203154 259200 203210 260000 6 instr_rdata_i[22]
port 368 nsew signal input
rlabel metal2 s 221462 259200 221518 260000 6 instr_rdata_i[23]
port 369 nsew signal input
rlabel metal3 s 0 206864 800 206984 6 instr_rdata_i[24]
port 370 nsew signal input
rlabel metal2 s 232410 259200 232466 260000 6 instr_rdata_i[25]
port 371 nsew signal input
rlabel metal3 s 0 214072 800 214192 6 instr_rdata_i[26]
port 372 nsew signal input
rlabel metal2 s 240690 0 240746 800 6 instr_rdata_i[27]
port 373 nsew signal input
rlabel metal2 s 247038 259200 247094 260000 6 instr_rdata_i[28]
port 374 nsew signal input
rlabel metal3 s 0 243448 800 243568 6 instr_rdata_i[29]
port 375 nsew signal input
rlabel metal2 s 63958 259200 64014 260000 6 instr_rdata_i[2]
port 376 nsew signal input
rlabel metal2 s 254398 259200 254454 260000 6 instr_rdata_i[30]
port 377 nsew signal input
rlabel metal3 s 0 258136 800 258256 6 instr_rdata_i[31]
port 378 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 instr_rdata_i[3]
port 379 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 instr_rdata_i[4]
port 380 nsew signal input
rlabel metal3 s 259200 76848 260000 76968 6 instr_rdata_i[5]
port 381 nsew signal input
rlabel metal3 s 259200 80248 260000 80368 6 instr_rdata_i[6]
port 382 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 instr_rdata_i[7]
port 383 nsew signal input
rlabel metal3 s 259200 90584 260000 90704 6 instr_rdata_i[8]
port 384 nsew signal input
rlabel metal3 s 0 96976 800 97096 6 instr_rdata_i[9]
port 385 nsew signal input
rlabel metal3 s 259200 11840 260000 11960 6 instr_req_o
port 386 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 instr_rvalid_i
port 387 nsew signal input
rlabel metal3 s 259200 15240 260000 15360 6 irq_ack_o
port 388 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 irq_i
port 389 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 irq_id_i[0]
port 390 nsew signal input
rlabel metal2 s 45650 259200 45706 260000 6 irq_id_i[1]
port 391 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 irq_id_i[2]
port 392 nsew signal input
rlabel metal3 s 259200 66648 260000 66768 6 irq_id_i[3]
port 393 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 irq_id_i[4]
port 394 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 irq_id_o[0]
port 395 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 irq_id_o[1]
port 396 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 irq_id_o[2]
port 397 nsew signal output
rlabel metal2 s 78586 259200 78642 260000 6 irq_id_o[3]
port 398 nsew signal output
rlabel metal3 s 259200 73448 260000 73568 6 irq_id_o[4]
port 399 nsew signal output
rlabel metal2 s 154026 0 154082 800 6 rst_ni
port 400 nsew signal input
rlabel metal3 s 259200 18640 260000 18760 6 test_en_i
port 401 nsew signal input
rlabel metal4 s 4208 2128 4528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 14208 2128 14528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 24208 2128 24528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 34208 2128 34528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 44208 2128 44528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 54208 2128 54528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 64208 2128 64528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 74208 2128 74528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 84208 2128 84528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 94208 2128 94528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 104208 2128 104528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 114208 2128 114528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 124208 2128 124528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 134208 2128 134528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 144208 2128 144528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 154208 2128 154528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 164208 2128 164528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 174208 2128 174528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 184208 2128 184528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 194208 2128 194528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 204208 2128 204528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 214208 2128 214528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 224208 2128 224528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 234208 2128 234528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 244208 2128 244528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 254208 2128 254528 257360 6 vccd1
port 402 nsew power input
rlabel metal4 s 9208 2128 9528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 19208 2128 19528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 29208 2128 29528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 39208 2128 39528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 49208 2128 49528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 59208 2128 59528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 69208 2128 69528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 79208 2128 79528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 89208 2128 89528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 99208 2128 99528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 109208 2128 109528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 119208 2128 119528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 129208 2128 129528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 139208 2128 139528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 149208 2128 149528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 159208 2128 159528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 169208 2128 169528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 179208 2128 179528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 189208 2128 189528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 199208 2128 199528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 209208 2128 209528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 219208 2128 219528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 229208 2128 229528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 239208 2128 239528 257360 6 vssd1
port 403 nsew ground input
rlabel metal4 s 249208 2128 249528 257360 6 vssd1
port 403 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 260000 260000
string LEFview TRUE
string GDS_FILE /project/openlane/flexbex_ibex_core/runs/flexbex_ibex_core/results/magic/flexbex_ibex_core.gds
string GDS_END 82620380
string GDS_START 1615266
<< end >>

