magic
tech sky130A
magscale 1 2
timestamp 1640351253
<< locali >>
rect 23121 27863 23155 28033
rect 23765 27387 23799 27489
rect 11529 26979 11563 27081
rect 24225 25143 24259 25245
rect 7849 22491 7883 22593
rect 16497 21403 16531 21505
rect 17233 20859 17267 20961
rect 5089 18615 5123 18717
rect 12173 18615 12207 18717
rect 15117 17731 15151 17833
rect 13461 17527 13495 17629
rect 8953 15351 8987 15589
rect 24685 15351 24719 15453
rect 17693 14943 17727 15113
rect 10701 14399 10735 14501
rect 24225 8823 24259 9061
rect 21189 8279 21223 8449
rect 3617 5695 3651 5797
rect 18981 5015 19015 5117
rect 17325 4471 17359 4573
rect 21833 4471 21867 4777
rect 29561 4131 29595 26469
rect 16129 3587 16163 3689
rect 16129 3383 16163 3553
<< viali >>
rect 20177 30277 20211 30311
rect 11805 30209 11839 30243
rect 12357 30209 12391 30243
rect 14933 30209 14967 30243
rect 19441 30209 19475 30243
rect 19827 30209 19861 30243
rect 19993 30209 20027 30243
rect 20729 30209 20763 30243
rect 22057 30209 22091 30243
rect 22201 30209 22235 30243
rect 22293 30209 22327 30243
rect 22477 30209 22511 30243
rect 22845 30209 22879 30243
rect 19625 30141 19659 30175
rect 19717 30141 19751 30175
rect 21557 30141 21591 30175
rect 11989 30073 12023 30107
rect 21925 30073 21959 30107
rect 12173 30005 12207 30039
rect 14749 30005 14783 30039
rect 19349 30005 19383 30039
rect 20545 30005 20579 30039
rect 22661 30005 22695 30039
rect 23029 30005 23063 30039
rect 19349 29801 19383 29835
rect 19625 29733 19659 29767
rect 3341 29665 3375 29699
rect 4629 29665 4663 29699
rect 7665 29665 7699 29699
rect 14197 29665 14231 29699
rect 15945 29665 15979 29699
rect 16681 29665 16715 29699
rect 18613 29665 18647 29699
rect 21097 29665 21131 29699
rect 5549 29597 5583 29631
rect 9045 29597 9079 29631
rect 11161 29597 11195 29631
rect 13277 29597 13311 29631
rect 18429 29597 18463 29631
rect 18705 29597 18739 29631
rect 18815 29597 18849 29631
rect 18981 29597 19015 29631
rect 21373 29597 21407 29631
rect 21833 29597 21867 29631
rect 5794 29529 5828 29563
rect 7573 29529 7607 29563
rect 9321 29529 9355 29563
rect 13001 29529 13035 29563
rect 15669 29529 15703 29563
rect 16948 29529 16982 29563
rect 18245 29529 18279 29563
rect 22109 29529 22143 29563
rect 6929 29461 6963 29495
rect 7113 29461 7147 29495
rect 7481 29461 7515 29495
rect 10793 29461 10827 29495
rect 10977 29461 11011 29495
rect 11529 29461 11563 29495
rect 18061 29461 18095 29495
rect 23581 29461 23615 29495
rect 5641 29257 5675 29291
rect 9321 29257 9355 29291
rect 10517 29257 10551 29291
rect 13478 29257 13512 29291
rect 15761 29257 15795 29291
rect 18613 29257 18647 29291
rect 20545 29257 20579 29291
rect 22845 29257 22879 29291
rect 7205 29189 7239 29223
rect 10149 29189 10183 29223
rect 12173 29189 12207 29223
rect 13182 29189 13216 29223
rect 13737 29189 13771 29223
rect 22201 29189 22235 29223
rect 22937 29189 22971 29223
rect 3433 29121 3467 29155
rect 3700 29121 3734 29155
rect 5825 29121 5859 29155
rect 5917 29121 5951 29155
rect 7297 29121 7331 29155
rect 9505 29121 9539 29155
rect 10701 29121 10735 29155
rect 11161 29121 11195 29155
rect 11621 29121 11655 29155
rect 11805 29121 11839 29155
rect 12449 29121 12483 29155
rect 12909 29121 12943 29155
rect 13093 29121 13127 29155
rect 13282 29121 13316 29155
rect 15945 29121 15979 29155
rect 16948 29121 16982 29155
rect 19726 29121 19760 29155
rect 19993 29121 20027 29155
rect 20729 29121 20763 29155
rect 22057 29121 22091 29155
rect 22293 29121 22327 29155
rect 22477 29121 22511 29155
rect 22661 29121 22695 29155
rect 6193 29053 6227 29087
rect 7389 29053 7423 29087
rect 10149 29053 10183 29087
rect 10241 29053 10275 29087
rect 12357 29053 12391 29087
rect 13829 29053 13863 29087
rect 15577 29053 15611 29087
rect 16681 29053 16715 29087
rect 4813 28985 4847 29019
rect 6101 28985 6135 29019
rect 6837 28985 6871 29019
rect 9689 28985 9723 29019
rect 11345 28985 11379 29019
rect 18061 28985 18095 29019
rect 21925 28985 21959 29019
rect 23213 28985 23247 29019
rect 14086 28917 14120 28951
rect 3985 28713 4019 28747
rect 4445 28713 4479 28747
rect 7297 28713 7331 28747
rect 13737 28713 13771 28747
rect 14841 28713 14875 28747
rect 15301 28713 15335 28747
rect 17233 28713 17267 28747
rect 23765 28713 23799 28747
rect 6561 28645 6595 28679
rect 17417 28645 17451 28679
rect 22201 28645 22235 28679
rect 5181 28577 5215 28611
rect 7389 28577 7423 28611
rect 17785 28577 17819 28611
rect 21741 28577 21775 28611
rect 4169 28509 4203 28543
rect 4261 28509 4295 28543
rect 4537 28509 4571 28543
rect 7021 28509 7055 28543
rect 7113 28509 7147 28543
rect 8585 28509 8619 28543
rect 10241 28509 10275 28543
rect 10885 28509 10919 28543
rect 11345 28509 11379 28543
rect 13185 28509 13219 28543
rect 13558 28509 13592 28543
rect 15025 28509 15059 28543
rect 15117 28509 15151 28543
rect 15761 28509 15795 28543
rect 17601 28509 17635 28543
rect 17877 28509 17911 28543
rect 17970 28509 18004 28543
rect 18153 28509 18187 28543
rect 22028 28509 22062 28543
rect 22333 28509 22367 28543
rect 22753 28509 22787 28543
rect 22845 28509 22879 28543
rect 23218 28509 23252 28543
rect 23581 28509 23615 28543
rect 24409 28509 24443 28543
rect 24869 28509 24903 28543
rect 5448 28441 5482 28475
rect 6837 28441 6871 28475
rect 13369 28441 13403 28475
rect 13461 28441 13495 28475
rect 22477 28441 22511 28475
rect 22569 28441 22603 28475
rect 23029 28441 23063 28475
rect 23121 28441 23155 28475
rect 8401 28373 8435 28407
rect 10057 28373 10091 28407
rect 11069 28373 11103 28407
rect 11161 28373 11195 28407
rect 14105 28373 14139 28407
rect 15945 28373 15979 28407
rect 20269 28373 20303 28407
rect 23414 28373 23448 28407
rect 23949 28373 23983 28407
rect 24593 28373 24627 28407
rect 24685 28373 24719 28407
rect 4445 28169 4479 28203
rect 7021 28169 7055 28203
rect 11253 28169 11287 28203
rect 18061 28169 18095 28203
rect 18889 28169 18923 28203
rect 20821 28169 20855 28203
rect 22477 28169 22511 28203
rect 22937 28169 22971 28203
rect 25053 28169 25087 28203
rect 4813 28101 4847 28135
rect 9781 28101 9815 28135
rect 23581 28101 23615 28135
rect 25513 28101 25547 28135
rect 6929 28033 6963 28067
rect 12449 28033 12483 28067
rect 14473 28033 14507 28067
rect 14749 28033 14783 28067
rect 14933 28033 14967 28067
rect 15301 28033 15335 28067
rect 17969 28033 18003 28067
rect 20002 28033 20036 28067
rect 20269 28033 20303 28067
rect 20637 28033 20671 28067
rect 22293 28033 22327 28067
rect 22753 28033 22787 28067
rect 23029 28033 23063 28067
rect 23121 28033 23155 28067
rect 25237 28033 25271 28067
rect 25421 28033 25455 28067
rect 25610 28033 25644 28067
rect 4905 27965 4939 27999
rect 5089 27965 5123 27999
rect 7113 27965 7147 27999
rect 9045 27965 9079 27999
rect 9321 27965 9355 27999
rect 9505 27965 9539 27999
rect 18245 27965 18279 27999
rect 15485 27897 15519 27931
rect 23305 27965 23339 27999
rect 25973 27897 26007 27931
rect 6561 27829 6595 27863
rect 7573 27829 7607 27863
rect 12633 27829 12667 27863
rect 14473 27829 14507 27863
rect 17601 27829 17635 27863
rect 22017 27829 22051 27863
rect 22569 27829 22603 27863
rect 23121 27829 23155 27863
rect 25789 27829 25823 27863
rect 10241 27625 10275 27659
rect 19349 27625 19383 27659
rect 23673 27625 23707 27659
rect 25316 27625 25350 27659
rect 4353 27557 4387 27591
rect 8125 27557 8159 27591
rect 9505 27557 9539 27591
rect 11713 27557 11747 27591
rect 17601 27557 17635 27591
rect 18429 27557 18463 27591
rect 23305 27557 23339 27591
rect 26801 27557 26835 27591
rect 8953 27489 8987 27523
rect 9689 27489 9723 27523
rect 10701 27489 10735 27523
rect 14197 27489 14231 27523
rect 18245 27489 18279 27523
rect 19625 27489 19659 27523
rect 23765 27489 23799 27523
rect 24133 27489 24167 27523
rect 4077 27421 4111 27455
rect 4169 27421 4203 27455
rect 4445 27421 4479 27455
rect 7941 27421 7975 27455
rect 8401 27421 8435 27455
rect 9137 27421 9171 27455
rect 9781 27421 9815 27455
rect 11529 27421 11563 27455
rect 13645 27421 13679 27455
rect 14105 27421 14139 27455
rect 14381 27421 14415 27455
rect 14565 27421 14599 27455
rect 14933 27421 14967 27455
rect 15669 27421 15703 27455
rect 17969 27421 18003 27455
rect 18613 27421 18647 27455
rect 18889 27421 18923 27455
rect 19441 27421 19475 27455
rect 19717 27421 19751 27455
rect 19827 27421 19861 27455
rect 19993 27421 20027 27455
rect 20453 27421 20487 27455
rect 22753 27421 22787 27455
rect 23029 27421 23063 27455
rect 23173 27421 23207 27455
rect 23489 27421 23523 27455
rect 23857 27421 23891 27455
rect 24777 27421 24811 27455
rect 25053 27421 25087 27455
rect 10793 27353 10827 27387
rect 13369 27353 13403 27387
rect 15936 27353 15970 27387
rect 22937 27353 22971 27387
rect 23765 27353 23799 27387
rect 3893 27285 3927 27319
rect 8217 27285 8251 27319
rect 10701 27285 10735 27319
rect 11897 27285 11931 27319
rect 15117 27285 15151 27319
rect 17049 27285 17083 27319
rect 18061 27285 18095 27319
rect 18705 27285 18739 27319
rect 20177 27285 20211 27319
rect 20361 27285 20395 27319
rect 20637 27285 20671 27319
rect 24041 27285 24075 27319
rect 24961 27285 24995 27319
rect 4169 27081 4203 27115
rect 4445 27081 4479 27115
rect 11161 27081 11195 27115
rect 11529 27081 11563 27115
rect 15669 27081 15703 27115
rect 16405 27081 16439 27115
rect 21649 27081 21683 27115
rect 21925 27081 21959 27115
rect 23857 27081 23891 27115
rect 25881 27081 25915 27115
rect 3056 27013 3090 27047
rect 8861 27013 8895 27047
rect 9781 27013 9815 27047
rect 12265 27013 12299 27047
rect 18521 27013 18555 27047
rect 23397 27013 23431 27047
rect 4629 26945 4663 26979
rect 4813 26945 4847 26979
rect 4905 26945 4939 26979
rect 5825 26945 5859 26979
rect 5917 26945 5951 26979
rect 6193 26945 6227 26979
rect 6837 26945 6871 26979
rect 9137 26945 9171 26979
rect 9413 26945 9447 26979
rect 10057 26945 10091 26979
rect 10517 26945 10551 26979
rect 11345 26945 11379 26979
rect 11529 26945 11563 26979
rect 11713 26945 11747 26979
rect 11897 26945 11931 26979
rect 12541 26945 12575 26979
rect 13553 26945 13587 26979
rect 14473 26945 14507 26979
rect 14657 26945 14691 26979
rect 14841 26945 14875 26979
rect 15117 26945 15151 26979
rect 15301 26945 15335 26979
rect 16681 26945 16715 26979
rect 16865 26945 16899 26979
rect 17234 26945 17268 26979
rect 17417 26945 17451 26979
rect 18981 26945 19015 26979
rect 19164 26945 19198 26979
rect 19533 26945 19567 26979
rect 19717 26945 19751 26979
rect 21014 26945 21048 26979
rect 21465 26945 21499 26979
rect 25697 26945 25731 26979
rect 2789 26877 2823 26911
rect 6929 26877 6963 26911
rect 7113 26877 7147 26911
rect 7389 26877 7423 26911
rect 9229 26877 9263 26911
rect 9965 26877 9999 26911
rect 12633 26877 12667 26911
rect 17049 26877 17083 26911
rect 17141 26877 17175 26911
rect 18613 26877 18647 26911
rect 18797 26877 18831 26911
rect 19257 26877 19291 26911
rect 19349 26877 19383 26911
rect 21281 26877 21315 26911
rect 23673 26877 23707 26911
rect 25329 26877 25363 26911
rect 25605 26877 25639 26911
rect 10333 26809 10367 26843
rect 13737 26809 13771 26843
rect 5089 26741 5123 26775
rect 5641 26741 5675 26775
rect 6101 26741 6135 26775
rect 6469 26741 6503 26775
rect 14381 26741 14415 26775
rect 15485 26741 15519 26775
rect 18153 26741 18187 26775
rect 19901 26741 19935 26775
rect 4077 26537 4111 26571
rect 6653 26537 6687 26571
rect 8309 26537 8343 26571
rect 10333 26537 10367 26571
rect 10793 26537 10827 26571
rect 12633 26537 12667 26571
rect 15577 26537 15611 26571
rect 16405 26537 16439 26571
rect 21649 26537 21683 26571
rect 22201 26537 22235 26571
rect 23765 26537 23799 26571
rect 14289 26469 14323 26503
rect 17509 26469 17543 26503
rect 19257 26469 19291 26503
rect 29561 26469 29595 26503
rect 5273 26401 5307 26435
rect 11345 26401 11379 26435
rect 16865 26401 16899 26435
rect 17049 26401 17083 26435
rect 18061 26401 18095 26435
rect 19901 26401 19935 26435
rect 2973 26333 3007 26367
rect 3249 26333 3283 26367
rect 4261 26333 4295 26367
rect 5540 26333 5574 26367
rect 8033 26333 8067 26367
rect 8125 26333 8159 26367
rect 10517 26333 10551 26367
rect 11161 26333 11195 26367
rect 12725 26333 12759 26367
rect 12909 26333 12943 26367
rect 13185 26333 13219 26367
rect 13461 26333 13495 26367
rect 14468 26333 14502 26367
rect 14841 26333 14875 26367
rect 15117 26333 15151 26367
rect 16773 26333 16807 26367
rect 17969 26333 18003 26367
rect 18889 26333 18923 26367
rect 19441 26333 19475 26367
rect 21833 26333 21867 26367
rect 22017 26333 22051 26367
rect 22293 26333 22327 26367
rect 23213 26333 23247 26367
rect 23489 26333 23523 26367
rect 23633 26333 23667 26367
rect 13645 26265 13679 26299
rect 14565 26265 14599 26299
rect 14657 26265 14691 26299
rect 15209 26265 15243 26299
rect 18705 26265 18739 26299
rect 19625 26265 19659 26299
rect 21557 26265 21591 26299
rect 23121 26265 23155 26299
rect 23397 26265 23431 26299
rect 3065 26197 3099 26231
rect 7849 26197 7883 26231
rect 11253 26197 11287 26231
rect 11621 26197 11655 26231
rect 12173 26197 12207 26231
rect 14933 26197 14967 26231
rect 17877 26197 17911 26231
rect 18613 26197 18647 26231
rect 19073 26197 19107 26231
rect 5365 25993 5399 26027
rect 10241 25993 10275 26027
rect 10609 25993 10643 26027
rect 14824 25993 14858 26027
rect 15577 25993 15611 26027
rect 26985 25993 27019 26027
rect 9413 25925 9447 25959
rect 11529 25925 11563 25959
rect 12817 25925 12851 25959
rect 15209 25925 15243 25959
rect 1777 25857 1811 25891
rect 2044 25857 2078 25891
rect 3617 25857 3651 25891
rect 3884 25857 3918 25891
rect 5181 25857 5215 25891
rect 6377 25857 6411 25891
rect 6653 25857 6687 25891
rect 6745 25857 6779 25891
rect 8401 25857 8435 25891
rect 11161 25857 11195 25891
rect 11805 25857 11839 25891
rect 12357 25857 12391 25891
rect 14565 25857 14599 25891
rect 15020 25857 15054 25891
rect 15117 25857 15151 25891
rect 15393 25857 15427 25891
rect 15761 25857 15795 25891
rect 15926 25860 15960 25894
rect 16037 25857 16071 25891
rect 16129 25857 16163 25891
rect 16313 25857 16347 25891
rect 16497 25857 16531 25891
rect 17886 25857 17920 25891
rect 18521 25857 18555 25891
rect 18704 25857 18738 25891
rect 19073 25857 19107 25891
rect 19257 25857 19291 25891
rect 20554 25857 20588 25891
rect 20821 25857 20855 25891
rect 22017 25857 22051 25891
rect 23305 25857 23339 25891
rect 27169 25857 27203 25891
rect 9413 25789 9447 25823
rect 9505 25789 9539 25823
rect 10701 25789 10735 25823
rect 10793 25789 10827 25823
rect 11713 25789 11747 25823
rect 13001 25789 13035 25823
rect 18153 25789 18187 25823
rect 18797 25789 18831 25823
rect 18889 25789 18923 25823
rect 24961 25789 24995 25823
rect 25237 25789 25271 25823
rect 26709 25789 26743 25823
rect 6469 25721 6503 25755
rect 8953 25721 8987 25755
rect 11345 25721 11379 25755
rect 13185 25721 13219 25755
rect 3157 25653 3191 25687
rect 4997 25653 5031 25687
rect 6929 25653 6963 25687
rect 8217 25653 8251 25687
rect 11805 25653 11839 25687
rect 11989 25653 12023 25687
rect 12265 25653 12299 25687
rect 12541 25653 12575 25687
rect 13369 25653 13403 25687
rect 14381 25653 14415 25687
rect 16773 25653 16807 25687
rect 19441 25653 19475 25687
rect 21833 25653 21867 25687
rect 23581 25653 23615 25687
rect 2697 25449 2731 25483
rect 3157 25449 3191 25483
rect 3893 25449 3927 25483
rect 6653 25449 6687 25483
rect 9965 25449 9999 25483
rect 11529 25449 11563 25483
rect 12173 25449 12207 25483
rect 12265 25449 12299 25483
rect 13921 25449 13955 25483
rect 16589 25449 16623 25483
rect 22569 25449 22603 25483
rect 25237 25449 25271 25483
rect 26065 25449 26099 25483
rect 8677 25381 8711 25415
rect 13461 25381 13495 25415
rect 14841 25381 14875 25415
rect 19257 25381 19291 25415
rect 23305 25381 23339 25415
rect 24041 25381 24075 25415
rect 24593 25381 24627 25415
rect 24685 25381 24719 25415
rect 5273 25313 5307 25347
rect 7297 25313 7331 25347
rect 7481 25313 7515 25347
rect 10609 25313 10643 25347
rect 11621 25313 11655 25347
rect 11989 25313 12023 25347
rect 12357 25313 12391 25347
rect 17049 25313 17083 25347
rect 17141 25313 17175 25347
rect 18429 25313 18463 25347
rect 19717 25313 19751 25347
rect 19809 25313 19843 25347
rect 20821 25313 20855 25347
rect 2881 25245 2915 25279
rect 2973 25245 3007 25279
rect 3249 25245 3283 25279
rect 4072 25245 4106 25279
rect 4261 25245 4295 25279
rect 4445 25245 4479 25279
rect 5540 25245 5574 25279
rect 8493 25245 8527 25279
rect 9137 25245 9171 25279
rect 10333 25245 10367 25279
rect 12265 25245 12299 25279
rect 12909 25245 12943 25279
rect 13282 25245 13316 25279
rect 13737 25245 13771 25279
rect 14197 25245 14231 25279
rect 15020 25245 15054 25279
rect 15393 25245 15427 25279
rect 15577 25245 15611 25279
rect 16497 25245 16531 25279
rect 18337 25245 18371 25279
rect 20453 25245 20487 25279
rect 22753 25245 22787 25279
rect 23126 25245 23160 25279
rect 23489 25245 23523 25279
rect 23862 25245 23896 25279
rect 24225 25245 24259 25279
rect 24409 25245 24443 25279
rect 24869 25245 24903 25279
rect 25392 25245 25426 25279
rect 25513 25245 25547 25279
rect 25789 25245 25823 25279
rect 25881 25245 25915 25279
rect 4169 25177 4203 25211
rect 8125 25177 8159 25211
rect 8309 25177 8343 25211
rect 13093 25177 13127 25211
rect 13185 25177 13219 25211
rect 15117 25177 15151 25211
rect 15209 25177 15243 25211
rect 21097 25177 21131 25211
rect 22937 25177 22971 25211
rect 23029 25177 23063 25211
rect 23673 25177 23707 25211
rect 23765 25177 23799 25211
rect 24961 25177 24995 25211
rect 25605 25177 25639 25211
rect 26157 25177 26191 25211
rect 6837 25109 6871 25143
rect 7205 25109 7239 25143
rect 8953 25109 8987 25143
rect 10425 25109 10459 25143
rect 11805 25109 11839 25143
rect 12633 25109 12667 25143
rect 14381 25109 14415 25143
rect 16313 25109 16347 25143
rect 16957 25109 16991 25143
rect 17877 25109 17911 25143
rect 18245 25109 18279 25143
rect 19625 25109 19659 25143
rect 20269 25109 20303 25143
rect 20637 25109 20671 25143
rect 24225 25109 24259 25143
rect 7205 24905 7239 24939
rect 9229 24905 9263 24939
rect 9689 24905 9723 24939
rect 10333 24905 10367 24939
rect 10885 24905 10919 24939
rect 15585 24905 15619 24939
rect 18061 24905 18095 24939
rect 22017 24905 22051 24939
rect 23305 24905 23339 24939
rect 2973 24837 3007 24871
rect 7757 24837 7791 24871
rect 10241 24837 10275 24871
rect 13369 24837 13403 24871
rect 15301 24837 15335 24871
rect 18613 24837 18647 24871
rect 19717 24837 19751 24871
rect 25513 24837 25547 24871
rect 2697 24769 2731 24803
rect 2881 24769 2915 24803
rect 4445 24769 4479 24803
rect 4813 24769 4847 24803
rect 6929 24769 6963 24803
rect 7389 24769 7423 24803
rect 9597 24769 9631 24803
rect 9781 24769 9815 24803
rect 10701 24769 10735 24803
rect 12173 24769 12207 24803
rect 12265 24769 12299 24803
rect 12357 24769 12391 24803
rect 12725 24769 12759 24803
rect 15025 24769 15059 24803
rect 15209 24769 15243 24803
rect 15445 24769 15479 24803
rect 17877 24769 17911 24803
rect 20545 24769 20579 24803
rect 21097 24769 21131 24803
rect 21833 24769 21867 24803
rect 22109 24769 22143 24803
rect 25237 24769 25271 24803
rect 25421 24769 25455 24803
rect 25657 24769 25691 24803
rect 26065 24769 26099 24803
rect 26341 24769 26375 24803
rect 7481 24701 7515 24735
rect 10517 24701 10551 24735
rect 11069 24701 11103 24735
rect 11805 24701 11839 24735
rect 13093 24701 13127 24735
rect 18705 24701 18739 24735
rect 18797 24701 18831 24735
rect 19809 24701 19843 24735
rect 19901 24701 19935 24735
rect 24777 24701 24811 24735
rect 25053 24701 25087 24735
rect 4261 24633 4295 24667
rect 12909 24633 12943 24667
rect 18245 24633 18279 24667
rect 26249 24633 26283 24667
rect 26985 24633 27019 24667
rect 2513 24565 2547 24599
rect 4629 24565 4663 24599
rect 7113 24565 7147 24599
rect 9873 24565 9907 24599
rect 11253 24565 11287 24599
rect 11529 24565 11563 24599
rect 11989 24565 12023 24599
rect 12541 24565 12575 24599
rect 14841 24565 14875 24599
rect 15853 24565 15887 24599
rect 19349 24565 19383 24599
rect 20729 24565 20763 24599
rect 21189 24565 21223 24599
rect 25789 24565 25823 24599
rect 26525 24565 26559 24599
rect 26709 24565 26743 24599
rect 2789 24361 2823 24395
rect 4721 24361 4755 24395
rect 10609 24361 10643 24395
rect 10793 24361 10827 24395
rect 10977 24361 11011 24395
rect 18245 24361 18279 24395
rect 19717 24361 19751 24395
rect 22753 24361 22787 24395
rect 19257 24293 19291 24327
rect 22477 24293 22511 24327
rect 1409 24225 1443 24259
rect 3065 24225 3099 24259
rect 3525 24225 3559 24259
rect 4169 24225 4203 24259
rect 4261 24225 4295 24259
rect 6929 24225 6963 24259
rect 9505 24225 9539 24259
rect 10057 24225 10091 24259
rect 10425 24225 10459 24259
rect 11437 24225 11471 24259
rect 25789 24225 25823 24259
rect 2973 24157 3007 24191
rect 3249 24157 3283 24191
rect 3341 24157 3375 24191
rect 4077 24157 4111 24191
rect 4353 24157 4387 24191
rect 4537 24157 4571 24191
rect 4813 24157 4847 24191
rect 5089 24157 5123 24191
rect 9597 24157 9631 24191
rect 14381 24157 14415 24191
rect 16865 24157 16899 24191
rect 21097 24157 21131 24191
rect 21925 24157 21959 24191
rect 22201 24157 22235 24191
rect 22345 24157 22379 24191
rect 23305 24157 23339 24191
rect 23581 24157 23615 24191
rect 23678 24157 23712 24191
rect 24409 24157 24443 24191
rect 25513 24157 25547 24191
rect 1676 24089 1710 24123
rect 5356 24089 5390 24123
rect 7205 24089 7239 24123
rect 9505 24089 9539 24123
rect 11713 24089 11747 24123
rect 17132 24089 17166 24123
rect 19073 24089 19107 24123
rect 19441 24089 19475 24123
rect 20830 24089 20864 24123
rect 22109 24089 22143 24123
rect 23489 24089 23523 24123
rect 3893 24021 3927 24055
rect 6469 24021 6503 24055
rect 8677 24021 8711 24055
rect 9027 24021 9061 24055
rect 10241 24021 10275 24055
rect 13185 24021 13219 24055
rect 14565 24021 14599 24055
rect 23121 24021 23155 24055
rect 23874 24021 23908 24055
rect 24593 24021 24627 24055
rect 27261 24021 27295 24055
rect 2513 23817 2547 23851
rect 2605 23817 2639 23851
rect 3341 23817 3375 23851
rect 3617 23817 3651 23851
rect 5549 23817 5583 23851
rect 6377 23817 6411 23851
rect 6745 23817 6779 23851
rect 7389 23817 7423 23851
rect 9873 23817 9907 23851
rect 11897 23817 11931 23851
rect 12725 23817 12759 23851
rect 17509 23817 17543 23851
rect 17785 23817 17819 23851
rect 19993 23817 20027 23851
rect 23673 23817 23707 23851
rect 25513 23817 25547 23851
rect 1961 23749 1995 23783
rect 2973 23749 3007 23783
rect 4721 23749 4755 23783
rect 6837 23749 6871 23783
rect 9965 23749 9999 23783
rect 24041 23749 24075 23783
rect 2145 23681 2179 23715
rect 2401 23681 2435 23715
rect 2789 23681 2823 23715
rect 3433 23681 3467 23715
rect 3709 23681 3743 23715
rect 4353 23681 4387 23715
rect 4537 23681 4571 23715
rect 4813 23681 4847 23715
rect 4957 23681 4991 23715
rect 5733 23681 5767 23715
rect 5825 23681 5859 23715
rect 7573 23681 7607 23715
rect 10149 23681 10183 23715
rect 10517 23681 10551 23715
rect 12081 23681 12115 23715
rect 12909 23681 12943 23715
rect 13185 23681 13219 23715
rect 15301 23681 15335 23715
rect 15853 23681 15887 23715
rect 16221 23681 16255 23715
rect 16865 23681 16899 23715
rect 17877 23681 17911 23715
rect 18015 23681 18049 23715
rect 18246 23681 18280 23715
rect 18429 23681 18463 23715
rect 18705 23681 18739 23715
rect 19349 23681 19383 23715
rect 19532 23681 19566 23715
rect 19901 23681 19935 23715
rect 22017 23681 22051 23715
rect 22753 23681 22787 23715
rect 23489 23681 23523 23715
rect 2697 23613 2731 23647
rect 3157 23613 3191 23647
rect 6101 23613 6135 23647
rect 6929 23613 6963 23647
rect 11713 23613 11747 23647
rect 13369 23613 13403 23647
rect 13737 23613 13771 23647
rect 15209 23613 15243 23647
rect 18153 23613 18187 23647
rect 19625 23613 19659 23647
rect 19717 23613 19751 23647
rect 23765 23613 23799 23647
rect 13001 23545 13035 23579
rect 16037 23545 16071 23579
rect 16405 23545 16439 23579
rect 20269 23545 20303 23579
rect 4169 23477 4203 23511
rect 5089 23477 5123 23511
rect 6009 23477 6043 23511
rect 10241 23477 10275 23511
rect 10977 23477 11011 23511
rect 11713 23477 11747 23511
rect 15485 23477 15519 23511
rect 16681 23477 16715 23511
rect 18521 23477 18555 23511
rect 21833 23477 21867 23511
rect 22569 23477 22603 23511
rect 9689 23273 9723 23307
rect 13553 23273 13587 23307
rect 14381 23273 14415 23307
rect 19257 23273 19291 23307
rect 21005 23273 21039 23307
rect 23305 23273 23339 23307
rect 24593 23273 24627 23307
rect 18613 23205 18647 23239
rect 23121 23205 23155 23239
rect 4077 23137 4111 23171
rect 10057 23137 10091 23171
rect 10149 23137 10183 23171
rect 10349 23137 10383 23171
rect 11161 23137 11195 23171
rect 15669 23137 15703 23171
rect 19809 23137 19843 23171
rect 22753 23137 22787 23171
rect 1961 23069 1995 23103
rect 3801 23069 3835 23103
rect 3893 23069 3927 23103
rect 6101 23069 6135 23103
rect 8217 23069 8251 23103
rect 9965 23069 9999 23103
rect 10885 23069 10919 23103
rect 11069 23069 11103 23103
rect 11529 23069 11563 23103
rect 13277 23069 13311 23103
rect 13369 23069 13403 23103
rect 14197 23069 14231 23103
rect 15117 23069 15151 23103
rect 15301 23069 15335 23103
rect 18429 23069 18463 23103
rect 22937 23069 22971 23103
rect 23213 23069 23247 23103
rect 23489 23069 23523 23103
rect 23862 23069 23896 23103
rect 5834 23001 5868 23035
rect 7941 23001 7975 23035
rect 9321 23001 9355 23035
rect 9735 23001 9769 23035
rect 10609 23001 10643 23035
rect 10793 23001 10827 23035
rect 11345 23001 11379 23035
rect 11713 23001 11747 23035
rect 12909 23001 12943 23035
rect 13093 23001 13127 23035
rect 17141 23001 17175 23035
rect 18705 23001 18739 23035
rect 22477 23001 22511 23035
rect 23673 23001 23707 23035
rect 23765 23001 23799 23035
rect 24501 23001 24535 23035
rect 1869 22933 1903 22967
rect 4261 22933 4295 22967
rect 4721 22933 4755 22967
rect 6469 22933 6503 22967
rect 8309 22933 8343 22967
rect 10241 22933 10275 22967
rect 14933 22933 14967 22967
rect 19625 22933 19659 22967
rect 19717 22933 19751 22967
rect 24058 22933 24092 22967
rect 2789 22729 2823 22763
rect 4537 22729 4571 22763
rect 7205 22729 7239 22763
rect 8844 22729 8878 22763
rect 9781 22729 9815 22763
rect 9873 22729 9907 22763
rect 13277 22729 13311 22763
rect 19625 22729 19659 22763
rect 21833 22729 21867 22763
rect 22753 22729 22787 22763
rect 3157 22661 3191 22695
rect 3341 22661 3375 22695
rect 9137 22661 9171 22695
rect 9229 22661 9263 22695
rect 9597 22661 9631 22695
rect 9965 22661 9999 22695
rect 11069 22661 11103 22695
rect 11161 22661 11195 22695
rect 1409 22593 1443 22627
rect 1676 22593 1710 22627
rect 3893 22593 3927 22627
rect 4077 22593 4111 22627
rect 4169 22593 4203 22627
rect 4905 22593 4939 22627
rect 7389 22593 7423 22627
rect 7481 22593 7515 22627
rect 7849 22593 7883 22627
rect 7941 22593 7975 22627
rect 8401 22593 8435 22627
rect 9040 22593 9074 22627
rect 9413 22593 9447 22627
rect 10333 22593 10367 22627
rect 10972 22593 11006 22627
rect 11345 22593 11379 22627
rect 11529 22593 11563 22627
rect 11989 22593 12023 22627
rect 13093 22593 13127 22627
rect 13553 22593 13587 22627
rect 14473 22593 14507 22627
rect 14933 22593 14967 22627
rect 15577 22593 15611 22627
rect 15853 22593 15887 22627
rect 17049 22593 17083 22627
rect 17316 22593 17350 22627
rect 18613 22593 18647 22627
rect 18797 22593 18831 22627
rect 18981 22593 19015 22627
rect 19166 22593 19200 22627
rect 19349 22593 19383 22627
rect 20738 22593 20772 22627
rect 21005 22593 21039 22627
rect 21097 22593 21131 22627
rect 22017 22593 22051 22627
rect 22109 22593 22143 22627
rect 22569 22593 22603 22627
rect 23029 22593 23063 22627
rect 23949 22593 23983 22627
rect 4261 22525 4295 22559
rect 12081 22525 12115 22559
rect 12265 22525 12299 22559
rect 19073 22525 19107 22559
rect 24225 22525 24259 22559
rect 3709 22457 3743 22491
rect 4721 22457 4755 22491
rect 7665 22457 7699 22491
rect 7849 22457 7883 22491
rect 8217 22457 8251 22491
rect 10149 22457 10183 22491
rect 11621 22457 11655 22491
rect 14657 22457 14691 22491
rect 21281 22457 21315 22491
rect 22845 22457 22879 22491
rect 3065 22389 3099 22423
rect 3893 22389 3927 22423
rect 4261 22389 4295 22423
rect 8125 22389 8159 22423
rect 10793 22389 10827 22423
rect 13369 22389 13403 22423
rect 14749 22389 14783 22423
rect 15761 22389 15795 22423
rect 16037 22389 16071 22423
rect 18429 22389 18463 22423
rect 22293 22389 22327 22423
rect 25697 22389 25731 22423
rect 3801 22185 3835 22219
rect 7192 22185 7226 22219
rect 9045 22185 9079 22219
rect 21268 22185 21302 22219
rect 11713 22117 11747 22151
rect 15117 22117 15151 22151
rect 23497 22117 23531 22151
rect 10793 22049 10827 22083
rect 11069 22049 11103 22083
rect 15577 22049 15611 22083
rect 18521 22049 18555 22083
rect 18613 22049 18647 22083
rect 19533 22049 19567 22083
rect 19993 22049 20027 22083
rect 24133 22049 24167 22083
rect 2881 21981 2915 22015
rect 3985 21981 4019 22015
rect 4077 21981 4111 22015
rect 4905 21981 4939 22015
rect 6929 21981 6963 22015
rect 9183 21981 9217 22015
rect 9321 21981 9355 22015
rect 9597 21981 9631 22015
rect 9965 21981 9999 22015
rect 10425 21981 10459 22015
rect 10701 21981 10735 22015
rect 11897 21981 11931 22015
rect 15025 21981 15059 22015
rect 15301 21981 15335 22015
rect 19257 21981 19291 22015
rect 19440 21981 19474 22015
rect 19625 21981 19659 22015
rect 19809 21981 19843 22015
rect 21005 21981 21039 22015
rect 22937 21981 22971 22015
rect 23310 21981 23344 22015
rect 23857 21981 23891 22015
rect 5172 21913 5206 21947
rect 9689 21913 9723 21947
rect 10241 21913 10275 21947
rect 10609 21913 10643 21947
rect 12173 21913 12207 21947
rect 15853 21913 15887 21947
rect 23121 21913 23155 21947
rect 23213 21913 23247 21947
rect 23765 21913 23799 21947
rect 3065 21845 3099 21879
rect 4169 21845 4203 21879
rect 6285 21845 6319 21879
rect 8677 21845 8711 21879
rect 9873 21845 9907 21879
rect 13645 21845 13679 21879
rect 14841 21845 14875 21879
rect 17325 21845 17359 21879
rect 18061 21845 18095 21879
rect 18429 21845 18463 21879
rect 20085 21845 20119 21879
rect 22753 21845 22787 21879
rect 24041 21845 24075 21879
rect 7389 21641 7423 21675
rect 7941 21641 7975 21675
rect 10057 21641 10091 21675
rect 10977 21641 11011 21675
rect 12449 21641 12483 21675
rect 12541 21641 12575 21675
rect 15853 21641 15887 21675
rect 16865 21641 16899 21675
rect 19441 21641 19475 21675
rect 22017 21641 22051 21675
rect 23213 21641 23247 21675
rect 4077 21573 4111 21607
rect 6561 21573 6595 21607
rect 7481 21573 7515 21607
rect 9045 21573 9079 21607
rect 9689 21573 9723 21607
rect 12173 21573 12207 21607
rect 12357 21573 12391 21607
rect 12728 21573 12762 21607
rect 19809 21573 19843 21607
rect 22477 21573 22511 21607
rect 23581 21573 23615 21607
rect 3433 21505 3467 21539
rect 3618 21505 3652 21539
rect 3709 21505 3743 21539
rect 3835 21505 3869 21539
rect 4629 21505 4663 21539
rect 4813 21505 4847 21539
rect 4905 21505 4939 21539
rect 6009 21505 6043 21539
rect 6193 21505 6227 21539
rect 6377 21505 6411 21539
rect 6837 21505 6871 21539
rect 7021 21505 7055 21539
rect 7665 21505 7699 21539
rect 8125 21505 8159 21539
rect 9229 21505 9263 21539
rect 9413 21505 9447 21539
rect 10241 21505 10275 21539
rect 10793 21505 10827 21539
rect 11069 21505 11103 21539
rect 11161 21505 11195 21539
rect 15393 21505 15427 21539
rect 15669 21505 15703 21539
rect 16129 21505 16163 21539
rect 16497 21505 16531 21539
rect 16681 21505 16715 21539
rect 20913 21505 20947 21539
rect 21833 21505 21867 21539
rect 22333 21505 22367 21539
rect 22569 21505 22603 21539
rect 22753 21505 22787 21539
rect 23029 21505 23063 21539
rect 9948 21437 9982 21471
rect 10149 21437 10183 21471
rect 10701 21437 10735 21471
rect 13277 21437 13311 21471
rect 13461 21437 13495 21471
rect 13737 21437 13771 21471
rect 23305 21437 23339 21471
rect 5089 21369 5123 21403
rect 6745 21369 6779 21403
rect 6929 21369 6963 21403
rect 11345 21369 11379 21403
rect 15209 21369 15243 21403
rect 16313 21369 16347 21403
rect 16497 21369 16531 21403
rect 19625 21369 19659 21403
rect 21097 21369 21131 21403
rect 22201 21369 22235 21403
rect 4537 21301 4571 21335
rect 6101 21301 6135 21335
rect 7849 21301 7883 21335
rect 9505 21301 9539 21335
rect 10425 21301 10459 21335
rect 10793 21301 10827 21335
rect 11529 21301 11563 21335
rect 15577 21301 15611 21335
rect 22845 21301 22879 21335
rect 25053 21301 25087 21335
rect 5365 21097 5399 21131
rect 7389 21097 7423 21131
rect 9505 21097 9539 21131
rect 12633 21097 12667 21131
rect 13829 21097 13863 21131
rect 17325 21097 17359 21131
rect 23029 21097 23063 21131
rect 16497 21029 16531 21063
rect 23949 21029 23983 21063
rect 2881 20961 2915 20995
rect 4721 20961 4755 20995
rect 17233 20961 17267 20995
rect 17877 20961 17911 20995
rect 18613 20961 18647 20995
rect 3157 20893 3191 20927
rect 3341 20893 3375 20927
rect 3433 20893 3467 20927
rect 3801 20893 3835 20927
rect 4097 20893 4131 20927
rect 4353 20893 4387 20927
rect 5457 20893 5491 20927
rect 5733 20893 5767 20927
rect 7205 20893 7239 20927
rect 7757 20893 7791 20927
rect 7941 20893 7975 20927
rect 9413 20893 9447 20927
rect 12633 20893 12667 20927
rect 12817 20893 12851 20927
rect 13553 20893 13587 20927
rect 13645 20893 13679 20927
rect 14565 20893 14599 20927
rect 14841 20893 14875 20927
rect 16313 20893 16347 20927
rect 16773 20893 16807 20927
rect 18153 20893 18187 20927
rect 18337 20893 18371 20927
rect 18502 20893 18536 20927
rect 18705 20893 18739 20927
rect 18889 20893 18923 20927
rect 20729 20893 20763 20927
rect 22293 20893 22327 20927
rect 22569 20893 22603 20927
rect 23397 20893 23431 20927
rect 23581 20893 23615 20927
rect 23817 20893 23851 20927
rect 2614 20825 2648 20859
rect 2973 20825 3007 20859
rect 4537 20825 4571 20859
rect 4997 20825 5031 20859
rect 9229 20825 9263 20859
rect 14473 20825 14507 20859
rect 16129 20825 16163 20859
rect 17233 20825 17267 20859
rect 19073 20825 19107 20859
rect 20462 20825 20496 20859
rect 22026 20825 22060 20859
rect 23673 20825 23707 20859
rect 24133 20825 24167 20859
rect 1501 20757 1535 20791
rect 3525 20757 3559 20791
rect 3893 20757 3927 20791
rect 3985 20757 4019 20791
rect 4905 20757 4939 20791
rect 5549 20757 5583 20791
rect 7573 20757 7607 20791
rect 8125 20757 8159 20791
rect 9781 20757 9815 20791
rect 13001 20757 13035 20791
rect 13461 20757 13495 20791
rect 16681 20757 16715 20791
rect 17693 20757 17727 20791
rect 17785 20757 17819 20791
rect 19349 20757 19383 20791
rect 20913 20757 20947 20791
rect 22385 20757 22419 20791
rect 23213 20757 23247 20791
rect 2421 20553 2455 20587
rect 2513 20553 2547 20587
rect 3985 20553 4019 20587
rect 6101 20553 6135 20587
rect 6469 20553 6503 20587
rect 6929 20553 6963 20587
rect 9597 20553 9631 20587
rect 9873 20553 9907 20587
rect 10241 20553 10275 20587
rect 13829 20553 13863 20587
rect 17325 20553 17359 20587
rect 17785 20553 17819 20587
rect 20453 20553 20487 20587
rect 21925 20553 21959 20587
rect 25605 20553 25639 20587
rect 1869 20485 1903 20519
rect 2053 20485 2087 20519
rect 7389 20485 7423 20519
rect 10333 20485 10367 20519
rect 14381 20485 14415 20519
rect 21465 20485 21499 20519
rect 21649 20485 21683 20519
rect 24133 20485 24167 20519
rect 2605 20417 2639 20451
rect 3617 20417 3651 20451
rect 4445 20417 4479 20451
rect 4988 20417 5022 20451
rect 6561 20417 6595 20451
rect 6837 20417 6871 20451
rect 10701 20417 10735 20451
rect 11161 20417 11195 20451
rect 11253 20417 11287 20451
rect 11529 20417 11563 20451
rect 11805 20417 11839 20451
rect 11989 20417 12023 20451
rect 12173 20417 12207 20451
rect 12541 20417 12575 20451
rect 12633 20417 12667 20451
rect 12909 20417 12943 20451
rect 13185 20417 13219 20451
rect 13461 20417 13495 20451
rect 14105 20417 14139 20451
rect 14565 20417 14599 20451
rect 14749 20417 14783 20451
rect 15301 20417 15335 20451
rect 15393 20417 15427 20451
rect 15669 20417 15703 20451
rect 15853 20417 15887 20451
rect 16129 20417 16163 20451
rect 16313 20417 16347 20451
rect 16681 20417 16715 20451
rect 16773 20417 16807 20451
rect 17693 20417 17727 20451
rect 18613 20417 18647 20451
rect 18889 20417 18923 20451
rect 19809 20417 19843 20451
rect 19992 20417 20026 20451
rect 20361 20417 20395 20451
rect 20637 20417 20671 20451
rect 23673 20417 23707 20451
rect 23857 20417 23891 20451
rect 2309 20349 2343 20383
rect 3341 20349 3375 20383
rect 3525 20349 3559 20383
rect 4721 20349 4755 20383
rect 7113 20349 7147 20383
rect 9505 20349 9539 20383
rect 9689 20349 9723 20383
rect 10517 20349 10551 20383
rect 13993 20349 14027 20383
rect 14473 20349 14507 20383
rect 15117 20349 15151 20383
rect 15945 20349 15979 20383
rect 17877 20349 17911 20383
rect 20085 20349 20119 20383
rect 20177 20349 20211 20383
rect 23397 20349 23431 20383
rect 9137 20281 9171 20315
rect 10793 20281 10827 20315
rect 11621 20281 11655 20315
rect 12633 20281 12667 20315
rect 15025 20281 15059 20315
rect 19073 20281 19107 20315
rect 1685 20213 1719 20247
rect 4353 20213 4387 20247
rect 6653 20213 6687 20247
rect 8861 20213 8895 20247
rect 16681 20213 16715 20247
rect 17049 20213 17083 20247
rect 18797 20213 18831 20247
rect 2513 20009 2547 20043
rect 2881 20009 2915 20043
rect 5273 20009 5307 20043
rect 7941 20009 7975 20043
rect 8217 20009 8251 20043
rect 9045 20009 9079 20043
rect 10977 20009 11011 20043
rect 14565 20009 14599 20043
rect 14933 20009 14967 20043
rect 15761 20009 15795 20043
rect 16589 20009 16623 20043
rect 18153 20009 18187 20043
rect 22385 20009 22419 20043
rect 23213 20009 23247 20043
rect 24409 20009 24443 20043
rect 25145 20009 25179 20043
rect 3433 19941 3467 19975
rect 24133 19941 24167 19975
rect 3893 19873 3927 19907
rect 4629 19873 4663 19907
rect 4813 19873 4847 19907
rect 11253 19873 11287 19907
rect 12633 19873 12667 19907
rect 15393 19873 15427 19907
rect 2697 19805 2731 19839
rect 3063 19805 3097 19839
rect 3525 19805 3559 19839
rect 3985 19805 4019 19839
rect 6837 19805 6871 19839
rect 7757 19805 7791 19839
rect 8309 19805 8343 19839
rect 11069 19805 11103 19839
rect 11345 19805 11379 19839
rect 11438 19805 11472 19839
rect 11621 19805 11655 19839
rect 13001 19805 13035 19839
rect 13369 19805 13403 19839
rect 14565 19805 14599 19839
rect 14749 19805 14783 19839
rect 15577 19805 15611 19839
rect 16681 19805 16715 19839
rect 16865 19805 16899 19839
rect 17969 19805 18003 19839
rect 18245 19805 18279 19839
rect 22201 19805 22235 19839
rect 22661 19805 22695 19839
rect 22937 19805 22971 19839
rect 23081 19805 23115 19839
rect 23581 19805 23615 19839
rect 23954 19805 23988 19839
rect 24961 19805 24995 19839
rect 6469 19737 6503 19771
rect 6653 19737 6687 19771
rect 12817 19737 12851 19771
rect 13185 19737 13219 19771
rect 13553 19737 13587 19771
rect 22845 19737 22879 19771
rect 23765 19737 23799 19771
rect 23857 19737 23891 19771
rect 3065 19669 3099 19703
rect 4905 19669 4939 19703
rect 6285 19669 6319 19703
rect 18429 19669 18463 19703
rect 20269 19669 20303 19703
rect 22569 19669 22603 19703
rect 2789 19465 2823 19499
rect 4353 19465 4387 19499
rect 4813 19465 4847 19499
rect 8309 19465 8343 19499
rect 10701 19465 10735 19499
rect 11989 19465 12023 19499
rect 13185 19465 13219 19499
rect 14657 19465 14691 19499
rect 16865 19465 16899 19499
rect 18337 19465 18371 19499
rect 19993 19465 20027 19499
rect 21557 19465 21591 19499
rect 24685 19465 24719 19499
rect 26525 19465 26559 19499
rect 5273 19397 5307 19431
rect 10425 19397 10459 19431
rect 25053 19397 25087 19431
rect 4445 19329 4479 19363
rect 5129 19329 5163 19363
rect 5365 19329 5399 19363
rect 5549 19329 5583 19363
rect 6377 19329 6411 19363
rect 8125 19329 8159 19363
rect 8585 19329 8619 19363
rect 10517 19329 10551 19363
rect 10885 19329 10919 19363
rect 11069 19329 11103 19363
rect 11161 19329 11195 19363
rect 11345 19329 11379 19363
rect 11529 19329 11563 19363
rect 12173 19329 12207 19363
rect 12541 19329 12575 19363
rect 12909 19329 12943 19363
rect 13047 19329 13081 19363
rect 14841 19329 14875 19363
rect 16681 19329 16715 19363
rect 17141 19329 17175 19363
rect 17785 19329 17819 19363
rect 17877 19329 17911 19363
rect 18705 19329 18739 19363
rect 19349 19329 19383 19363
rect 19532 19332 19566 19366
rect 19901 19329 19935 19363
rect 20177 19329 20211 19363
rect 20433 19329 20467 19363
rect 24501 19329 24535 19363
rect 24777 19329 24811 19363
rect 2881 19261 2915 19295
rect 3065 19261 3099 19295
rect 4169 19261 4203 19295
rect 12633 19261 12667 19295
rect 18797 19261 18831 19295
rect 18981 19261 19015 19295
rect 19625 19261 19659 19295
rect 19717 19261 19751 19295
rect 4997 19193 5031 19227
rect 10977 19193 11011 19227
rect 2421 19125 2455 19159
rect 5641 19125 5675 19159
rect 6561 19125 6595 19159
rect 8769 19125 8803 19159
rect 11713 19125 11747 19159
rect 17325 19125 17359 19159
rect 7481 18921 7515 18955
rect 13921 18921 13955 18955
rect 19073 18921 19107 18955
rect 19993 18921 20027 18955
rect 22293 18921 22327 18955
rect 22569 18921 22603 18955
rect 23765 18921 23799 18955
rect 25973 18921 26007 18955
rect 11989 18853 12023 18887
rect 12909 18853 12943 18887
rect 23397 18853 23431 18887
rect 24041 18853 24075 18887
rect 24869 18853 24903 18887
rect 25513 18853 25547 18887
rect 2312 18785 2346 18819
rect 2605 18785 2639 18819
rect 7757 18785 7791 18819
rect 7849 18785 7883 18819
rect 9873 18785 9907 18819
rect 11345 18785 11379 18819
rect 11621 18785 11655 18819
rect 11805 18785 11839 18819
rect 14473 18785 14507 18819
rect 14933 18785 14967 18819
rect 16037 18785 16071 18819
rect 16497 18785 16531 18819
rect 18521 18785 18555 18819
rect 19349 18785 19383 18819
rect 20361 18785 20395 18819
rect 20453 18785 20487 18819
rect 20913 18785 20947 18819
rect 2053 18717 2087 18751
rect 5089 18717 5123 18751
rect 5365 18717 5399 18751
rect 5641 18717 5675 18751
rect 5825 18717 5859 18751
rect 7665 18717 7699 18751
rect 7941 18717 7975 18751
rect 8125 18717 8159 18751
rect 8309 18717 8343 18751
rect 8401 18717 8435 18751
rect 9597 18717 9631 18751
rect 9781 18717 9815 18751
rect 10057 18717 10091 18751
rect 10241 18717 10275 18751
rect 10425 18717 10459 18751
rect 11161 18717 11195 18751
rect 11437 18717 11471 18751
rect 12081 18717 12115 18751
rect 12173 18717 12207 18751
rect 12541 18717 12575 18751
rect 12725 18717 12759 18751
rect 13001 18717 13035 18751
rect 13369 18717 13403 18751
rect 13461 18717 13495 18751
rect 13737 18717 13771 18751
rect 14197 18717 14231 18751
rect 14362 18717 14396 18751
rect 14565 18717 14599 18751
rect 14749 18717 14783 18751
rect 15209 18717 15243 18751
rect 15485 18717 15519 18751
rect 15669 18717 15703 18751
rect 15853 18717 15887 18751
rect 16129 18717 16163 18751
rect 16313 18717 16347 18751
rect 18889 18717 18923 18751
rect 19625 18717 19659 18751
rect 20085 18717 20119 18751
rect 20268 18717 20302 18751
rect 20637 18717 20671 18751
rect 22753 18717 22787 18751
rect 22845 18717 22879 18751
rect 23029 18717 23063 18751
rect 23265 18717 23299 18751
rect 23581 18717 23615 18751
rect 24685 18717 24719 18751
rect 25145 18717 25179 18751
rect 25329 18717 25363 18751
rect 25789 18717 25823 18751
rect 1869 18649 1903 18683
rect 5733 18649 5767 18683
rect 6070 18649 6104 18683
rect 10977 18649 11011 18683
rect 12449 18649 12483 18683
rect 15117 18649 15151 18683
rect 16773 18649 16807 18683
rect 18705 18649 18739 18683
rect 20821 18649 20855 18683
rect 21158 18649 21192 18683
rect 23121 18649 23155 18683
rect 23857 18649 23891 18683
rect 2421 18581 2455 18615
rect 2513 18581 2547 18615
rect 2697 18581 2731 18615
rect 3801 18581 3835 18615
rect 5089 18581 5123 18615
rect 5273 18581 5307 18615
rect 7205 18581 7239 18615
rect 10517 18581 10551 18615
rect 12173 18581 12207 18615
rect 15301 18581 15335 18615
rect 18245 18581 18279 18615
rect 19533 18581 19567 18615
rect 24961 18581 24995 18615
rect 1869 18377 1903 18411
rect 1961 18377 1995 18411
rect 3617 18377 3651 18411
rect 3985 18377 4019 18411
rect 7481 18377 7515 18411
rect 9965 18377 9999 18411
rect 13001 18377 13035 18411
rect 17049 18377 17083 18411
rect 24869 18377 24903 18411
rect 2421 18309 2455 18343
rect 3065 18309 3099 18343
rect 3157 18309 3191 18343
rect 8309 18309 8343 18343
rect 11161 18309 11195 18343
rect 13829 18309 13863 18343
rect 15393 18309 15427 18343
rect 15761 18309 15795 18343
rect 2605 18241 2639 18275
rect 2789 18241 2823 18275
rect 2881 18241 2915 18275
rect 3301 18241 3335 18275
rect 4629 18241 4663 18275
rect 6009 18241 6043 18275
rect 7573 18241 7607 18275
rect 7757 18241 7791 18275
rect 8033 18241 8067 18275
rect 11345 18241 11379 18275
rect 11529 18241 11563 18275
rect 12357 18241 12391 18275
rect 12725 18241 12759 18275
rect 13737 18241 13771 18275
rect 14013 18241 14047 18275
rect 14289 18241 14323 18275
rect 14749 18241 14783 18275
rect 15025 18241 15059 18275
rect 15577 18241 15611 18275
rect 16681 18241 16715 18275
rect 18705 18241 18739 18275
rect 19717 18241 19751 18275
rect 22661 18241 22695 18275
rect 23121 18241 23155 18275
rect 2145 18173 2179 18207
rect 4077 18173 4111 18207
rect 4169 18173 4203 18207
rect 9781 18173 9815 18207
rect 12541 18173 12575 18207
rect 12633 18173 12667 18207
rect 12817 18173 12851 18207
rect 16773 18173 16807 18207
rect 19809 18173 19843 18207
rect 19901 18173 19935 18207
rect 23397 18173 23431 18207
rect 4445 18105 4479 18139
rect 7849 18105 7883 18139
rect 14105 18105 14139 18139
rect 14841 18105 14875 18139
rect 19349 18105 19383 18139
rect 1501 18037 1535 18071
rect 3433 18037 3467 18071
rect 5917 18037 5951 18071
rect 11069 18037 11103 18071
rect 11713 18037 11747 18071
rect 13553 18037 13587 18071
rect 15209 18037 15243 18071
rect 16681 18037 16715 18071
rect 18889 18037 18923 18071
rect 20913 18037 20947 18071
rect 22753 18037 22787 18071
rect 9229 17833 9263 17867
rect 11989 17833 12023 17867
rect 12449 17833 12483 17867
rect 13369 17833 13403 17867
rect 15117 17833 15151 17867
rect 17877 17833 17911 17867
rect 20085 17833 20119 17867
rect 6653 17765 6687 17799
rect 7113 17765 7147 17799
rect 10977 17765 11011 17799
rect 12173 17765 12207 17799
rect 14197 17765 14231 17799
rect 16681 17765 16715 17799
rect 17417 17765 17451 17799
rect 13553 17697 13587 17731
rect 15117 17697 15151 17731
rect 15485 17697 15519 17731
rect 15669 17697 15703 17731
rect 15945 17697 15979 17731
rect 19441 17697 19475 17731
rect 20453 17697 20487 17731
rect 22477 17697 22511 17731
rect 24593 17697 24627 17731
rect 1409 17629 1443 17663
rect 3893 17629 3927 17663
rect 6469 17629 6503 17663
rect 6561 17629 6595 17663
rect 6745 17629 6779 17663
rect 6929 17629 6963 17663
rect 7849 17629 7883 17663
rect 8125 17629 8159 17663
rect 9781 17629 9815 17663
rect 10793 17629 10827 17663
rect 10885 17629 10919 17663
rect 11161 17629 11195 17663
rect 11529 17629 11563 17663
rect 11805 17629 11839 17663
rect 11989 17629 12023 17663
rect 12541 17629 12575 17663
rect 12725 17629 12759 17663
rect 13277 17629 13311 17663
rect 13369 17629 13403 17663
rect 13461 17629 13495 17663
rect 14105 17629 14139 17663
rect 15577 17629 15611 17663
rect 16037 17629 16071 17663
rect 16773 17629 16807 17663
rect 17233 17629 17267 17663
rect 18245 17629 18279 17663
rect 18429 17629 18463 17663
rect 18521 17629 18555 17663
rect 1654 17561 1688 17595
rect 4138 17561 4172 17595
rect 9597 17561 9631 17595
rect 9965 17561 9999 17595
rect 18649 17626 18683 17660
rect 18797 17629 18831 17663
rect 20177 17629 20211 17663
rect 20360 17629 20394 17663
rect 20545 17629 20579 17663
rect 20729 17629 20763 17663
rect 22937 17629 22971 17663
rect 23213 17629 23247 17663
rect 15209 17561 15243 17595
rect 19625 17561 19659 17595
rect 20913 17561 20947 17595
rect 22210 17561 22244 17595
rect 24869 17561 24903 17595
rect 2789 17493 2823 17527
rect 3065 17493 3099 17527
rect 5273 17493 5307 17527
rect 6285 17493 6319 17527
rect 8125 17493 8159 17527
rect 11253 17493 11287 17527
rect 11713 17493 11747 17527
rect 13001 17493 13035 17527
rect 13461 17493 13495 17527
rect 16221 17493 16255 17527
rect 18153 17493 18187 17527
rect 19717 17493 19751 17527
rect 21097 17493 21131 17527
rect 23121 17493 23155 17527
rect 23397 17493 23431 17527
rect 26341 17493 26375 17527
rect 2237 17289 2271 17323
rect 2605 17289 2639 17323
rect 4169 17289 4203 17323
rect 7573 17289 7607 17323
rect 8861 17289 8895 17323
rect 10793 17289 10827 17323
rect 11621 17289 11655 17323
rect 12633 17289 12667 17323
rect 15025 17289 15059 17323
rect 17049 17289 17083 17323
rect 17693 17289 17727 17323
rect 19625 17289 19659 17323
rect 21097 17289 21131 17323
rect 25513 17289 25547 17323
rect 25789 17289 25823 17323
rect 4997 17221 5031 17255
rect 6837 17221 6871 17255
rect 6929 17221 6963 17255
rect 13737 17221 13771 17255
rect 18490 17221 18524 17255
rect 24777 17221 24811 17255
rect 25605 17221 25639 17255
rect 3065 17153 3099 17187
rect 3250 17153 3284 17187
rect 3617 17153 3651 17187
rect 3709 17153 3743 17187
rect 5181 17153 5215 17187
rect 6561 17153 6595 17187
rect 7205 17153 7239 17187
rect 7461 17153 7495 17187
rect 7849 17153 7883 17187
rect 8217 17153 8251 17187
rect 8677 17153 8711 17187
rect 9321 17153 9355 17187
rect 9413 17153 9447 17187
rect 9680 17153 9714 17187
rect 11529 17153 11563 17187
rect 12725 17153 12759 17187
rect 12909 17153 12943 17187
rect 13093 17153 13127 17187
rect 13369 17153 13403 17187
rect 13553 17153 13587 17187
rect 15577 17153 15611 17187
rect 15853 17153 15887 17187
rect 16129 17153 16163 17187
rect 16313 17153 16347 17187
rect 16681 17153 16715 17187
rect 17417 17153 17451 17187
rect 17509 17153 17543 17187
rect 17969 17153 18003 17187
rect 18245 17153 18279 17187
rect 24501 17153 24535 17187
rect 24685 17153 24719 17187
rect 24921 17153 24955 17187
rect 25329 17153 25363 17187
rect 2697 17085 2731 17119
rect 2881 17085 2915 17119
rect 4261 17085 4295 17119
rect 4445 17085 4479 17119
rect 6745 17085 6779 17119
rect 7665 17085 7699 17119
rect 7757 17085 7791 17119
rect 8401 17085 8435 17119
rect 9045 17085 9079 17119
rect 13277 17085 13311 17119
rect 15945 17085 15979 17119
rect 16773 17085 16807 17119
rect 22661 17085 22695 17119
rect 24133 17085 24167 17119
rect 24409 17085 24443 17119
rect 7941 17017 7975 17051
rect 17233 17017 17267 17051
rect 25053 17017 25087 17051
rect 3801 16949 3835 16983
rect 4905 16949 4939 16983
rect 7205 16949 7239 16983
rect 8493 16949 8527 16983
rect 9229 16949 9263 16983
rect 16681 16949 16715 16983
rect 17785 16949 17819 16983
rect 2697 16745 2731 16779
rect 7573 16745 7607 16779
rect 8585 16745 8619 16779
rect 13001 16745 13035 16779
rect 13277 16745 13311 16779
rect 13553 16745 13587 16779
rect 14749 16745 14783 16779
rect 22661 16745 22695 16779
rect 23397 16745 23431 16779
rect 23857 16745 23891 16779
rect 25145 16745 25179 16779
rect 7021 16677 7055 16711
rect 7297 16677 7331 16711
rect 8401 16677 8435 16711
rect 9965 16677 9999 16711
rect 18521 16677 18555 16711
rect 4813 16609 4847 16643
rect 5365 16609 5399 16643
rect 7665 16609 7699 16643
rect 9321 16609 9355 16643
rect 9505 16609 9539 16643
rect 10057 16609 10091 16643
rect 11529 16609 11563 16643
rect 13277 16609 13311 16643
rect 15117 16609 15151 16643
rect 20269 16609 20303 16643
rect 20361 16609 20395 16643
rect 22293 16609 22327 16643
rect 2789 16541 2823 16575
rect 4629 16541 4663 16575
rect 5632 16541 5666 16575
rect 7389 16541 7423 16575
rect 7941 16541 7975 16575
rect 8677 16541 8711 16575
rect 9229 16541 9263 16575
rect 9597 16541 9631 16575
rect 11253 16541 11287 16575
rect 11437 16541 11471 16575
rect 11713 16541 11747 16575
rect 11989 16541 12023 16575
rect 12357 16541 12391 16575
rect 12633 16541 12667 16575
rect 13369 16541 13403 16575
rect 13461 16541 13495 16575
rect 14381 16541 14415 16575
rect 14841 16541 14875 16575
rect 17601 16541 17635 16575
rect 18061 16541 18095 16575
rect 18337 16541 18371 16575
rect 19993 16541 20027 16575
rect 20176 16541 20210 16575
rect 20545 16541 20579 16575
rect 22845 16541 22879 16575
rect 23121 16541 23155 16575
rect 23265 16541 23299 16575
rect 23581 16541 23615 16575
rect 24041 16541 24075 16575
rect 24409 16541 24443 16575
rect 24961 16541 24995 16575
rect 25697 16541 25731 16575
rect 26065 16541 26099 16575
rect 2973 16473 3007 16507
rect 8033 16473 8067 16507
rect 8217 16473 8251 16507
rect 12725 16473 12759 16507
rect 15393 16473 15427 16507
rect 20729 16473 20763 16507
rect 22026 16473 22060 16507
rect 23029 16473 23063 16507
rect 4261 16405 4295 16439
rect 4721 16405 4755 16439
rect 6745 16405 6779 16439
rect 14473 16405 14507 16439
rect 16865 16405 16899 16439
rect 17417 16405 17451 16439
rect 18245 16405 18279 16439
rect 20913 16405 20947 16439
rect 23765 16405 23799 16439
rect 24133 16405 24167 16439
rect 24593 16405 24627 16439
rect 25881 16405 25915 16439
rect 26249 16405 26283 16439
rect 3893 16201 3927 16235
rect 4629 16201 4663 16235
rect 7205 16201 7239 16235
rect 8401 16201 8435 16235
rect 9413 16201 9447 16235
rect 16129 16201 16163 16235
rect 18153 16201 18187 16235
rect 18981 16201 19015 16235
rect 19441 16201 19475 16235
rect 21097 16201 21131 16235
rect 3157 16133 3191 16167
rect 7849 16133 7883 16167
rect 8585 16133 8619 16167
rect 14749 16133 14783 16167
rect 18521 16133 18555 16167
rect 18613 16133 18647 16167
rect 2145 16065 2179 16099
rect 3433 16065 3467 16099
rect 3709 16065 3743 16099
rect 4779 16065 4813 16099
rect 5089 16065 5123 16099
rect 5549 16065 5583 16099
rect 5825 16065 5859 16099
rect 7389 16065 7423 16099
rect 8033 16065 8067 16099
rect 8217 16065 8251 16099
rect 8861 16065 8895 16099
rect 9505 16065 9539 16099
rect 15393 16065 15427 16099
rect 15945 16065 15979 16099
rect 17969 16065 18003 16099
rect 19349 16065 19383 16099
rect 19993 16065 20027 16099
rect 20176 16068 20210 16102
rect 20407 16065 20441 16099
rect 20545 16065 20579 16099
rect 24961 16065 24995 16099
rect 2237 15997 2271 16031
rect 2421 15997 2455 16031
rect 3525 15997 3559 16031
rect 5181 15997 5215 16031
rect 5733 15997 5767 16031
rect 8677 15997 8711 16031
rect 15025 15997 15059 16031
rect 18797 15997 18831 16031
rect 19625 15997 19659 16031
rect 20269 15997 20303 16031
rect 25237 15997 25271 16031
rect 2881 15929 2915 15963
rect 9045 15929 9079 15963
rect 20821 15929 20855 15963
rect 1777 15861 1811 15895
rect 2697 15861 2731 15895
rect 3433 15861 3467 15895
rect 5365 15861 5399 15895
rect 6653 15861 6687 15895
rect 7665 15861 7699 15895
rect 8217 15861 8251 15895
rect 8769 15861 8803 15895
rect 9689 15861 9723 15895
rect 13277 15861 13311 15895
rect 15209 15861 15243 15895
rect 17785 15861 17819 15895
rect 20637 15861 20671 15895
rect 26709 15861 26743 15895
rect 2145 15657 2179 15691
rect 2973 15657 3007 15691
rect 3157 15657 3191 15691
rect 5365 15657 5399 15691
rect 8401 15657 8435 15691
rect 10793 15657 10827 15691
rect 12725 15657 12759 15691
rect 14657 15657 14691 15691
rect 17509 15657 17543 15691
rect 18521 15657 18555 15691
rect 20269 15657 20303 15691
rect 24593 15657 24627 15691
rect 25329 15657 25363 15691
rect 4169 15589 4203 15623
rect 8953 15589 8987 15623
rect 24133 15589 24167 15623
rect 3893 15521 3927 15555
rect 7297 15521 7331 15555
rect 2329 15453 2363 15487
rect 2789 15453 2823 15487
rect 2973 15453 3007 15487
rect 6745 15453 6779 15487
rect 7021 15453 7055 15487
rect 7205 15453 7239 15487
rect 7390 15453 7424 15487
rect 7573 15453 7607 15487
rect 7757 15453 7791 15487
rect 7932 15453 7966 15487
rect 8033 15453 8067 15487
rect 8217 15453 8251 15487
rect 8309 15453 8343 15487
rect 8585 15453 8619 15487
rect 6500 15385 6534 15419
rect 6837 15385 6871 15419
rect 9045 15521 9079 15555
rect 10977 15521 11011 15555
rect 11253 15521 11287 15555
rect 17969 15521 18003 15555
rect 14841 15453 14875 15487
rect 16129 15453 16163 15487
rect 17693 15453 17727 15487
rect 17858 15453 17892 15487
rect 18061 15453 18095 15487
rect 18245 15453 18279 15487
rect 18705 15453 18739 15487
rect 21382 15453 21416 15487
rect 21649 15453 21683 15487
rect 21741 15453 21775 15487
rect 23581 15453 23615 15487
rect 23765 15453 23799 15487
rect 23857 15453 23891 15487
rect 24001 15453 24035 15487
rect 24409 15453 24443 15487
rect 24685 15453 24719 15487
rect 24777 15453 24811 15487
rect 25150 15453 25184 15487
rect 9321 15385 9355 15419
rect 13369 15385 13403 15419
rect 16396 15385 16430 15419
rect 22008 15385 22042 15419
rect 24961 15385 24995 15419
rect 25053 15385 25087 15419
rect 4353 15317 4387 15351
rect 8677 15317 8711 15351
rect 8953 15317 8987 15351
rect 18337 15317 18371 15351
rect 23121 15317 23155 15351
rect 24685 15317 24719 15351
rect 25513 15317 25547 15351
rect 2789 15113 2823 15147
rect 3341 15113 3375 15147
rect 4353 15113 4387 15147
rect 4813 15113 4847 15147
rect 6469 15113 6503 15147
rect 7757 15113 7791 15147
rect 8217 15113 8251 15147
rect 10609 15113 10643 15147
rect 11713 15113 11747 15147
rect 16405 15113 16439 15147
rect 17325 15113 17359 15147
rect 17693 15113 17727 15147
rect 19257 15113 19291 15147
rect 19809 15113 19843 15147
rect 23857 15113 23891 15147
rect 24317 15113 24351 15147
rect 1676 15045 1710 15079
rect 4445 15045 4479 15079
rect 7113 15045 7147 15079
rect 7205 15045 7239 15079
rect 4997 14977 5031 15011
rect 6561 14977 6595 15011
rect 7849 14977 7883 15011
rect 8033 14977 8067 15011
rect 8677 14977 8711 15011
rect 8769 14977 8803 15011
rect 9045 14977 9079 15011
rect 9321 14977 9355 15011
rect 9505 14977 9539 15011
rect 9689 14977 9723 15011
rect 10057 14977 10091 15011
rect 10793 14977 10827 15011
rect 11069 14977 11103 15011
rect 11529 14977 11563 15011
rect 12449 14977 12483 15011
rect 12633 14977 12667 15011
rect 12725 14977 12759 15011
rect 12822 14977 12856 15011
rect 15485 14977 15519 15011
rect 15577 14977 15611 15011
rect 16681 14977 16715 15011
rect 16846 14977 16880 15011
rect 17049 14977 17083 15011
rect 17233 14977 17267 15011
rect 18144 15045 18178 15079
rect 25053 15045 25087 15079
rect 17877 14977 17911 15011
rect 20922 14977 20956 15011
rect 22733 14977 22767 15011
rect 24225 14977 24259 15011
rect 24501 14977 24535 15011
rect 24777 14977 24811 15011
rect 1409 14909 1443 14943
rect 3433 14909 3467 14943
rect 3617 14909 3651 14943
rect 4537 14909 4571 14943
rect 7297 14909 7331 14943
rect 9229 14909 9263 14943
rect 13369 14909 13403 14943
rect 13645 14909 13679 14943
rect 16957 14909 16991 14943
rect 17693 14909 17727 14943
rect 21189 14909 21223 14943
rect 22477 14909 22511 14943
rect 2973 14841 3007 14875
rect 8953 14841 8987 14875
rect 9689 14841 9723 14875
rect 11253 14841 11287 14875
rect 13001 14841 13035 14875
rect 15301 14841 15335 14875
rect 24041 14841 24075 14875
rect 3985 14773 4019 14807
rect 6745 14773 6779 14807
rect 8493 14773 8527 14807
rect 13277 14773 13311 14807
rect 15117 14773 15151 14807
rect 15761 14773 15795 14807
rect 17509 14773 17543 14807
rect 24685 14773 24719 14807
rect 26525 14773 26559 14807
rect 3065 14569 3099 14603
rect 4537 14569 4571 14603
rect 5641 14569 5675 14603
rect 10793 14569 10827 14603
rect 11161 14569 11195 14603
rect 16497 14569 16531 14603
rect 18981 14569 19015 14603
rect 22017 14569 22051 14603
rect 25605 14569 25639 14603
rect 10701 14501 10735 14535
rect 16773 14501 16807 14535
rect 22385 14501 22419 14535
rect 5089 14433 5123 14467
rect 13553 14433 13587 14467
rect 18613 14433 18647 14467
rect 19533 14433 19567 14467
rect 20177 14433 20211 14467
rect 2513 14365 2547 14399
rect 2933 14365 2967 14399
rect 3249 14365 3283 14399
rect 5549 14365 5583 14399
rect 7113 14365 7147 14399
rect 8309 14365 8343 14399
rect 8401 14365 8435 14399
rect 10425 14365 10459 14399
rect 10701 14365 10735 14399
rect 10977 14365 11011 14399
rect 13829 14365 13863 14399
rect 15117 14365 15151 14399
rect 16313 14365 16347 14399
rect 16589 14365 16623 14399
rect 17417 14365 17451 14399
rect 17877 14365 17911 14399
rect 18337 14365 18371 14399
rect 18502 14365 18536 14399
rect 18705 14365 18739 14399
rect 18889 14365 18923 14399
rect 19257 14365 19291 14399
rect 19440 14365 19474 14399
rect 19625 14365 19659 14399
rect 19809 14365 19843 14399
rect 21465 14365 21499 14399
rect 21838 14365 21872 14399
rect 25421 14365 25455 14399
rect 2697 14297 2731 14331
rect 2789 14297 2823 14331
rect 4905 14297 4939 14331
rect 5365 14297 5399 14331
rect 13277 14297 13311 14331
rect 19993 14297 20027 14331
rect 21649 14297 21683 14331
rect 21741 14297 21775 14331
rect 3341 14229 3375 14263
rect 4997 14229 5031 14263
rect 7021 14229 7055 14263
rect 7941 14229 7975 14263
rect 8217 14229 8251 14263
rect 10609 14229 10643 14263
rect 11805 14229 11839 14263
rect 13645 14229 13679 14263
rect 14933 14229 14967 14263
rect 17601 14229 17635 14263
rect 17693 14229 17727 14263
rect 18153 14229 18187 14263
rect 22293 14229 22327 14263
rect 3433 14025 3467 14059
rect 4997 14025 5031 14059
rect 5733 14025 5767 14059
rect 6653 14025 6687 14059
rect 9321 14025 9355 14059
rect 10057 14025 10091 14059
rect 10149 14025 10183 14059
rect 10793 14025 10827 14059
rect 12374 14025 12408 14059
rect 13553 14025 13587 14059
rect 14105 14025 14139 14059
rect 16405 14025 16439 14059
rect 18705 14025 18739 14059
rect 19809 14025 19843 14059
rect 3065 13957 3099 13991
rect 3249 13957 3283 13991
rect 3884 13957 3918 13991
rect 7389 13957 7423 13991
rect 8208 13957 8242 13991
rect 12633 13957 12667 13991
rect 19073 13957 19107 13991
rect 20922 13957 20956 13991
rect 2513 13889 2547 13923
rect 2697 13889 2731 13923
rect 2789 13889 2823 13923
rect 2881 13889 2915 13923
rect 3341 13889 3375 13923
rect 5181 13889 5215 13923
rect 5583 13889 5617 13923
rect 6745 13889 6779 13923
rect 7021 13889 7055 13923
rect 7114 13889 7148 13923
rect 7297 13889 7331 13923
rect 9873 13889 9907 13923
rect 10333 13889 10367 13923
rect 10609 13889 10643 13923
rect 11805 13889 11839 13923
rect 11989 13889 12023 13923
rect 12081 13889 12115 13923
rect 12225 13889 12259 13923
rect 13369 13889 13403 13923
rect 14013 13889 14047 13923
rect 14289 13889 14323 13923
rect 15025 13889 15059 13923
rect 15292 13889 15326 13923
rect 16865 13889 16899 13923
rect 17141 13889 17175 13923
rect 17408 13889 17442 13923
rect 22100 13889 22134 13923
rect 23664 13889 23698 13923
rect 24961 13889 24995 13923
rect 25217 13889 25251 13923
rect 3617 13821 3651 13855
rect 5273 13821 5307 13855
rect 6929 13821 6963 13855
rect 7941 13821 7975 13855
rect 19165 13821 19199 13855
rect 19257 13821 19291 13855
rect 21189 13821 21223 13855
rect 21833 13821 21867 13855
rect 23397 13821 23431 13855
rect 13829 13753 13863 13787
rect 2329 13685 2363 13719
rect 10425 13685 10459 13719
rect 16681 13685 16715 13719
rect 18521 13685 18555 13719
rect 23213 13685 23247 13719
rect 24777 13685 24811 13719
rect 26341 13685 26375 13719
rect 2237 13481 2271 13515
rect 8309 13481 8343 13515
rect 10995 13481 11029 13515
rect 11437 13481 11471 13515
rect 17141 13481 17175 13515
rect 19901 13481 19935 13515
rect 20913 13481 20947 13515
rect 21649 13481 21683 13515
rect 22385 13481 22419 13515
rect 23857 13481 23891 13515
rect 24133 13481 24167 13515
rect 24961 13481 24995 13515
rect 9505 13413 9539 13447
rect 12725 13413 12759 13447
rect 15577 13413 15611 13447
rect 17325 13413 17359 13447
rect 25329 13413 25363 13447
rect 2697 13345 2731 13379
rect 2881 13345 2915 13379
rect 6929 13345 6963 13379
rect 11253 13345 11287 13379
rect 15209 13345 15243 13379
rect 17693 13345 17727 13379
rect 22569 13345 22603 13379
rect 5365 13277 5399 13311
rect 5632 13277 5666 13311
rect 7196 13277 7230 13311
rect 11616 13277 11650 13311
rect 11989 13277 12023 13311
rect 12173 13277 12207 13311
rect 12449 13277 12483 13311
rect 12593 13277 12627 13311
rect 14841 13277 14875 13311
rect 15006 13274 15040 13308
rect 15117 13277 15151 13311
rect 15393 13277 15427 13311
rect 15853 13277 15887 13311
rect 17509 13277 17543 13311
rect 17785 13277 17819 13311
rect 17878 13277 17912 13311
rect 18061 13277 18095 13311
rect 21097 13277 21131 13311
rect 21517 13277 21551 13311
rect 21833 13277 21867 13311
rect 22017 13277 22051 13311
rect 22206 13277 22240 13311
rect 23305 13277 23339 13311
rect 23581 13277 23615 13311
rect 23725 13277 23759 13311
rect 24409 13277 24443 13311
rect 24782 13277 24816 13311
rect 11713 13209 11747 13243
rect 11805 13209 11839 13243
rect 12357 13209 12391 13243
rect 18337 13209 18371 13243
rect 20821 13209 20855 13243
rect 21281 13209 21315 13243
rect 21373 13209 21407 13243
rect 22109 13209 22143 13243
rect 23489 13209 23523 13243
rect 24593 13209 24627 13243
rect 24685 13209 24719 13243
rect 25145 13209 25179 13243
rect 2605 13141 2639 13175
rect 6745 13141 6779 13175
rect 13001 13141 13035 13175
rect 14657 13141 14691 13175
rect 15669 13141 15703 13175
rect 18245 13141 18279 13175
rect 22753 13141 22787 13175
rect 23213 13141 23247 13175
rect 3985 12937 4019 12971
rect 8677 12937 8711 12971
rect 12541 12937 12575 12971
rect 14381 12937 14415 12971
rect 17601 12937 17635 12971
rect 18061 12937 18095 12971
rect 18613 12937 18647 12971
rect 20269 12937 20303 12971
rect 22293 12937 22327 12971
rect 22845 12937 22879 12971
rect 2697 12869 2731 12903
rect 6745 12869 6779 12903
rect 6929 12869 6963 12903
rect 10609 12869 10643 12903
rect 10793 12869 10827 12903
rect 20177 12869 20211 12903
rect 22109 12869 22143 12903
rect 23765 12869 23799 12903
rect 24133 12869 24167 12903
rect 24225 12869 24259 12903
rect 4077 12801 4111 12835
rect 6653 12801 6687 12835
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 7573 12801 7607 12835
rect 7699 12801 7733 12835
rect 10425 12801 10459 12835
rect 11800 12801 11834 12835
rect 11897 12801 11931 12835
rect 11989 12801 12023 12835
rect 12173 12801 12207 12835
rect 12265 12801 12299 12835
rect 12633 12801 12667 12835
rect 14749 12801 14783 12835
rect 17969 12801 18003 12835
rect 19726 12801 19760 12835
rect 20729 12801 20763 12835
rect 22017 12801 22051 12835
rect 22661 12801 22695 12835
rect 23949 12801 23983 12835
rect 24369 12801 24403 12835
rect 24869 12801 24903 12835
rect 3893 12733 3927 12767
rect 10149 12733 10183 12767
rect 12909 12733 12943 12767
rect 18245 12733 18279 12767
rect 19993 12733 20027 12767
rect 2421 12665 2455 12699
rect 7941 12665 7975 12699
rect 11621 12665 11655 12699
rect 24685 12665 24719 12699
rect 2237 12597 2271 12631
rect 4445 12597 4479 12631
rect 6561 12597 6595 12631
rect 14565 12597 14599 12631
rect 20545 12597 20579 12631
rect 21833 12597 21867 12631
rect 24501 12597 24535 12631
rect 2789 12393 2823 12427
rect 5273 12393 5307 12427
rect 8677 12393 8711 12427
rect 9505 12393 9539 12427
rect 12817 12393 12851 12427
rect 14105 12393 14139 12427
rect 18429 12393 18463 12427
rect 21465 12393 21499 12427
rect 3433 12325 3467 12359
rect 11253 12325 11287 12359
rect 12449 12325 12483 12359
rect 1409 12257 1443 12291
rect 3065 12257 3099 12291
rect 14657 12257 14691 12291
rect 15117 12257 15151 12291
rect 18153 12257 18187 12291
rect 19441 12257 19475 12291
rect 24593 12257 24627 12291
rect 3893 12189 3927 12223
rect 5457 12189 5491 12223
rect 6193 12189 6227 12223
rect 6377 12189 6411 12223
rect 7297 12189 7331 12223
rect 7564 12189 7598 12223
rect 9229 12189 9263 12223
rect 9689 12189 9723 12223
rect 11069 12189 11103 12223
rect 11437 12189 11471 12223
rect 11897 12189 11931 12223
rect 12270 12189 12304 12223
rect 12633 12189 12667 12223
rect 14289 12189 14323 12223
rect 14841 12189 14875 12223
rect 15006 12189 15040 12223
rect 15209 12189 15243 12223
rect 15393 12189 15427 12223
rect 15669 12189 15703 12223
rect 17785 12189 17819 12223
rect 17968 12189 18002 12223
rect 18061 12189 18095 12223
rect 18310 12189 18344 12223
rect 22845 12189 22879 12223
rect 23121 12189 23155 12223
rect 23305 12189 23339 12223
rect 23581 12189 23615 12223
rect 23857 12189 23891 12223
rect 24001 12189 24035 12223
rect 1676 12121 1710 12155
rect 4160 12121 4194 12155
rect 12081 12121 12115 12155
rect 12173 12121 12207 12155
rect 13001 12121 13035 12155
rect 15577 12121 15611 12155
rect 15914 12121 15948 12155
rect 19717 12121 19751 12155
rect 22578 12121 22612 12155
rect 23765 12121 23799 12155
rect 24150 12121 24184 12155
rect 24838 12121 24872 12155
rect 3525 12053 3559 12087
rect 5549 12053 5583 12087
rect 6009 12053 6043 12087
rect 6377 12053 6411 12087
rect 9413 12053 9447 12087
rect 11621 12053 11655 12087
rect 13185 12053 13219 12087
rect 17049 12053 17083 12087
rect 17601 12053 17635 12087
rect 21189 12053 21223 12087
rect 22937 12053 22971 12087
rect 23489 12053 23523 12087
rect 24501 12053 24535 12087
rect 25973 12053 26007 12087
rect 1961 11849 1995 11883
rect 2329 11849 2363 11883
rect 2789 11849 2823 11883
rect 3985 11849 4019 11883
rect 9321 11849 9355 11883
rect 17417 11849 17451 11883
rect 19441 11849 19475 11883
rect 21557 11849 21591 11883
rect 4997 11781 5031 11815
rect 8861 11781 8895 11815
rect 9045 11781 9079 11815
rect 19809 11781 19843 11815
rect 22109 11781 22143 11815
rect 24746 11781 24780 11815
rect 2421 11713 2455 11747
rect 2973 11713 3007 11747
rect 3801 11713 3835 11747
rect 4517 11713 4551 11747
rect 4629 11713 4663 11747
rect 4905 11713 4939 11747
rect 5641 11713 5675 11747
rect 6633 11713 6667 11747
rect 10057 11713 10091 11747
rect 10425 11713 10459 11747
rect 10972 11713 11006 11747
rect 11069 11713 11103 11747
rect 11161 11713 11195 11747
rect 11345 11713 11379 11747
rect 12173 11713 12207 11747
rect 12357 11713 12391 11747
rect 12449 11713 12483 11747
rect 12593 11713 12627 11747
rect 12909 11713 12943 11747
rect 15117 11713 15151 11747
rect 15300 11713 15334 11747
rect 15393 11713 15427 11747
rect 15669 11713 15703 11747
rect 17785 11713 17819 11747
rect 21833 11713 21867 11747
rect 22017 11713 22051 11747
rect 22206 11713 22240 11747
rect 22569 11713 22603 11747
rect 22836 11713 22870 11747
rect 24501 11713 24535 11747
rect 2605 11645 2639 11679
rect 6377 11645 6411 11679
rect 11621 11645 11655 11679
rect 13185 11645 13219 11679
rect 14933 11645 14967 11679
rect 15485 11645 15519 11679
rect 17877 11645 17911 11679
rect 17969 11645 18003 11679
rect 19901 11645 19935 11679
rect 19993 11645 20027 11679
rect 4353 11577 4387 11611
rect 10241 11577 10275 11611
rect 12725 11577 12759 11611
rect 22385 11577 22419 11611
rect 5549 11509 5583 11543
rect 7757 11509 7791 11543
rect 10609 11509 10643 11543
rect 10793 11509 10827 11543
rect 14657 11509 14691 11543
rect 15761 11509 15795 11543
rect 18337 11509 18371 11543
rect 21373 11509 21407 11543
rect 23949 11509 23983 11543
rect 25881 11509 25915 11543
rect 2605 11305 2639 11339
rect 4997 11305 5031 11339
rect 6745 11305 6779 11339
rect 7113 11305 7147 11339
rect 10044 11305 10078 11339
rect 12173 11305 12207 11339
rect 13921 11305 13955 11339
rect 17141 11305 17175 11339
rect 20637 11305 20671 11339
rect 7481 11237 7515 11271
rect 9137 11237 9171 11271
rect 9505 11237 9539 11271
rect 13185 11237 13219 11271
rect 14105 11237 14139 11271
rect 9781 11169 9815 11203
rect 11529 11169 11563 11203
rect 15209 11169 15243 11203
rect 15301 11169 15335 11203
rect 15761 11169 15795 11203
rect 17601 11169 17635 11203
rect 18429 11169 18463 11203
rect 18521 11169 18555 11203
rect 19257 11169 19291 11203
rect 2237 11101 2271 11135
rect 3801 11101 3835 11135
rect 3985 11101 4019 11135
rect 5181 11101 5215 11135
rect 5549 11101 5583 11135
rect 5733 11101 5767 11135
rect 6745 11101 6779 11135
rect 6837 11101 6871 11135
rect 7297 11101 7331 11135
rect 8953 11101 8987 11135
rect 9413 11101 9447 11135
rect 9689 11101 9723 11135
rect 12357 11101 12391 11135
rect 13737 11101 13771 11135
rect 14289 11101 14323 11135
rect 14933 11101 14967 11135
rect 15098 11101 15132 11135
rect 15485 11101 15519 11135
rect 17325 11101 17359 11135
rect 17473 11101 17507 11135
rect 17693 11101 17727 11135
rect 17877 11101 17911 11135
rect 18153 11101 18187 11135
rect 18336 11101 18370 11135
rect 18705 11101 18739 11135
rect 2053 11033 2087 11067
rect 2421 11033 2455 11067
rect 14749 11033 14783 11067
rect 16006 11033 16040 11067
rect 18889 11033 18923 11067
rect 19502 11033 19536 11067
rect 4077 10965 4111 10999
rect 5733 10965 5767 10999
rect 9229 10965 9263 10999
rect 13001 10965 13035 10999
rect 15577 10965 15611 10999
rect 17969 10965 18003 10999
rect 1593 10761 1627 10795
rect 2145 10761 2179 10795
rect 2513 10761 2547 10795
rect 2881 10761 2915 10795
rect 5549 10761 5583 10795
rect 12265 10761 12299 10795
rect 16405 10761 16439 10795
rect 18797 10761 18831 10795
rect 22661 10761 22695 10795
rect 2053 10693 2087 10727
rect 5641 10693 5675 10727
rect 6469 10693 6503 10727
rect 9965 10693 9999 10727
rect 17684 10693 17718 10727
rect 1409 10625 1443 10659
rect 2697 10625 2731 10659
rect 3994 10625 4028 10659
rect 4629 10625 4663 10659
rect 4905 10625 4939 10659
rect 6377 10625 6411 10659
rect 7573 10625 7607 10659
rect 9729 10625 9763 10659
rect 9873 10625 9907 10659
rect 10149 10625 10183 10659
rect 10425 10625 10459 10659
rect 12357 10625 12391 10659
rect 12633 10625 12667 10659
rect 12909 10625 12943 10659
rect 13645 10625 13679 10659
rect 15025 10625 15059 10659
rect 15292 10625 15326 10659
rect 20177 10625 20211 10659
rect 20444 10625 20478 10659
rect 21925 10625 21959 10659
rect 22109 10625 22143 10659
rect 22247 10625 22281 10659
rect 22569 10625 22603 10659
rect 22937 10625 22971 10659
rect 23121 10625 23155 10659
rect 23397 10625 23431 10659
rect 23581 10625 23615 10659
rect 23949 10625 23983 10659
rect 24961 10625 24995 10659
rect 25053 10625 25087 10659
rect 2237 10557 2271 10591
rect 4261 10557 4295 10591
rect 4537 10557 4571 10591
rect 5457 10557 5491 10591
rect 7849 10557 7883 10591
rect 17417 10557 17451 10591
rect 22385 10557 22419 10591
rect 22477 10557 22511 10591
rect 23213 10557 23247 10591
rect 24685 10557 24719 10591
rect 9597 10489 9631 10523
rect 21557 10489 21591 10523
rect 23857 10489 23891 10523
rect 1685 10421 1719 10455
rect 6009 10421 6043 10455
rect 6193 10421 6227 10455
rect 9321 10421 9355 10455
rect 10241 10421 10275 10455
rect 10609 10421 10643 10455
rect 12449 10421 12483 10455
rect 12725 10421 12759 10455
rect 13461 10421 13495 10455
rect 17141 10421 17175 10455
rect 24777 10421 24811 10455
rect 25237 10421 25271 10455
rect 2329 10217 2363 10251
rect 3801 10217 3835 10251
rect 14197 10217 14231 10251
rect 14933 10217 14967 10251
rect 15301 10217 15335 10251
rect 19349 10217 19383 10251
rect 22293 10217 22327 10251
rect 22845 10217 22879 10251
rect 24133 10217 24167 10251
rect 24777 10217 24811 10251
rect 24593 10149 24627 10183
rect 4261 10081 4295 10115
rect 4445 10081 4479 10115
rect 5825 10081 5859 10115
rect 13921 10081 13955 10115
rect 14473 10081 14507 10115
rect 14657 10081 14691 10115
rect 14749 10081 14783 10115
rect 25053 10081 25087 10115
rect 2421 10013 2455 10047
rect 3065 10013 3099 10047
rect 9137 10013 9171 10047
rect 14381 10013 14415 10047
rect 14933 10013 14967 10047
rect 15117 10013 15151 10047
rect 21925 10013 21959 10047
rect 22201 10013 22235 10047
rect 23024 10013 23058 10047
rect 23213 10013 23247 10047
rect 23397 10013 23431 10047
rect 23673 10013 23707 10047
rect 24041 10013 24075 10047
rect 2605 9945 2639 9979
rect 6070 9945 6104 9979
rect 11529 9945 11563 9979
rect 13645 9945 13679 9979
rect 14841 9945 14875 9979
rect 23121 9945 23155 9979
rect 23489 9945 23523 9979
rect 23857 9945 23891 9979
rect 24961 9945 24995 9979
rect 25298 9945 25332 9979
rect 3157 9877 3191 9911
rect 4169 9877 4203 9911
rect 4721 9877 4755 9911
rect 7205 9877 7239 9911
rect 8953 9877 8987 9911
rect 12173 9877 12207 9911
rect 22109 9877 22143 9911
rect 24777 9877 24811 9911
rect 26433 9877 26467 9911
rect 2789 9673 2823 9707
rect 4169 9673 4203 9707
rect 6469 9673 6503 9707
rect 6653 9673 6687 9707
rect 11713 9673 11747 9707
rect 13461 9673 13495 9707
rect 14013 9673 14047 9707
rect 15025 9673 15059 9707
rect 16129 9673 16163 9707
rect 19165 9673 19199 9707
rect 23581 9673 23615 9707
rect 25513 9673 25547 9707
rect 1676 9605 1710 9639
rect 3065 9605 3099 9639
rect 10149 9605 10183 9639
rect 15209 9605 15243 9639
rect 15761 9605 15795 9639
rect 19441 9605 19475 9639
rect 20177 9605 20211 9639
rect 21833 9605 21867 9639
rect 3249 9537 3283 9571
rect 3341 9537 3375 9571
rect 3617 9537 3651 9571
rect 3709 9537 3743 9571
rect 3985 9537 4019 9571
rect 4721 9537 4755 9571
rect 4813 9537 4847 9571
rect 5181 9537 5215 9571
rect 5273 9537 5307 9571
rect 5549 9537 5583 9571
rect 6651 9537 6685 9571
rect 7113 9537 7147 9571
rect 7389 9537 7423 9571
rect 10005 9537 10039 9571
rect 10241 9537 10275 9571
rect 10425 9537 10459 9571
rect 10701 9537 10735 9571
rect 10885 9537 10919 9571
rect 10977 9537 11011 9571
rect 11121 9537 11155 9571
rect 11529 9537 11563 9571
rect 11989 9537 12023 9571
rect 12081 9537 12115 9571
rect 12265 9537 12299 9571
rect 12357 9537 12391 9571
rect 12495 9537 12529 9571
rect 13645 9537 13679 9571
rect 14841 9537 14875 9571
rect 15117 9537 15151 9571
rect 15393 9537 15427 9571
rect 15853 9537 15887 9571
rect 15945 9537 15979 9571
rect 17776 9537 17810 9571
rect 20085 9537 20119 9571
rect 20913 9537 20947 9571
rect 21005 9537 21039 9571
rect 21557 9537 21591 9571
rect 23121 9537 23155 9571
rect 23397 9537 23431 9571
rect 23489 9537 23523 9571
rect 24593 9537 24627 9571
rect 24777 9537 24811 9571
rect 25053 9537 25087 9571
rect 25329 9537 25363 9571
rect 25605 9537 25639 9571
rect 1409 9469 1443 9503
rect 3525 9469 3559 9503
rect 3801 9469 3835 9503
rect 4997 9469 5031 9503
rect 9413 9469 9447 9503
rect 9689 9469 9723 9503
rect 12909 9469 12943 9503
rect 15577 9469 15611 9503
rect 17509 9469 17543 9503
rect 20269 9469 20303 9503
rect 21097 9469 21131 9503
rect 23305 9469 23339 9503
rect 24961 9469 24995 9503
rect 7021 9401 7055 9435
rect 9873 9401 9907 9435
rect 10609 9401 10643 9435
rect 12633 9401 12667 9435
rect 19257 9401 19291 9435
rect 21373 9401 21407 9435
rect 22937 9401 22971 9435
rect 3709 9333 3743 9367
rect 4353 9333 4387 9367
rect 5733 9333 5767 9367
rect 7205 9333 7239 9367
rect 7941 9333 7975 9367
rect 11253 9333 11287 9367
rect 11805 9333 11839 9367
rect 14657 9333 14691 9367
rect 18889 9333 18923 9367
rect 19717 9333 19751 9367
rect 20545 9333 20579 9367
rect 23121 9333 23155 9367
rect 3893 9129 3927 9163
rect 4997 9129 5031 9163
rect 6285 9129 6319 9163
rect 9137 9129 9171 9163
rect 13093 9129 13127 9163
rect 15025 9129 15059 9163
rect 15209 9129 15243 9163
rect 18245 9129 18279 9163
rect 22293 9129 22327 9163
rect 20453 9061 20487 9095
rect 22753 9061 22787 9095
rect 24225 9061 24259 9095
rect 6653 8993 6687 9027
rect 11713 8993 11747 9027
rect 18061 8993 18095 9027
rect 18797 8993 18831 9027
rect 19901 8993 19935 9027
rect 21005 8993 21039 9027
rect 23121 8993 23155 9027
rect 23765 8993 23799 9027
rect 3157 8925 3191 8959
rect 3341 8925 3375 8959
rect 3985 8925 4019 8959
rect 5089 8925 5123 8959
rect 6469 8925 6503 8959
rect 8217 8925 8251 8959
rect 8953 8925 8987 8959
rect 11989 8925 12023 8959
rect 13737 8925 13771 8959
rect 17233 8925 17267 8959
rect 19349 8925 19383 8959
rect 19809 8925 19843 8959
rect 20177 8925 20211 8959
rect 20361 8925 20395 8959
rect 20821 8925 20855 8959
rect 21373 8925 21407 8959
rect 21649 8925 21683 8959
rect 21741 8925 21775 8959
rect 22017 8925 22051 8959
rect 22201 8925 22235 8959
rect 22661 8925 22695 8959
rect 22845 8925 22879 8959
rect 22937 8925 22971 8959
rect 23305 8925 23339 8959
rect 23581 8925 23615 8959
rect 23857 8925 23891 8959
rect 24041 8925 24075 8959
rect 3525 8857 3559 8891
rect 7950 8857 7984 8891
rect 12909 8857 12943 8891
rect 16988 8857 17022 8891
rect 17785 8857 17819 8891
rect 19441 8857 19475 8891
rect 22385 8857 22419 8891
rect 25881 8925 25915 8959
rect 25614 8857 25648 8891
rect 6837 8789 6871 8823
rect 10241 8789 10275 8823
rect 13921 8789 13955 8823
rect 15853 8789 15887 8823
rect 17417 8789 17451 8823
rect 17877 8789 17911 8823
rect 18613 8789 18647 8823
rect 18705 8789 18739 8823
rect 20913 8789 20947 8823
rect 24225 8789 24259 8823
rect 24501 8789 24535 8823
rect 5273 8585 5307 8619
rect 6101 8585 6135 8619
rect 7113 8585 7147 8619
rect 7573 8585 7607 8619
rect 11529 8585 11563 8619
rect 15025 8585 15059 8619
rect 16681 8585 16715 8619
rect 19165 8585 19199 8619
rect 19349 8585 19383 8619
rect 24041 8585 24075 8619
rect 7205 8517 7239 8551
rect 9229 8517 9263 8551
rect 12357 8517 12391 8551
rect 15209 8517 15243 8551
rect 17601 8517 17635 8551
rect 17785 8517 17819 8551
rect 2329 8449 2363 8483
rect 5273 8449 5307 8483
rect 5733 8449 5767 8483
rect 5825 8449 5859 8483
rect 6561 8449 6595 8483
rect 8769 8449 8803 8483
rect 9684 8449 9718 8483
rect 9781 8449 9815 8483
rect 9873 8449 9907 8483
rect 10057 8449 10091 8483
rect 10373 8449 10407 8483
rect 10517 8449 10551 8483
rect 10609 8449 10643 8483
rect 10793 8449 10827 8483
rect 10885 8449 10919 8483
rect 11161 8449 11195 8483
rect 12081 8449 12115 8483
rect 12265 8449 12299 8483
rect 12501 8449 12535 8483
rect 12817 8449 12851 8483
rect 15301 8449 15335 8483
rect 15485 8449 15519 8483
rect 15945 8449 15979 8483
rect 16221 8449 16255 8483
rect 17049 8449 17083 8483
rect 17969 8449 18003 8483
rect 18429 8449 18463 8483
rect 18797 8449 18831 8483
rect 19533 8449 19567 8483
rect 19625 8449 19659 8483
rect 19901 8449 19935 8483
rect 21189 8449 21223 8483
rect 21281 8449 21315 8483
rect 21465 8449 21499 8483
rect 21833 8449 21867 8483
rect 22017 8449 22051 8483
rect 22201 8449 22235 8483
rect 22293 8449 22327 8483
rect 24133 8449 24167 8483
rect 25329 8449 25363 8483
rect 5089 8381 5123 8415
rect 5641 8381 5675 8415
rect 6745 8381 6779 8415
rect 7021 8381 7055 8415
rect 13093 8381 13127 8415
rect 14565 8381 14599 8415
rect 16037 8381 16071 8415
rect 17141 8381 17175 8415
rect 17325 8381 17359 8415
rect 18521 8381 18555 8415
rect 18705 8381 18739 8415
rect 19809 8381 19843 8415
rect 9045 8313 9079 8347
rect 11069 8313 11103 8347
rect 11345 8313 11379 8347
rect 15669 8313 15703 8347
rect 16405 8313 16439 8347
rect 18613 8313 18647 8347
rect 21649 8381 21683 8415
rect 22477 8313 22511 8347
rect 25421 8313 25455 8347
rect 2145 8245 2179 8279
rect 5733 8245 5767 8279
rect 6469 8245 6503 8279
rect 8953 8245 8987 8279
rect 9505 8245 9539 8279
rect 10241 8245 10275 8279
rect 11805 8245 11839 8279
rect 12633 8245 12667 8279
rect 14841 8245 14875 8279
rect 15025 8245 15059 8279
rect 15853 8245 15887 8279
rect 21189 8245 21223 8279
rect 6377 8041 6411 8075
rect 9413 8041 9447 8075
rect 12817 8041 12851 8075
rect 13737 8041 13771 8075
rect 15025 8041 15059 8075
rect 16681 8041 16715 8075
rect 17141 8041 17175 8075
rect 21373 8041 21407 8075
rect 21741 8041 21775 8075
rect 5733 7973 5767 8007
rect 13185 7973 13219 8007
rect 13921 7973 13955 8007
rect 16129 7973 16163 8007
rect 17785 7973 17819 8007
rect 24409 7973 24443 8007
rect 7389 7905 7423 7939
rect 10057 7905 10091 7939
rect 14197 7905 14231 7939
rect 15577 7905 15611 7939
rect 16773 7905 16807 7939
rect 23029 7905 23063 7939
rect 24961 7905 24995 7939
rect 1501 7837 1535 7871
rect 3893 7837 3927 7871
rect 5457 7837 5491 7871
rect 5641 7837 5675 7871
rect 6101 7837 6135 7871
rect 6285 7837 6319 7871
rect 7941 7837 7975 7871
rect 9137 7837 9171 7871
rect 12265 7837 12299 7871
rect 12541 7837 12575 7871
rect 12638 7837 12672 7871
rect 13001 7837 13035 7871
rect 13277 7837 13311 7871
rect 13553 7837 13587 7871
rect 14933 7837 14967 7871
rect 15209 7837 15243 7871
rect 15945 7837 15979 7871
rect 16221 7837 16255 7871
rect 16957 7837 16991 7871
rect 17509 7837 17543 7871
rect 17969 7837 18003 7871
rect 20637 7837 20671 7871
rect 21189 7837 21223 7871
rect 21649 7837 21683 7871
rect 23213 7837 23247 7871
rect 24869 7837 24903 7871
rect 1768 7769 1802 7803
rect 4160 7769 4194 7803
rect 6469 7769 6503 7803
rect 7573 7769 7607 7803
rect 10333 7769 10367 7803
rect 12449 7769 12483 7803
rect 15393 7769 15427 7803
rect 16681 7769 16715 7803
rect 20821 7769 20855 7803
rect 2881 7701 2915 7735
rect 5273 7701 5307 7735
rect 7757 7701 7791 7735
rect 8953 7701 8987 7735
rect 11805 7701 11839 7735
rect 13461 7701 13495 7735
rect 14749 7701 14783 7735
rect 16405 7701 16439 7735
rect 17601 7701 17635 7735
rect 23397 7701 23431 7735
rect 24777 7701 24811 7735
rect 1777 7497 1811 7531
rect 2237 7497 2271 7531
rect 3801 7497 3835 7531
rect 6837 7497 6871 7531
rect 7297 7497 7331 7531
rect 19073 7497 19107 7531
rect 24777 7497 24811 7531
rect 4261 7429 4295 7463
rect 4905 7429 4939 7463
rect 10977 7429 11011 7463
rect 12541 7429 12575 7463
rect 17509 7429 17543 7463
rect 17693 7429 17727 7463
rect 21925 7429 21959 7463
rect 2145 7361 2179 7395
rect 2789 7361 2823 7395
rect 2973 7361 3007 7395
rect 3215 7361 3249 7395
rect 3525 7361 3559 7395
rect 3985 7361 4019 7395
rect 4353 7361 4387 7395
rect 5089 7361 5123 7395
rect 6009 7361 6043 7395
rect 6561 7361 6595 7395
rect 6653 7361 6687 7395
rect 7389 7361 7423 7395
rect 17233 7361 17267 7395
rect 17325 7361 17359 7395
rect 18061 7361 18095 7395
rect 18245 7361 18279 7395
rect 18429 7361 18463 7395
rect 18705 7361 18739 7395
rect 18889 7361 18923 7395
rect 19349 7361 19383 7395
rect 19441 7361 19475 7395
rect 19533 7361 19567 7395
rect 19993 7361 20027 7395
rect 20361 7361 20395 7395
rect 21005 7361 21039 7395
rect 21097 7361 21131 7395
rect 22293 7361 22327 7395
rect 23213 7361 23247 7395
rect 23397 7361 23431 7395
rect 23673 7361 23707 7395
rect 23857 7361 23891 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 24501 7361 24535 7395
rect 24593 7361 24627 7395
rect 25789 7361 25823 7395
rect 2329 7293 2363 7327
rect 3617 7293 3651 7327
rect 4077 7293 4111 7327
rect 4445 7293 4479 7327
rect 7113 7293 7147 7327
rect 9597 7293 9631 7327
rect 9873 7293 9907 7327
rect 12265 7293 12299 7327
rect 20085 7293 20119 7327
rect 20269 7293 20303 7327
rect 21281 7293 21315 7327
rect 22477 7293 22511 7327
rect 23489 7293 23523 7327
rect 2605 7225 2639 7259
rect 6193 7225 6227 7259
rect 17877 7225 17911 7259
rect 19625 7225 19659 7259
rect 20637 7225 20671 7259
rect 22201 7225 22235 7259
rect 4169 7157 4203 7191
rect 4353 7157 4387 7191
rect 4721 7157 4755 7191
rect 5181 7157 5215 7191
rect 7757 7157 7791 7191
rect 8125 7157 8159 7191
rect 11069 7157 11103 7191
rect 14013 7157 14047 7191
rect 17693 7157 17727 7191
rect 18705 7157 18739 7191
rect 25973 7157 26007 7191
rect 2697 6953 2731 6987
rect 5641 6953 5675 6987
rect 15669 6953 15703 6987
rect 18613 6953 18647 6987
rect 19533 6953 19567 6987
rect 20269 6953 20303 6987
rect 25789 6953 25823 6987
rect 19349 6885 19383 6919
rect 23213 6885 23247 6919
rect 2145 6817 2179 6851
rect 4445 6817 4479 6851
rect 12541 6817 12575 6851
rect 12725 6817 12759 6851
rect 15025 6817 15059 6851
rect 17785 6817 17819 6851
rect 19625 6817 19659 6851
rect 20729 6817 20763 6851
rect 20913 6817 20947 6851
rect 21373 6817 21407 6851
rect 21741 6817 21775 6851
rect 22477 6817 22511 6851
rect 24961 6817 24995 6851
rect 2329 6749 2363 6783
rect 2513 6749 2547 6783
rect 4043 6749 4077 6783
rect 4353 6749 4387 6783
rect 4721 6749 4755 6783
rect 4905 6749 4939 6783
rect 5089 6749 5123 6783
rect 5734 6749 5768 6783
rect 6101 6749 6135 6783
rect 6193 6749 6227 6783
rect 6929 6749 6963 6783
rect 8226 6749 8260 6783
rect 8493 6749 8527 6783
rect 9505 6749 9539 6783
rect 9597 6749 9631 6783
rect 11989 6749 12023 6783
rect 17049 6749 17083 6783
rect 17509 6749 17543 6783
rect 18797 6749 18831 6783
rect 19717 6749 19751 6783
rect 21557 6749 21591 6783
rect 21925 6749 21959 6783
rect 22385 6749 22419 6783
rect 22753 6749 22787 6783
rect 22845 6749 22879 6783
rect 23213 6749 23247 6783
rect 24685 6749 24719 6783
rect 24869 6749 24903 6783
rect 25145 6749 25179 6783
rect 25329 6749 25363 6783
rect 25973 6749 26007 6783
rect 9321 6681 9355 6715
rect 11744 6681 11778 6715
rect 16804 6681 16838 6715
rect 22017 6681 22051 6715
rect 25513 6681 25547 6715
rect 25697 6681 25731 6715
rect 26218 6681 26252 6715
rect 3893 6613 3927 6647
rect 7113 6613 7147 6647
rect 9137 6613 9171 6647
rect 10609 6613 10643 6647
rect 12081 6613 12115 6647
rect 12449 6613 12483 6647
rect 14473 6613 14507 6647
rect 14841 6613 14875 6647
rect 14933 6613 14967 6647
rect 17141 6613 17175 6647
rect 17601 6613 17635 6647
rect 20177 6613 20211 6647
rect 20637 6613 20671 6647
rect 27353 6613 27387 6647
rect 2881 6409 2915 6443
rect 5549 6409 5583 6443
rect 11989 6409 12023 6443
rect 12265 6409 12299 6443
rect 15853 6409 15887 6443
rect 18889 6409 18923 6443
rect 22477 6409 22511 6443
rect 22569 6409 22603 6443
rect 22937 6409 22971 6443
rect 24777 6409 24811 6443
rect 25145 6409 25179 6443
rect 25513 6409 25547 6443
rect 25881 6409 25915 6443
rect 6009 6341 6043 6375
rect 14464 6341 14498 6375
rect 18061 6341 18095 6375
rect 20637 6341 20671 6375
rect 21005 6341 21039 6375
rect 1768 6273 1802 6307
rect 3249 6273 3283 6307
rect 4353 6273 4387 6307
rect 4812 6273 4846 6307
rect 5733 6273 5767 6307
rect 6377 6273 6411 6307
rect 8861 6273 8895 6307
rect 9137 6273 9171 6307
rect 9404 6273 9438 6307
rect 11805 6273 11839 6307
rect 11989 6273 12023 6307
rect 12173 6273 12207 6307
rect 12900 6273 12934 6307
rect 14197 6273 14231 6307
rect 15853 6273 15887 6307
rect 16037 6273 16071 6307
rect 17969 6273 18003 6307
rect 18521 6273 18555 6307
rect 18613 6273 18647 6307
rect 19901 6273 19935 6307
rect 20821 6273 20855 6307
rect 23305 6273 23339 6307
rect 25421 6273 25455 6307
rect 1501 6205 1535 6239
rect 4445 6205 4479 6239
rect 5825 6205 5859 6239
rect 6469 6205 6503 6239
rect 12633 6205 12667 6239
rect 17877 6205 17911 6239
rect 22661 6205 22695 6239
rect 23397 6205 23431 6239
rect 23489 6205 23523 6239
rect 24501 6205 24535 6239
rect 24685 6205 24719 6239
rect 25329 6205 25363 6239
rect 25973 6205 26007 6239
rect 26065 6205 26099 6239
rect 6745 6137 6779 6171
rect 18429 6137 18463 6171
rect 3065 6069 3099 6103
rect 4905 6069 4939 6103
rect 5733 6069 5767 6103
rect 6377 6069 6411 6103
rect 9045 6069 9079 6103
rect 10517 6069 10551 6103
rect 14013 6069 14047 6103
rect 15577 6069 15611 6103
rect 18705 6069 18739 6103
rect 19717 6069 19751 6103
rect 22109 6069 22143 6103
rect 2237 5865 2271 5899
rect 4905 5865 4939 5899
rect 9321 5865 9355 5899
rect 15393 5865 15427 5899
rect 18705 5865 18739 5899
rect 20637 5865 20671 5899
rect 20913 5865 20947 5899
rect 21097 5865 21131 5899
rect 21649 5865 21683 5899
rect 24133 5865 24167 5899
rect 24593 5865 24627 5899
rect 3617 5797 3651 5831
rect 7205 5797 7239 5831
rect 19625 5797 19659 5831
rect 22661 5797 22695 5831
rect 2881 5729 2915 5763
rect 3985 5729 4019 5763
rect 5365 5729 5399 5763
rect 9781 5729 9815 5763
rect 9873 5729 9907 5763
rect 15117 5729 15151 5763
rect 2605 5661 2639 5695
rect 3341 5661 3375 5695
rect 3525 5661 3559 5695
rect 3617 5661 3651 5695
rect 4169 5661 4203 5695
rect 5273 5661 5307 5695
rect 5457 5661 5491 5695
rect 5824 5661 5858 5695
rect 6101 5661 6135 5695
rect 6193 5661 6227 5695
rect 6503 5661 6537 5695
rect 6745 5661 6779 5695
rect 6837 5661 6871 5695
rect 8585 5661 8619 5695
rect 11253 5661 11287 5695
rect 11529 5661 11563 5695
rect 13001 5661 13035 5695
rect 13553 5661 13587 5695
rect 14657 5661 14691 5695
rect 14841 5661 14875 5695
rect 15209 5661 15243 5695
rect 15485 5661 15519 5695
rect 17601 5661 17635 5695
rect 17785 5661 17819 5695
rect 18521 5661 18555 5695
rect 18613 5661 18647 5695
rect 18705 5661 18739 5695
rect 19257 5661 19291 5695
rect 19533 5661 19567 5695
rect 19717 5661 19751 5695
rect 20085 5661 20119 5695
rect 20269 5661 20303 5695
rect 20361 5661 20395 5695
rect 20821 5661 20855 5695
rect 21281 5661 21315 5695
rect 21373 5661 21407 5695
rect 21833 5661 21867 5695
rect 22385 5661 22419 5695
rect 22661 5661 22695 5695
rect 23949 5661 23983 5695
rect 24133 5661 24167 5695
rect 24409 5661 24443 5695
rect 25329 5661 25363 5695
rect 4629 5593 4663 5627
rect 4813 5593 4847 5627
rect 6009 5593 6043 5627
rect 8318 5593 8352 5627
rect 11621 5593 11655 5627
rect 20545 5593 20579 5627
rect 25513 5593 25547 5627
rect 25697 5593 25731 5627
rect 2697 5525 2731 5559
rect 3157 5525 3191 5559
rect 3893 5525 3927 5559
rect 4353 5525 4387 5559
rect 5089 5525 5123 5559
rect 7021 5525 7055 5559
rect 9689 5525 9723 5559
rect 13185 5525 13219 5559
rect 13369 5525 13403 5559
rect 17693 5525 17727 5559
rect 18429 5525 18463 5559
rect 18981 5525 19015 5559
rect 21557 5525 21591 5559
rect 23765 5525 23799 5559
rect 2605 5321 2639 5355
rect 4261 5321 4295 5355
rect 4353 5321 4387 5355
rect 4721 5321 4755 5355
rect 7481 5321 7515 5355
rect 8033 5321 8067 5355
rect 11713 5321 11747 5355
rect 12817 5321 12851 5355
rect 13277 5321 13311 5355
rect 15301 5321 15335 5355
rect 17325 5321 17359 5355
rect 17969 5321 18003 5355
rect 19625 5321 19659 5355
rect 19993 5321 20027 5355
rect 20637 5321 20671 5355
rect 24041 5321 24075 5355
rect 25421 5321 25455 5355
rect 25881 5321 25915 5355
rect 26249 5321 26283 5355
rect 27537 5321 27571 5355
rect 5825 5253 5859 5287
rect 6009 5253 6043 5287
rect 6193 5253 6227 5287
rect 11253 5253 11287 5287
rect 12633 5253 12667 5287
rect 13829 5253 13863 5287
rect 16773 5253 16807 5287
rect 17877 5253 17911 5287
rect 18429 5253 18463 5287
rect 23121 5253 23155 5287
rect 24317 5253 24351 5287
rect 27905 5253 27939 5287
rect 2789 5185 2823 5219
rect 4905 5185 4939 5219
rect 6653 5185 6687 5219
rect 6837 5185 6871 5219
rect 7573 5185 7607 5219
rect 8217 5185 8251 5219
rect 9137 5185 9171 5219
rect 9689 5185 9723 5219
rect 10885 5185 10919 5219
rect 11069 5185 11103 5219
rect 11161 5185 11195 5219
rect 11713 5185 11747 5219
rect 12081 5185 12115 5219
rect 12173 5185 12207 5219
rect 12357 5185 12391 5219
rect 12725 5185 12759 5219
rect 13185 5185 13219 5219
rect 14071 5185 14105 5219
rect 14841 5185 14875 5219
rect 15025 5185 15059 5219
rect 15301 5185 15335 5219
rect 15485 5185 15519 5219
rect 17049 5185 17083 5219
rect 18337 5185 18371 5219
rect 20085 5185 20119 5219
rect 20821 5185 20855 5219
rect 21925 5185 21959 5219
rect 22109 5185 22143 5219
rect 22385 5185 22419 5219
rect 22569 5185 22603 5219
rect 23581 5185 23615 5219
rect 23765 5185 23799 5219
rect 23857 5185 23891 5219
rect 24409 5185 24443 5219
rect 24593 5185 24627 5219
rect 24777 5185 24811 5219
rect 25053 5185 25087 5219
rect 25237 5185 25271 5219
rect 25789 5185 25823 5219
rect 26433 5185 26467 5219
rect 27169 5185 27203 5219
rect 27425 5185 27459 5219
rect 27721 5185 27755 5219
rect 27813 5185 27847 5219
rect 4537 5117 4571 5151
rect 4997 5117 5031 5151
rect 7297 5117 7331 5151
rect 8769 5117 8803 5151
rect 9321 5117 9355 5151
rect 10701 5117 10735 5151
rect 11529 5117 11563 5151
rect 13461 5117 13495 5151
rect 14381 5117 14415 5151
rect 14473 5117 14507 5151
rect 16681 5117 16715 5151
rect 17161 5117 17195 5151
rect 18061 5117 18095 5151
rect 18981 5117 19015 5151
rect 19073 5117 19107 5151
rect 19349 5117 19383 5151
rect 19533 5117 19567 5151
rect 20177 5117 20211 5151
rect 22201 5117 22235 5151
rect 23213 5117 23247 5151
rect 23305 5117 23339 5151
rect 24869 5117 24903 5151
rect 25973 5117 26007 5151
rect 27629 5117 27663 5151
rect 7021 5049 7055 5083
rect 7941 5049 7975 5083
rect 9505 5049 9539 5083
rect 22753 5049 22787 5083
rect 3893 4981 3927 5015
rect 8953 4981 8987 5015
rect 17509 4981 17543 5015
rect 18981 4981 19015 5015
rect 20913 4981 20947 5015
rect 23581 4981 23615 5015
rect 26985 4981 27019 5015
rect 5181 4777 5215 4811
rect 10609 4777 10643 4811
rect 11253 4777 11287 4811
rect 12909 4777 12943 4811
rect 15393 4777 15427 4811
rect 15853 4777 15887 4811
rect 21833 4777 21867 4811
rect 22845 4777 22879 4811
rect 25605 4777 25639 4811
rect 26433 4777 26467 4811
rect 10333 4709 10367 4743
rect 14565 4709 14599 4743
rect 8953 4641 8987 4675
rect 11069 4641 11103 4675
rect 11345 4641 11379 4675
rect 12633 4641 12667 4675
rect 15209 4641 15243 4675
rect 19717 4641 19751 4675
rect 19809 4641 19843 4675
rect 21557 4641 21591 4675
rect 1869 4573 1903 4607
rect 3801 4573 3835 4607
rect 4057 4573 4091 4607
rect 6009 4573 6043 4607
rect 8585 4573 8619 4607
rect 10702 4573 10736 4607
rect 11161 4573 11195 4607
rect 11253 4573 11287 4607
rect 11529 4573 11563 4607
rect 13093 4573 13127 4607
rect 13277 4573 13311 4607
rect 13553 4573 13587 4607
rect 14197 4573 14231 4607
rect 15393 4573 15427 4607
rect 17233 4573 17267 4607
rect 17325 4573 17359 4607
rect 17509 4573 17543 4607
rect 17785 4573 17819 4607
rect 19625 4573 19659 4607
rect 21373 4573 21407 4607
rect 9198 4505 9232 4539
rect 12265 4505 12299 4539
rect 12449 4505 12483 4539
rect 14381 4505 14415 4539
rect 15117 4505 15151 4539
rect 16988 4505 17022 4539
rect 27353 4709 27387 4743
rect 22293 4641 22327 4675
rect 23397 4641 23431 4675
rect 23581 4641 23615 4675
rect 24501 4641 24535 4675
rect 26157 4641 26191 4675
rect 26893 4641 26927 4675
rect 26985 4641 27019 4675
rect 22109 4573 22143 4607
rect 22569 4573 22603 4607
rect 22661 4573 22695 4607
rect 23673 4573 23707 4607
rect 24685 4573 24719 4607
rect 26801 4573 26835 4607
rect 27261 4573 27295 4607
rect 27537 4573 27571 4607
rect 21925 4505 21959 4539
rect 24777 4505 24811 4539
rect 26065 4505 26099 4539
rect 27721 4505 27755 4539
rect 1409 4437 1443 4471
rect 6193 4437 6227 4471
rect 7021 4437 7055 4471
rect 8769 4437 8803 4471
rect 11713 4437 11747 4471
rect 13369 4437 13403 4471
rect 15577 4437 15611 4471
rect 17325 4437 17359 4471
rect 17693 4437 17727 4471
rect 19257 4437 19291 4471
rect 21005 4437 21039 4471
rect 21465 4437 21499 4471
rect 21833 4437 21867 4471
rect 22477 4437 22511 4471
rect 24041 4437 24075 4471
rect 25145 4437 25179 4471
rect 25973 4437 26007 4471
rect 6745 4233 6779 4267
rect 8953 4233 8987 4267
rect 9413 4233 9447 4267
rect 18705 4233 18739 4267
rect 20361 4233 20395 4267
rect 21557 4233 21591 4267
rect 23765 4233 23799 4267
rect 27261 4233 27295 4267
rect 9321 4165 9355 4199
rect 11253 4165 11287 4199
rect 13369 4165 13403 4199
rect 15301 4165 15335 4199
rect 17785 4165 17819 4199
rect 18429 4165 18463 4199
rect 18613 4165 18647 4199
rect 24860 4165 24894 4199
rect 26801 4165 26835 4199
rect 5926 4097 5960 4131
rect 6193 4097 6227 4131
rect 7481 4097 7515 4131
rect 7757 4097 7791 4131
rect 11069 4097 11103 4131
rect 12357 4097 12391 4131
rect 13553 4097 13587 4131
rect 13737 4097 13771 4131
rect 15485 4097 15519 4131
rect 16773 4097 16807 4131
rect 16957 4097 16991 4131
rect 17601 4097 17635 4131
rect 18889 4097 18923 4131
rect 19165 4097 19199 4131
rect 20729 4097 20763 4131
rect 21373 4097 21407 4131
rect 23857 4097 23891 4131
rect 26433 4097 26467 4131
rect 26617 4097 26651 4131
rect 26985 4097 27019 4131
rect 29561 4097 29595 4131
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 7665 4029 7699 4063
rect 9505 4029 9539 4063
rect 16681 4029 16715 4063
rect 17969 4029 18003 4063
rect 20821 4029 20855 4063
rect 20913 4029 20947 4063
rect 24593 4029 24627 4063
rect 18245 3961 18279 3995
rect 25973 3961 26007 3995
rect 4813 3893 4847 3927
rect 6377 3893 6411 3927
rect 7297 3893 7331 3927
rect 10977 3893 11011 3927
rect 12173 3893 12207 3927
rect 12725 3893 12759 3927
rect 15209 3893 15243 3927
rect 18981 3893 19015 3927
rect 6653 3689 6687 3723
rect 9505 3689 9539 3723
rect 13185 3689 13219 3723
rect 15577 3689 15611 3723
rect 15761 3689 15795 3723
rect 16129 3689 16163 3723
rect 17601 3689 17635 3723
rect 21281 3689 21315 3723
rect 22477 3689 22511 3723
rect 23213 3689 23247 3723
rect 26617 3689 26651 3723
rect 12909 3621 12943 3655
rect 20637 3621 20671 3655
rect 10057 3553 10091 3587
rect 11161 3553 11195 3587
rect 13737 3553 13771 3587
rect 16129 3553 16163 3587
rect 16313 3553 16347 3587
rect 16497 3553 16531 3587
rect 17141 3553 17175 3587
rect 18245 3553 18279 3587
rect 18429 3553 18463 3587
rect 21445 3553 21479 3587
rect 23765 3553 23799 3587
rect 6469 3485 6503 3519
rect 9873 3485 9907 3519
rect 10333 3485 10367 3519
rect 10517 3485 10551 3519
rect 10759 3485 10793 3519
rect 11069 3485 11103 3519
rect 11529 3485 11563 3519
rect 13278 3485 13312 3519
rect 13645 3485 13679 3519
rect 14289 3485 14323 3519
rect 14991 3485 15025 3519
rect 15301 3485 15335 3519
rect 15393 3485 15427 3519
rect 15761 3485 15795 3519
rect 15853 3485 15887 3519
rect 9689 3417 9723 3451
rect 11796 3417 11830 3451
rect 14749 3417 14783 3451
rect 16037 3417 16071 3451
rect 17049 3485 17083 3519
rect 17325 3485 17359 3519
rect 17417 3485 17451 3519
rect 17969 3485 18003 3519
rect 18521 3485 18555 3519
rect 19257 3485 19291 3519
rect 21557 3485 21591 3519
rect 21833 3485 21867 3519
rect 22017 3485 22051 3519
rect 22293 3485 22327 3519
rect 24041 3485 24075 3519
rect 26525 3485 26559 3519
rect 16589 3417 16623 3451
rect 17877 3417 17911 3451
rect 19524 3417 19558 3451
rect 21925 3417 21959 3451
rect 24133 3417 24167 3451
rect 10149 3349 10183 3383
rect 14105 3349 14139 3383
rect 16129 3349 16163 3383
rect 16957 3349 16991 3383
rect 18889 3349 18923 3383
rect 22109 3349 22143 3383
rect 23581 3349 23615 3383
rect 23673 3349 23707 3383
rect 10701 3145 10735 3179
rect 11713 3145 11747 3179
rect 12081 3145 12115 3179
rect 12541 3145 12575 3179
rect 13185 3145 13219 3179
rect 13645 3145 13679 3179
rect 15117 3145 15151 3179
rect 18337 3145 18371 3179
rect 21281 3145 21315 3179
rect 23581 3145 23615 3179
rect 25421 3145 25455 3179
rect 25881 3145 25915 3179
rect 26433 3145 26467 3179
rect 13982 3077 14016 3111
rect 15577 3077 15611 3111
rect 15761 3077 15795 3111
rect 15945 3077 15979 3111
rect 16948 3077 16982 3111
rect 19450 3077 19484 3111
rect 9045 3009 9079 3043
rect 9321 3009 9355 3043
rect 9588 3009 9622 3043
rect 12173 3009 12207 3043
rect 12725 3009 12759 3043
rect 13277 3009 13311 3043
rect 13737 3009 13771 3043
rect 16681 3009 16715 3043
rect 19717 3009 19751 3043
rect 19901 3009 19935 3043
rect 20168 3009 20202 3043
rect 21925 3009 21959 3043
rect 22192 3009 22226 3043
rect 23673 3009 23707 3043
rect 23857 3009 23891 3043
rect 24124 3009 24158 3043
rect 25789 3009 25823 3043
rect 26433 3009 26467 3043
rect 26801 3009 26835 3043
rect 2973 2941 3007 2975
rect 7849 2941 7883 2975
rect 12265 2941 12299 2975
rect 13001 2941 13035 2975
rect 25973 2941 26007 2975
rect 26249 2941 26283 2975
rect 18061 2873 18095 2907
rect 23305 2873 23339 2907
rect 9229 2805 9263 2839
rect 25237 2805 25271 2839
rect 9597 2601 9631 2635
rect 12081 2601 12115 2635
rect 13369 2601 13403 2635
rect 13829 2601 13863 2635
rect 17509 2601 17543 2635
rect 25697 2601 25731 2635
rect 26157 2601 26191 2635
rect 23673 2533 23707 2567
rect 10057 2465 10091 2499
rect 10149 2465 10183 2499
rect 11621 2465 11655 2499
rect 11713 2465 11747 2499
rect 13461 2465 13495 2499
rect 9965 2397 9999 2431
rect 11897 2397 11931 2431
rect 13645 2397 13679 2431
rect 14473 2397 14507 2431
rect 17601 2397 17635 2431
rect 21833 2397 21867 2431
rect 22017 2397 22051 2431
rect 23489 2397 23523 2431
rect 23765 2397 23799 2431
rect 24041 2397 24075 2431
rect 25605 2397 25639 2431
rect 26065 2397 26099 2431
rect 22201 2329 22235 2363
rect 23857 2329 23891 2363
rect 24225 2329 24259 2363
rect 25881 2329 25915 2363
rect 14289 2261 14323 2295
rect 23305 2261 23339 2295
<< metal1 >>
rect 4062 30540 4068 30592
rect 4120 30580 4126 30592
rect 19610 30580 19616 30592
rect 4120 30552 19616 30580
rect 4120 30540 4126 30552
rect 19610 30540 19616 30552
rect 19668 30540 19674 30592
rect 1104 30490 29440 30512
rect 1104 30438 10395 30490
rect 10447 30438 10459 30490
rect 10511 30438 10523 30490
rect 10575 30438 10587 30490
rect 10639 30438 10651 30490
rect 10703 30438 19840 30490
rect 19892 30438 19904 30490
rect 19956 30438 19968 30490
rect 20020 30438 20032 30490
rect 20084 30438 20096 30490
rect 20148 30438 29440 30490
rect 1104 30416 29440 30438
rect 3970 30336 3976 30388
rect 4028 30376 4034 30388
rect 22186 30376 22192 30388
rect 4028 30348 22192 30376
rect 4028 30336 4034 30348
rect 22186 30336 22192 30348
rect 22244 30336 22250 30388
rect 20165 30311 20223 30317
rect 20165 30308 20177 30311
rect 19904 30280 20177 30308
rect 11146 30200 11152 30252
rect 11204 30240 11210 30252
rect 11793 30243 11851 30249
rect 11793 30240 11805 30243
rect 11204 30212 11805 30240
rect 11204 30200 11210 30212
rect 11793 30209 11805 30212
rect 11839 30209 11851 30243
rect 12345 30243 12403 30249
rect 12345 30240 12357 30243
rect 11793 30203 11851 30209
rect 11992 30212 12357 30240
rect 11992 30113 12020 30212
rect 12345 30209 12357 30212
rect 12391 30209 12403 30243
rect 14918 30240 14924 30252
rect 14879 30212 14924 30240
rect 12345 30203 12403 30209
rect 14918 30200 14924 30212
rect 14976 30200 14982 30252
rect 18598 30200 18604 30252
rect 18656 30240 18662 30252
rect 19429 30243 19487 30249
rect 19429 30240 19441 30243
rect 18656 30212 19441 30240
rect 18656 30200 18662 30212
rect 19429 30209 19441 30212
rect 19475 30209 19487 30243
rect 19429 30203 19487 30209
rect 19815 30243 19873 30249
rect 19815 30209 19827 30243
rect 19861 30240 19873 30243
rect 19904 30240 19932 30280
rect 20165 30277 20177 30280
rect 20211 30308 20223 30311
rect 26234 30308 26240 30320
rect 20211 30280 26240 30308
rect 20211 30277 20223 30280
rect 20165 30271 20223 30277
rect 26234 30268 26240 30280
rect 26292 30268 26298 30320
rect 19861 30212 19932 30240
rect 19981 30243 20039 30249
rect 19861 30209 19873 30212
rect 19815 30203 19873 30209
rect 19981 30209 19993 30243
rect 20027 30240 20039 30243
rect 20346 30240 20352 30252
rect 20027 30212 20352 30240
rect 20027 30209 20039 30212
rect 19981 30203 20039 30209
rect 20346 30200 20352 30212
rect 20404 30200 20410 30252
rect 20714 30240 20720 30252
rect 20675 30212 20720 30240
rect 20714 30200 20720 30212
rect 20772 30200 20778 30252
rect 22002 30200 22008 30252
rect 22060 30249 22066 30252
rect 22060 30243 22103 30249
rect 22091 30209 22103 30243
rect 22060 30203 22103 30209
rect 22189 30243 22247 30249
rect 22189 30209 22201 30243
rect 22235 30209 22247 30243
rect 22189 30203 22247 30209
rect 22281 30243 22339 30249
rect 22281 30209 22293 30243
rect 22327 30209 22339 30243
rect 22462 30240 22468 30252
rect 22423 30212 22468 30240
rect 22281 30203 22339 30209
rect 22060 30200 22066 30203
rect 18690 30132 18696 30184
rect 18748 30172 18754 30184
rect 19613 30175 19671 30181
rect 19613 30172 19625 30175
rect 18748 30144 19625 30172
rect 18748 30132 18754 30144
rect 19613 30141 19625 30144
rect 19659 30141 19671 30175
rect 19613 30135 19671 30141
rect 19705 30175 19763 30181
rect 19705 30141 19717 30175
rect 19751 30141 19763 30175
rect 21545 30175 21603 30181
rect 21545 30172 21557 30175
rect 19705 30135 19763 30141
rect 20364 30144 21557 30172
rect 11977 30107 12035 30113
rect 11977 30073 11989 30107
rect 12023 30073 12035 30107
rect 11977 30067 12035 30073
rect 19058 30064 19064 30116
rect 19116 30104 19122 30116
rect 19720 30104 19748 30135
rect 19116 30076 19748 30104
rect 19116 30064 19122 30076
rect 12161 30039 12219 30045
rect 12161 30005 12173 30039
rect 12207 30036 12219 30039
rect 12250 30036 12256 30048
rect 12207 30008 12256 30036
rect 12207 30005 12219 30008
rect 12161 29999 12219 30005
rect 12250 29996 12256 30008
rect 12308 29996 12314 30048
rect 14642 29996 14648 30048
rect 14700 30036 14706 30048
rect 14737 30039 14795 30045
rect 14737 30036 14749 30039
rect 14700 30008 14749 30036
rect 14700 29996 14706 30008
rect 14737 30005 14749 30008
rect 14783 30005 14795 30039
rect 19334 30036 19340 30048
rect 19295 30008 19340 30036
rect 14737 29999 14795 30005
rect 19334 29996 19340 30008
rect 19392 29996 19398 30048
rect 19610 29996 19616 30048
rect 19668 30036 19674 30048
rect 20364 30036 20392 30144
rect 21545 30141 21557 30144
rect 21591 30172 21603 30175
rect 21726 30172 21732 30184
rect 21591 30144 21732 30172
rect 21591 30141 21603 30144
rect 21545 30135 21603 30141
rect 21726 30132 21732 30144
rect 21784 30132 21790 30184
rect 21082 30064 21088 30116
rect 21140 30104 21146 30116
rect 21913 30107 21971 30113
rect 21913 30104 21925 30107
rect 21140 30076 21925 30104
rect 21140 30064 21146 30076
rect 21913 30073 21925 30076
rect 21959 30073 21971 30107
rect 21913 30067 21971 30073
rect 20530 30036 20536 30048
rect 19668 30008 20392 30036
rect 20491 30008 20536 30036
rect 19668 29996 19674 30008
rect 20530 29996 20536 30008
rect 20588 29996 20594 30048
rect 21726 29996 21732 30048
rect 21784 30036 21790 30048
rect 22204 30036 22232 30203
rect 22296 30172 22324 30203
rect 22462 30200 22468 30212
rect 22520 30200 22526 30252
rect 22830 30240 22836 30252
rect 22791 30212 22836 30240
rect 22830 30200 22836 30212
rect 22888 30200 22894 30252
rect 22296 30144 22692 30172
rect 22664 30048 22692 30144
rect 22646 30036 22652 30048
rect 21784 30008 22232 30036
rect 22607 30008 22652 30036
rect 21784 29996 21790 30008
rect 22646 29996 22652 30008
rect 22704 29996 22710 30048
rect 23017 30039 23075 30045
rect 23017 30005 23029 30039
rect 23063 30036 23075 30039
rect 23106 30036 23112 30048
rect 23063 30008 23112 30036
rect 23063 30005 23075 30008
rect 23017 29999 23075 30005
rect 23106 29996 23112 30008
rect 23164 29996 23170 30048
rect 1104 29946 29440 29968
rect 1104 29894 5672 29946
rect 5724 29894 5736 29946
rect 5788 29894 5800 29946
rect 5852 29894 5864 29946
rect 5916 29894 5928 29946
rect 5980 29894 15118 29946
rect 15170 29894 15182 29946
rect 15234 29894 15246 29946
rect 15298 29894 15310 29946
rect 15362 29894 15374 29946
rect 15426 29894 24563 29946
rect 24615 29894 24627 29946
rect 24679 29894 24691 29946
rect 24743 29894 24755 29946
rect 24807 29894 24819 29946
rect 24871 29894 29440 29946
rect 1104 29872 29440 29894
rect 4062 29792 4068 29844
rect 4120 29832 4126 29844
rect 17034 29832 17040 29844
rect 4120 29804 17040 29832
rect 4120 29792 4126 29804
rect 17034 29792 17040 29804
rect 17092 29792 17098 29844
rect 19337 29835 19395 29841
rect 19337 29801 19349 29835
rect 19383 29832 19395 29835
rect 26142 29832 26148 29844
rect 19383 29804 26148 29832
rect 19383 29801 19395 29804
rect 19337 29795 19395 29801
rect 18690 29764 18696 29776
rect 18616 29736 18696 29764
rect 3234 29656 3240 29708
rect 3292 29696 3298 29708
rect 3329 29699 3387 29705
rect 3329 29696 3341 29699
rect 3292 29668 3341 29696
rect 3292 29656 3298 29668
rect 3329 29665 3341 29668
rect 3375 29665 3387 29699
rect 4614 29696 4620 29708
rect 4575 29668 4620 29696
rect 3329 29659 3387 29665
rect 4614 29656 4620 29668
rect 4672 29656 4678 29708
rect 7098 29656 7104 29708
rect 7156 29696 7162 29708
rect 7653 29699 7711 29705
rect 7653 29696 7665 29699
rect 7156 29668 7665 29696
rect 7156 29656 7162 29668
rect 7653 29665 7665 29668
rect 7699 29665 7711 29699
rect 7653 29659 7711 29665
rect 12526 29656 12532 29708
rect 12584 29696 12590 29708
rect 14185 29699 14243 29705
rect 14185 29696 14197 29699
rect 12584 29668 14197 29696
rect 12584 29656 12590 29668
rect 14185 29665 14197 29668
rect 14231 29665 14243 29699
rect 14185 29659 14243 29665
rect 15654 29656 15660 29708
rect 15712 29696 15718 29708
rect 15933 29699 15991 29705
rect 15933 29696 15945 29699
rect 15712 29668 15945 29696
rect 15712 29656 15718 29668
rect 15933 29665 15945 29668
rect 15979 29696 15991 29699
rect 16669 29699 16727 29705
rect 16669 29696 16681 29699
rect 15979 29668 16681 29696
rect 15979 29665 15991 29668
rect 15933 29659 15991 29665
rect 16669 29665 16681 29668
rect 16715 29665 16727 29699
rect 16669 29659 16727 29665
rect 17954 29656 17960 29708
rect 18012 29696 18018 29708
rect 18616 29705 18644 29736
rect 18690 29724 18696 29736
rect 18748 29724 18754 29776
rect 18601 29699 18659 29705
rect 18012 29668 18552 29696
rect 18012 29656 18018 29668
rect 5166 29588 5172 29640
rect 5224 29628 5230 29640
rect 5537 29631 5595 29637
rect 5537 29628 5549 29631
rect 5224 29600 5549 29628
rect 5224 29588 5230 29600
rect 5537 29597 5549 29600
rect 5583 29628 5595 29631
rect 9033 29631 9091 29637
rect 9033 29628 9045 29631
rect 5583 29600 9045 29628
rect 5583 29597 5595 29600
rect 5537 29591 5595 29597
rect 9033 29597 9045 29600
rect 9079 29597 9091 29631
rect 11146 29628 11152 29640
rect 11107 29600 11152 29628
rect 9033 29591 9091 29597
rect 11146 29588 11152 29600
rect 11204 29588 11210 29640
rect 13265 29631 13323 29637
rect 13265 29597 13277 29631
rect 13311 29628 13323 29631
rect 13630 29628 13636 29640
rect 13311 29600 13636 29628
rect 13311 29597 13323 29600
rect 13265 29591 13323 29597
rect 13630 29588 13636 29600
rect 13688 29588 13694 29640
rect 18417 29631 18475 29637
rect 18417 29597 18429 29631
rect 18463 29597 18475 29631
rect 18524 29628 18552 29668
rect 18601 29665 18613 29699
rect 18647 29665 18659 29699
rect 19352 29696 19380 29795
rect 26142 29792 26148 29804
rect 26200 29792 26206 29844
rect 19610 29764 19616 29776
rect 19571 29736 19616 29764
rect 19610 29724 19616 29736
rect 19668 29724 19674 29776
rect 20346 29696 20352 29708
rect 18601 29659 18659 29665
rect 18892 29668 19380 29696
rect 19536 29668 20352 29696
rect 18693 29631 18751 29637
rect 18693 29628 18705 29631
rect 18524 29600 18705 29628
rect 18417 29591 18475 29597
rect 18693 29597 18705 29600
rect 18739 29597 18751 29631
rect 18693 29591 18751 29597
rect 18803 29631 18861 29637
rect 18803 29597 18815 29631
rect 18849 29628 18861 29631
rect 18892 29628 18920 29668
rect 18849 29600 18920 29628
rect 18849 29597 18861 29600
rect 18803 29591 18861 29597
rect 5626 29520 5632 29572
rect 5684 29560 5690 29572
rect 5782 29563 5840 29569
rect 5782 29560 5794 29563
rect 5684 29532 5794 29560
rect 5684 29520 5690 29532
rect 5782 29529 5794 29532
rect 5828 29529 5840 29563
rect 7561 29563 7619 29569
rect 7561 29560 7573 29563
rect 5782 29523 5840 29529
rect 6932 29532 7573 29560
rect 6932 29504 6960 29532
rect 7561 29529 7573 29532
rect 7607 29529 7619 29563
rect 9306 29560 9312 29572
rect 9267 29532 9312 29560
rect 7561 29523 7619 29529
rect 9306 29520 9312 29532
rect 9364 29520 9370 29572
rect 10318 29520 10324 29572
rect 10376 29520 10382 29572
rect 10612 29532 11560 29560
rect 6914 29492 6920 29504
rect 6875 29464 6920 29492
rect 6914 29452 6920 29464
rect 6972 29452 6978 29504
rect 7101 29495 7159 29501
rect 7101 29461 7113 29495
rect 7147 29492 7159 29495
rect 7374 29492 7380 29504
rect 7147 29464 7380 29492
rect 7147 29461 7159 29464
rect 7101 29455 7159 29461
rect 7374 29452 7380 29464
rect 7432 29452 7438 29504
rect 7469 29495 7527 29501
rect 7469 29461 7481 29495
rect 7515 29492 7527 29495
rect 10612 29492 10640 29532
rect 10778 29492 10784 29504
rect 7515 29464 10640 29492
rect 10739 29464 10784 29492
rect 7515 29461 7527 29464
rect 7469 29455 7527 29461
rect 10778 29452 10784 29464
rect 10836 29452 10842 29504
rect 10962 29492 10968 29504
rect 10923 29464 10968 29492
rect 10962 29452 10968 29464
rect 11020 29452 11026 29504
rect 11532 29501 11560 29532
rect 12250 29520 12256 29572
rect 12308 29520 12314 29572
rect 12986 29560 12992 29572
rect 12947 29532 12992 29560
rect 12986 29520 12992 29532
rect 13044 29520 13050 29572
rect 14642 29520 14648 29572
rect 14700 29520 14706 29572
rect 15378 29520 15384 29572
rect 15436 29560 15442 29572
rect 15657 29563 15715 29569
rect 15657 29560 15669 29563
rect 15436 29532 15669 29560
rect 15436 29520 15442 29532
rect 15657 29529 15669 29532
rect 15703 29529 15715 29563
rect 15657 29523 15715 29529
rect 16936 29563 16994 29569
rect 16936 29529 16948 29563
rect 16982 29560 16994 29563
rect 18233 29563 18291 29569
rect 18233 29560 18245 29563
rect 16982 29532 18245 29560
rect 16982 29529 16994 29532
rect 16936 29523 16994 29529
rect 18233 29529 18245 29532
rect 18279 29529 18291 29563
rect 18233 29523 18291 29529
rect 11517 29495 11575 29501
rect 11517 29461 11529 29495
rect 11563 29492 11575 29495
rect 11606 29492 11612 29504
rect 11563 29464 11612 29492
rect 11563 29461 11575 29464
rect 11517 29455 11575 29461
rect 11606 29452 11612 29464
rect 11664 29452 11670 29504
rect 14366 29452 14372 29504
rect 14424 29492 14430 29504
rect 15838 29492 15844 29504
rect 14424 29464 15844 29492
rect 14424 29452 14430 29464
rect 15838 29452 15844 29464
rect 15896 29452 15902 29504
rect 18049 29495 18107 29501
rect 18049 29461 18061 29495
rect 18095 29492 18107 29495
rect 18138 29492 18144 29504
rect 18095 29464 18144 29492
rect 18095 29461 18107 29464
rect 18049 29455 18107 29461
rect 18138 29452 18144 29464
rect 18196 29492 18202 29504
rect 18432 29492 18460 29591
rect 18708 29560 18736 29591
rect 18966 29588 18972 29640
rect 19024 29628 19030 29640
rect 19536 29628 19564 29668
rect 20346 29656 20352 29668
rect 20404 29656 20410 29708
rect 21082 29696 21088 29708
rect 21043 29668 21088 29696
rect 21082 29656 21088 29668
rect 21140 29656 21146 29708
rect 19024 29600 19564 29628
rect 21361 29631 21419 29637
rect 19024 29588 19030 29600
rect 21361 29597 21373 29631
rect 21407 29628 21419 29631
rect 21726 29628 21732 29640
rect 21407 29600 21732 29628
rect 21407 29597 21419 29600
rect 21361 29591 21419 29597
rect 21726 29588 21732 29600
rect 21784 29628 21790 29640
rect 21821 29631 21879 29637
rect 21821 29628 21833 29631
rect 21784 29600 21833 29628
rect 21784 29588 21790 29600
rect 21821 29597 21833 29600
rect 21867 29597 21879 29631
rect 21821 29591 21879 29597
rect 19058 29560 19064 29572
rect 18708 29532 19064 29560
rect 19058 29520 19064 29532
rect 19116 29520 19122 29572
rect 20530 29520 20536 29572
rect 20588 29520 20594 29572
rect 22094 29520 22100 29572
rect 22152 29560 22158 29572
rect 22152 29532 22197 29560
rect 22152 29520 22158 29532
rect 23106 29520 23112 29572
rect 23164 29520 23170 29572
rect 18196 29464 18460 29492
rect 18196 29452 18202 29464
rect 22922 29452 22928 29504
rect 22980 29492 22986 29504
rect 23569 29495 23627 29501
rect 23569 29492 23581 29495
rect 22980 29464 23581 29492
rect 22980 29452 22986 29464
rect 23569 29461 23581 29464
rect 23615 29461 23627 29495
rect 23569 29455 23627 29461
rect 1104 29402 29440 29424
rect 1104 29350 10395 29402
rect 10447 29350 10459 29402
rect 10511 29350 10523 29402
rect 10575 29350 10587 29402
rect 10639 29350 10651 29402
rect 10703 29350 19840 29402
rect 19892 29350 19904 29402
rect 19956 29350 19968 29402
rect 20020 29350 20032 29402
rect 20084 29350 20096 29402
rect 20148 29350 29440 29402
rect 1104 29328 29440 29350
rect 5626 29288 5632 29300
rect 5587 29260 5632 29288
rect 5626 29248 5632 29260
rect 5684 29248 5690 29300
rect 9306 29288 9312 29300
rect 9267 29260 9312 29288
rect 9306 29248 9312 29260
rect 9364 29248 9370 29300
rect 10318 29248 10324 29300
rect 10376 29288 10382 29300
rect 10505 29291 10563 29297
rect 10505 29288 10517 29291
rect 10376 29260 10517 29288
rect 10376 29248 10382 29260
rect 10505 29257 10517 29260
rect 10551 29257 10563 29291
rect 10505 29251 10563 29257
rect 12526 29248 12532 29300
rect 12584 29288 12590 29300
rect 13466 29291 13524 29297
rect 12584 29260 13124 29288
rect 12584 29248 12590 29260
rect 5166 29220 5172 29232
rect 3436 29192 5172 29220
rect 3436 29161 3464 29192
rect 5166 29180 5172 29192
rect 5224 29180 5230 29232
rect 6914 29220 6920 29232
rect 5828 29192 6920 29220
rect 3421 29155 3479 29161
rect 3421 29121 3433 29155
rect 3467 29121 3479 29155
rect 3421 29115 3479 29121
rect 3688 29155 3746 29161
rect 3688 29121 3700 29155
rect 3734 29152 3746 29155
rect 3970 29152 3976 29164
rect 3734 29124 3976 29152
rect 3734 29121 3746 29124
rect 3688 29115 3746 29121
rect 3970 29112 3976 29124
rect 4028 29112 4034 29164
rect 5828 29161 5856 29192
rect 6914 29180 6920 29192
rect 6972 29180 6978 29232
rect 7193 29223 7251 29229
rect 7193 29189 7205 29223
rect 7239 29220 7251 29223
rect 10137 29223 10195 29229
rect 10137 29220 10149 29223
rect 7239 29192 10149 29220
rect 7239 29189 7251 29192
rect 7193 29183 7251 29189
rect 10137 29189 10149 29192
rect 10183 29220 10195 29223
rect 10778 29220 10784 29232
rect 10183 29192 10784 29220
rect 10183 29189 10195 29192
rect 10137 29183 10195 29189
rect 10778 29180 10784 29192
rect 10836 29180 10842 29232
rect 12161 29223 12219 29229
rect 12161 29189 12173 29223
rect 12207 29220 12219 29223
rect 12986 29220 12992 29232
rect 12207 29192 12992 29220
rect 12207 29189 12219 29192
rect 12161 29183 12219 29189
rect 12986 29180 12992 29192
rect 13044 29180 13050 29232
rect 13096 29220 13124 29260
rect 13466 29257 13478 29291
rect 13512 29288 13524 29291
rect 15378 29288 15384 29300
rect 13512 29260 15384 29288
rect 13512 29257 13524 29260
rect 13466 29251 13524 29257
rect 15378 29248 15384 29260
rect 15436 29248 15442 29300
rect 15749 29291 15807 29297
rect 15749 29257 15761 29291
rect 15795 29257 15807 29291
rect 18598 29288 18604 29300
rect 18559 29260 18604 29288
rect 15749 29251 15807 29257
rect 13170 29223 13228 29229
rect 13170 29220 13182 29223
rect 13096 29192 13182 29220
rect 13170 29189 13182 29192
rect 13216 29189 13228 29223
rect 13170 29183 13228 29189
rect 13725 29223 13783 29229
rect 13725 29189 13737 29223
rect 13771 29220 13783 29223
rect 14366 29220 14372 29232
rect 13771 29192 14372 29220
rect 13771 29189 13783 29192
rect 13725 29183 13783 29189
rect 5813 29155 5871 29161
rect 5813 29121 5825 29155
rect 5859 29121 5871 29155
rect 5813 29115 5871 29121
rect 5902 29112 5908 29164
rect 5960 29152 5966 29164
rect 7285 29155 7343 29161
rect 7285 29152 7297 29155
rect 5960 29124 6005 29152
rect 6104 29124 7297 29152
rect 5960 29112 5966 29124
rect 6104 29084 6132 29124
rect 7285 29121 7297 29124
rect 7331 29121 7343 29155
rect 7285 29115 7343 29121
rect 9493 29155 9551 29161
rect 9493 29121 9505 29155
rect 9539 29152 9551 29155
rect 10689 29155 10747 29161
rect 9539 29124 9720 29152
rect 9539 29121 9551 29124
rect 9493 29115 9551 29121
rect 4816 29056 6132 29084
rect 6181 29087 6239 29093
rect 4816 29025 4844 29056
rect 6181 29053 6193 29087
rect 6227 29084 6239 29087
rect 6227 29056 6868 29084
rect 6227 29053 6239 29056
rect 6181 29047 6239 29053
rect 4801 29019 4859 29025
rect 4801 28985 4813 29019
rect 4847 28985 4859 29019
rect 4801 28979 4859 28985
rect 4154 28908 4160 28960
rect 4212 28948 4218 28960
rect 4816 28948 4844 28979
rect 6086 28976 6092 29028
rect 6144 29016 6150 29028
rect 6840 29025 6868 29056
rect 7098 29044 7104 29096
rect 7156 29084 7162 29096
rect 7377 29087 7435 29093
rect 7377 29084 7389 29087
rect 7156 29056 7389 29084
rect 7156 29044 7162 29056
rect 7377 29053 7389 29056
rect 7423 29053 7435 29087
rect 7377 29047 7435 29053
rect 9692 29025 9720 29124
rect 10689 29121 10701 29155
rect 10735 29152 10747 29155
rect 10962 29152 10968 29164
rect 10735 29124 10968 29152
rect 10735 29121 10747 29124
rect 10689 29115 10747 29121
rect 10962 29112 10968 29124
rect 11020 29112 11026 29164
rect 11149 29155 11207 29161
rect 11149 29121 11161 29155
rect 11195 29121 11207 29155
rect 11606 29152 11612 29164
rect 11567 29124 11612 29152
rect 11149 29115 11207 29121
rect 10134 29084 10140 29096
rect 10095 29056 10140 29084
rect 10134 29044 10140 29056
rect 10192 29044 10198 29096
rect 10229 29087 10287 29093
rect 10229 29053 10241 29087
rect 10275 29084 10287 29087
rect 10870 29084 10876 29096
rect 10275 29056 10876 29084
rect 10275 29053 10287 29056
rect 10229 29047 10287 29053
rect 10870 29044 10876 29056
rect 10928 29084 10934 29096
rect 11164 29084 11192 29115
rect 11606 29112 11612 29124
rect 11664 29112 11670 29164
rect 11793 29155 11851 29161
rect 11793 29121 11805 29155
rect 11839 29152 11851 29155
rect 12437 29155 12495 29161
rect 11839 29124 12204 29152
rect 11839 29121 11851 29124
rect 11793 29115 11851 29121
rect 10928 29056 11192 29084
rect 10928 29044 10934 29056
rect 6825 29019 6883 29025
rect 6144 28988 6189 29016
rect 6144 28976 6150 28988
rect 6825 28985 6837 29019
rect 6871 28985 6883 29019
rect 6825 28979 6883 28985
rect 9677 29019 9735 29025
rect 9677 28985 9689 29019
rect 9723 28985 9735 29019
rect 9677 28979 9735 28985
rect 11333 29019 11391 29025
rect 11333 28985 11345 29019
rect 11379 29016 11391 29019
rect 11808 29016 11836 29115
rect 12176 29096 12204 29124
rect 12437 29121 12449 29155
rect 12483 29152 12495 29155
rect 12526 29152 12532 29164
rect 12483 29124 12532 29152
rect 12483 29121 12495 29124
rect 12437 29115 12495 29121
rect 12526 29112 12532 29124
rect 12584 29112 12590 29164
rect 12894 29152 12900 29164
rect 12855 29124 12900 29152
rect 12894 29112 12900 29124
rect 12952 29112 12958 29164
rect 13081 29155 13139 29161
rect 13081 29121 13093 29155
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 12158 29044 12164 29096
rect 12216 29084 12222 29096
rect 12345 29087 12403 29093
rect 12345 29084 12357 29087
rect 12216 29056 12357 29084
rect 12216 29044 12222 29056
rect 12345 29053 12357 29056
rect 12391 29053 12403 29087
rect 13096 29084 13124 29115
rect 13262 29112 13268 29164
rect 13320 29161 13326 29164
rect 13320 29152 13328 29161
rect 13740 29152 13768 29183
rect 14366 29180 14372 29192
rect 14424 29180 14430 29232
rect 15764 29220 15792 29251
rect 18598 29248 18604 29260
rect 18656 29248 18662 29300
rect 20533 29291 20591 29297
rect 20533 29257 20545 29291
rect 20579 29288 20591 29291
rect 20714 29288 20720 29300
rect 20579 29260 20720 29288
rect 20579 29257 20591 29260
rect 20533 29251 20591 29257
rect 20714 29248 20720 29260
rect 20772 29248 20778 29300
rect 22830 29288 22836 29300
rect 22791 29260 22836 29288
rect 22830 29248 22836 29260
rect 22888 29248 22894 29300
rect 22186 29220 22192 29232
rect 15318 29192 15792 29220
rect 16684 29192 20024 29220
rect 22147 29192 22192 29220
rect 15930 29152 15936 29164
rect 13320 29124 13365 29152
rect 13464 29124 13768 29152
rect 15891 29124 15936 29152
rect 13320 29115 13328 29124
rect 13320 29112 13326 29115
rect 13464 29084 13492 29124
rect 15930 29112 15936 29124
rect 15988 29112 15994 29164
rect 13096 29056 13492 29084
rect 12345 29047 12403 29053
rect 13630 29044 13636 29096
rect 13688 29084 13694 29096
rect 13817 29087 13875 29093
rect 13817 29084 13829 29087
rect 13688 29056 13829 29084
rect 13688 29044 13694 29056
rect 13817 29053 13829 29056
rect 13863 29053 13875 29087
rect 13817 29047 13875 29053
rect 14090 29044 14096 29096
rect 14148 29084 14154 29096
rect 15565 29087 15623 29093
rect 15565 29084 15577 29087
rect 14148 29056 15577 29084
rect 14148 29044 14154 29056
rect 15565 29053 15577 29056
rect 15611 29053 15623 29087
rect 15565 29047 15623 29053
rect 15654 29044 15660 29096
rect 15712 29084 15718 29096
rect 16684 29093 16712 29192
rect 16936 29155 16994 29161
rect 16936 29121 16948 29155
rect 16982 29152 16994 29155
rect 17402 29152 17408 29164
rect 16982 29124 17408 29152
rect 16982 29121 16994 29124
rect 16936 29115 16994 29121
rect 17402 29112 17408 29124
rect 17460 29112 17466 29164
rect 19334 29112 19340 29164
rect 19392 29152 19398 29164
rect 19996 29161 20024 29192
rect 22186 29180 22192 29192
rect 22244 29220 22250 29232
rect 22922 29220 22928 29232
rect 22244 29192 22928 29220
rect 22244 29180 22250 29192
rect 22922 29180 22928 29192
rect 22980 29180 22986 29232
rect 19714 29155 19772 29161
rect 19714 29152 19726 29155
rect 19392 29124 19726 29152
rect 19392 29112 19398 29124
rect 19714 29121 19726 29124
rect 19760 29121 19772 29155
rect 19714 29115 19772 29121
rect 19981 29155 20039 29161
rect 19981 29121 19993 29155
rect 20027 29152 20039 29155
rect 20254 29152 20260 29164
rect 20027 29124 20260 29152
rect 20027 29121 20039 29124
rect 19981 29115 20039 29121
rect 20254 29112 20260 29124
rect 20312 29112 20318 29164
rect 20346 29112 20352 29164
rect 20404 29152 20410 29164
rect 20530 29152 20536 29164
rect 20404 29124 20536 29152
rect 20404 29112 20410 29124
rect 20530 29112 20536 29124
rect 20588 29112 20594 29164
rect 20714 29152 20720 29164
rect 20675 29124 20720 29152
rect 20714 29112 20720 29124
rect 20772 29112 20778 29164
rect 22002 29112 22008 29164
rect 22060 29161 22066 29164
rect 22060 29155 22103 29161
rect 22091 29152 22103 29155
rect 22281 29155 22339 29161
rect 22091 29124 22232 29152
rect 22091 29121 22103 29124
rect 22060 29115 22103 29121
rect 22060 29112 22066 29115
rect 22204 29096 22232 29124
rect 22281 29121 22293 29155
rect 22327 29121 22339 29155
rect 22281 29115 22339 29121
rect 22465 29155 22523 29161
rect 22465 29121 22477 29155
rect 22511 29152 22523 29155
rect 22554 29152 22560 29164
rect 22511 29124 22560 29152
rect 22511 29121 22523 29124
rect 22465 29115 22523 29121
rect 16669 29087 16727 29093
rect 16669 29084 16681 29087
rect 15712 29056 16681 29084
rect 15712 29044 15718 29056
rect 16669 29053 16681 29056
rect 16715 29053 16727 29087
rect 16669 29047 16727 29053
rect 22186 29044 22192 29096
rect 22244 29044 22250 29096
rect 11379 28988 11836 29016
rect 18049 29019 18107 29025
rect 11379 28985 11391 28988
rect 11333 28979 11391 28985
rect 18049 28985 18061 29019
rect 18095 29016 18107 29019
rect 18230 29016 18236 29028
rect 18095 28988 18236 29016
rect 18095 28985 18107 28988
rect 18049 28979 18107 28985
rect 18230 28976 18236 28988
rect 18288 28976 18294 29028
rect 21913 29019 21971 29025
rect 21913 28985 21925 29019
rect 21959 29016 21971 29019
rect 22094 29016 22100 29028
rect 21959 28988 22100 29016
rect 21959 28985 21971 28988
rect 21913 28979 21971 28985
rect 22094 28976 22100 28988
rect 22152 28976 22158 29028
rect 22296 29016 22324 29115
rect 22554 29112 22560 29124
rect 22612 29112 22618 29164
rect 22649 29155 22707 29161
rect 22649 29121 22661 29155
rect 22695 29152 22707 29155
rect 22738 29152 22744 29164
rect 22695 29124 22744 29152
rect 22695 29121 22707 29124
rect 22649 29115 22707 29121
rect 22738 29112 22744 29124
rect 22796 29152 22802 29164
rect 24394 29152 24400 29164
rect 22796 29124 24400 29152
rect 22796 29112 22802 29124
rect 24394 29112 24400 29124
rect 24452 29112 24458 29164
rect 23201 29019 23259 29025
rect 23201 29016 23213 29019
rect 22296 28988 23213 29016
rect 23201 28985 23213 28988
rect 23247 29016 23259 29019
rect 23842 29016 23848 29028
rect 23247 28988 23848 29016
rect 23247 28985 23259 28988
rect 23201 28979 23259 28985
rect 23842 28976 23848 28988
rect 23900 28976 23906 29028
rect 4212 28920 4844 28948
rect 4212 28908 4218 28920
rect 13722 28908 13728 28960
rect 13780 28948 13786 28960
rect 14074 28951 14132 28957
rect 14074 28948 14086 28951
rect 13780 28920 14086 28948
rect 13780 28908 13786 28920
rect 14074 28917 14086 28920
rect 14120 28917 14132 28951
rect 14074 28911 14132 28917
rect 19242 28908 19248 28960
rect 19300 28948 19306 28960
rect 20806 28948 20812 28960
rect 19300 28920 20812 28948
rect 19300 28908 19306 28920
rect 20806 28908 20812 28920
rect 20864 28908 20870 28960
rect 23934 28908 23940 28960
rect 23992 28948 23998 28960
rect 25866 28948 25872 28960
rect 23992 28920 25872 28948
rect 23992 28908 23998 28920
rect 25866 28908 25872 28920
rect 25924 28908 25930 28960
rect 1104 28858 29440 28880
rect 1104 28806 5672 28858
rect 5724 28806 5736 28858
rect 5788 28806 5800 28858
rect 5852 28806 5864 28858
rect 5916 28806 5928 28858
rect 5980 28806 15118 28858
rect 15170 28806 15182 28858
rect 15234 28806 15246 28858
rect 15298 28806 15310 28858
rect 15362 28806 15374 28858
rect 15426 28806 24563 28858
rect 24615 28806 24627 28858
rect 24679 28806 24691 28858
rect 24743 28806 24755 28858
rect 24807 28806 24819 28858
rect 24871 28806 29440 28858
rect 1104 28784 29440 28806
rect 3970 28744 3976 28756
rect 3931 28716 3976 28744
rect 3970 28704 3976 28716
rect 4028 28704 4034 28756
rect 4338 28704 4344 28756
rect 4396 28744 4402 28756
rect 4433 28747 4491 28753
rect 4433 28744 4445 28747
rect 4396 28716 4445 28744
rect 4396 28704 4402 28716
rect 4433 28713 4445 28716
rect 4479 28744 4491 28747
rect 6086 28744 6092 28756
rect 4479 28716 6092 28744
rect 4479 28713 4491 28716
rect 4433 28707 4491 28713
rect 6086 28704 6092 28716
rect 6144 28744 6150 28756
rect 7285 28747 7343 28753
rect 7285 28744 7297 28747
rect 6144 28716 7297 28744
rect 6144 28704 6150 28716
rect 7285 28713 7297 28716
rect 7331 28713 7343 28747
rect 13722 28744 13728 28756
rect 13683 28716 13728 28744
rect 7285 28707 7343 28713
rect 13722 28704 13728 28716
rect 13780 28704 13786 28756
rect 14829 28747 14887 28753
rect 14829 28713 14841 28747
rect 14875 28744 14887 28747
rect 14918 28744 14924 28756
rect 14875 28716 14924 28744
rect 14875 28713 14887 28716
rect 14829 28707 14887 28713
rect 14918 28704 14924 28716
rect 14976 28704 14982 28756
rect 15289 28747 15347 28753
rect 15289 28713 15301 28747
rect 15335 28744 15347 28747
rect 15930 28744 15936 28756
rect 15335 28716 15936 28744
rect 15335 28713 15347 28716
rect 15289 28707 15347 28713
rect 15930 28704 15936 28716
rect 15988 28704 15994 28756
rect 17034 28704 17040 28756
rect 17092 28744 17098 28756
rect 17221 28747 17279 28753
rect 17221 28744 17233 28747
rect 17092 28716 17233 28744
rect 17092 28704 17098 28716
rect 17221 28713 17233 28716
rect 17267 28744 17279 28747
rect 18046 28744 18052 28756
rect 17267 28716 18052 28744
rect 17267 28713 17279 28716
rect 17221 28707 17279 28713
rect 18046 28704 18052 28716
rect 18104 28704 18110 28756
rect 23753 28747 23811 28753
rect 23753 28713 23765 28747
rect 23799 28744 23811 28747
rect 25222 28744 25228 28756
rect 23799 28716 25228 28744
rect 23799 28713 23811 28716
rect 23753 28707 23811 28713
rect 25222 28704 25228 28716
rect 25280 28704 25286 28756
rect 6549 28679 6607 28685
rect 6549 28645 6561 28679
rect 6595 28645 6607 28679
rect 6549 28639 6607 28645
rect 5166 28608 5172 28620
rect 5127 28580 5172 28608
rect 5166 28568 5172 28580
rect 5224 28568 5230 28620
rect 4154 28540 4160 28552
rect 4115 28512 4160 28540
rect 4154 28500 4160 28512
rect 4212 28500 4218 28552
rect 4246 28500 4252 28552
rect 4304 28540 4310 28552
rect 4522 28540 4528 28552
rect 4304 28512 4349 28540
rect 4483 28512 4528 28540
rect 4304 28500 4310 28512
rect 4522 28500 4528 28512
rect 4580 28500 4586 28552
rect 6564 28540 6592 28639
rect 15470 28636 15476 28688
rect 15528 28676 15534 28688
rect 16206 28676 16212 28688
rect 15528 28648 16212 28676
rect 15528 28636 15534 28648
rect 16206 28636 16212 28648
rect 16264 28636 16270 28688
rect 17402 28676 17408 28688
rect 17363 28648 17408 28676
rect 17402 28636 17408 28648
rect 17460 28636 17466 28688
rect 22189 28679 22247 28685
rect 22189 28676 22201 28679
rect 22066 28648 22201 28676
rect 7374 28568 7380 28620
rect 7432 28608 7438 28620
rect 11146 28608 11152 28620
rect 7432 28580 7477 28608
rect 10888 28580 11152 28608
rect 7432 28568 7438 28580
rect 7006 28540 7012 28552
rect 6564 28512 7012 28540
rect 7006 28500 7012 28512
rect 7064 28500 7070 28552
rect 7101 28543 7159 28549
rect 7101 28509 7113 28543
rect 7147 28509 7159 28543
rect 8570 28540 8576 28552
rect 8531 28512 8576 28540
rect 7101 28503 7159 28509
rect 5436 28475 5494 28481
rect 5436 28441 5448 28475
rect 5482 28472 5494 28475
rect 6825 28475 6883 28481
rect 6825 28472 6837 28475
rect 5482 28444 6837 28472
rect 5482 28441 5494 28444
rect 5436 28435 5494 28441
rect 6825 28441 6837 28444
rect 6871 28441 6883 28475
rect 6825 28435 6883 28441
rect 5994 28364 6000 28416
rect 6052 28404 6058 28416
rect 7116 28404 7144 28503
rect 8570 28500 8576 28512
rect 8628 28500 8634 28552
rect 10226 28540 10232 28552
rect 10187 28512 10232 28540
rect 10226 28500 10232 28512
rect 10284 28500 10290 28552
rect 10888 28549 10916 28580
rect 11146 28568 11152 28580
rect 11204 28568 11210 28620
rect 11238 28568 11244 28620
rect 11296 28608 11302 28620
rect 11974 28608 11980 28620
rect 11296 28580 11980 28608
rect 11296 28568 11302 28580
rect 11974 28568 11980 28580
rect 12032 28568 12038 28620
rect 17773 28611 17831 28617
rect 17773 28577 17785 28611
rect 17819 28608 17831 28611
rect 18690 28608 18696 28620
rect 17819 28580 18696 28608
rect 17819 28577 17831 28580
rect 17773 28571 17831 28577
rect 18690 28568 18696 28580
rect 18748 28568 18754 28620
rect 21729 28611 21787 28617
rect 21729 28577 21741 28611
rect 21775 28608 21787 28611
rect 22066 28608 22094 28648
rect 22189 28645 22201 28648
rect 22235 28645 22247 28679
rect 29822 28676 29828 28688
rect 22189 28639 22247 28645
rect 22296 28648 29828 28676
rect 22296 28608 22324 28648
rect 29822 28636 29828 28648
rect 29880 28636 29886 28688
rect 21775 28580 22094 28608
rect 22204 28580 22324 28608
rect 21775 28577 21787 28580
rect 21729 28571 21787 28577
rect 10873 28543 10931 28549
rect 10873 28509 10885 28543
rect 10919 28509 10931 28543
rect 11333 28543 11391 28549
rect 11333 28540 11345 28543
rect 10873 28503 10931 28509
rect 11072 28512 11345 28540
rect 8386 28404 8392 28416
rect 6052 28376 7144 28404
rect 8347 28376 8392 28404
rect 6052 28364 6058 28376
rect 8386 28364 8392 28376
rect 8444 28364 8450 28416
rect 9766 28364 9772 28416
rect 9824 28404 9830 28416
rect 11072 28413 11100 28512
rect 11333 28509 11345 28512
rect 11379 28509 11391 28543
rect 11333 28503 11391 28509
rect 12894 28500 12900 28552
rect 12952 28540 12958 28552
rect 13173 28543 13231 28549
rect 13173 28540 13185 28543
rect 12952 28512 13185 28540
rect 12952 28500 12958 28512
rect 13173 28509 13185 28512
rect 13219 28509 13231 28543
rect 13173 28503 13231 28509
rect 13262 28500 13268 28552
rect 13320 28540 13326 28552
rect 13546 28543 13604 28549
rect 13546 28540 13558 28543
rect 13320 28512 13558 28540
rect 13320 28500 13326 28512
rect 13546 28509 13558 28512
rect 13592 28509 13604 28543
rect 13546 28503 13604 28509
rect 15013 28543 15071 28549
rect 15013 28509 15025 28543
rect 15059 28540 15071 28543
rect 15105 28543 15163 28549
rect 15105 28540 15117 28543
rect 15059 28512 15117 28540
rect 15059 28509 15071 28512
rect 15013 28503 15071 28509
rect 15105 28509 15117 28512
rect 15151 28540 15163 28543
rect 15470 28540 15476 28552
rect 15151 28512 15476 28540
rect 15151 28509 15163 28512
rect 15105 28503 15163 28509
rect 15470 28500 15476 28512
rect 15528 28540 15534 28552
rect 15749 28543 15807 28549
rect 15749 28540 15761 28543
rect 15528 28512 15761 28540
rect 15528 28500 15534 28512
rect 15749 28509 15761 28512
rect 15795 28509 15807 28543
rect 15749 28503 15807 28509
rect 17589 28543 17647 28549
rect 17589 28509 17601 28543
rect 17635 28509 17647 28543
rect 17862 28540 17868 28552
rect 17823 28512 17868 28540
rect 17589 28503 17647 28509
rect 13357 28475 13415 28481
rect 13357 28441 13369 28475
rect 13403 28441 13415 28475
rect 13357 28435 13415 28441
rect 13449 28475 13507 28481
rect 13449 28441 13461 28475
rect 13495 28472 13507 28475
rect 13906 28472 13912 28484
rect 13495 28444 13912 28472
rect 13495 28441 13507 28444
rect 13449 28435 13507 28441
rect 10045 28407 10103 28413
rect 10045 28404 10057 28407
rect 9824 28376 10057 28404
rect 9824 28364 9830 28376
rect 10045 28373 10057 28376
rect 10091 28373 10103 28407
rect 10045 28367 10103 28373
rect 11057 28407 11115 28413
rect 11057 28373 11069 28407
rect 11103 28373 11115 28407
rect 11057 28367 11115 28373
rect 11146 28364 11152 28416
rect 11204 28404 11210 28416
rect 13372 28404 13400 28435
rect 13906 28432 13912 28444
rect 13964 28432 13970 28484
rect 17604 28472 17632 28503
rect 17862 28500 17868 28512
rect 17920 28500 17926 28552
rect 17958 28543 18016 28549
rect 17958 28509 17970 28543
rect 18004 28540 18016 28543
rect 18046 28540 18052 28552
rect 18004 28512 18052 28540
rect 18004 28509 18016 28512
rect 17958 28503 18016 28509
rect 18046 28500 18052 28512
rect 18104 28500 18110 28552
rect 18141 28543 18199 28549
rect 18141 28509 18153 28543
rect 18187 28540 18199 28543
rect 18966 28540 18972 28552
rect 18187 28512 18972 28540
rect 18187 28509 18199 28512
rect 18141 28503 18199 28509
rect 18966 28500 18972 28512
rect 19024 28500 19030 28552
rect 22016 28543 22074 28549
rect 22016 28509 22028 28543
rect 22062 28540 22074 28543
rect 22062 28509 22094 28540
rect 22016 28503 22094 28509
rect 18230 28472 18236 28484
rect 17604 28444 18236 28472
rect 18230 28432 18236 28444
rect 18288 28432 18294 28484
rect 20714 28432 20720 28484
rect 20772 28432 20778 28484
rect 21726 28432 21732 28484
rect 21784 28472 21790 28484
rect 22066 28472 22094 28503
rect 21784 28444 22094 28472
rect 22204 28472 22232 28580
rect 22462 28568 22468 28620
rect 22520 28608 22526 28620
rect 22520 28580 22784 28608
rect 22520 28568 22526 28580
rect 22278 28500 22284 28552
rect 22336 28549 22342 28552
rect 22756 28549 22784 28580
rect 22336 28543 22379 28549
rect 22367 28509 22379 28543
rect 22336 28503 22379 28509
rect 22741 28543 22799 28549
rect 22741 28509 22753 28543
rect 22787 28540 22799 28543
rect 22833 28543 22891 28549
rect 22833 28540 22845 28543
rect 22787 28512 22845 28540
rect 22787 28509 22799 28512
rect 22741 28503 22799 28509
rect 22833 28509 22845 28512
rect 22879 28509 22891 28543
rect 22833 28503 22891 28509
rect 22336 28500 22342 28503
rect 23198 28500 23204 28552
rect 23256 28549 23262 28552
rect 23256 28540 23264 28549
rect 23256 28512 23301 28540
rect 23256 28503 23264 28512
rect 23256 28500 23262 28503
rect 23382 28500 23388 28552
rect 23440 28540 23446 28552
rect 23569 28543 23627 28549
rect 23569 28540 23581 28543
rect 23440 28512 23581 28540
rect 23440 28500 23446 28512
rect 23569 28509 23581 28512
rect 23615 28509 23627 28543
rect 24394 28540 24400 28552
rect 24355 28512 24400 28540
rect 23569 28503 23627 28509
rect 24394 28500 24400 28512
rect 24452 28500 24458 28552
rect 24857 28543 24915 28549
rect 24857 28540 24869 28543
rect 24596 28512 24869 28540
rect 22465 28475 22523 28481
rect 22465 28472 22477 28475
rect 22204 28444 22477 28472
rect 21784 28432 21790 28444
rect 13998 28404 14004 28416
rect 11204 28376 11249 28404
rect 13372 28376 14004 28404
rect 11204 28364 11210 28376
rect 13998 28364 14004 28376
rect 14056 28404 14062 28416
rect 14093 28407 14151 28413
rect 14093 28404 14105 28407
rect 14056 28376 14105 28404
rect 14056 28364 14062 28376
rect 14093 28373 14105 28376
rect 14139 28373 14151 28407
rect 15930 28404 15936 28416
rect 15891 28376 15936 28404
rect 14093 28367 14151 28373
rect 15930 28364 15936 28376
rect 15988 28364 15994 28416
rect 20257 28407 20315 28413
rect 20257 28373 20269 28407
rect 20303 28404 20315 28407
rect 22204 28404 22232 28444
rect 22465 28441 22477 28444
rect 22511 28441 22523 28475
rect 22465 28435 22523 28441
rect 22554 28432 22560 28484
rect 22612 28472 22618 28484
rect 22612 28444 22657 28472
rect 22612 28432 22618 28444
rect 22922 28432 22928 28484
rect 22980 28472 22986 28484
rect 23017 28475 23075 28481
rect 23017 28472 23029 28475
rect 22980 28444 23029 28472
rect 22980 28432 22986 28444
rect 23017 28441 23029 28444
rect 23063 28441 23075 28475
rect 23017 28435 23075 28441
rect 23109 28475 23167 28481
rect 23109 28441 23121 28475
rect 23155 28472 23167 28475
rect 23658 28472 23664 28484
rect 23155 28444 23664 28472
rect 23155 28441 23167 28444
rect 23109 28435 23167 28441
rect 23658 28432 23664 28444
rect 23716 28432 23722 28484
rect 20303 28376 22232 28404
rect 20303 28373 20315 28376
rect 20257 28367 20315 28373
rect 22278 28364 22284 28416
rect 22336 28404 22342 28416
rect 23198 28404 23204 28416
rect 22336 28376 23204 28404
rect 22336 28364 22342 28376
rect 23198 28364 23204 28376
rect 23256 28364 23262 28416
rect 23402 28407 23460 28413
rect 23402 28373 23414 28407
rect 23448 28404 23460 28407
rect 23566 28404 23572 28416
rect 23448 28376 23572 28404
rect 23448 28373 23460 28376
rect 23402 28367 23460 28373
rect 23566 28364 23572 28376
rect 23624 28364 23630 28416
rect 23937 28407 23995 28413
rect 23937 28373 23949 28407
rect 23983 28404 23995 28407
rect 24026 28404 24032 28416
rect 23983 28376 24032 28404
rect 23983 28373 23995 28376
rect 23937 28367 23995 28373
rect 24026 28364 24032 28376
rect 24084 28364 24090 28416
rect 24596 28413 24624 28512
rect 24857 28509 24869 28512
rect 24903 28509 24915 28543
rect 24857 28503 24915 28509
rect 24581 28407 24639 28413
rect 24581 28373 24593 28407
rect 24627 28373 24639 28407
rect 24581 28367 24639 28373
rect 24670 28364 24676 28416
rect 24728 28404 24734 28416
rect 24728 28376 24773 28404
rect 24728 28364 24734 28376
rect 1104 28314 29440 28336
rect 1104 28262 10395 28314
rect 10447 28262 10459 28314
rect 10511 28262 10523 28314
rect 10575 28262 10587 28314
rect 10639 28262 10651 28314
rect 10703 28262 19840 28314
rect 19892 28262 19904 28314
rect 19956 28262 19968 28314
rect 20020 28262 20032 28314
rect 20084 28262 20096 28314
rect 20148 28262 29440 28314
rect 1104 28240 29440 28262
rect 4433 28203 4491 28209
rect 4433 28169 4445 28203
rect 4479 28200 4491 28203
rect 4522 28200 4528 28212
rect 4479 28172 4528 28200
rect 4479 28169 4491 28172
rect 4433 28163 4491 28169
rect 4522 28160 4528 28172
rect 4580 28160 4586 28212
rect 7006 28200 7012 28212
rect 6967 28172 7012 28200
rect 7006 28160 7012 28172
rect 7064 28160 7070 28212
rect 10042 28200 10048 28212
rect 7760 28172 10048 28200
rect 4801 28135 4859 28141
rect 4801 28101 4813 28135
rect 4847 28132 4859 28135
rect 7760 28132 7788 28172
rect 10042 28160 10048 28172
rect 10100 28200 10106 28212
rect 11241 28203 11299 28209
rect 11241 28200 11253 28203
rect 10100 28172 11253 28200
rect 10100 28160 10106 28172
rect 11241 28169 11253 28172
rect 11287 28169 11299 28203
rect 11241 28163 11299 28169
rect 18049 28203 18107 28209
rect 18049 28169 18061 28203
rect 18095 28200 18107 28203
rect 18877 28203 18935 28209
rect 18877 28200 18889 28203
rect 18095 28172 18889 28200
rect 18095 28169 18107 28172
rect 18049 28163 18107 28169
rect 18877 28169 18889 28172
rect 18923 28200 18935 28203
rect 19242 28200 19248 28212
rect 18923 28172 19248 28200
rect 18923 28169 18935 28172
rect 18877 28163 18935 28169
rect 19242 28160 19248 28172
rect 19300 28160 19306 28212
rect 20714 28160 20720 28212
rect 20772 28200 20778 28212
rect 20809 28203 20867 28209
rect 20809 28200 20821 28203
rect 20772 28172 20821 28200
rect 20772 28160 20778 28172
rect 20809 28169 20821 28172
rect 20855 28169 20867 28203
rect 22462 28200 22468 28212
rect 22423 28172 22468 28200
rect 20809 28163 20867 28169
rect 22462 28160 22468 28172
rect 22520 28160 22526 28212
rect 22925 28203 22983 28209
rect 22925 28169 22937 28203
rect 22971 28200 22983 28203
rect 23382 28200 23388 28212
rect 22971 28172 23388 28200
rect 22971 28169 22983 28172
rect 22925 28163 22983 28169
rect 4847 28104 7788 28132
rect 4847 28101 4859 28104
rect 4801 28095 4859 28101
rect 8386 28092 8392 28144
rect 8444 28092 8450 28144
rect 9766 28132 9772 28144
rect 9727 28104 9772 28132
rect 9766 28092 9772 28104
rect 9824 28092 9830 28144
rect 11146 28132 11152 28144
rect 10994 28104 11152 28132
rect 11146 28092 11152 28104
rect 11204 28092 11210 28144
rect 13814 28092 13820 28144
rect 13872 28132 13878 28144
rect 13872 28104 15240 28132
rect 13872 28092 13878 28104
rect 6917 28067 6975 28073
rect 6917 28033 6929 28067
rect 6963 28064 6975 28067
rect 6963 28036 7604 28064
rect 6963 28033 6975 28036
rect 6917 28027 6975 28033
rect 4246 27956 4252 28008
rect 4304 27996 4310 28008
rect 4893 27999 4951 28005
rect 4893 27996 4905 27999
rect 4304 27968 4905 27996
rect 4304 27956 4310 27968
rect 4893 27965 4905 27968
rect 4939 27965 4951 27999
rect 4893 27959 4951 27965
rect 5077 27999 5135 28005
rect 5077 27965 5089 27999
rect 5123 27996 5135 27999
rect 7098 27996 7104 28008
rect 5123 27968 7104 27996
rect 5123 27965 5135 27968
rect 5077 27959 5135 27965
rect 7098 27956 7104 27968
rect 7156 27956 7162 28008
rect 6546 27860 6552 27872
rect 6507 27832 6552 27860
rect 6546 27820 6552 27832
rect 6604 27820 6610 27872
rect 7576 27869 7604 28036
rect 12434 28024 12440 28076
rect 12492 28064 12498 28076
rect 12492 28036 12537 28064
rect 12492 28024 12498 28036
rect 14090 28024 14096 28076
rect 14148 28064 14154 28076
rect 14752 28073 14780 28104
rect 14461 28067 14519 28073
rect 14461 28064 14473 28067
rect 14148 28036 14473 28064
rect 14148 28024 14154 28036
rect 14461 28033 14473 28036
rect 14507 28033 14519 28067
rect 14461 28027 14519 28033
rect 14737 28067 14795 28073
rect 14737 28033 14749 28067
rect 14783 28033 14795 28067
rect 14737 28027 14795 28033
rect 14921 28067 14979 28073
rect 14921 28033 14933 28067
rect 14967 28033 14979 28067
rect 14921 28027 14979 28033
rect 9030 27996 9036 28008
rect 8991 27968 9036 27996
rect 9030 27956 9036 27968
rect 9088 27956 9094 28008
rect 9306 27996 9312 28008
rect 9267 27968 9312 27996
rect 9306 27956 9312 27968
rect 9364 27996 9370 28008
rect 9493 27999 9551 28005
rect 9493 27996 9505 27999
rect 9364 27968 9505 27996
rect 9364 27956 9370 27968
rect 9493 27965 9505 27968
rect 9539 27965 9551 27999
rect 9493 27959 9551 27965
rect 14550 27888 14556 27940
rect 14608 27928 14614 27940
rect 14936 27928 14964 28027
rect 15212 27996 15240 28104
rect 15930 28092 15936 28144
rect 15988 28132 15994 28144
rect 22940 28132 22968 28163
rect 23382 28160 23388 28172
rect 23440 28160 23446 28212
rect 23658 28160 23664 28212
rect 23716 28200 23722 28212
rect 25041 28203 25099 28209
rect 25041 28200 25053 28203
rect 23716 28172 25053 28200
rect 23716 28160 23722 28172
rect 25041 28169 25053 28172
rect 25087 28200 25099 28203
rect 28534 28200 28540 28212
rect 25087 28172 28540 28200
rect 25087 28169 25099 28172
rect 25041 28163 25099 28169
rect 28534 28160 28540 28172
rect 28592 28160 28598 28212
rect 23566 28132 23572 28144
rect 15988 28104 20668 28132
rect 15988 28092 15994 28104
rect 15289 28067 15347 28073
rect 15289 28033 15301 28067
rect 15335 28064 15347 28067
rect 16390 28064 16396 28076
rect 15335 28036 16396 28064
rect 15335 28033 15347 28036
rect 15289 28027 15347 28033
rect 16390 28024 16396 28036
rect 16448 28024 16454 28076
rect 17954 28064 17960 28076
rect 17915 28036 17960 28064
rect 17954 28024 17960 28036
rect 18012 28024 18018 28076
rect 19426 28024 19432 28076
rect 19484 28064 19490 28076
rect 19990 28067 20048 28073
rect 19990 28064 20002 28067
rect 19484 28036 20002 28064
rect 19484 28024 19490 28036
rect 19990 28033 20002 28036
rect 20036 28033 20048 28067
rect 20254 28064 20260 28076
rect 20215 28036 20260 28064
rect 19990 28027 20048 28033
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 20640 28073 20668 28104
rect 22296 28104 22968 28132
rect 23527 28104 23572 28132
rect 20625 28067 20683 28073
rect 20625 28033 20637 28067
rect 20671 28033 20683 28067
rect 22186 28064 22192 28076
rect 20625 28027 20683 28033
rect 20732 28036 22192 28064
rect 15212 27968 15516 27996
rect 15488 27937 15516 27968
rect 16574 27956 16580 28008
rect 16632 27996 16638 28008
rect 17586 27996 17592 28008
rect 16632 27968 17592 27996
rect 16632 27956 16638 27968
rect 17586 27956 17592 27968
rect 17644 27956 17650 28008
rect 18233 27999 18291 28005
rect 18233 27965 18245 27999
rect 18279 27996 18291 27999
rect 18322 27996 18328 28008
rect 18279 27968 18328 27996
rect 18279 27965 18291 27968
rect 18233 27959 18291 27965
rect 18322 27956 18328 27968
rect 18380 27956 18386 28008
rect 14608 27900 14964 27928
rect 15473 27931 15531 27937
rect 14608 27888 14614 27900
rect 15473 27897 15485 27931
rect 15519 27928 15531 27931
rect 15519 27900 17724 27928
rect 15519 27897 15531 27900
rect 15473 27891 15531 27897
rect 7561 27863 7619 27869
rect 7561 27829 7573 27863
rect 7607 27860 7619 27863
rect 8938 27860 8944 27872
rect 7607 27832 8944 27860
rect 7607 27829 7619 27832
rect 7561 27823 7619 27829
rect 8938 27820 8944 27832
rect 8996 27820 9002 27872
rect 12618 27860 12624 27872
rect 12579 27832 12624 27860
rect 12618 27820 12624 27832
rect 12676 27820 12682 27872
rect 14458 27860 14464 27872
rect 14419 27832 14464 27860
rect 14458 27820 14464 27832
rect 14516 27820 14522 27872
rect 15746 27820 15752 27872
rect 15804 27860 15810 27872
rect 17589 27863 17647 27869
rect 17589 27860 17601 27863
rect 15804 27832 17601 27860
rect 15804 27820 15810 27832
rect 17589 27829 17601 27832
rect 17635 27829 17647 27863
rect 17696 27860 17724 27900
rect 20732 27860 20760 28036
rect 22186 28024 22192 28036
rect 22244 28024 22250 28076
rect 22296 28073 22324 28104
rect 23566 28092 23572 28104
rect 23624 28092 23630 28144
rect 25501 28135 25559 28141
rect 25501 28101 25513 28135
rect 25547 28132 25559 28135
rect 26786 28132 26792 28144
rect 25547 28104 26792 28132
rect 25547 28101 25559 28104
rect 25501 28095 25559 28101
rect 26786 28092 26792 28104
rect 26844 28092 26850 28144
rect 22281 28067 22339 28073
rect 22281 28033 22293 28067
rect 22327 28033 22339 28067
rect 22281 28027 22339 28033
rect 22741 28067 22799 28073
rect 22741 28033 22753 28067
rect 22787 28064 22799 28067
rect 23017 28067 23075 28073
rect 23017 28064 23029 28067
rect 22787 28036 23029 28064
rect 22787 28033 22799 28036
rect 22741 28027 22799 28033
rect 23017 28033 23029 28036
rect 23063 28064 23075 28067
rect 23109 28067 23167 28073
rect 23109 28064 23121 28067
rect 23063 28036 23121 28064
rect 23063 28033 23075 28036
rect 23017 28027 23075 28033
rect 23109 28033 23121 28036
rect 23155 28033 23167 28067
rect 23109 28027 23167 28033
rect 24670 28024 24676 28076
rect 24728 28024 24734 28076
rect 25222 28064 25228 28076
rect 25183 28036 25228 28064
rect 25222 28024 25228 28036
rect 25280 28024 25286 28076
rect 25406 28064 25412 28076
rect 25367 28036 25412 28064
rect 25406 28024 25412 28036
rect 25464 28024 25470 28076
rect 25598 28067 25656 28073
rect 25598 28033 25610 28067
rect 25644 28033 25656 28067
rect 25598 28027 25656 28033
rect 21266 27956 21272 28008
rect 21324 27996 21330 28008
rect 21726 27996 21732 28008
rect 21324 27968 21732 27996
rect 21324 27956 21330 27968
rect 21726 27956 21732 27968
rect 21784 27996 21790 28008
rect 23293 27999 23351 28005
rect 23293 27996 23305 27999
rect 21784 27968 23305 27996
rect 21784 27956 21790 27968
rect 23293 27965 23305 27968
rect 23339 27965 23351 27999
rect 23293 27959 23351 27965
rect 23658 27956 23664 28008
rect 23716 27996 23722 28008
rect 25613 27996 25641 28027
rect 23716 27968 25641 27996
rect 23716 27956 23722 27968
rect 21818 27888 21824 27940
rect 21876 27928 21882 27940
rect 22462 27928 22468 27940
rect 21876 27900 22468 27928
rect 21876 27888 21882 27900
rect 22462 27888 22468 27900
rect 22520 27888 22526 27940
rect 25406 27888 25412 27940
rect 25464 27928 25470 27940
rect 25961 27931 26019 27937
rect 25961 27928 25973 27931
rect 25464 27900 25973 27928
rect 25464 27888 25470 27900
rect 25961 27897 25973 27900
rect 26007 27897 26019 27931
rect 25961 27891 26019 27897
rect 22002 27860 22008 27872
rect 17696 27832 20760 27860
rect 21963 27832 22008 27860
rect 17589 27823 17647 27829
rect 22002 27820 22008 27832
rect 22060 27820 22066 27872
rect 22278 27820 22284 27872
rect 22336 27860 22342 27872
rect 22557 27863 22615 27869
rect 22557 27860 22569 27863
rect 22336 27832 22569 27860
rect 22336 27820 22342 27832
rect 22557 27829 22569 27832
rect 22603 27829 22615 27863
rect 22557 27823 22615 27829
rect 23109 27863 23167 27869
rect 23109 27829 23121 27863
rect 23155 27860 23167 27863
rect 23382 27860 23388 27872
rect 23155 27832 23388 27860
rect 23155 27829 23167 27832
rect 23109 27823 23167 27829
rect 23382 27820 23388 27832
rect 23440 27820 23446 27872
rect 25774 27860 25780 27872
rect 25735 27832 25780 27860
rect 25774 27820 25780 27832
rect 25832 27820 25838 27872
rect 1104 27770 29440 27792
rect 1104 27718 5672 27770
rect 5724 27718 5736 27770
rect 5788 27718 5800 27770
rect 5852 27718 5864 27770
rect 5916 27718 5928 27770
rect 5980 27718 15118 27770
rect 15170 27718 15182 27770
rect 15234 27718 15246 27770
rect 15298 27718 15310 27770
rect 15362 27718 15374 27770
rect 15426 27718 24563 27770
rect 24615 27718 24627 27770
rect 24679 27718 24691 27770
rect 24743 27718 24755 27770
rect 24807 27718 24819 27770
rect 24871 27718 29440 27770
rect 1104 27696 29440 27718
rect 4062 27616 4068 27668
rect 4120 27656 4126 27668
rect 10226 27656 10232 27668
rect 4120 27628 10088 27656
rect 10187 27628 10232 27656
rect 4120 27616 4126 27628
rect 4338 27588 4344 27600
rect 4299 27560 4344 27588
rect 4338 27548 4344 27560
rect 4396 27548 4402 27600
rect 8113 27591 8171 27597
rect 8113 27557 8125 27591
rect 8159 27588 8171 27591
rect 8570 27588 8576 27600
rect 8159 27560 8576 27588
rect 8159 27557 8171 27560
rect 8113 27551 8171 27557
rect 8570 27548 8576 27560
rect 8628 27548 8634 27600
rect 9030 27548 9036 27600
rect 9088 27588 9094 27600
rect 9493 27591 9551 27597
rect 9493 27588 9505 27591
rect 9088 27560 9505 27588
rect 9088 27548 9094 27560
rect 9493 27557 9505 27560
rect 9539 27557 9551 27591
rect 10060 27588 10088 27628
rect 10226 27616 10232 27628
rect 10284 27616 10290 27668
rect 16298 27656 16304 27668
rect 10352 27628 16304 27656
rect 10352 27588 10380 27628
rect 16298 27616 16304 27628
rect 16356 27656 16362 27668
rect 17218 27656 17224 27668
rect 16356 27628 17224 27656
rect 16356 27616 16362 27628
rect 17218 27616 17224 27628
rect 17276 27616 17282 27668
rect 17770 27616 17776 27668
rect 17828 27656 17834 27668
rect 19337 27659 19395 27665
rect 17828 27628 19288 27656
rect 17828 27616 17834 27628
rect 11330 27588 11336 27600
rect 9493 27551 9551 27557
rect 9600 27560 9812 27588
rect 10060 27560 10380 27588
rect 10428 27560 11336 27588
rect 4246 27520 4252 27532
rect 4080 27492 4252 27520
rect 4080 27461 4108 27492
rect 4246 27480 4252 27492
rect 4304 27480 4310 27532
rect 8938 27520 8944 27532
rect 8899 27492 8944 27520
rect 8938 27480 8944 27492
rect 8996 27480 9002 27532
rect 9306 27480 9312 27532
rect 9364 27520 9370 27532
rect 9600 27520 9628 27560
rect 9364 27492 9628 27520
rect 9677 27523 9735 27529
rect 9364 27480 9370 27492
rect 9677 27489 9689 27523
rect 9723 27489 9735 27523
rect 9784 27520 9812 27560
rect 10428 27520 10456 27560
rect 11330 27548 11336 27560
rect 11388 27548 11394 27600
rect 11701 27591 11759 27597
rect 11701 27557 11713 27591
rect 11747 27588 11759 27591
rect 12342 27588 12348 27600
rect 11747 27560 12348 27588
rect 11747 27557 11759 27560
rect 11701 27551 11759 27557
rect 12342 27548 12348 27560
rect 12400 27548 12406 27600
rect 17589 27591 17647 27597
rect 17589 27557 17601 27591
rect 17635 27557 17647 27591
rect 17589 27551 17647 27557
rect 18417 27591 18475 27597
rect 18417 27557 18429 27591
rect 18463 27588 18475 27591
rect 18690 27588 18696 27600
rect 18463 27560 18696 27588
rect 18463 27557 18475 27560
rect 18417 27551 18475 27557
rect 9784 27492 10456 27520
rect 10689 27523 10747 27529
rect 9677 27483 9735 27489
rect 10689 27489 10701 27523
rect 10735 27520 10747 27523
rect 10778 27520 10784 27532
rect 10735 27492 10784 27520
rect 10735 27489 10747 27492
rect 10689 27483 10747 27489
rect 4065 27455 4123 27461
rect 4065 27421 4077 27455
rect 4111 27421 4123 27455
rect 4065 27415 4123 27421
rect 4154 27412 4160 27464
rect 4212 27452 4218 27464
rect 4430 27452 4436 27464
rect 4212 27424 4257 27452
rect 4391 27424 4436 27452
rect 4212 27412 4218 27424
rect 4430 27412 4436 27424
rect 4488 27412 4494 27464
rect 7834 27412 7840 27464
rect 7892 27452 7898 27464
rect 7929 27455 7987 27461
rect 7929 27452 7941 27455
rect 7892 27424 7941 27452
rect 7892 27412 7898 27424
rect 7929 27421 7941 27424
rect 7975 27421 7987 27455
rect 7929 27415 7987 27421
rect 8294 27412 8300 27464
rect 8352 27452 8358 27464
rect 8389 27455 8447 27461
rect 8389 27452 8401 27455
rect 8352 27424 8401 27452
rect 8352 27412 8358 27424
rect 8389 27421 8401 27424
rect 8435 27421 8447 27455
rect 8389 27415 8447 27421
rect 9125 27455 9183 27461
rect 9125 27421 9137 27455
rect 9171 27452 9183 27455
rect 9398 27452 9404 27464
rect 9171 27424 9404 27452
rect 9171 27421 9183 27424
rect 9125 27415 9183 27421
rect 9398 27412 9404 27424
rect 9456 27452 9462 27464
rect 9692 27452 9720 27483
rect 10778 27480 10784 27492
rect 10836 27480 10842 27532
rect 11238 27480 11244 27532
rect 11296 27520 11302 27532
rect 11296 27492 11560 27520
rect 11296 27480 11302 27492
rect 11532 27461 11560 27492
rect 12710 27480 12716 27532
rect 12768 27520 12774 27532
rect 14185 27523 14243 27529
rect 14185 27520 14197 27523
rect 12768 27492 14197 27520
rect 12768 27480 12774 27492
rect 14185 27489 14197 27492
rect 14231 27489 14243 27523
rect 14185 27483 14243 27489
rect 9456 27424 9720 27452
rect 9769 27455 9827 27461
rect 9456 27412 9462 27424
rect 9769 27421 9781 27455
rect 9815 27421 9827 27455
rect 11517 27455 11575 27461
rect 9769 27415 9827 27421
rect 10704 27424 11468 27452
rect 9784 27384 9812 27415
rect 10704 27384 10732 27424
rect 9784 27356 10732 27384
rect 10781 27387 10839 27393
rect 10781 27353 10793 27387
rect 10827 27384 10839 27387
rect 10870 27384 10876 27396
rect 10827 27356 10876 27384
rect 10827 27353 10839 27356
rect 10781 27347 10839 27353
rect 10870 27344 10876 27356
rect 10928 27344 10934 27396
rect 11440 27384 11468 27424
rect 11517 27421 11529 27455
rect 11563 27421 11575 27455
rect 11517 27415 11575 27421
rect 13630 27412 13636 27464
rect 13688 27452 13694 27464
rect 14090 27452 14096 27464
rect 13688 27424 13781 27452
rect 14051 27424 14096 27452
rect 13688 27412 13694 27424
rect 14090 27412 14096 27424
rect 14148 27412 14154 27464
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27421 14427 27455
rect 14550 27452 14556 27464
rect 14511 27424 14556 27452
rect 14369 27415 14427 27421
rect 11440 27356 12020 27384
rect 3878 27316 3884 27328
rect 3839 27288 3884 27316
rect 3878 27276 3884 27288
rect 3936 27276 3942 27328
rect 8202 27276 8208 27328
rect 8260 27316 8266 27328
rect 8260 27288 8305 27316
rect 8260 27276 8266 27288
rect 10042 27276 10048 27328
rect 10100 27316 10106 27328
rect 10689 27319 10747 27325
rect 10689 27316 10701 27319
rect 10100 27288 10701 27316
rect 10100 27276 10106 27288
rect 10689 27285 10701 27288
rect 10735 27285 10747 27319
rect 10689 27279 10747 27285
rect 11606 27276 11612 27328
rect 11664 27316 11670 27328
rect 11885 27319 11943 27325
rect 11885 27316 11897 27319
rect 11664 27288 11897 27316
rect 11664 27276 11670 27288
rect 11885 27285 11897 27288
rect 11931 27285 11943 27319
rect 11992 27316 12020 27356
rect 12618 27344 12624 27396
rect 12676 27344 12682 27396
rect 13354 27384 13360 27396
rect 13315 27356 13360 27384
rect 13354 27344 13360 27356
rect 13412 27344 13418 27396
rect 12986 27316 12992 27328
rect 11992 27288 12992 27316
rect 11885 27279 11943 27285
rect 12986 27276 12992 27288
rect 13044 27276 13050 27328
rect 13078 27276 13084 27328
rect 13136 27316 13142 27328
rect 13648 27316 13676 27412
rect 13722 27344 13728 27396
rect 13780 27384 13786 27396
rect 14384 27384 14412 27415
rect 14550 27412 14556 27424
rect 14608 27412 14614 27464
rect 14921 27455 14979 27461
rect 14921 27421 14933 27455
rect 14967 27421 14979 27455
rect 15654 27452 15660 27464
rect 15615 27424 15660 27452
rect 14921 27415 14979 27421
rect 14936 27384 14964 27415
rect 15654 27412 15660 27424
rect 15712 27412 15718 27464
rect 17604 27452 17632 27551
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 19260 27588 19288 27628
rect 19337 27625 19349 27659
rect 19383 27656 19395 27659
rect 19426 27656 19432 27668
rect 19383 27628 19432 27656
rect 19383 27625 19395 27628
rect 19337 27619 19395 27625
rect 19426 27616 19432 27628
rect 19484 27616 19490 27668
rect 21542 27656 21548 27668
rect 19536 27628 21548 27656
rect 19536 27588 19564 27628
rect 21542 27616 21548 27628
rect 21600 27616 21606 27668
rect 23658 27656 23664 27668
rect 23619 27628 23664 27656
rect 23658 27616 23664 27628
rect 23716 27616 23722 27668
rect 25304 27659 25362 27665
rect 25304 27625 25316 27659
rect 25350 27656 25362 27659
rect 25774 27656 25780 27668
rect 25350 27628 25780 27656
rect 25350 27625 25362 27628
rect 25304 27619 25362 27625
rect 25774 27616 25780 27628
rect 25832 27616 25838 27668
rect 19260 27560 19564 27588
rect 19702 27548 19708 27600
rect 19760 27588 19766 27600
rect 22002 27588 22008 27600
rect 19760 27560 22008 27588
rect 19760 27548 19766 27560
rect 22002 27548 22008 27560
rect 22060 27588 22066 27600
rect 22554 27588 22560 27600
rect 22060 27560 22560 27588
rect 22060 27548 22066 27560
rect 22554 27548 22560 27560
rect 22612 27588 22618 27600
rect 22922 27588 22928 27600
rect 22612 27560 22928 27588
rect 22612 27548 22618 27560
rect 22922 27548 22928 27560
rect 22980 27548 22986 27600
rect 23290 27588 23296 27600
rect 23251 27560 23296 27588
rect 23290 27548 23296 27560
rect 23348 27548 23354 27600
rect 26786 27588 26792 27600
rect 26747 27560 26792 27588
rect 26786 27548 26792 27560
rect 26844 27548 26850 27600
rect 18233 27523 18291 27529
rect 18233 27489 18245 27523
rect 18279 27520 18291 27523
rect 18322 27520 18328 27532
rect 18279 27492 18328 27520
rect 18279 27489 18291 27492
rect 18233 27483 18291 27489
rect 15764 27424 17632 27452
rect 17957 27455 18015 27461
rect 15764 27384 15792 27424
rect 17957 27421 17969 27455
rect 18003 27452 18015 27455
rect 18046 27452 18052 27464
rect 18003 27424 18052 27452
rect 18003 27421 18015 27424
rect 17957 27415 18015 27421
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 13780 27356 14504 27384
rect 14936 27356 15792 27384
rect 15924 27387 15982 27393
rect 13780 27344 13786 27356
rect 13136 27288 13676 27316
rect 14476 27316 14504 27356
rect 15924 27353 15936 27387
rect 15970 27384 15982 27387
rect 16666 27384 16672 27396
rect 15970 27356 16672 27384
rect 15970 27353 15982 27356
rect 15924 27347 15982 27353
rect 16666 27344 16672 27356
rect 16724 27344 16730 27396
rect 17862 27384 17868 27396
rect 16776 27356 17868 27384
rect 15105 27319 15163 27325
rect 15105 27316 15117 27319
rect 14476 27288 15117 27316
rect 13136 27276 13142 27288
rect 15105 27285 15117 27288
rect 15151 27316 15163 27319
rect 16776 27316 16804 27356
rect 17862 27344 17868 27356
rect 17920 27344 17926 27396
rect 18248 27384 18276 27483
rect 18322 27480 18328 27492
rect 18380 27480 18386 27532
rect 18708 27520 18736 27548
rect 19613 27523 19671 27529
rect 19613 27520 19625 27523
rect 18708 27492 19625 27520
rect 19613 27489 19625 27492
rect 19659 27489 19671 27523
rect 23658 27520 23664 27532
rect 19613 27483 19671 27489
rect 19904 27492 20208 27520
rect 18414 27412 18420 27464
rect 18472 27452 18478 27464
rect 18601 27455 18659 27461
rect 18601 27452 18613 27455
rect 18472 27424 18613 27452
rect 18472 27412 18478 27424
rect 18601 27421 18613 27424
rect 18647 27421 18659 27455
rect 18601 27415 18659 27421
rect 18690 27412 18696 27464
rect 18748 27412 18754 27464
rect 18877 27455 18935 27461
rect 18877 27421 18889 27455
rect 18923 27452 18935 27455
rect 18966 27452 18972 27464
rect 18923 27424 18972 27452
rect 18923 27421 18935 27424
rect 18877 27415 18935 27421
rect 18966 27412 18972 27424
rect 19024 27412 19030 27464
rect 19242 27412 19248 27464
rect 19300 27452 19306 27464
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 19300 27424 19441 27452
rect 19300 27412 19306 27424
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 19705 27455 19763 27461
rect 19705 27421 19717 27455
rect 19751 27421 19763 27455
rect 19705 27415 19763 27421
rect 19815 27455 19873 27461
rect 19815 27421 19827 27455
rect 19861 27452 19873 27455
rect 19904 27452 19932 27492
rect 19861 27424 19932 27452
rect 19981 27455 20039 27461
rect 19861 27421 19873 27424
rect 19815 27415 19873 27421
rect 19981 27421 19993 27455
rect 20027 27421 20039 27455
rect 19981 27415 20039 27421
rect 18708 27384 18736 27412
rect 19720 27384 19748 27415
rect 18248 27356 18736 27384
rect 19076 27356 19748 27384
rect 19076 27328 19104 27356
rect 15151 27288 16804 27316
rect 15151 27285 15163 27288
rect 15105 27279 15163 27285
rect 16850 27276 16856 27328
rect 16908 27316 16914 27328
rect 17037 27319 17095 27325
rect 17037 27316 17049 27319
rect 16908 27288 17049 27316
rect 16908 27276 16914 27288
rect 17037 27285 17049 27288
rect 17083 27285 17095 27319
rect 17037 27279 17095 27285
rect 18049 27319 18107 27325
rect 18049 27285 18061 27319
rect 18095 27316 18107 27319
rect 18138 27316 18144 27328
rect 18095 27288 18144 27316
rect 18095 27285 18107 27288
rect 18049 27279 18107 27285
rect 18138 27276 18144 27288
rect 18196 27276 18202 27328
rect 18693 27319 18751 27325
rect 18693 27285 18705 27319
rect 18739 27316 18751 27319
rect 19058 27316 19064 27328
rect 18739 27288 19064 27316
rect 18739 27285 18751 27288
rect 18693 27279 18751 27285
rect 19058 27276 19064 27288
rect 19116 27276 19122 27328
rect 19334 27276 19340 27328
rect 19392 27316 19398 27328
rect 19996 27316 20024 27415
rect 20180 27328 20208 27492
rect 23313 27492 23664 27520
rect 20441 27455 20499 27461
rect 20441 27452 20453 27455
rect 20364 27424 20453 27452
rect 20364 27328 20392 27424
rect 20441 27421 20453 27424
rect 20487 27421 20499 27455
rect 22738 27452 22744 27464
rect 22699 27424 22744 27452
rect 20441 27415 20499 27421
rect 22738 27412 22744 27424
rect 22796 27412 22802 27464
rect 23014 27412 23020 27464
rect 23072 27452 23078 27464
rect 23161 27455 23219 27461
rect 23072 27424 23117 27452
rect 23072 27412 23078 27424
rect 23161 27421 23173 27455
rect 23207 27452 23219 27455
rect 23313 27452 23341 27492
rect 23658 27480 23664 27492
rect 23716 27480 23722 27532
rect 23753 27523 23811 27529
rect 23753 27489 23765 27523
rect 23799 27520 23811 27523
rect 24026 27520 24032 27532
rect 23799 27492 24032 27520
rect 23799 27489 23811 27492
rect 23753 27483 23811 27489
rect 24026 27480 24032 27492
rect 24084 27520 24090 27532
rect 24121 27523 24179 27529
rect 24121 27520 24133 27523
rect 24084 27492 24133 27520
rect 24084 27480 24090 27492
rect 24121 27489 24133 27492
rect 24167 27489 24179 27523
rect 24121 27483 24179 27489
rect 23474 27452 23480 27464
rect 23207 27424 23341 27452
rect 23435 27424 23480 27452
rect 23207 27421 23219 27424
rect 23161 27415 23219 27421
rect 23474 27412 23480 27424
rect 23532 27412 23538 27464
rect 23566 27412 23572 27464
rect 23624 27452 23630 27464
rect 23845 27455 23903 27461
rect 23845 27452 23857 27455
rect 23624 27424 23857 27452
rect 23624 27412 23630 27424
rect 23845 27421 23857 27424
rect 23891 27421 23903 27455
rect 23845 27415 23903 27421
rect 24765 27455 24823 27461
rect 24765 27421 24777 27455
rect 24811 27421 24823 27455
rect 24765 27415 24823 27421
rect 21450 27344 21456 27396
rect 21508 27384 21514 27396
rect 22554 27384 22560 27396
rect 21508 27356 22560 27384
rect 21508 27344 21514 27356
rect 22554 27344 22560 27356
rect 22612 27384 22618 27396
rect 22830 27384 22836 27396
rect 22612 27356 22836 27384
rect 22612 27344 22618 27356
rect 22830 27344 22836 27356
rect 22888 27384 22894 27396
rect 22925 27387 22983 27393
rect 22925 27384 22937 27387
rect 22888 27356 22937 27384
rect 22888 27344 22894 27356
rect 22925 27353 22937 27356
rect 22971 27384 22983 27387
rect 23753 27387 23811 27393
rect 23753 27384 23765 27387
rect 22971 27356 23765 27384
rect 22971 27353 22983 27356
rect 22925 27347 22983 27353
rect 23753 27353 23765 27356
rect 23799 27353 23811 27387
rect 24394 27384 24400 27396
rect 23753 27347 23811 27353
rect 23877 27356 24400 27384
rect 20162 27316 20168 27328
rect 19392 27288 20024 27316
rect 20123 27288 20168 27316
rect 19392 27276 19398 27288
rect 20162 27276 20168 27288
rect 20220 27276 20226 27328
rect 20346 27316 20352 27328
rect 20307 27288 20352 27316
rect 20346 27276 20352 27288
rect 20404 27276 20410 27328
rect 20625 27319 20683 27325
rect 20625 27285 20637 27319
rect 20671 27316 20683 27319
rect 23877 27316 23905 27356
rect 24394 27344 24400 27356
rect 24452 27384 24458 27396
rect 24780 27384 24808 27415
rect 24946 27412 24952 27464
rect 25004 27452 25010 27464
rect 25041 27455 25099 27461
rect 25041 27452 25053 27455
rect 25004 27424 25053 27452
rect 25004 27412 25010 27424
rect 25041 27421 25053 27424
rect 25087 27421 25099 27455
rect 25041 27415 25099 27421
rect 24452 27356 24808 27384
rect 24452 27344 24458 27356
rect 25866 27344 25872 27396
rect 25924 27344 25930 27396
rect 24026 27316 24032 27328
rect 20671 27288 23905 27316
rect 23987 27288 24032 27316
rect 20671 27285 20683 27288
rect 20625 27279 20683 27285
rect 24026 27276 24032 27288
rect 24084 27276 24090 27328
rect 24949 27319 25007 27325
rect 24949 27285 24961 27319
rect 24995 27316 25007 27319
rect 25682 27316 25688 27328
rect 24995 27288 25688 27316
rect 24995 27285 25007 27288
rect 24949 27279 25007 27285
rect 25682 27276 25688 27288
rect 25740 27276 25746 27328
rect 1104 27226 29440 27248
rect 1104 27174 10395 27226
rect 10447 27174 10459 27226
rect 10511 27174 10523 27226
rect 10575 27174 10587 27226
rect 10639 27174 10651 27226
rect 10703 27174 19840 27226
rect 19892 27174 19904 27226
rect 19956 27174 19968 27226
rect 20020 27174 20032 27226
rect 20084 27174 20096 27226
rect 20148 27174 29440 27226
rect 1104 27152 29440 27174
rect 4157 27115 4215 27121
rect 4157 27081 4169 27115
rect 4203 27112 4215 27115
rect 4246 27112 4252 27124
rect 4203 27084 4252 27112
rect 4203 27081 4215 27084
rect 4157 27075 4215 27081
rect 4246 27072 4252 27084
rect 4304 27072 4310 27124
rect 4430 27112 4436 27124
rect 4391 27084 4436 27112
rect 4430 27072 4436 27084
rect 4488 27072 4494 27124
rect 11149 27115 11207 27121
rect 4816 27084 11100 27112
rect 3044 27047 3102 27053
rect 3044 27013 3056 27047
rect 3090 27044 3102 27047
rect 3878 27044 3884 27056
rect 3090 27016 3884 27044
rect 3090 27013 3102 27016
rect 3044 27007 3102 27013
rect 3878 27004 3884 27016
rect 3936 27004 3942 27056
rect 3326 26936 3332 26988
rect 3384 26976 3390 26988
rect 4816 26985 4844 27084
rect 8202 27004 8208 27056
rect 8260 27004 8266 27056
rect 8849 27047 8907 27053
rect 8849 27013 8861 27047
rect 8895 27044 8907 27047
rect 9769 27047 9827 27053
rect 9769 27044 9781 27047
rect 8895 27016 9781 27044
rect 8895 27013 8907 27016
rect 8849 27007 8907 27013
rect 9769 27013 9781 27016
rect 9815 27013 9827 27047
rect 10962 27044 10968 27056
rect 9769 27007 9827 27013
rect 10244 27016 10968 27044
rect 4617 26979 4675 26985
rect 4617 26976 4629 26979
rect 3384 26948 4629 26976
rect 3384 26936 3390 26948
rect 4617 26945 4629 26948
rect 4663 26945 4675 26979
rect 4617 26939 4675 26945
rect 4801 26979 4859 26985
rect 4801 26945 4813 26979
rect 4847 26945 4859 26979
rect 4801 26939 4859 26945
rect 4893 26979 4951 26985
rect 4893 26945 4905 26979
rect 4939 26976 4951 26979
rect 4982 26976 4988 26988
rect 4939 26948 4988 26976
rect 4939 26945 4951 26948
rect 4893 26939 4951 26945
rect 4982 26936 4988 26948
rect 5040 26936 5046 26988
rect 5813 26979 5871 26985
rect 5813 26945 5825 26979
rect 5859 26945 5871 26979
rect 5813 26939 5871 26945
rect 5905 26979 5963 26985
rect 5905 26945 5917 26979
rect 5951 26976 5963 26979
rect 5994 26976 6000 26988
rect 5951 26948 6000 26976
rect 5951 26945 5963 26948
rect 5905 26939 5963 26945
rect 2682 26868 2688 26920
rect 2740 26908 2746 26920
rect 2777 26911 2835 26917
rect 2777 26908 2789 26911
rect 2740 26880 2789 26908
rect 2740 26868 2746 26880
rect 2777 26877 2789 26880
rect 2823 26877 2835 26911
rect 5828 26908 5856 26939
rect 5994 26936 6000 26948
rect 6052 26936 6058 26988
rect 6181 26979 6239 26985
rect 6181 26945 6193 26979
rect 6227 26976 6239 26979
rect 6546 26976 6552 26988
rect 6227 26948 6552 26976
rect 6227 26945 6239 26948
rect 6181 26939 6239 26945
rect 6546 26936 6552 26948
rect 6604 26936 6610 26988
rect 6825 26979 6883 26985
rect 6825 26945 6837 26979
rect 6871 26976 6883 26979
rect 9125 26979 9183 26985
rect 6871 26948 7420 26976
rect 6871 26945 6883 26948
rect 6825 26939 6883 26945
rect 6638 26908 6644 26920
rect 5828 26880 6644 26908
rect 2777 26871 2835 26877
rect 6638 26868 6644 26880
rect 6696 26908 6702 26920
rect 6917 26911 6975 26917
rect 6917 26908 6929 26911
rect 6696 26880 6929 26908
rect 6696 26868 6702 26880
rect 6917 26877 6929 26880
rect 6963 26877 6975 26911
rect 6917 26871 6975 26877
rect 7098 26868 7104 26920
rect 7156 26908 7162 26920
rect 7392 26917 7420 26948
rect 9125 26945 9137 26979
rect 9171 26976 9183 26979
rect 9306 26976 9312 26988
rect 9171 26948 9312 26976
rect 9171 26945 9183 26948
rect 9125 26939 9183 26945
rect 9306 26936 9312 26948
rect 9364 26936 9370 26988
rect 9398 26936 9404 26988
rect 9456 26976 9462 26988
rect 10045 26979 10103 26985
rect 9456 26948 9996 26976
rect 9456 26936 9462 26948
rect 9968 26917 9996 26948
rect 10045 26945 10057 26979
rect 10091 26976 10103 26979
rect 10244 26976 10272 27016
rect 10962 27004 10968 27016
rect 11020 27004 11026 27056
rect 11072 27044 11100 27084
rect 11149 27081 11161 27115
rect 11195 27112 11207 27115
rect 11238 27112 11244 27124
rect 11195 27084 11244 27112
rect 11195 27081 11207 27084
rect 11149 27075 11207 27081
rect 11238 27072 11244 27084
rect 11296 27072 11302 27124
rect 11517 27115 11575 27121
rect 11517 27081 11529 27115
rect 11563 27112 11575 27115
rect 12618 27112 12624 27124
rect 11563 27084 12624 27112
rect 11563 27081 11575 27084
rect 11517 27075 11575 27081
rect 12618 27072 12624 27084
rect 12676 27072 12682 27124
rect 12728 27084 12940 27112
rect 11606 27044 11612 27056
rect 11072 27016 11612 27044
rect 11606 27004 11612 27016
rect 11664 27004 11670 27056
rect 12253 27047 12311 27053
rect 12253 27013 12265 27047
rect 12299 27044 12311 27047
rect 12728 27044 12756 27084
rect 12299 27016 12756 27044
rect 12912 27044 12940 27084
rect 12986 27072 12992 27124
rect 13044 27112 13050 27124
rect 14458 27112 14464 27124
rect 13044 27084 14464 27112
rect 13044 27072 13050 27084
rect 14458 27072 14464 27084
rect 14516 27072 14522 27124
rect 14550 27072 14556 27124
rect 14608 27112 14614 27124
rect 14608 27084 14872 27112
rect 14608 27072 14614 27084
rect 13354 27044 13360 27056
rect 12912 27016 13360 27044
rect 12299 27013 12311 27016
rect 12253 27007 12311 27013
rect 13354 27004 13360 27016
rect 13412 27004 13418 27056
rect 10091 26948 10272 26976
rect 10091 26945 10103 26948
rect 10045 26939 10103 26945
rect 10318 26936 10324 26988
rect 10376 26976 10382 26988
rect 10505 26979 10563 26985
rect 10505 26976 10517 26979
rect 10376 26948 10517 26976
rect 10376 26936 10382 26948
rect 10505 26945 10517 26948
rect 10551 26976 10563 26979
rect 10870 26976 10876 26988
rect 10551 26948 10876 26976
rect 10551 26945 10563 26948
rect 10505 26939 10563 26945
rect 10870 26936 10876 26948
rect 10928 26936 10934 26988
rect 11054 26936 11060 26988
rect 11112 26976 11118 26988
rect 11333 26979 11391 26985
rect 11333 26976 11345 26979
rect 11112 26948 11345 26976
rect 11112 26936 11118 26948
rect 11333 26945 11345 26948
rect 11379 26976 11391 26979
rect 11517 26979 11575 26985
rect 11517 26976 11529 26979
rect 11379 26948 11529 26976
rect 11379 26945 11391 26948
rect 11333 26939 11391 26945
rect 11517 26945 11529 26948
rect 11563 26945 11575 26979
rect 11624 26976 11652 27004
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11624 26948 11713 26976
rect 11517 26939 11575 26945
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26976 11943 26979
rect 12158 26976 12164 26988
rect 11931 26948 12164 26976
rect 11931 26945 11943 26948
rect 11885 26939 11943 26945
rect 12158 26936 12164 26948
rect 12216 26976 12222 26988
rect 12529 26979 12587 26985
rect 12360 26976 12480 26979
rect 12216 26951 12480 26976
rect 12216 26948 12388 26951
rect 12216 26936 12222 26948
rect 7377 26911 7435 26917
rect 7156 26880 7249 26908
rect 7156 26868 7162 26880
rect 7377 26877 7389 26911
rect 7423 26908 7435 26911
rect 9217 26911 9275 26917
rect 9217 26908 9229 26911
rect 7423 26880 9229 26908
rect 7423 26877 7435 26880
rect 7377 26871 7435 26877
rect 9217 26877 9229 26880
rect 9263 26877 9275 26911
rect 9217 26871 9275 26877
rect 9953 26911 10011 26917
rect 9953 26877 9965 26911
rect 9999 26908 10011 26911
rect 12452 26908 12480 26951
rect 12529 26945 12541 26979
rect 12575 26976 12587 26979
rect 12710 26976 12716 26988
rect 12575 26948 12716 26976
rect 12575 26945 12587 26948
rect 12529 26939 12587 26945
rect 12710 26936 12716 26948
rect 12768 26936 12774 26988
rect 13538 26976 13544 26988
rect 13499 26948 13544 26976
rect 13538 26936 13544 26948
rect 13596 26936 13602 26988
rect 14090 26936 14096 26988
rect 14148 26936 14154 26988
rect 14458 26936 14464 26988
rect 14516 26976 14522 26988
rect 14844 26985 14872 27084
rect 14918 27072 14924 27124
rect 14976 27112 14982 27124
rect 15657 27115 15715 27121
rect 15657 27112 15669 27115
rect 14976 27084 15669 27112
rect 14976 27072 14982 27084
rect 15657 27081 15669 27084
rect 15703 27112 15715 27115
rect 15703 27084 15884 27112
rect 15703 27081 15715 27084
rect 15657 27075 15715 27081
rect 15746 27044 15752 27056
rect 15120 27016 15752 27044
rect 15120 26985 15148 27016
rect 15746 27004 15752 27016
rect 15804 27004 15810 27056
rect 15856 27044 15884 27084
rect 16298 27072 16304 27124
rect 16356 27112 16362 27124
rect 16393 27115 16451 27121
rect 16393 27112 16405 27115
rect 16356 27084 16405 27112
rect 16356 27072 16362 27084
rect 16393 27081 16405 27084
rect 16439 27081 16451 27115
rect 21450 27112 21456 27124
rect 16393 27075 16451 27081
rect 16500 27084 21456 27112
rect 16500 27044 16528 27084
rect 21450 27072 21456 27084
rect 21508 27072 21514 27124
rect 21637 27115 21695 27121
rect 21637 27081 21649 27115
rect 21683 27081 21695 27115
rect 21637 27075 21695 27081
rect 21913 27115 21971 27121
rect 21913 27081 21925 27115
rect 21959 27112 21971 27115
rect 23014 27112 23020 27124
rect 21959 27084 23020 27112
rect 21959 27081 21971 27084
rect 21913 27075 21971 27081
rect 15856 27016 16528 27044
rect 18506 27004 18512 27056
rect 18564 27044 18570 27056
rect 18564 27016 18609 27044
rect 18564 27004 18570 27016
rect 18782 27004 18788 27056
rect 18840 27044 18846 27056
rect 19334 27044 19340 27056
rect 18840 27016 19340 27044
rect 18840 27004 18846 27016
rect 19334 27004 19340 27016
rect 19392 27004 19398 27056
rect 21652 27044 21680 27075
rect 23014 27072 23020 27084
rect 23072 27072 23078 27124
rect 23474 27072 23480 27124
rect 23532 27112 23538 27124
rect 23845 27115 23903 27121
rect 23845 27112 23857 27115
rect 23532 27084 23857 27112
rect 23532 27072 23538 27084
rect 23845 27081 23857 27084
rect 23891 27112 23903 27115
rect 24486 27112 24492 27124
rect 23891 27084 24492 27112
rect 23891 27081 23903 27084
rect 23845 27075 23903 27081
rect 24486 27072 24492 27084
rect 24544 27072 24550 27124
rect 25866 27112 25872 27124
rect 25827 27084 25872 27112
rect 25866 27072 25872 27084
rect 25924 27072 25930 27124
rect 21652 27016 22218 27044
rect 23290 27004 23296 27056
rect 23348 27044 23354 27056
rect 23385 27047 23443 27053
rect 23385 27044 23397 27047
rect 23348 27016 23397 27044
rect 23348 27004 23354 27016
rect 23385 27013 23397 27016
rect 23431 27013 23443 27047
rect 23385 27007 23443 27013
rect 24026 27004 24032 27056
rect 24084 27044 24090 27056
rect 24084 27016 24150 27044
rect 24084 27004 24090 27016
rect 14645 26979 14703 26985
rect 14516 26948 14561 26976
rect 14516 26936 14522 26948
rect 14645 26945 14657 26979
rect 14691 26945 14703 26979
rect 14645 26939 14703 26945
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26945 14887 26979
rect 14829 26939 14887 26945
rect 15105 26979 15163 26985
rect 15105 26945 15117 26979
rect 15151 26945 15163 26979
rect 15105 26939 15163 26945
rect 12621 26911 12679 26917
rect 12621 26908 12633 26911
rect 9999 26880 10364 26908
rect 12452 26880 12633 26908
rect 9999 26877 10011 26880
rect 9953 26871 10011 26877
rect 4062 26800 4068 26852
rect 4120 26840 4126 26852
rect 7116 26840 7144 26868
rect 7558 26840 7564 26852
rect 4120 26812 6592 26840
rect 7116 26812 7564 26840
rect 4120 26800 4126 26812
rect 4338 26732 4344 26784
rect 4396 26772 4402 26784
rect 5077 26775 5135 26781
rect 5077 26772 5089 26775
rect 4396 26744 5089 26772
rect 4396 26732 4402 26744
rect 5077 26741 5089 26744
rect 5123 26741 5135 26775
rect 5077 26735 5135 26741
rect 5534 26732 5540 26784
rect 5592 26772 5598 26784
rect 5629 26775 5687 26781
rect 5629 26772 5641 26775
rect 5592 26744 5641 26772
rect 5592 26732 5598 26744
rect 5629 26741 5641 26744
rect 5675 26741 5687 26775
rect 6086 26772 6092 26784
rect 6047 26744 6092 26772
rect 5629 26735 5687 26741
rect 6086 26732 6092 26744
rect 6144 26732 6150 26784
rect 6454 26772 6460 26784
rect 6415 26744 6460 26772
rect 6454 26732 6460 26744
rect 6512 26732 6518 26784
rect 6564 26772 6592 26812
rect 7558 26800 7564 26812
rect 7616 26800 7622 26852
rect 10336 26849 10364 26880
rect 12621 26877 12633 26880
rect 12667 26877 12679 26911
rect 14108 26908 14136 26936
rect 14476 26908 14504 26936
rect 12621 26871 12679 26877
rect 13740 26880 14504 26908
rect 13740 26849 13768 26880
rect 10321 26843 10379 26849
rect 10321 26809 10333 26843
rect 10367 26809 10379 26843
rect 10321 26803 10379 26809
rect 13725 26843 13783 26849
rect 13725 26809 13737 26843
rect 13771 26809 13783 26843
rect 13725 26803 13783 26809
rect 14090 26800 14096 26852
rect 14148 26840 14154 26852
rect 14660 26840 14688 26939
rect 15194 26936 15200 26988
rect 15252 26976 15258 26988
rect 15289 26979 15347 26985
rect 15289 26976 15301 26979
rect 15252 26948 15301 26976
rect 15252 26936 15258 26948
rect 15289 26945 15301 26948
rect 15335 26976 15347 26979
rect 16022 26976 16028 26988
rect 15335 26948 16028 26976
rect 15335 26945 15347 26948
rect 15289 26939 15347 26945
rect 16022 26936 16028 26948
rect 16080 26936 16086 26988
rect 16666 26976 16672 26988
rect 16627 26948 16672 26976
rect 16666 26936 16672 26948
rect 16724 26936 16730 26988
rect 16758 26936 16764 26988
rect 16816 26976 16822 26988
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16816 26948 16865 26976
rect 16816 26936 16822 26948
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 17218 26936 17224 26988
rect 17276 26976 17282 26988
rect 17276 26948 17321 26976
rect 17276 26936 17282 26948
rect 17402 26936 17408 26988
rect 17460 26976 17466 26988
rect 18969 26979 19027 26985
rect 17460 26948 17505 26976
rect 17460 26936 17466 26948
rect 18969 26945 18981 26979
rect 19015 26945 19027 26979
rect 19150 26976 19156 26988
rect 19111 26948 19156 26976
rect 18969 26939 19027 26945
rect 17034 26908 17040 26920
rect 16995 26880 17040 26908
rect 17034 26868 17040 26880
rect 17092 26868 17098 26920
rect 17126 26868 17132 26920
rect 17184 26908 17190 26920
rect 17184 26880 17229 26908
rect 17184 26868 17190 26880
rect 18598 26868 18604 26920
rect 18656 26908 18662 26920
rect 18785 26911 18843 26917
rect 18656 26880 18701 26908
rect 18656 26868 18662 26880
rect 18785 26877 18797 26911
rect 18831 26877 18843 26911
rect 18984 26908 19012 26939
rect 19150 26936 19156 26948
rect 19208 26936 19214 26988
rect 19518 26976 19524 26988
rect 19479 26948 19524 26976
rect 19518 26936 19524 26948
rect 19576 26936 19582 26988
rect 19705 26979 19763 26985
rect 19705 26945 19717 26979
rect 19751 26976 19763 26979
rect 21002 26979 21060 26985
rect 21002 26976 21014 26979
rect 19751 26948 21014 26976
rect 19751 26945 19763 26948
rect 19705 26939 19763 26945
rect 21002 26945 21014 26948
rect 21048 26945 21060 26979
rect 21002 26939 21060 26945
rect 21453 26979 21511 26985
rect 21453 26945 21465 26979
rect 21499 26976 21511 26979
rect 21634 26976 21640 26988
rect 21499 26948 21640 26976
rect 21499 26945 21511 26948
rect 21453 26939 21511 26945
rect 21634 26936 21640 26948
rect 21692 26936 21698 26988
rect 25682 26976 25688 26988
rect 25643 26948 25688 26976
rect 25682 26936 25688 26948
rect 25740 26936 25746 26988
rect 19058 26908 19064 26920
rect 18984 26880 19064 26908
rect 18785 26871 18843 26877
rect 14918 26840 14924 26852
rect 14148 26812 14924 26840
rect 14148 26800 14154 26812
rect 14918 26800 14924 26812
rect 14976 26800 14982 26852
rect 15746 26800 15752 26852
rect 15804 26840 15810 26852
rect 15804 26812 18276 26840
rect 15804 26800 15810 26812
rect 10042 26772 10048 26784
rect 6564 26744 10048 26772
rect 10042 26732 10048 26744
rect 10100 26732 10106 26784
rect 12526 26732 12532 26784
rect 12584 26772 12590 26784
rect 14369 26775 14427 26781
rect 14369 26772 14381 26775
rect 12584 26744 14381 26772
rect 12584 26732 12590 26744
rect 14369 26741 14381 26744
rect 14415 26741 14427 26775
rect 14369 26735 14427 26741
rect 14458 26732 14464 26784
rect 14516 26772 14522 26784
rect 14826 26772 14832 26784
rect 14516 26744 14832 26772
rect 14516 26732 14522 26744
rect 14826 26732 14832 26744
rect 14884 26732 14890 26784
rect 15470 26772 15476 26784
rect 15431 26744 15476 26772
rect 15470 26732 15476 26744
rect 15528 26732 15534 26784
rect 16482 26732 16488 26784
rect 16540 26772 16546 26784
rect 18141 26775 18199 26781
rect 18141 26772 18153 26775
rect 16540 26744 18153 26772
rect 16540 26732 16546 26744
rect 18141 26741 18153 26744
rect 18187 26741 18199 26775
rect 18248 26772 18276 26812
rect 18690 26800 18696 26852
rect 18748 26840 18754 26852
rect 18800 26840 18828 26871
rect 19058 26868 19064 26880
rect 19116 26868 19122 26920
rect 19242 26908 19248 26920
rect 19203 26880 19248 26908
rect 19242 26868 19248 26880
rect 19300 26868 19306 26920
rect 19337 26911 19395 26917
rect 19337 26877 19349 26911
rect 19383 26877 19395 26911
rect 21266 26908 21272 26920
rect 21227 26880 21272 26908
rect 19337 26871 19395 26877
rect 18748 26812 18828 26840
rect 18748 26800 18754 26812
rect 18874 26800 18880 26852
rect 18932 26840 18938 26852
rect 19352 26840 19380 26871
rect 21266 26868 21272 26880
rect 21324 26868 21330 26920
rect 23661 26911 23719 26917
rect 23661 26877 23673 26911
rect 23707 26908 23719 26911
rect 24946 26908 24952 26920
rect 23707 26880 24952 26908
rect 23707 26877 23719 26880
rect 23661 26871 23719 26877
rect 24946 26868 24952 26880
rect 25004 26868 25010 26920
rect 25314 26908 25320 26920
rect 25275 26880 25320 26908
rect 25314 26868 25320 26880
rect 25372 26868 25378 26920
rect 25593 26911 25651 26917
rect 25593 26877 25605 26911
rect 25639 26877 25651 26911
rect 25593 26871 25651 26877
rect 18932 26812 19380 26840
rect 19443 26812 20024 26840
rect 18932 26800 18938 26812
rect 19443 26772 19471 26812
rect 18248 26744 19471 26772
rect 18141 26735 18199 26741
rect 19518 26732 19524 26784
rect 19576 26772 19582 26784
rect 19889 26775 19947 26781
rect 19889 26772 19901 26775
rect 19576 26744 19901 26772
rect 19576 26732 19582 26744
rect 19889 26741 19901 26744
rect 19935 26741 19947 26775
rect 19996 26772 20024 26812
rect 22646 26772 22652 26784
rect 19996 26744 22652 26772
rect 19889 26735 19947 26741
rect 22646 26732 22652 26744
rect 22704 26772 22710 26784
rect 23014 26772 23020 26784
rect 22704 26744 23020 26772
rect 22704 26732 22710 26744
rect 23014 26732 23020 26744
rect 23072 26732 23078 26784
rect 24946 26732 24952 26784
rect 25004 26772 25010 26784
rect 25608 26772 25636 26871
rect 25004 26744 25636 26772
rect 25004 26732 25010 26744
rect 1104 26682 29440 26704
rect 1104 26630 5672 26682
rect 5724 26630 5736 26682
rect 5788 26630 5800 26682
rect 5852 26630 5864 26682
rect 5916 26630 5928 26682
rect 5980 26630 15118 26682
rect 15170 26630 15182 26682
rect 15234 26630 15246 26682
rect 15298 26630 15310 26682
rect 15362 26630 15374 26682
rect 15426 26630 24563 26682
rect 24615 26630 24627 26682
rect 24679 26630 24691 26682
rect 24743 26630 24755 26682
rect 24807 26630 24819 26682
rect 24871 26630 29440 26682
rect 1104 26608 29440 26630
rect 4065 26571 4123 26577
rect 4065 26537 4077 26571
rect 4111 26568 4123 26571
rect 4154 26568 4160 26580
rect 4111 26540 4160 26568
rect 4111 26537 4123 26540
rect 4065 26531 4123 26537
rect 4154 26528 4160 26540
rect 4212 26528 4218 26580
rect 6638 26568 6644 26580
rect 6599 26540 6644 26568
rect 6638 26528 6644 26540
rect 6696 26528 6702 26580
rect 8294 26568 8300 26580
rect 8255 26540 8300 26568
rect 8294 26528 8300 26540
rect 8352 26528 8358 26580
rect 10318 26568 10324 26580
rect 10279 26540 10324 26568
rect 10318 26528 10324 26540
rect 10376 26528 10382 26580
rect 10778 26568 10784 26580
rect 10739 26540 10784 26568
rect 10778 26528 10784 26540
rect 10836 26528 10842 26580
rect 10962 26528 10968 26580
rect 11020 26568 11026 26580
rect 12621 26571 12679 26577
rect 12621 26568 12633 26571
rect 11020 26540 12633 26568
rect 11020 26528 11026 26540
rect 12621 26537 12633 26540
rect 12667 26537 12679 26571
rect 12621 26531 12679 26537
rect 13170 26528 13176 26580
rect 13228 26568 13234 26580
rect 14550 26568 14556 26580
rect 13228 26540 14556 26568
rect 13228 26528 13234 26540
rect 14550 26528 14556 26540
rect 14608 26528 14614 26580
rect 15565 26571 15623 26577
rect 15565 26537 15577 26571
rect 15611 26568 15623 26571
rect 15746 26568 15752 26580
rect 15611 26540 15752 26568
rect 15611 26537 15623 26540
rect 15565 26531 15623 26537
rect 15746 26528 15752 26540
rect 15804 26528 15810 26580
rect 16390 26568 16396 26580
rect 16351 26540 16396 26568
rect 16390 26528 16396 26540
rect 16448 26528 16454 26580
rect 21634 26568 21640 26580
rect 21595 26540 21640 26568
rect 21634 26528 21640 26540
rect 21692 26528 21698 26580
rect 22189 26571 22247 26577
rect 22189 26537 22201 26571
rect 22235 26568 22247 26571
rect 23566 26568 23572 26580
rect 22235 26540 23572 26568
rect 22235 26537 22247 26540
rect 22189 26531 22247 26537
rect 23566 26528 23572 26540
rect 23624 26528 23630 26580
rect 23753 26571 23811 26577
rect 23753 26537 23765 26571
rect 23799 26568 23811 26571
rect 25314 26568 25320 26580
rect 23799 26540 25320 26568
rect 23799 26537 23811 26540
rect 23753 26531 23811 26537
rect 25314 26528 25320 26540
rect 25372 26528 25378 26580
rect 14277 26503 14335 26509
rect 14277 26500 14289 26503
rect 11164 26472 14289 26500
rect 5166 26392 5172 26444
rect 5224 26432 5230 26444
rect 5261 26435 5319 26441
rect 5261 26432 5273 26435
rect 5224 26404 5273 26432
rect 5224 26392 5230 26404
rect 5261 26401 5273 26404
rect 5307 26401 5319 26435
rect 11054 26432 11060 26444
rect 5261 26395 5319 26401
rect 8036 26404 11060 26432
rect 8036 26376 8064 26404
rect 11054 26392 11060 26404
rect 11112 26392 11118 26444
rect 2774 26324 2780 26376
rect 2832 26364 2838 26376
rect 2961 26367 3019 26373
rect 2961 26364 2973 26367
rect 2832 26336 2973 26364
rect 2832 26324 2838 26336
rect 2961 26333 2973 26336
rect 3007 26333 3019 26367
rect 2961 26327 3019 26333
rect 3237 26367 3295 26373
rect 3237 26333 3249 26367
rect 3283 26364 3295 26367
rect 3326 26364 3332 26376
rect 3283 26336 3332 26364
rect 3283 26333 3295 26336
rect 3237 26327 3295 26333
rect 3326 26324 3332 26336
rect 3384 26324 3390 26376
rect 4249 26367 4307 26373
rect 4249 26333 4261 26367
rect 4295 26364 4307 26367
rect 4890 26364 4896 26376
rect 4295 26336 4896 26364
rect 4295 26333 4307 26336
rect 4249 26327 4307 26333
rect 4890 26324 4896 26336
rect 4948 26324 4954 26376
rect 5534 26373 5540 26376
rect 5528 26364 5540 26373
rect 5495 26336 5540 26364
rect 5528 26327 5540 26336
rect 5534 26324 5540 26327
rect 5592 26324 5598 26376
rect 8018 26364 8024 26376
rect 7979 26336 8024 26364
rect 8018 26324 8024 26336
rect 8076 26324 8082 26376
rect 8113 26367 8171 26373
rect 8113 26333 8125 26367
rect 8159 26333 8171 26367
rect 8113 26327 8171 26333
rect 8128 26296 8156 26327
rect 9582 26324 9588 26376
rect 9640 26364 9646 26376
rect 11164 26373 11192 26472
rect 14277 26469 14289 26472
rect 14323 26469 14335 26503
rect 14918 26500 14924 26512
rect 14277 26463 14335 26469
rect 14384 26472 14924 26500
rect 11333 26435 11391 26441
rect 11333 26432 11345 26435
rect 11256 26404 11345 26432
rect 10505 26367 10563 26373
rect 10505 26364 10517 26367
rect 9640 26336 10517 26364
rect 9640 26324 9646 26336
rect 10505 26333 10517 26336
rect 10551 26333 10563 26367
rect 10505 26327 10563 26333
rect 11149 26367 11207 26373
rect 11149 26333 11161 26367
rect 11195 26333 11207 26367
rect 11149 26327 11207 26333
rect 7852 26268 8156 26296
rect 7852 26240 7880 26268
rect 10962 26256 10968 26308
rect 11020 26296 11026 26308
rect 11256 26296 11284 26404
rect 11333 26401 11345 26404
rect 11379 26401 11391 26435
rect 13538 26432 13544 26444
rect 11333 26395 11391 26401
rect 12728 26404 13544 26432
rect 12728 26373 12756 26404
rect 13538 26392 13544 26404
rect 13596 26392 13602 26444
rect 12713 26367 12771 26373
rect 12713 26333 12725 26367
rect 12759 26333 12771 26367
rect 12713 26327 12771 26333
rect 12897 26367 12955 26373
rect 12897 26333 12909 26367
rect 12943 26333 12955 26367
rect 13170 26364 13176 26376
rect 13131 26336 13176 26364
rect 12897 26327 12955 26333
rect 12912 26296 12940 26327
rect 13170 26324 13176 26336
rect 13228 26324 13234 26376
rect 13449 26367 13507 26373
rect 13449 26333 13461 26367
rect 13495 26364 13507 26367
rect 14384 26364 14412 26472
rect 14918 26460 14924 26472
rect 14976 26460 14982 26512
rect 15010 26460 15016 26512
rect 15068 26500 15074 26512
rect 17497 26503 17555 26509
rect 17497 26500 17509 26503
rect 15068 26472 17509 26500
rect 15068 26460 15074 26472
rect 17497 26469 17509 26472
rect 17543 26469 17555 26503
rect 18690 26500 18696 26512
rect 17497 26463 17555 26469
rect 17788 26472 18696 26500
rect 16482 26432 16488 26444
rect 14752 26404 16488 26432
rect 13495 26336 14412 26364
rect 14456 26367 14514 26373
rect 13495 26333 13507 26336
rect 13449 26327 13507 26333
rect 14456 26333 14468 26367
rect 14502 26364 14514 26367
rect 14752 26364 14780 26404
rect 16482 26392 16488 26404
rect 16540 26392 16546 26444
rect 16850 26432 16856 26444
rect 16811 26404 16856 26432
rect 16850 26392 16856 26404
rect 16908 26392 16914 26444
rect 17037 26435 17095 26441
rect 17037 26401 17049 26435
rect 17083 26432 17095 26435
rect 17218 26432 17224 26444
rect 17083 26404 17224 26432
rect 17083 26401 17095 26404
rect 17037 26395 17095 26401
rect 17218 26392 17224 26404
rect 17276 26432 17282 26444
rect 17788 26432 17816 26472
rect 18064 26441 18092 26472
rect 18690 26460 18696 26472
rect 18748 26460 18754 26512
rect 18782 26460 18788 26512
rect 18840 26500 18846 26512
rect 19242 26500 19248 26512
rect 18840 26472 19248 26500
rect 18840 26460 18846 26472
rect 19242 26460 19248 26472
rect 19300 26460 19306 26512
rect 20162 26460 20168 26512
rect 20220 26500 20226 26512
rect 29549 26503 29607 26509
rect 29549 26500 29561 26503
rect 20220 26472 29561 26500
rect 20220 26460 20226 26472
rect 29549 26469 29561 26472
rect 29595 26469 29607 26503
rect 29549 26463 29607 26469
rect 17276 26404 17816 26432
rect 18049 26435 18107 26441
rect 17276 26392 17282 26404
rect 18049 26401 18061 26435
rect 18095 26401 18107 26435
rect 18049 26395 18107 26401
rect 18598 26392 18604 26444
rect 18656 26432 18662 26444
rect 18966 26432 18972 26444
rect 18656 26404 18972 26432
rect 18656 26392 18662 26404
rect 18966 26392 18972 26404
rect 19024 26392 19030 26444
rect 19150 26392 19156 26444
rect 19208 26432 19214 26444
rect 19889 26435 19947 26441
rect 19889 26432 19901 26435
rect 19208 26404 19901 26432
rect 19208 26392 19214 26404
rect 19889 26401 19901 26404
rect 19935 26432 19947 26435
rect 23934 26432 23940 26444
rect 19935 26404 23940 26432
rect 19935 26401 19947 26404
rect 19889 26395 19947 26401
rect 23934 26392 23940 26404
rect 23992 26392 23998 26444
rect 14502 26336 14780 26364
rect 14502 26333 14514 26336
rect 14456 26327 14514 26333
rect 14826 26324 14832 26376
rect 14884 26364 14890 26376
rect 15105 26367 15163 26373
rect 14884 26336 14929 26364
rect 14884 26324 14890 26336
rect 15105 26333 15117 26367
rect 15151 26364 15163 26367
rect 15470 26364 15476 26376
rect 15151 26336 15476 26364
rect 15151 26333 15163 26336
rect 15105 26327 15163 26333
rect 15470 26324 15476 26336
rect 15528 26324 15534 26376
rect 16761 26367 16819 26373
rect 16761 26333 16773 26367
rect 16807 26364 16819 26367
rect 17310 26364 17316 26376
rect 16807 26336 17316 26364
rect 16807 26333 16819 26336
rect 16761 26327 16819 26333
rect 17310 26324 17316 26336
rect 17368 26324 17374 26376
rect 17957 26367 18015 26373
rect 17957 26333 17969 26367
rect 18003 26364 18015 26367
rect 18138 26364 18144 26376
rect 18003 26336 18144 26364
rect 18003 26333 18015 26336
rect 17957 26327 18015 26333
rect 18138 26324 18144 26336
rect 18196 26324 18202 26376
rect 18414 26324 18420 26376
rect 18472 26364 18478 26376
rect 18877 26367 18935 26373
rect 18877 26364 18889 26367
rect 18472 26336 18889 26364
rect 18472 26324 18478 26336
rect 18877 26333 18889 26336
rect 18923 26333 18935 26367
rect 18984 26364 19012 26392
rect 19429 26367 19487 26373
rect 19429 26364 19441 26367
rect 18984 26336 19441 26364
rect 18877 26327 18935 26333
rect 19429 26333 19441 26336
rect 19475 26333 19487 26367
rect 19429 26327 19487 26333
rect 21821 26367 21879 26373
rect 21821 26333 21833 26367
rect 21867 26364 21879 26367
rect 22005 26367 22063 26373
rect 22005 26364 22017 26367
rect 21867 26336 22017 26364
rect 21867 26333 21879 26336
rect 21821 26327 21879 26333
rect 22005 26333 22017 26336
rect 22051 26364 22063 26367
rect 22281 26367 22339 26373
rect 22281 26364 22293 26367
rect 22051 26336 22293 26364
rect 22051 26333 22063 26336
rect 22005 26327 22063 26333
rect 22281 26333 22293 26336
rect 22327 26333 22339 26367
rect 22281 26327 22339 26333
rect 13633 26299 13691 26305
rect 13633 26296 13645 26299
rect 11020 26268 11284 26296
rect 12406 26268 13645 26296
rect 11020 26256 11026 26268
rect 3050 26228 3056 26240
rect 3011 26200 3056 26228
rect 3050 26188 3056 26200
rect 3108 26188 3114 26240
rect 7834 26228 7840 26240
rect 7795 26200 7840 26228
rect 7834 26188 7840 26200
rect 7892 26188 7898 26240
rect 11241 26231 11299 26237
rect 11241 26197 11253 26231
rect 11287 26228 11299 26231
rect 11422 26228 11428 26240
rect 11287 26200 11428 26228
rect 11287 26197 11299 26200
rect 11241 26191 11299 26197
rect 11422 26188 11428 26200
rect 11480 26228 11486 26240
rect 11609 26231 11667 26237
rect 11609 26228 11621 26231
rect 11480 26200 11621 26228
rect 11480 26188 11486 26200
rect 11609 26197 11621 26200
rect 11655 26197 11667 26231
rect 12158 26228 12164 26240
rect 12119 26200 12164 26228
rect 11609 26191 11667 26197
rect 12158 26188 12164 26200
rect 12216 26228 12222 26240
rect 12406 26228 12434 26268
rect 13633 26265 13645 26268
rect 13679 26265 13691 26299
rect 14550 26296 14556 26308
rect 14511 26268 14556 26296
rect 13633 26259 13691 26265
rect 12216 26200 12434 26228
rect 13648 26228 13676 26259
rect 14550 26256 14556 26268
rect 14608 26256 14614 26308
rect 14645 26299 14703 26305
rect 14645 26265 14657 26299
rect 14691 26296 14703 26299
rect 15197 26299 15255 26305
rect 15197 26296 15209 26299
rect 14691 26268 15209 26296
rect 14691 26265 14703 26268
rect 14645 26259 14703 26265
rect 15197 26265 15209 26268
rect 15243 26265 15255 26299
rect 15197 26259 15255 26265
rect 13998 26228 14004 26240
rect 13648 26200 14004 26228
rect 12216 26188 12222 26200
rect 13998 26188 14004 26200
rect 14056 26188 14062 26240
rect 14458 26188 14464 26240
rect 14516 26228 14522 26240
rect 14660 26228 14688 26259
rect 15654 26256 15660 26308
rect 15712 26296 15718 26308
rect 18690 26296 18696 26308
rect 15712 26268 18184 26296
rect 18651 26268 18696 26296
rect 15712 26256 15718 26268
rect 18156 26240 18184 26268
rect 18690 26256 18696 26268
rect 18748 26256 18754 26308
rect 19610 26296 19616 26308
rect 19571 26268 19616 26296
rect 19610 26256 19616 26268
rect 19668 26256 19674 26308
rect 21545 26299 21603 26305
rect 21545 26265 21557 26299
rect 21591 26296 21603 26299
rect 21726 26296 21732 26308
rect 21591 26268 21732 26296
rect 21591 26265 21603 26268
rect 21545 26259 21603 26265
rect 21726 26256 21732 26268
rect 21784 26296 21790 26308
rect 21836 26296 21864 26327
rect 22738 26324 22744 26376
rect 22796 26364 22802 26376
rect 23198 26364 23204 26376
rect 22796 26336 23204 26364
rect 22796 26324 22802 26336
rect 23198 26324 23204 26336
rect 23256 26324 23262 26376
rect 23474 26364 23480 26376
rect 23435 26336 23480 26364
rect 23474 26324 23480 26336
rect 23532 26324 23538 26376
rect 23658 26373 23664 26376
rect 23621 26367 23664 26373
rect 23621 26333 23633 26367
rect 23621 26327 23664 26333
rect 23658 26324 23664 26327
rect 23716 26324 23722 26376
rect 23106 26296 23112 26308
rect 21784 26268 21864 26296
rect 23067 26268 23112 26296
rect 21784 26256 21790 26268
rect 23106 26256 23112 26268
rect 23164 26296 23170 26308
rect 23385 26299 23443 26305
rect 23385 26296 23397 26299
rect 23164 26268 23397 26296
rect 23164 26256 23170 26268
rect 23385 26265 23397 26268
rect 23431 26265 23443 26299
rect 23385 26259 23443 26265
rect 14516 26200 14688 26228
rect 14516 26188 14522 26200
rect 14734 26188 14740 26240
rect 14792 26228 14798 26240
rect 14921 26231 14979 26237
rect 14921 26228 14933 26231
rect 14792 26200 14933 26228
rect 14792 26188 14798 26200
rect 14921 26197 14933 26200
rect 14967 26197 14979 26231
rect 17862 26228 17868 26240
rect 17823 26200 17868 26228
rect 14921 26191 14979 26197
rect 17862 26188 17868 26200
rect 17920 26188 17926 26240
rect 18138 26188 18144 26240
rect 18196 26228 18202 26240
rect 18601 26231 18659 26237
rect 18601 26228 18613 26231
rect 18196 26200 18613 26228
rect 18196 26188 18202 26200
rect 18601 26197 18613 26200
rect 18647 26197 18659 26231
rect 18601 26191 18659 26197
rect 18874 26188 18880 26240
rect 18932 26228 18938 26240
rect 19061 26231 19119 26237
rect 19061 26228 19073 26231
rect 18932 26200 19073 26228
rect 18932 26188 18938 26200
rect 19061 26197 19073 26200
rect 19107 26197 19119 26231
rect 19061 26191 19119 26197
rect 1104 26138 29440 26160
rect 1104 26086 10395 26138
rect 10447 26086 10459 26138
rect 10511 26086 10523 26138
rect 10575 26086 10587 26138
rect 10639 26086 10651 26138
rect 10703 26086 19840 26138
rect 19892 26086 19904 26138
rect 19956 26086 19968 26138
rect 20020 26086 20032 26138
rect 20084 26086 20096 26138
rect 20148 26086 29440 26138
rect 1104 26064 29440 26086
rect 5166 25984 5172 26036
rect 5224 25984 5230 26036
rect 5353 26027 5411 26033
rect 5353 25993 5365 26027
rect 5399 26024 5411 26027
rect 5994 26024 6000 26036
rect 5399 25996 6000 26024
rect 5399 25993 5411 25996
rect 5353 25987 5411 25993
rect 5994 25984 6000 25996
rect 6052 26024 6058 26036
rect 6052 25996 6684 26024
rect 6052 25984 6058 25996
rect 2682 25956 2688 25968
rect 1780 25928 2688 25956
rect 1394 25848 1400 25900
rect 1452 25888 1458 25900
rect 1780 25897 1808 25928
rect 2682 25916 2688 25928
rect 2740 25956 2746 25968
rect 5184 25956 5212 25984
rect 2740 25928 5212 25956
rect 2740 25916 2746 25928
rect 1765 25891 1823 25897
rect 1765 25888 1777 25891
rect 1452 25860 1777 25888
rect 1452 25848 1458 25860
rect 1765 25857 1777 25860
rect 1811 25857 1823 25891
rect 1765 25851 1823 25857
rect 2032 25891 2090 25897
rect 2032 25857 2044 25891
rect 2078 25888 2090 25891
rect 2590 25888 2596 25900
rect 2078 25860 2596 25888
rect 2078 25857 2090 25860
rect 2032 25851 2090 25857
rect 2590 25848 2596 25860
rect 2648 25848 2654 25900
rect 3620 25897 3648 25928
rect 3878 25897 3884 25900
rect 3605 25891 3663 25897
rect 3605 25857 3617 25891
rect 3651 25857 3663 25891
rect 3872 25888 3884 25897
rect 3839 25860 3884 25888
rect 3605 25851 3663 25857
rect 3872 25851 3884 25860
rect 3878 25848 3884 25851
rect 3936 25848 3942 25900
rect 4890 25848 4896 25900
rect 4948 25888 4954 25900
rect 5169 25891 5227 25897
rect 5169 25888 5181 25891
rect 4948 25860 5181 25888
rect 4948 25848 4954 25860
rect 5169 25857 5181 25860
rect 5215 25857 5227 25891
rect 5169 25851 5227 25857
rect 6365 25891 6423 25897
rect 6365 25857 6377 25891
rect 6411 25888 6423 25891
rect 6454 25888 6460 25900
rect 6411 25860 6460 25888
rect 6411 25857 6423 25860
rect 6365 25851 6423 25857
rect 6454 25848 6460 25860
rect 6512 25848 6518 25900
rect 6656 25897 6684 25996
rect 10134 25984 10140 26036
rect 10192 26024 10198 26036
rect 10229 26027 10287 26033
rect 10229 26024 10241 26027
rect 10192 25996 10241 26024
rect 10192 25984 10198 25996
rect 10229 25993 10241 25996
rect 10275 25993 10287 26027
rect 10229 25987 10287 25993
rect 10597 26027 10655 26033
rect 10597 25993 10609 26027
rect 10643 26024 10655 26027
rect 14812 26027 14870 26033
rect 14812 26024 14824 26027
rect 10643 25996 14824 26024
rect 10643 25993 10655 25996
rect 10597 25987 10655 25993
rect 14812 25993 14824 25996
rect 14858 25993 14870 26027
rect 15562 26024 15568 26036
rect 15523 25996 15568 26024
rect 14812 25987 14870 25993
rect 15562 25984 15568 25996
rect 15620 25984 15626 26036
rect 17126 26024 17132 26036
rect 16040 25996 17132 26024
rect 9214 25916 9220 25968
rect 9272 25956 9278 25968
rect 9401 25959 9459 25965
rect 9401 25956 9413 25959
rect 9272 25928 9413 25956
rect 9272 25916 9278 25928
rect 9401 25925 9413 25928
rect 9447 25925 9459 25959
rect 9401 25919 9459 25925
rect 11517 25959 11575 25965
rect 11517 25925 11529 25959
rect 11563 25956 11575 25959
rect 12158 25956 12164 25968
rect 11563 25928 12164 25956
rect 11563 25925 11575 25928
rect 11517 25919 11575 25925
rect 12158 25916 12164 25928
rect 12216 25916 12222 25968
rect 12805 25959 12863 25965
rect 12805 25956 12817 25959
rect 12268 25928 12817 25956
rect 6641 25891 6699 25897
rect 6641 25857 6653 25891
rect 6687 25857 6699 25891
rect 6641 25851 6699 25857
rect 6730 25848 6736 25900
rect 6788 25888 6794 25900
rect 8389 25891 8447 25897
rect 6788 25860 6833 25888
rect 6788 25848 6794 25860
rect 8389 25857 8401 25891
rect 8435 25888 8447 25891
rect 8435 25860 8984 25888
rect 8435 25857 8447 25860
rect 8389 25851 8447 25857
rect 6086 25712 6092 25764
rect 6144 25752 6150 25764
rect 8956 25761 8984 25860
rect 10870 25848 10876 25900
rect 10928 25888 10934 25900
rect 11149 25891 11207 25897
rect 11149 25888 11161 25891
rect 10928 25860 11161 25888
rect 10928 25848 10934 25860
rect 11149 25857 11161 25860
rect 11195 25857 11207 25891
rect 11790 25888 11796 25900
rect 11703 25860 11796 25888
rect 11149 25851 11207 25857
rect 11790 25848 11796 25860
rect 11848 25888 11854 25900
rect 12268 25888 12296 25928
rect 12805 25925 12817 25928
rect 12851 25956 12863 25959
rect 15197 25959 15255 25965
rect 15197 25956 15209 25959
rect 12851 25928 15209 25956
rect 12851 25925 12863 25928
rect 12805 25919 12863 25925
rect 15197 25925 15209 25928
rect 15243 25956 15255 25959
rect 15470 25956 15476 25968
rect 15243 25928 15476 25956
rect 15243 25925 15255 25928
rect 15197 25919 15255 25925
rect 15470 25916 15476 25928
rect 15528 25916 15534 25968
rect 15580 25956 15608 25984
rect 15580 25928 15957 25956
rect 15929 25900 15957 25928
rect 11848 25860 12296 25888
rect 12345 25891 12403 25897
rect 11848 25848 11854 25860
rect 12345 25857 12357 25891
rect 12391 25888 12403 25891
rect 12526 25888 12532 25900
rect 12391 25860 12532 25888
rect 12391 25857 12403 25860
rect 12345 25851 12403 25857
rect 12526 25848 12532 25860
rect 12584 25888 12590 25900
rect 14458 25888 14464 25900
rect 12584 25860 14464 25888
rect 12584 25848 12590 25860
rect 14458 25848 14464 25860
rect 14516 25848 14522 25900
rect 14553 25891 14611 25897
rect 14553 25857 14565 25891
rect 14599 25888 14611 25891
rect 14734 25888 14740 25900
rect 14599 25860 14740 25888
rect 14599 25857 14611 25860
rect 14553 25851 14611 25857
rect 14734 25848 14740 25860
rect 14792 25848 14798 25900
rect 15010 25897 15016 25900
rect 15008 25888 15016 25897
rect 14971 25860 15016 25888
rect 15008 25851 15016 25860
rect 15010 25848 15016 25851
rect 15068 25848 15074 25900
rect 15102 25848 15108 25900
rect 15160 25888 15166 25900
rect 15381 25891 15439 25897
rect 15160 25860 15205 25888
rect 15160 25848 15166 25860
rect 15381 25857 15393 25891
rect 15427 25857 15439 25891
rect 15746 25888 15752 25900
rect 15707 25860 15752 25888
rect 15381 25851 15439 25857
rect 9398 25820 9404 25832
rect 9359 25792 9404 25820
rect 9398 25780 9404 25792
rect 9456 25780 9462 25832
rect 9493 25823 9551 25829
rect 9493 25789 9505 25823
rect 9539 25820 9551 25823
rect 9582 25820 9588 25832
rect 9539 25792 9588 25820
rect 9539 25789 9551 25792
rect 9493 25783 9551 25789
rect 9582 25780 9588 25792
rect 9640 25780 9646 25832
rect 10134 25780 10140 25832
rect 10192 25820 10198 25832
rect 10689 25823 10747 25829
rect 10689 25820 10701 25823
rect 10192 25792 10701 25820
rect 10192 25780 10198 25792
rect 10689 25789 10701 25792
rect 10735 25789 10747 25823
rect 10689 25783 10747 25789
rect 10781 25823 10839 25829
rect 10781 25789 10793 25823
rect 10827 25820 10839 25823
rect 10962 25820 10968 25832
rect 10827 25792 10968 25820
rect 10827 25789 10839 25792
rect 10781 25783 10839 25789
rect 10962 25780 10968 25792
rect 11020 25780 11026 25832
rect 11698 25820 11704 25832
rect 11659 25792 11704 25820
rect 11698 25780 11704 25792
rect 11756 25780 11762 25832
rect 12989 25823 13047 25829
rect 12989 25789 13001 25823
rect 13035 25820 13047 25823
rect 14090 25820 14096 25832
rect 13035 25792 14096 25820
rect 13035 25789 13047 25792
rect 12989 25783 13047 25789
rect 6457 25755 6515 25761
rect 6457 25752 6469 25755
rect 6144 25724 6469 25752
rect 6144 25712 6150 25724
rect 6457 25721 6469 25724
rect 6503 25721 6515 25755
rect 6457 25715 6515 25721
rect 8941 25755 8999 25761
rect 8941 25721 8953 25755
rect 8987 25721 8999 25755
rect 11330 25752 11336 25764
rect 11291 25724 11336 25752
rect 8941 25715 8999 25721
rect 11330 25712 11336 25724
rect 11388 25712 11394 25764
rect 13004 25752 13032 25783
rect 14090 25780 14096 25792
rect 14148 25780 14154 25832
rect 14826 25780 14832 25832
rect 14884 25820 14890 25832
rect 15396 25820 15424 25851
rect 15746 25848 15752 25860
rect 15804 25848 15810 25900
rect 15914 25894 15972 25900
rect 16040 25897 16068 25996
rect 17126 25984 17132 25996
rect 17184 26024 17190 26036
rect 18782 26024 18788 26036
rect 17184 25996 18788 26024
rect 17184 25984 17190 25996
rect 18782 25984 18788 25996
rect 18840 25984 18846 26036
rect 19610 25984 19616 26036
rect 19668 26024 19674 26036
rect 26234 26024 26240 26036
rect 19668 25996 26240 26024
rect 19668 25984 19674 25996
rect 26234 25984 26240 25996
rect 26292 25984 26298 26036
rect 26973 26027 27031 26033
rect 26973 25993 26985 26027
rect 27019 25993 27031 26027
rect 26973 25987 27031 25993
rect 17034 25956 17040 25968
rect 16132 25928 17040 25956
rect 16132 25897 16160 25928
rect 17034 25916 17040 25928
rect 17092 25956 17098 25968
rect 19628 25956 19656 25984
rect 17092 25928 18644 25956
rect 17092 25916 17098 25928
rect 15914 25860 15926 25894
rect 15960 25860 15972 25894
rect 15914 25854 15972 25860
rect 16025 25891 16083 25897
rect 16025 25857 16037 25891
rect 16071 25857 16083 25891
rect 16025 25851 16083 25857
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25857 16175 25891
rect 16117 25851 16175 25857
rect 16301 25891 16359 25897
rect 16301 25857 16313 25891
rect 16347 25857 16359 25891
rect 16301 25851 16359 25857
rect 16485 25891 16543 25897
rect 16485 25857 16497 25891
rect 16531 25888 16543 25891
rect 17874 25891 17932 25897
rect 17874 25888 17886 25891
rect 16531 25860 17886 25888
rect 16531 25857 16543 25860
rect 16485 25851 16543 25857
rect 17874 25857 17886 25860
rect 17920 25857 17932 25891
rect 17874 25851 17932 25857
rect 18509 25891 18567 25897
rect 18509 25857 18521 25891
rect 18555 25857 18567 25891
rect 18509 25851 18567 25857
rect 14884 25792 15424 25820
rect 16316 25820 16344 25851
rect 18138 25820 18144 25832
rect 16316 25792 16804 25820
rect 18099 25792 18144 25820
rect 14884 25780 14890 25792
rect 13170 25752 13176 25764
rect 11808 25724 13032 25752
rect 13083 25724 13176 25752
rect 2774 25644 2780 25696
rect 2832 25684 2838 25696
rect 3145 25687 3203 25693
rect 3145 25684 3157 25687
rect 2832 25656 3157 25684
rect 2832 25644 2838 25656
rect 3145 25653 3157 25656
rect 3191 25653 3203 25687
rect 3145 25647 3203 25653
rect 3970 25644 3976 25696
rect 4028 25684 4034 25696
rect 4985 25687 5043 25693
rect 4985 25684 4997 25687
rect 4028 25656 4997 25684
rect 4028 25644 4034 25656
rect 4985 25653 4997 25656
rect 5031 25653 5043 25687
rect 6914 25684 6920 25696
rect 6875 25656 6920 25684
rect 4985 25647 5043 25653
rect 6914 25644 6920 25656
rect 6972 25644 6978 25696
rect 7742 25644 7748 25696
rect 7800 25684 7806 25696
rect 11808 25693 11836 25724
rect 13170 25712 13176 25724
rect 13228 25752 13234 25764
rect 13814 25752 13820 25764
rect 13228 25724 13820 25752
rect 13228 25712 13234 25724
rect 13814 25712 13820 25724
rect 13872 25712 13878 25764
rect 14550 25712 14556 25764
rect 14608 25752 14614 25764
rect 15010 25752 15016 25764
rect 14608 25724 15016 25752
rect 14608 25712 14614 25724
rect 15010 25712 15016 25724
rect 15068 25712 15074 25764
rect 16776 25696 16804 25792
rect 18138 25780 18144 25792
rect 18196 25780 18202 25832
rect 8205 25687 8263 25693
rect 8205 25684 8217 25687
rect 7800 25656 8217 25684
rect 7800 25644 7806 25656
rect 8205 25653 8217 25656
rect 8251 25653 8263 25687
rect 8205 25647 8263 25653
rect 11793 25687 11851 25693
rect 11793 25653 11805 25687
rect 11839 25653 11851 25687
rect 11793 25647 11851 25653
rect 11977 25687 12035 25693
rect 11977 25653 11989 25687
rect 12023 25684 12035 25687
rect 12066 25684 12072 25696
rect 12023 25656 12072 25684
rect 12023 25653 12035 25656
rect 11977 25647 12035 25653
rect 12066 25644 12072 25656
rect 12124 25644 12130 25696
rect 12250 25684 12256 25696
rect 12211 25656 12256 25684
rect 12250 25644 12256 25656
rect 12308 25644 12314 25696
rect 12526 25684 12532 25696
rect 12487 25656 12532 25684
rect 12526 25644 12532 25656
rect 12584 25644 12590 25696
rect 12986 25644 12992 25696
rect 13044 25684 13050 25696
rect 13357 25687 13415 25693
rect 13357 25684 13369 25687
rect 13044 25656 13369 25684
rect 13044 25644 13050 25656
rect 13357 25653 13369 25656
rect 13403 25684 13415 25687
rect 13630 25684 13636 25696
rect 13403 25656 13636 25684
rect 13403 25653 13415 25656
rect 13357 25647 13415 25653
rect 13630 25644 13636 25656
rect 13688 25644 13694 25696
rect 14366 25684 14372 25696
rect 14327 25656 14372 25684
rect 14366 25644 14372 25656
rect 14424 25644 14430 25696
rect 16758 25684 16764 25696
rect 16719 25656 16764 25684
rect 16758 25644 16764 25656
rect 16816 25644 16822 25696
rect 18524 25684 18552 25851
rect 18616 25752 18644 25928
rect 18800 25928 19656 25956
rect 18692 25891 18750 25897
rect 18692 25857 18704 25891
rect 18738 25888 18750 25891
rect 18800 25888 18828 25928
rect 20254 25916 20260 25968
rect 20312 25956 20318 25968
rect 26988 25956 27016 25987
rect 20312 25928 20852 25956
rect 26450 25928 27016 25956
rect 20312 25916 20318 25928
rect 20824 25897 20852 25928
rect 18738 25860 18828 25888
rect 19061 25891 19119 25897
rect 18738 25857 18750 25860
rect 18692 25851 18750 25857
rect 19061 25857 19073 25891
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 19245 25891 19303 25897
rect 19245 25857 19257 25891
rect 19291 25888 19303 25891
rect 20542 25891 20600 25897
rect 20542 25888 20554 25891
rect 19291 25860 20554 25888
rect 19291 25857 19303 25860
rect 19245 25851 19303 25857
rect 20542 25857 20554 25860
rect 20588 25857 20600 25891
rect 20542 25851 20600 25857
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25857 20867 25891
rect 22002 25888 22008 25900
rect 21963 25860 22008 25888
rect 20809 25851 20867 25857
rect 18782 25820 18788 25832
rect 18743 25792 18788 25820
rect 18782 25780 18788 25792
rect 18840 25780 18846 25832
rect 18874 25780 18880 25832
rect 18932 25820 18938 25832
rect 19076 25820 19104 25851
rect 22002 25848 22008 25860
rect 22060 25848 22066 25900
rect 23290 25888 23296 25900
rect 23251 25860 23296 25888
rect 23290 25848 23296 25860
rect 23348 25848 23354 25900
rect 27154 25888 27160 25900
rect 27115 25860 27160 25888
rect 27154 25848 27160 25860
rect 27212 25848 27218 25900
rect 24946 25820 24952 25832
rect 18932 25792 19025 25820
rect 19076 25792 19472 25820
rect 24907 25792 24952 25820
rect 18932 25780 18938 25792
rect 18892 25752 18920 25780
rect 19334 25752 19340 25764
rect 18616 25724 18920 25752
rect 19306 25712 19340 25752
rect 19392 25712 19398 25764
rect 19306 25684 19334 25712
rect 19444 25696 19472 25792
rect 24946 25780 24952 25792
rect 25004 25780 25010 25832
rect 25222 25820 25228 25832
rect 25183 25792 25228 25820
rect 25222 25780 25228 25792
rect 25280 25780 25286 25832
rect 26697 25823 26755 25829
rect 26697 25789 26709 25823
rect 26743 25820 26755 25823
rect 27062 25820 27068 25832
rect 26743 25792 27068 25820
rect 26743 25789 26755 25792
rect 26697 25783 26755 25789
rect 27062 25780 27068 25792
rect 27120 25780 27126 25832
rect 19426 25684 19432 25696
rect 18524 25656 19334 25684
rect 19387 25656 19432 25684
rect 19426 25644 19432 25656
rect 19484 25644 19490 25696
rect 21818 25684 21824 25696
rect 21779 25656 21824 25684
rect 21818 25644 21824 25656
rect 21876 25644 21882 25696
rect 22186 25644 22192 25696
rect 22244 25684 22250 25696
rect 22646 25684 22652 25696
rect 22244 25656 22652 25684
rect 22244 25644 22250 25656
rect 22646 25644 22652 25656
rect 22704 25684 22710 25696
rect 23569 25687 23627 25693
rect 23569 25684 23581 25687
rect 22704 25656 23581 25684
rect 22704 25644 22710 25656
rect 23569 25653 23581 25656
rect 23615 25684 23627 25687
rect 25406 25684 25412 25696
rect 23615 25656 25412 25684
rect 23615 25653 23627 25656
rect 23569 25647 23627 25653
rect 25406 25644 25412 25656
rect 25464 25644 25470 25696
rect 1104 25594 29440 25616
rect 1104 25542 5672 25594
rect 5724 25542 5736 25594
rect 5788 25542 5800 25594
rect 5852 25542 5864 25594
rect 5916 25542 5928 25594
rect 5980 25542 15118 25594
rect 15170 25542 15182 25594
rect 15234 25542 15246 25594
rect 15298 25542 15310 25594
rect 15362 25542 15374 25594
rect 15426 25542 24563 25594
rect 24615 25542 24627 25594
rect 24679 25542 24691 25594
rect 24743 25542 24755 25594
rect 24807 25542 24819 25594
rect 24871 25542 29440 25594
rect 1104 25520 29440 25542
rect 2590 25440 2596 25492
rect 2648 25480 2654 25492
rect 2685 25483 2743 25489
rect 2685 25480 2697 25483
rect 2648 25452 2697 25480
rect 2648 25440 2654 25452
rect 2685 25449 2697 25452
rect 2731 25449 2743 25483
rect 2685 25443 2743 25449
rect 3050 25440 3056 25492
rect 3108 25480 3114 25492
rect 3145 25483 3203 25489
rect 3145 25480 3157 25483
rect 3108 25452 3157 25480
rect 3108 25440 3114 25452
rect 3145 25449 3157 25452
rect 3191 25449 3203 25483
rect 3878 25480 3884 25492
rect 3839 25452 3884 25480
rect 3145 25443 3203 25449
rect 3878 25440 3884 25452
rect 3936 25440 3942 25492
rect 6641 25483 6699 25489
rect 6641 25449 6653 25483
rect 6687 25480 6699 25483
rect 6730 25480 6736 25492
rect 6687 25452 6736 25480
rect 6687 25449 6699 25452
rect 6641 25443 6699 25449
rect 6730 25440 6736 25452
rect 6788 25480 6794 25492
rect 6788 25452 7328 25480
rect 6788 25440 6794 25452
rect 4982 25412 4988 25424
rect 3252 25384 4988 25412
rect 2774 25236 2780 25288
rect 2832 25276 2838 25288
rect 3252 25285 3280 25384
rect 4982 25372 4988 25384
rect 5040 25372 5046 25424
rect 4154 25344 4160 25356
rect 3712 25316 4160 25344
rect 2869 25279 2927 25285
rect 2869 25276 2881 25279
rect 2832 25248 2881 25276
rect 2832 25236 2838 25248
rect 2869 25245 2881 25248
rect 2915 25245 2927 25279
rect 2869 25239 2927 25245
rect 2961 25279 3019 25285
rect 2961 25245 2973 25279
rect 3007 25245 3019 25279
rect 2961 25239 3019 25245
rect 3237 25279 3295 25285
rect 3237 25245 3249 25279
rect 3283 25245 3295 25279
rect 3237 25239 3295 25245
rect 2976 25208 3004 25239
rect 3712 25208 3740 25316
rect 4154 25304 4160 25316
rect 4212 25344 4218 25356
rect 4212 25316 4292 25344
rect 4212 25304 4218 25316
rect 4062 25285 4068 25288
rect 4060 25276 4068 25285
rect 4023 25248 4068 25276
rect 4060 25239 4068 25248
rect 4062 25236 4068 25239
rect 4120 25236 4126 25288
rect 4264 25285 4292 25316
rect 5166 25304 5172 25356
rect 5224 25344 5230 25356
rect 7300 25353 7328 25452
rect 9398 25440 9404 25492
rect 9456 25480 9462 25492
rect 9953 25483 10011 25489
rect 9953 25480 9965 25483
rect 9456 25452 9965 25480
rect 9456 25440 9462 25452
rect 9953 25449 9965 25452
rect 9999 25449 10011 25483
rect 9953 25443 10011 25449
rect 11517 25483 11575 25489
rect 11517 25449 11529 25483
rect 11563 25480 11575 25483
rect 11790 25480 11796 25492
rect 11563 25452 11796 25480
rect 11563 25449 11575 25452
rect 11517 25443 11575 25449
rect 8665 25415 8723 25421
rect 8665 25381 8677 25415
rect 8711 25381 8723 25415
rect 8665 25375 8723 25381
rect 5261 25347 5319 25353
rect 5261 25344 5273 25347
rect 5224 25316 5273 25344
rect 5224 25304 5230 25316
rect 5261 25313 5273 25316
rect 5307 25313 5319 25347
rect 5261 25307 5319 25313
rect 7285 25347 7343 25353
rect 7285 25313 7297 25347
rect 7331 25313 7343 25347
rect 7285 25307 7343 25313
rect 7469 25347 7527 25353
rect 7469 25313 7481 25347
rect 7515 25344 7527 25347
rect 7558 25344 7564 25356
rect 7515 25316 7564 25344
rect 7515 25313 7527 25316
rect 7469 25307 7527 25313
rect 7558 25304 7564 25316
rect 7616 25304 7622 25356
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25245 4307 25279
rect 4430 25276 4436 25288
rect 4391 25248 4436 25276
rect 4249 25239 4307 25245
rect 4430 25236 4436 25248
rect 4488 25236 4494 25288
rect 5528 25279 5586 25285
rect 5528 25245 5540 25279
rect 5574 25276 5586 25279
rect 6914 25276 6920 25288
rect 5574 25248 6920 25276
rect 5574 25245 5586 25248
rect 5528 25239 5586 25245
rect 6914 25236 6920 25248
rect 6972 25236 6978 25288
rect 7834 25276 7840 25288
rect 7392 25248 7840 25276
rect 7392 25220 7420 25248
rect 7834 25236 7840 25248
rect 7892 25276 7898 25288
rect 8481 25279 8539 25285
rect 8481 25276 8493 25279
rect 7892 25248 8493 25276
rect 7892 25236 7898 25248
rect 8481 25245 8493 25248
rect 8527 25245 8539 25279
rect 8680 25276 8708 25375
rect 10597 25347 10655 25353
rect 10597 25313 10609 25347
rect 10643 25344 10655 25347
rect 10962 25344 10968 25356
rect 10643 25316 10968 25344
rect 10643 25313 10655 25316
rect 10597 25307 10655 25313
rect 10962 25304 10968 25316
rect 11020 25304 11026 25356
rect 11624 25353 11652 25452
rect 11790 25440 11796 25452
rect 11848 25440 11854 25492
rect 12161 25483 12219 25489
rect 12161 25449 12173 25483
rect 12207 25480 12219 25483
rect 12250 25480 12256 25492
rect 12207 25452 12256 25480
rect 12207 25449 12219 25452
rect 12161 25443 12219 25449
rect 12250 25440 12256 25452
rect 12308 25440 12314 25492
rect 13909 25483 13967 25489
rect 13909 25449 13921 25483
rect 13955 25480 13967 25483
rect 14734 25480 14740 25492
rect 13955 25452 14740 25480
rect 13955 25449 13967 25452
rect 13909 25443 13967 25449
rect 14734 25440 14740 25452
rect 14792 25440 14798 25492
rect 14918 25440 14924 25492
rect 14976 25480 14982 25492
rect 16577 25483 16635 25489
rect 16577 25480 16589 25483
rect 14976 25452 16589 25480
rect 14976 25440 14982 25452
rect 16577 25449 16589 25452
rect 16623 25449 16635 25483
rect 16577 25443 16635 25449
rect 17862 25440 17868 25492
rect 17920 25480 17926 25492
rect 19058 25480 19064 25492
rect 17920 25452 19064 25480
rect 17920 25440 17926 25452
rect 19058 25440 19064 25452
rect 19116 25440 19122 25492
rect 22462 25440 22468 25492
rect 22520 25480 22526 25492
rect 22557 25483 22615 25489
rect 22557 25480 22569 25483
rect 22520 25452 22569 25480
rect 22520 25440 22526 25452
rect 22557 25449 22569 25452
rect 22603 25480 22615 25483
rect 23014 25480 23020 25492
rect 22603 25452 23020 25480
rect 22603 25449 22615 25452
rect 22557 25443 22615 25449
rect 23014 25440 23020 25452
rect 23072 25440 23078 25492
rect 25038 25480 25044 25492
rect 23676 25452 25044 25480
rect 12986 25412 12992 25424
rect 12360 25384 12992 25412
rect 12360 25353 12388 25384
rect 12986 25372 12992 25384
rect 13044 25372 13050 25424
rect 13446 25412 13452 25424
rect 13407 25384 13452 25412
rect 13446 25372 13452 25384
rect 13504 25372 13510 25424
rect 14829 25415 14887 25421
rect 14829 25381 14841 25415
rect 14875 25381 14887 25415
rect 19245 25415 19303 25421
rect 19245 25412 19257 25415
rect 14829 25375 14887 25381
rect 15304 25384 19257 25412
rect 11609 25347 11667 25353
rect 11609 25313 11621 25347
rect 11655 25313 11667 25347
rect 11609 25307 11667 25313
rect 11977 25347 12035 25353
rect 11977 25313 11989 25347
rect 12023 25344 12035 25347
rect 12345 25347 12403 25353
rect 12345 25344 12357 25347
rect 12023 25316 12357 25344
rect 12023 25313 12035 25316
rect 11977 25307 12035 25313
rect 12345 25313 12357 25316
rect 12391 25313 12403 25347
rect 14844 25344 14872 25375
rect 12345 25307 12403 25313
rect 13004 25316 14872 25344
rect 9125 25279 9183 25285
rect 9125 25276 9137 25279
rect 8680 25248 9137 25276
rect 8481 25239 8539 25245
rect 9125 25245 9137 25248
rect 9171 25245 9183 25279
rect 9125 25239 9183 25245
rect 10321 25279 10379 25285
rect 10321 25245 10333 25279
rect 10367 25276 10379 25279
rect 10367 25248 11376 25276
rect 10367 25245 10379 25248
rect 10321 25239 10379 25245
rect 4157 25211 4215 25217
rect 4157 25208 4169 25211
rect 2976 25180 3740 25208
rect 3988 25180 4169 25208
rect 3988 25152 4016 25180
rect 4157 25177 4169 25180
rect 4203 25177 4215 25211
rect 4157 25171 4215 25177
rect 7374 25168 7380 25220
rect 7432 25168 7438 25220
rect 7466 25168 7472 25220
rect 7524 25208 7530 25220
rect 8113 25211 8171 25217
rect 8113 25208 8125 25211
rect 7524 25180 8125 25208
rect 7524 25168 7530 25180
rect 8113 25177 8125 25180
rect 8159 25177 8171 25211
rect 8113 25171 8171 25177
rect 8297 25211 8355 25217
rect 8297 25177 8309 25211
rect 8343 25208 8355 25211
rect 10870 25208 10876 25220
rect 8343 25180 10876 25208
rect 8343 25177 8355 25180
rect 8297 25171 8355 25177
rect 10870 25168 10876 25180
rect 10928 25168 10934 25220
rect 11348 25208 11376 25248
rect 12066 25236 12072 25288
rect 12124 25276 12130 25288
rect 12253 25279 12311 25285
rect 12253 25276 12265 25279
rect 12124 25248 12265 25276
rect 12124 25236 12130 25248
rect 12253 25245 12265 25248
rect 12299 25245 12311 25279
rect 12253 25239 12311 25245
rect 12710 25236 12716 25288
rect 12768 25276 12774 25288
rect 12897 25279 12955 25285
rect 12897 25276 12909 25279
rect 12768 25248 12909 25276
rect 12768 25236 12774 25248
rect 12897 25245 12909 25248
rect 12943 25245 12955 25279
rect 12897 25239 12955 25245
rect 13004 25208 13032 25316
rect 13262 25236 13268 25288
rect 13320 25285 13326 25288
rect 13320 25276 13328 25285
rect 13320 25248 13365 25276
rect 13320 25239 13328 25248
rect 13320 25236 13326 25239
rect 13630 25236 13636 25288
rect 13688 25276 13694 25288
rect 13725 25279 13783 25285
rect 13725 25276 13737 25279
rect 13688 25248 13737 25276
rect 13688 25236 13694 25248
rect 13725 25245 13737 25248
rect 13771 25245 13783 25279
rect 13725 25239 13783 25245
rect 14185 25279 14243 25285
rect 14185 25245 14197 25279
rect 14231 25276 14243 25279
rect 14274 25276 14280 25288
rect 14231 25248 14280 25276
rect 14231 25245 14243 25248
rect 14185 25239 14243 25245
rect 11348 25180 13032 25208
rect 13081 25211 13139 25217
rect 13081 25177 13093 25211
rect 13127 25177 13139 25211
rect 13081 25171 13139 25177
rect 13173 25211 13231 25217
rect 13173 25177 13185 25211
rect 13219 25208 13231 25211
rect 14200 25208 14228 25239
rect 14274 25236 14280 25248
rect 14332 25236 14338 25288
rect 15008 25279 15066 25285
rect 15008 25245 15020 25279
rect 15054 25276 15066 25279
rect 15304 25276 15332 25384
rect 19245 25381 19257 25384
rect 19291 25381 19303 25415
rect 23293 25415 23351 25421
rect 19245 25375 19303 25381
rect 19352 25384 19840 25412
rect 15396 25316 15700 25344
rect 15396 25285 15424 25316
rect 15054 25248 15332 25276
rect 15381 25279 15439 25285
rect 15054 25245 15066 25248
rect 15008 25239 15066 25245
rect 15381 25245 15393 25279
rect 15427 25245 15439 25279
rect 15562 25276 15568 25288
rect 15523 25248 15568 25276
rect 15381 25239 15439 25245
rect 15562 25236 15568 25248
rect 15620 25236 15626 25288
rect 15102 25208 15108 25220
rect 13219 25180 14228 25208
rect 15063 25180 15108 25208
rect 13219 25177 13231 25180
rect 13173 25171 13231 25177
rect 3970 25100 3976 25152
rect 4028 25100 4034 25152
rect 6822 25140 6828 25152
rect 6783 25112 6828 25140
rect 6822 25100 6828 25112
rect 6880 25100 6886 25152
rect 7193 25143 7251 25149
rect 7193 25109 7205 25143
rect 7239 25140 7251 25143
rect 8386 25140 8392 25152
rect 7239 25112 8392 25140
rect 7239 25109 7251 25112
rect 7193 25103 7251 25109
rect 8386 25100 8392 25112
rect 8444 25100 8450 25152
rect 8754 25100 8760 25152
rect 8812 25140 8818 25152
rect 8941 25143 8999 25149
rect 8941 25140 8953 25143
rect 8812 25112 8953 25140
rect 8812 25100 8818 25112
rect 8941 25109 8953 25112
rect 8987 25109 8999 25143
rect 8941 25103 8999 25109
rect 10318 25100 10324 25152
rect 10376 25140 10382 25152
rect 10413 25143 10471 25149
rect 10413 25140 10425 25143
rect 10376 25112 10425 25140
rect 10376 25100 10382 25112
rect 10413 25109 10425 25112
rect 10459 25109 10471 25143
rect 11790 25140 11796 25152
rect 11751 25112 11796 25140
rect 10413 25103 10471 25109
rect 11790 25100 11796 25112
rect 11848 25100 11854 25152
rect 12618 25140 12624 25152
rect 12579 25112 12624 25140
rect 12618 25100 12624 25112
rect 12676 25100 12682 25152
rect 12802 25100 12808 25152
rect 12860 25140 12866 25152
rect 13096 25140 13124 25171
rect 15102 25168 15108 25180
rect 15160 25168 15166 25220
rect 15197 25211 15255 25217
rect 15197 25177 15209 25211
rect 15243 25208 15255 25211
rect 15580 25208 15608 25236
rect 15243 25180 15608 25208
rect 15243 25177 15255 25180
rect 15197 25171 15255 25177
rect 14369 25143 14427 25149
rect 14369 25140 14381 25143
rect 12860 25112 14381 25140
rect 12860 25100 12866 25112
rect 14369 25109 14381 25112
rect 14415 25140 14427 25143
rect 14642 25140 14648 25152
rect 14415 25112 14648 25140
rect 14415 25109 14427 25112
rect 14369 25103 14427 25109
rect 14642 25100 14648 25112
rect 14700 25100 14706 25152
rect 14826 25100 14832 25152
rect 14884 25140 14890 25152
rect 15672 25140 15700 25316
rect 16758 25304 16764 25356
rect 16816 25344 16822 25356
rect 17037 25347 17095 25353
rect 17037 25344 17049 25347
rect 16816 25316 17049 25344
rect 16816 25304 16822 25316
rect 17037 25313 17049 25316
rect 17083 25313 17095 25347
rect 17037 25307 17095 25313
rect 17126 25304 17132 25356
rect 17184 25344 17190 25356
rect 18417 25347 18475 25353
rect 18417 25344 18429 25347
rect 17184 25316 18429 25344
rect 17184 25304 17190 25316
rect 18417 25313 18429 25316
rect 18463 25344 18475 25347
rect 19352 25344 19380 25384
rect 18463 25316 19380 25344
rect 18463 25313 18475 25316
rect 18417 25307 18475 25313
rect 19426 25304 19432 25356
rect 19484 25344 19490 25356
rect 19812 25353 19840 25384
rect 23293 25381 23305 25415
rect 23339 25381 23351 25415
rect 23293 25375 23351 25381
rect 19705 25347 19763 25353
rect 19705 25344 19717 25347
rect 19484 25316 19717 25344
rect 19484 25304 19490 25316
rect 19705 25313 19717 25316
rect 19751 25313 19763 25347
rect 19705 25307 19763 25313
rect 19797 25347 19855 25353
rect 19797 25313 19809 25347
rect 19843 25313 19855 25347
rect 19797 25307 19855 25313
rect 20254 25304 20260 25356
rect 20312 25344 20318 25356
rect 20809 25347 20867 25353
rect 20809 25344 20821 25347
rect 20312 25316 20821 25344
rect 20312 25304 20318 25316
rect 20809 25313 20821 25316
rect 20855 25313 20867 25347
rect 23308 25344 23336 25375
rect 20809 25307 20867 25313
rect 22480 25316 23336 25344
rect 16298 25236 16304 25288
rect 16356 25276 16362 25288
rect 16485 25279 16543 25285
rect 16485 25276 16497 25279
rect 16356 25248 16497 25276
rect 16356 25236 16362 25248
rect 16485 25245 16497 25248
rect 16531 25245 16543 25279
rect 16485 25239 16543 25245
rect 18325 25279 18383 25285
rect 18325 25245 18337 25279
rect 18371 25276 18383 25279
rect 19518 25276 19524 25288
rect 18371 25248 19524 25276
rect 18371 25245 18383 25248
rect 18325 25239 18383 25245
rect 19518 25236 19524 25248
rect 19576 25236 19582 25288
rect 20346 25276 20352 25288
rect 20259 25248 20352 25276
rect 15746 25168 15752 25220
rect 15804 25208 15810 25220
rect 19334 25208 19340 25220
rect 15804 25180 19340 25208
rect 15804 25168 15810 25180
rect 16316 25149 16344 25180
rect 19334 25168 19340 25180
rect 19392 25168 19398 25220
rect 14884 25112 15700 25140
rect 16301 25143 16359 25149
rect 14884 25100 14890 25112
rect 16301 25109 16313 25143
rect 16347 25109 16359 25143
rect 16942 25140 16948 25152
rect 16903 25112 16948 25140
rect 16301 25103 16359 25109
rect 16942 25100 16948 25112
rect 17000 25100 17006 25152
rect 17034 25100 17040 25152
rect 17092 25140 17098 25152
rect 17865 25143 17923 25149
rect 17865 25140 17877 25143
rect 17092 25112 17877 25140
rect 17092 25100 17098 25112
rect 17865 25109 17877 25112
rect 17911 25109 17923 25143
rect 18230 25140 18236 25152
rect 18191 25112 18236 25140
rect 17865 25103 17923 25109
rect 18230 25100 18236 25112
rect 18288 25100 18294 25152
rect 19518 25100 19524 25152
rect 19576 25140 19582 25152
rect 19613 25143 19671 25149
rect 19613 25140 19625 25143
rect 19576 25112 19625 25140
rect 19576 25100 19582 25112
rect 19613 25109 19625 25112
rect 19659 25109 19671 25143
rect 19613 25103 19671 25109
rect 19702 25100 19708 25152
rect 19760 25140 19766 25152
rect 20272 25149 20300 25248
rect 20346 25236 20352 25248
rect 20404 25276 20410 25288
rect 20441 25279 20499 25285
rect 20441 25276 20453 25279
rect 20404 25248 20453 25276
rect 20404 25236 20410 25248
rect 20441 25245 20453 25248
rect 20487 25245 20499 25279
rect 20441 25239 20499 25245
rect 21085 25211 21143 25217
rect 21085 25177 21097 25211
rect 21131 25177 21143 25211
rect 21085 25171 21143 25177
rect 20257 25143 20315 25149
rect 20257 25140 20269 25143
rect 19760 25112 20269 25140
rect 19760 25100 19766 25112
rect 20257 25109 20269 25112
rect 20303 25109 20315 25143
rect 20622 25140 20628 25152
rect 20583 25112 20628 25140
rect 20257 25103 20315 25109
rect 20622 25100 20628 25112
rect 20680 25100 20686 25152
rect 21100 25140 21128 25171
rect 21818 25168 21824 25220
rect 21876 25168 21882 25220
rect 22480 25140 22508 25316
rect 22738 25276 22744 25288
rect 22699 25248 22744 25276
rect 22738 25236 22744 25248
rect 22796 25236 22802 25288
rect 22830 25236 22836 25288
rect 22888 25276 22894 25288
rect 23114 25279 23172 25285
rect 23114 25276 23126 25279
rect 22888 25248 23126 25276
rect 22888 25236 22894 25248
rect 23114 25245 23126 25248
rect 23160 25245 23172 25279
rect 23114 25239 23172 25245
rect 23477 25279 23535 25285
rect 23477 25245 23489 25279
rect 23523 25276 23535 25279
rect 23676 25276 23704 25452
rect 25038 25440 25044 25452
rect 25096 25440 25102 25492
rect 25222 25480 25228 25492
rect 25183 25452 25228 25480
rect 25222 25440 25228 25452
rect 25280 25440 25286 25492
rect 26053 25483 26111 25489
rect 26053 25449 26065 25483
rect 26099 25480 26111 25483
rect 27154 25480 27160 25492
rect 26099 25452 27160 25480
rect 26099 25449 26111 25452
rect 26053 25443 26111 25449
rect 27154 25440 27160 25452
rect 27212 25440 27218 25492
rect 24026 25412 24032 25424
rect 23987 25384 24032 25412
rect 24026 25372 24032 25384
rect 24084 25372 24090 25424
rect 24581 25415 24639 25421
rect 24581 25412 24593 25415
rect 24504 25384 24593 25412
rect 23750 25304 23756 25356
rect 23808 25344 23814 25356
rect 23808 25316 23893 25344
rect 23808 25304 23814 25316
rect 23865 25285 23893 25316
rect 23523 25248 23704 25276
rect 23850 25279 23908 25285
rect 23523 25245 23535 25248
rect 23477 25239 23535 25245
rect 23850 25245 23862 25279
rect 23896 25276 23908 25279
rect 24213 25279 24271 25285
rect 24213 25276 24225 25279
rect 23896 25248 24225 25276
rect 23896 25245 23908 25248
rect 23850 25239 23908 25245
rect 24213 25245 24225 25248
rect 24259 25245 24271 25279
rect 24394 25276 24400 25288
rect 24355 25248 24400 25276
rect 24213 25239 24271 25245
rect 24394 25236 24400 25248
rect 24452 25236 24458 25288
rect 24504 25276 24532 25384
rect 24581 25381 24593 25384
rect 24627 25381 24639 25415
rect 24581 25375 24639 25381
rect 24670 25372 24676 25424
rect 24728 25412 24734 25424
rect 25056 25412 25084 25440
rect 25774 25412 25780 25424
rect 24728 25384 24773 25412
rect 25056 25384 25780 25412
rect 24728 25372 24734 25384
rect 25774 25372 25780 25384
rect 25832 25372 25838 25424
rect 27062 25344 27068 25356
rect 25516 25316 27068 25344
rect 25516 25285 25544 25316
rect 27062 25304 27068 25316
rect 27120 25304 27126 25356
rect 24857 25279 24915 25285
rect 24857 25276 24869 25279
rect 24504 25248 24869 25276
rect 24857 25245 24869 25248
rect 24903 25245 24915 25279
rect 25380 25279 25438 25285
rect 25380 25276 25392 25279
rect 24857 25239 24915 25245
rect 25378 25245 25392 25276
rect 25426 25245 25438 25279
rect 25378 25239 25438 25245
rect 25501 25279 25559 25285
rect 25501 25245 25513 25279
rect 25547 25245 25559 25279
rect 25774 25276 25780 25288
rect 25735 25248 25780 25276
rect 25501 25239 25559 25245
rect 22646 25168 22652 25220
rect 22704 25208 22710 25220
rect 22925 25211 22983 25217
rect 22925 25208 22937 25211
rect 22704 25180 22937 25208
rect 22704 25168 22710 25180
rect 22925 25177 22937 25180
rect 22971 25177 22983 25211
rect 22925 25171 22983 25177
rect 23014 25168 23020 25220
rect 23072 25208 23078 25220
rect 23072 25180 23117 25208
rect 23072 25168 23078 25180
rect 23382 25168 23388 25220
rect 23440 25208 23446 25220
rect 23661 25211 23719 25217
rect 23661 25208 23673 25211
rect 23440 25180 23673 25208
rect 23440 25168 23446 25180
rect 23661 25177 23673 25180
rect 23707 25177 23719 25211
rect 23661 25171 23719 25177
rect 21100 25112 22508 25140
rect 23676 25140 23704 25171
rect 23750 25168 23756 25220
rect 23808 25208 23814 25220
rect 24949 25211 25007 25217
rect 24949 25208 24961 25211
rect 23808 25180 23853 25208
rect 23952 25180 24961 25208
rect 23808 25168 23814 25180
rect 23952 25140 23980 25180
rect 24949 25177 24961 25180
rect 24995 25177 25007 25211
rect 24949 25171 25007 25177
rect 23676 25112 23980 25140
rect 24213 25143 24271 25149
rect 24213 25109 24225 25143
rect 24259 25140 24271 25143
rect 25378 25140 25406 25239
rect 25774 25236 25780 25248
rect 25832 25236 25838 25288
rect 25866 25236 25872 25288
rect 25924 25276 25930 25288
rect 25924 25248 25969 25276
rect 25924 25236 25930 25248
rect 25590 25208 25596 25220
rect 25503 25180 25596 25208
rect 25590 25168 25596 25180
rect 25648 25208 25654 25220
rect 26145 25211 26203 25217
rect 26145 25208 26157 25211
rect 25648 25180 26157 25208
rect 25648 25168 25654 25180
rect 26145 25177 26157 25180
rect 26191 25177 26203 25211
rect 26145 25171 26203 25177
rect 25682 25140 25688 25152
rect 24259 25112 25688 25140
rect 24259 25109 24271 25112
rect 24213 25103 24271 25109
rect 25682 25100 25688 25112
rect 25740 25100 25746 25152
rect 1104 25050 29440 25072
rect 1104 24998 10395 25050
rect 10447 24998 10459 25050
rect 10511 24998 10523 25050
rect 10575 24998 10587 25050
rect 10639 24998 10651 25050
rect 10703 24998 19840 25050
rect 19892 24998 19904 25050
rect 19956 24998 19968 25050
rect 20020 24998 20032 25050
rect 20084 24998 20096 25050
rect 20148 24998 29440 25050
rect 1104 24976 29440 24998
rect 7193 24939 7251 24945
rect 7193 24905 7205 24939
rect 7239 24905 7251 24939
rect 7193 24899 7251 24905
rect 2774 24828 2780 24880
rect 2832 24868 2838 24880
rect 2961 24871 3019 24877
rect 2961 24868 2973 24871
rect 2832 24840 2973 24868
rect 2832 24828 2838 24840
rect 2961 24837 2973 24840
rect 3007 24837 3019 24871
rect 2961 24831 3019 24837
rect 2685 24803 2743 24809
rect 2685 24769 2697 24803
rect 2731 24769 2743 24803
rect 2866 24800 2872 24812
rect 2827 24772 2872 24800
rect 2685 24763 2743 24769
rect 2700 24732 2728 24763
rect 2866 24760 2872 24772
rect 2924 24760 2930 24812
rect 4433 24803 4491 24809
rect 4433 24769 4445 24803
rect 4479 24800 4491 24803
rect 4706 24800 4712 24812
rect 4479 24772 4712 24800
rect 4479 24769 4491 24772
rect 4433 24763 4491 24769
rect 4706 24760 4712 24772
rect 4764 24760 4770 24812
rect 4801 24803 4859 24809
rect 4801 24769 4813 24803
rect 4847 24800 4859 24803
rect 4890 24800 4896 24812
rect 4847 24772 4896 24800
rect 4847 24769 4859 24772
rect 4801 24763 4859 24769
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 6917 24803 6975 24809
rect 6917 24769 6929 24803
rect 6963 24800 6975 24803
rect 7208 24800 7236 24899
rect 8386 24896 8392 24948
rect 8444 24936 8450 24948
rect 9214 24936 9220 24948
rect 8444 24908 9220 24936
rect 8444 24896 8450 24908
rect 9214 24896 9220 24908
rect 9272 24896 9278 24948
rect 9677 24939 9735 24945
rect 9677 24905 9689 24939
rect 9723 24936 9735 24939
rect 10321 24939 10379 24945
rect 10321 24936 10333 24939
rect 9723 24908 10333 24936
rect 9723 24905 9735 24908
rect 9677 24899 9735 24905
rect 10321 24905 10333 24908
rect 10367 24905 10379 24939
rect 10873 24939 10931 24945
rect 10873 24936 10885 24939
rect 10321 24899 10379 24905
rect 10520 24908 10885 24936
rect 7742 24868 7748 24880
rect 7703 24840 7748 24868
rect 7742 24828 7748 24840
rect 7800 24828 7806 24880
rect 8754 24828 8760 24880
rect 8812 24828 8818 24880
rect 10229 24871 10287 24877
rect 10229 24837 10241 24871
rect 10275 24868 10287 24871
rect 10410 24868 10416 24880
rect 10275 24840 10416 24868
rect 10275 24837 10287 24840
rect 10229 24831 10287 24837
rect 10410 24828 10416 24840
rect 10468 24828 10474 24880
rect 7374 24800 7380 24812
rect 6963 24772 7236 24800
rect 7335 24772 7380 24800
rect 6963 24769 6975 24772
rect 6917 24763 6975 24769
rect 7374 24760 7380 24772
rect 7432 24760 7438 24812
rect 9585 24803 9643 24809
rect 9585 24769 9597 24803
rect 9631 24769 9643 24803
rect 9766 24800 9772 24812
rect 9727 24772 9772 24800
rect 9585 24763 9643 24769
rect 3234 24732 3240 24744
rect 2700 24704 3240 24732
rect 3234 24692 3240 24704
rect 3292 24692 3298 24744
rect 5166 24692 5172 24744
rect 5224 24732 5230 24744
rect 7466 24732 7472 24744
rect 5224 24704 7472 24732
rect 5224 24692 5230 24704
rect 6932 24676 6960 24704
rect 7466 24692 7472 24704
rect 7524 24692 7530 24744
rect 9600 24732 9628 24763
rect 9766 24760 9772 24772
rect 9824 24800 9830 24812
rect 10520 24800 10548 24908
rect 10873 24905 10885 24908
rect 10919 24905 10931 24939
rect 15573 24939 15631 24945
rect 15573 24936 15585 24939
rect 10873 24899 10931 24905
rect 12406 24908 15585 24936
rect 10594 24828 10600 24880
rect 10652 24868 10658 24880
rect 12406 24868 12434 24908
rect 15573 24905 15585 24908
rect 15619 24905 15631 24939
rect 15573 24899 15631 24905
rect 18049 24939 18107 24945
rect 18049 24905 18061 24939
rect 18095 24936 18107 24939
rect 18966 24936 18972 24948
rect 18095 24908 18972 24936
rect 18095 24905 18107 24908
rect 18049 24899 18107 24905
rect 18966 24896 18972 24908
rect 19024 24896 19030 24948
rect 22002 24936 22008 24948
rect 21963 24908 22008 24936
rect 22002 24896 22008 24908
rect 22060 24896 22066 24948
rect 23290 24936 23296 24948
rect 23251 24908 23296 24936
rect 23290 24896 23296 24908
rect 23348 24896 23354 24948
rect 24394 24936 24400 24948
rect 23492 24908 24400 24936
rect 10652 24840 12434 24868
rect 10652 24828 10658 24840
rect 12526 24828 12532 24880
rect 12584 24868 12590 24880
rect 13262 24868 13268 24880
rect 12584 24840 13268 24868
rect 12584 24828 12590 24840
rect 13262 24828 13268 24840
rect 13320 24828 13326 24880
rect 13357 24871 13415 24877
rect 13357 24837 13369 24871
rect 13403 24868 13415 24871
rect 13446 24868 13452 24880
rect 13403 24840 13452 24868
rect 13403 24837 13415 24840
rect 13357 24831 13415 24837
rect 13446 24828 13452 24840
rect 13504 24828 13510 24880
rect 14366 24828 14372 24880
rect 14424 24828 14430 24880
rect 14642 24828 14648 24880
rect 14700 24868 14706 24880
rect 14700 24840 15240 24868
rect 14700 24828 14706 24840
rect 9824 24772 10548 24800
rect 10689 24803 10747 24809
rect 9824 24760 9830 24772
rect 10689 24769 10701 24803
rect 10735 24800 10747 24803
rect 10778 24800 10784 24812
rect 10735 24772 10784 24800
rect 10735 24769 10747 24772
rect 10689 24763 10747 24769
rect 10778 24760 10784 24772
rect 10836 24800 10842 24812
rect 12158 24800 12164 24812
rect 10836 24772 11836 24800
rect 12119 24772 12164 24800
rect 10836 24760 10842 24772
rect 10134 24732 10140 24744
rect 9600 24704 10140 24732
rect 10134 24692 10140 24704
rect 10192 24692 10198 24744
rect 10505 24735 10563 24741
rect 10505 24701 10517 24735
rect 10551 24732 10563 24735
rect 10962 24732 10968 24744
rect 10551 24704 10968 24732
rect 10551 24701 10563 24704
rect 10505 24695 10563 24701
rect 10962 24692 10968 24704
rect 11020 24692 11026 24744
rect 11057 24735 11115 24741
rect 11057 24701 11069 24735
rect 11103 24732 11115 24735
rect 11514 24732 11520 24744
rect 11103 24704 11520 24732
rect 11103 24701 11115 24704
rect 11057 24695 11115 24701
rect 11514 24692 11520 24704
rect 11572 24692 11578 24744
rect 11808 24741 11836 24772
rect 12158 24760 12164 24772
rect 12216 24800 12222 24812
rect 12253 24803 12311 24809
rect 12253 24800 12265 24803
rect 12216 24772 12265 24800
rect 12216 24760 12222 24772
rect 12253 24769 12265 24772
rect 12299 24769 12311 24803
rect 12253 24763 12311 24769
rect 12345 24803 12403 24809
rect 12345 24769 12357 24803
rect 12391 24800 12403 24803
rect 12710 24800 12716 24812
rect 12391 24772 12716 24800
rect 12391 24769 12403 24772
rect 12345 24763 12403 24769
rect 12710 24760 12716 24772
rect 12768 24760 12774 24812
rect 14826 24760 14832 24812
rect 14884 24800 14890 24812
rect 15212 24809 15240 24840
rect 15286 24828 15292 24880
rect 15344 24868 15350 24880
rect 16114 24868 16120 24880
rect 15344 24840 16120 24868
rect 15344 24828 15350 24840
rect 16114 24828 16120 24840
rect 16172 24828 16178 24880
rect 18601 24871 18659 24877
rect 18601 24837 18613 24871
rect 18647 24868 18659 24871
rect 18874 24868 18880 24880
rect 18647 24840 18880 24868
rect 18647 24837 18659 24840
rect 18601 24831 18659 24837
rect 18874 24828 18880 24840
rect 18932 24828 18938 24880
rect 19705 24871 19763 24877
rect 19705 24837 19717 24871
rect 19751 24868 19763 24871
rect 20254 24868 20260 24880
rect 19751 24840 20260 24868
rect 19751 24837 19763 24840
rect 19705 24831 19763 24837
rect 20254 24828 20260 24840
rect 20312 24828 20318 24880
rect 20622 24868 20628 24880
rect 20535 24840 20628 24868
rect 15013 24803 15071 24809
rect 15013 24800 15025 24803
rect 14884 24772 15025 24800
rect 14884 24760 14890 24772
rect 15013 24769 15025 24772
rect 15059 24769 15071 24803
rect 15013 24763 15071 24769
rect 15197 24803 15255 24809
rect 15197 24769 15209 24803
rect 15243 24769 15255 24803
rect 15197 24763 15255 24769
rect 15433 24803 15491 24809
rect 15433 24769 15445 24803
rect 15479 24800 15491 24803
rect 17034 24800 17040 24812
rect 15479 24772 17040 24800
rect 15479 24769 15491 24772
rect 15433 24763 15491 24769
rect 11793 24735 11851 24741
rect 11793 24701 11805 24735
rect 11839 24732 11851 24735
rect 12802 24732 12808 24744
rect 11839 24704 12808 24732
rect 11839 24701 11851 24704
rect 11793 24695 11851 24701
rect 12802 24692 12808 24704
rect 12860 24692 12866 24744
rect 13078 24732 13084 24744
rect 13039 24704 13084 24732
rect 13078 24692 13084 24704
rect 13136 24692 13142 24744
rect 15212 24732 15240 24763
rect 17034 24760 17040 24772
rect 17092 24760 17098 24812
rect 20548 24809 20576 24840
rect 20622 24828 20628 24840
rect 20680 24868 20686 24880
rect 23492 24868 23520 24908
rect 24394 24896 24400 24908
rect 24452 24936 24458 24948
rect 25866 24936 25872 24948
rect 24452 24908 25872 24936
rect 24452 24896 24458 24908
rect 25866 24896 25872 24908
rect 25924 24896 25930 24948
rect 24670 24868 24676 24880
rect 20680 24840 23520 24868
rect 24334 24840 24676 24868
rect 20680 24828 20686 24840
rect 24670 24828 24676 24840
rect 24728 24828 24734 24880
rect 25501 24871 25559 24877
rect 25501 24837 25513 24871
rect 25547 24868 25559 24871
rect 26694 24868 26700 24880
rect 25547 24840 26700 24868
rect 25547 24837 25559 24840
rect 25501 24831 25559 24837
rect 26694 24828 26700 24840
rect 26752 24828 26758 24880
rect 17865 24803 17923 24809
rect 17865 24769 17877 24803
rect 17911 24800 17923 24803
rect 20533 24803 20591 24809
rect 17911 24772 18000 24800
rect 17911 24769 17923 24772
rect 17865 24763 17923 24769
rect 15212 24704 15884 24732
rect 4062 24624 4068 24676
rect 4120 24664 4126 24676
rect 4249 24667 4307 24673
rect 4249 24664 4261 24667
rect 4120 24636 4261 24664
rect 4120 24624 4126 24636
rect 4249 24633 4261 24636
rect 4295 24664 4307 24667
rect 6086 24664 6092 24676
rect 4295 24636 6092 24664
rect 4295 24633 4307 24636
rect 4249 24627 4307 24633
rect 6086 24624 6092 24636
rect 6144 24624 6150 24676
rect 6914 24624 6920 24676
rect 6972 24624 6978 24676
rect 12618 24664 12624 24676
rect 11256 24636 12624 24664
rect 2501 24599 2559 24605
rect 2501 24565 2513 24599
rect 2547 24596 2559 24599
rect 2590 24596 2596 24608
rect 2547 24568 2596 24596
rect 2547 24565 2559 24568
rect 2501 24559 2559 24565
rect 2590 24556 2596 24568
rect 2648 24556 2654 24608
rect 4338 24556 4344 24608
rect 4396 24596 4402 24608
rect 4617 24599 4675 24605
rect 4617 24596 4629 24599
rect 4396 24568 4629 24596
rect 4396 24556 4402 24568
rect 4617 24565 4629 24568
rect 4663 24565 4675 24599
rect 4617 24559 4675 24565
rect 7101 24599 7159 24605
rect 7101 24565 7113 24599
rect 7147 24596 7159 24599
rect 7282 24596 7288 24608
rect 7147 24568 7288 24596
rect 7147 24565 7159 24568
rect 7101 24559 7159 24565
rect 7282 24556 7288 24568
rect 7340 24556 7346 24608
rect 9490 24556 9496 24608
rect 9548 24596 9554 24608
rect 9861 24599 9919 24605
rect 9861 24596 9873 24599
rect 9548 24568 9873 24596
rect 9548 24556 9554 24568
rect 9861 24565 9873 24568
rect 9907 24565 9919 24599
rect 9861 24559 9919 24565
rect 10410 24556 10416 24608
rect 10468 24596 10474 24608
rect 11256 24605 11284 24636
rect 12618 24624 12624 24636
rect 12676 24624 12682 24676
rect 12894 24664 12900 24676
rect 12855 24636 12900 24664
rect 12894 24624 12900 24636
rect 12952 24624 12958 24676
rect 15856 24608 15884 24704
rect 11241 24599 11299 24605
rect 11241 24596 11253 24599
rect 10468 24568 11253 24596
rect 10468 24556 10474 24568
rect 11241 24565 11253 24568
rect 11287 24565 11299 24599
rect 11514 24596 11520 24608
rect 11475 24568 11520 24596
rect 11241 24559 11299 24565
rect 11514 24556 11520 24568
rect 11572 24556 11578 24608
rect 11977 24599 12035 24605
rect 11977 24565 11989 24599
rect 12023 24596 12035 24599
rect 12434 24596 12440 24608
rect 12023 24568 12440 24596
rect 12023 24565 12035 24568
rect 11977 24559 12035 24565
rect 12434 24556 12440 24568
rect 12492 24556 12498 24608
rect 12529 24599 12587 24605
rect 12529 24565 12541 24599
rect 12575 24596 12587 24599
rect 12986 24596 12992 24608
rect 12575 24568 12992 24596
rect 12575 24565 12587 24568
rect 12529 24559 12587 24565
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 14366 24556 14372 24608
rect 14424 24596 14430 24608
rect 14829 24599 14887 24605
rect 14829 24596 14841 24599
rect 14424 24568 14841 24596
rect 14424 24556 14430 24568
rect 14829 24565 14841 24568
rect 14875 24565 14887 24599
rect 15838 24596 15844 24608
rect 15799 24568 15844 24596
rect 14829 24559 14887 24565
rect 15838 24556 15844 24568
rect 15896 24556 15902 24608
rect 16298 24556 16304 24608
rect 16356 24596 16362 24608
rect 17972 24596 18000 24772
rect 18800 24772 19932 24800
rect 18800 24744 18828 24772
rect 18046 24692 18052 24744
rect 18104 24732 18110 24744
rect 18104 24704 18276 24732
rect 18104 24692 18110 24704
rect 18248 24673 18276 24704
rect 18322 24692 18328 24744
rect 18380 24732 18386 24744
rect 18693 24735 18751 24741
rect 18693 24732 18705 24735
rect 18380 24704 18705 24732
rect 18380 24692 18386 24704
rect 18693 24701 18705 24704
rect 18739 24701 18751 24735
rect 18693 24695 18751 24701
rect 18782 24692 18788 24744
rect 18840 24732 18846 24744
rect 18840 24704 18885 24732
rect 18840 24692 18846 24704
rect 19702 24692 19708 24744
rect 19760 24732 19766 24744
rect 19904 24741 19932 24772
rect 20533 24769 20545 24803
rect 20579 24769 20591 24803
rect 20533 24763 20591 24769
rect 21085 24803 21143 24809
rect 21085 24769 21097 24803
rect 21131 24769 21143 24803
rect 21085 24763 21143 24769
rect 19797 24735 19855 24741
rect 19797 24732 19809 24735
rect 19760 24704 19809 24732
rect 19760 24692 19766 24704
rect 19797 24701 19809 24704
rect 19843 24701 19855 24735
rect 19797 24695 19855 24701
rect 19889 24735 19947 24741
rect 19889 24701 19901 24735
rect 19935 24701 19947 24735
rect 19889 24695 19947 24701
rect 18233 24667 18291 24673
rect 18233 24633 18245 24667
rect 18279 24633 18291 24667
rect 19150 24664 19156 24676
rect 18233 24627 18291 24633
rect 18340 24636 19156 24664
rect 18340 24596 18368 24636
rect 19150 24624 19156 24636
rect 19208 24624 19214 24676
rect 19242 24624 19248 24676
rect 19300 24664 19306 24676
rect 21100 24664 21128 24763
rect 21726 24760 21732 24812
rect 21784 24800 21790 24812
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 21784 24772 21833 24800
rect 21784 24760 21790 24772
rect 21821 24769 21833 24772
rect 21867 24800 21879 24803
rect 22097 24803 22155 24809
rect 22097 24800 22109 24803
rect 21867 24772 22109 24800
rect 21867 24769 21879 24772
rect 21821 24763 21879 24769
rect 22097 24769 22109 24772
rect 22143 24769 22155 24803
rect 22097 24763 22155 24769
rect 25130 24760 25136 24812
rect 25188 24800 25194 24812
rect 25682 24809 25688 24812
rect 25225 24803 25283 24809
rect 25225 24800 25237 24803
rect 25188 24772 25237 24800
rect 25188 24760 25194 24772
rect 25225 24769 25237 24772
rect 25271 24769 25283 24803
rect 25409 24803 25467 24809
rect 25409 24800 25421 24803
rect 25225 24763 25283 24769
rect 25332 24772 25421 24800
rect 24026 24692 24032 24744
rect 24084 24732 24090 24744
rect 24765 24735 24823 24741
rect 24765 24732 24777 24735
rect 24084 24704 24777 24732
rect 24084 24692 24090 24704
rect 24765 24701 24777 24704
rect 24811 24701 24823 24735
rect 25038 24732 25044 24744
rect 24999 24704 25044 24732
rect 24765 24695 24823 24701
rect 25038 24692 25044 24704
rect 25096 24692 25102 24744
rect 19300 24636 21128 24664
rect 25332 24664 25360 24772
rect 25409 24769 25421 24772
rect 25455 24769 25467 24803
rect 25409 24763 25467 24769
rect 25645 24803 25688 24809
rect 25645 24769 25657 24803
rect 25645 24763 25688 24769
rect 25682 24760 25688 24763
rect 25740 24760 25746 24812
rect 25866 24760 25872 24812
rect 25924 24800 25930 24812
rect 26053 24803 26111 24809
rect 26053 24800 26065 24803
rect 25924 24772 26065 24800
rect 25924 24760 25930 24772
rect 26053 24769 26065 24772
rect 26099 24769 26111 24803
rect 26329 24803 26387 24809
rect 26329 24800 26341 24803
rect 26053 24763 26111 24769
rect 26252 24772 26341 24800
rect 26252 24673 26280 24772
rect 26329 24769 26341 24772
rect 26375 24769 26387 24803
rect 26329 24763 26387 24769
rect 26237 24667 26295 24673
rect 25332 24636 25912 24664
rect 19300 24624 19306 24636
rect 16356 24568 18368 24596
rect 16356 24556 16362 24568
rect 19058 24556 19064 24608
rect 19116 24596 19122 24608
rect 19337 24599 19395 24605
rect 19337 24596 19349 24599
rect 19116 24568 19349 24596
rect 19116 24556 19122 24568
rect 19337 24565 19349 24568
rect 19383 24565 19395 24599
rect 19337 24559 19395 24565
rect 20717 24599 20775 24605
rect 20717 24565 20729 24599
rect 20763 24596 20775 24599
rect 20898 24596 20904 24608
rect 20763 24568 20904 24596
rect 20763 24565 20775 24568
rect 20717 24559 20775 24565
rect 20898 24556 20904 24568
rect 20956 24556 20962 24608
rect 20990 24556 20996 24608
rect 21048 24596 21054 24608
rect 21177 24599 21235 24605
rect 21177 24596 21189 24599
rect 21048 24568 21189 24596
rect 21048 24556 21054 24568
rect 21177 24565 21189 24568
rect 21223 24596 21235 24599
rect 21266 24596 21272 24608
rect 21223 24568 21272 24596
rect 21223 24565 21235 24568
rect 21177 24559 21235 24565
rect 21266 24556 21272 24568
rect 21324 24556 21330 24608
rect 24118 24556 24124 24608
rect 24176 24596 24182 24608
rect 25332 24596 25360 24636
rect 25774 24596 25780 24608
rect 24176 24568 25360 24596
rect 25735 24568 25780 24596
rect 24176 24556 24182 24568
rect 25774 24556 25780 24568
rect 25832 24556 25838 24608
rect 25884 24596 25912 24636
rect 26237 24633 26249 24667
rect 26283 24633 26295 24667
rect 26973 24667 27031 24673
rect 26973 24664 26985 24667
rect 26237 24627 26295 24633
rect 26344 24636 26985 24664
rect 26344 24596 26372 24636
rect 26973 24633 26985 24636
rect 27019 24633 27031 24667
rect 26973 24627 27031 24633
rect 26510 24596 26516 24608
rect 25884 24568 26372 24596
rect 26471 24568 26516 24596
rect 26510 24556 26516 24568
rect 26568 24556 26574 24608
rect 26694 24596 26700 24608
rect 26655 24568 26700 24596
rect 26694 24556 26700 24568
rect 26752 24556 26758 24608
rect 1104 24506 29440 24528
rect 1104 24454 5672 24506
rect 5724 24454 5736 24506
rect 5788 24454 5800 24506
rect 5852 24454 5864 24506
rect 5916 24454 5928 24506
rect 5980 24454 15118 24506
rect 15170 24454 15182 24506
rect 15234 24454 15246 24506
rect 15298 24454 15310 24506
rect 15362 24454 15374 24506
rect 15426 24454 24563 24506
rect 24615 24454 24627 24506
rect 24679 24454 24691 24506
rect 24743 24454 24755 24506
rect 24807 24454 24819 24506
rect 24871 24454 29440 24506
rect 1104 24432 29440 24454
rect 2777 24395 2835 24401
rect 2777 24361 2789 24395
rect 2823 24392 2835 24395
rect 2866 24392 2872 24404
rect 2823 24364 2872 24392
rect 2823 24361 2835 24364
rect 2777 24355 2835 24361
rect 2866 24352 2872 24364
rect 2924 24352 2930 24404
rect 4706 24392 4712 24404
rect 4667 24364 4712 24392
rect 4706 24352 4712 24364
rect 4764 24352 4770 24404
rect 10597 24395 10655 24401
rect 10597 24361 10609 24395
rect 10643 24392 10655 24395
rect 10778 24392 10784 24404
rect 10643 24364 10784 24392
rect 10643 24361 10655 24364
rect 10597 24355 10655 24361
rect 10778 24352 10784 24364
rect 10836 24352 10842 24404
rect 10965 24395 11023 24401
rect 10965 24361 10977 24395
rect 11011 24392 11023 24395
rect 11514 24392 11520 24404
rect 11011 24364 11520 24392
rect 11011 24361 11023 24364
rect 10965 24355 11023 24361
rect 1394 24256 1400 24268
rect 1355 24228 1400 24256
rect 1394 24216 1400 24228
rect 1452 24216 1458 24268
rect 3050 24256 3056 24268
rect 3011 24228 3056 24256
rect 3050 24216 3056 24228
rect 3108 24216 3114 24268
rect 3513 24259 3571 24265
rect 3513 24225 3525 24259
rect 3559 24256 3571 24259
rect 4157 24259 4215 24265
rect 4157 24256 4169 24259
rect 3559 24228 4169 24256
rect 3559 24225 3571 24228
rect 3513 24219 3571 24225
rect 4157 24225 4169 24228
rect 4203 24225 4215 24259
rect 4157 24219 4215 24225
rect 4246 24216 4252 24268
rect 4304 24256 4310 24268
rect 4724 24256 4752 24352
rect 10980 24324 11008 24355
rect 11514 24352 11520 24364
rect 11572 24392 11578 24404
rect 15562 24392 15568 24404
rect 11572 24364 15568 24392
rect 11572 24352 11578 24364
rect 15562 24352 15568 24364
rect 15620 24352 15626 24404
rect 15838 24352 15844 24404
rect 15896 24392 15902 24404
rect 15896 24364 17816 24392
rect 15896 24352 15902 24364
rect 10060 24296 11008 24324
rect 17788 24324 17816 24364
rect 17862 24352 17868 24404
rect 17920 24392 17926 24404
rect 18233 24395 18291 24401
rect 18233 24392 18245 24395
rect 17920 24364 18245 24392
rect 17920 24352 17926 24364
rect 18233 24361 18245 24364
rect 18279 24392 18291 24395
rect 18322 24392 18328 24404
rect 18279 24364 18328 24392
rect 18279 24361 18291 24364
rect 18233 24355 18291 24361
rect 18322 24352 18328 24364
rect 18380 24352 18386 24404
rect 19702 24392 19708 24404
rect 19663 24364 19708 24392
rect 19702 24352 19708 24364
rect 19760 24352 19766 24404
rect 22646 24352 22652 24404
rect 22704 24392 22710 24404
rect 22741 24395 22799 24401
rect 22741 24392 22753 24395
rect 22704 24364 22753 24392
rect 22704 24352 22710 24364
rect 22741 24361 22753 24364
rect 22787 24392 22799 24395
rect 23382 24392 23388 24404
rect 22787 24364 23388 24392
rect 22787 24361 22799 24364
rect 22741 24355 22799 24361
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 26234 24392 26240 24404
rect 23584 24364 26240 24392
rect 17788 24296 18276 24324
rect 6914 24256 6920 24268
rect 4304 24228 4752 24256
rect 6875 24228 6920 24256
rect 4304 24216 4310 24228
rect 6914 24216 6920 24228
rect 6972 24216 6978 24268
rect 9490 24256 9496 24268
rect 9451 24228 9496 24256
rect 9490 24216 9496 24228
rect 9548 24216 9554 24268
rect 10060 24265 10088 24296
rect 10045 24259 10103 24265
rect 10045 24225 10057 24259
rect 10091 24225 10103 24259
rect 10410 24256 10416 24268
rect 10371 24228 10416 24256
rect 10045 24219 10103 24225
rect 10410 24216 10416 24228
rect 10468 24216 10474 24268
rect 11330 24216 11336 24268
rect 11388 24256 11394 24268
rect 11425 24259 11483 24265
rect 11425 24256 11437 24259
rect 11388 24228 11437 24256
rect 11388 24216 11394 24228
rect 11425 24225 11437 24228
rect 11471 24256 11483 24259
rect 13078 24256 13084 24268
rect 11471 24228 13084 24256
rect 11471 24225 11483 24228
rect 11425 24219 11483 24225
rect 13078 24216 13084 24228
rect 13136 24216 13142 24268
rect 2961 24191 3019 24197
rect 2961 24157 2973 24191
rect 3007 24157 3019 24191
rect 3234 24188 3240 24200
rect 3195 24160 3240 24188
rect 2961 24151 3019 24157
rect 1664 24123 1722 24129
rect 1664 24089 1676 24123
rect 1710 24120 1722 24123
rect 1946 24120 1952 24132
rect 1710 24092 1952 24120
rect 1710 24089 1722 24092
rect 1664 24083 1722 24089
rect 1946 24080 1952 24092
rect 2004 24080 2010 24132
rect 2976 24120 3004 24151
rect 3234 24148 3240 24160
rect 3292 24148 3298 24200
rect 3329 24191 3387 24197
rect 3329 24157 3341 24191
rect 3375 24157 3387 24191
rect 3329 24151 3387 24157
rect 3142 24120 3148 24132
rect 2976 24092 3148 24120
rect 3142 24080 3148 24092
rect 3200 24080 3206 24132
rect 3344 24120 3372 24151
rect 3418 24148 3424 24200
rect 3476 24188 3482 24200
rect 4065 24191 4123 24197
rect 4065 24188 4077 24191
rect 3476 24160 4077 24188
rect 3476 24148 3482 24160
rect 4065 24157 4077 24160
rect 4111 24157 4123 24191
rect 4338 24188 4344 24200
rect 4299 24160 4344 24188
rect 4065 24151 4123 24157
rect 4338 24148 4344 24160
rect 4396 24148 4402 24200
rect 4525 24191 4583 24197
rect 4525 24157 4537 24191
rect 4571 24157 4583 24191
rect 4525 24151 4583 24157
rect 4801 24191 4859 24197
rect 4801 24157 4813 24191
rect 4847 24188 4859 24191
rect 4890 24188 4896 24200
rect 4847 24160 4896 24188
rect 4847 24157 4859 24160
rect 4801 24151 4859 24157
rect 3602 24120 3608 24132
rect 3344 24092 3608 24120
rect 3602 24080 3608 24092
rect 3660 24120 3666 24132
rect 4540 24120 4568 24151
rect 4890 24148 4896 24160
rect 4948 24148 4954 24200
rect 5077 24191 5135 24197
rect 5077 24157 5089 24191
rect 5123 24188 5135 24191
rect 5166 24188 5172 24200
rect 5123 24160 5172 24188
rect 5123 24157 5135 24160
rect 5077 24151 5135 24157
rect 5166 24148 5172 24160
rect 5224 24148 5230 24200
rect 9582 24188 9588 24200
rect 9495 24160 9588 24188
rect 9582 24148 9588 24160
rect 9640 24188 9646 24200
rect 11146 24188 11152 24200
rect 9640 24160 11152 24188
rect 9640 24148 9646 24160
rect 11146 24148 11152 24160
rect 11204 24148 11210 24200
rect 14366 24188 14372 24200
rect 14327 24160 14372 24188
rect 14366 24148 14372 24160
rect 14424 24148 14430 24200
rect 16850 24188 16856 24200
rect 16811 24160 16856 24188
rect 16850 24148 16856 24160
rect 16908 24188 16914 24200
rect 18138 24188 18144 24200
rect 16908 24160 18144 24188
rect 16908 24148 16914 24160
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18248 24188 18276 24296
rect 18690 24284 18696 24336
rect 18748 24324 18754 24336
rect 19242 24324 19248 24336
rect 18748 24296 19248 24324
rect 18748 24284 18754 24296
rect 19242 24284 19248 24296
rect 19300 24284 19306 24336
rect 22462 24324 22468 24336
rect 22423 24296 22468 24324
rect 22462 24284 22468 24296
rect 22520 24284 22526 24336
rect 22738 24256 22744 24268
rect 22066 24228 22744 24256
rect 20346 24188 20352 24200
rect 18248 24160 20352 24188
rect 20346 24148 20352 24160
rect 20404 24148 20410 24200
rect 20990 24148 20996 24200
rect 21048 24188 21054 24200
rect 21085 24191 21143 24197
rect 21085 24188 21097 24191
rect 21048 24160 21097 24188
rect 21048 24148 21054 24160
rect 21085 24157 21097 24160
rect 21131 24157 21143 24191
rect 21085 24151 21143 24157
rect 21913 24191 21971 24197
rect 21913 24157 21925 24191
rect 21959 24188 21971 24191
rect 22066 24188 22094 24228
rect 22738 24216 22744 24228
rect 22796 24256 22802 24268
rect 22922 24256 22928 24268
rect 22796 24228 22928 24256
rect 22796 24216 22802 24228
rect 22922 24216 22928 24228
rect 22980 24216 22986 24268
rect 21959 24160 22094 24188
rect 21959 24157 21971 24160
rect 21913 24151 21971 24157
rect 22186 24148 22192 24200
rect 22244 24188 22250 24200
rect 22333 24191 22391 24197
rect 22244 24160 22289 24188
rect 22244 24148 22250 24160
rect 22333 24157 22345 24191
rect 22379 24188 22391 24191
rect 22830 24188 22836 24200
rect 22379 24160 22836 24188
rect 22379 24157 22391 24160
rect 22333 24151 22391 24157
rect 22830 24148 22836 24160
rect 22888 24148 22894 24200
rect 23198 24148 23204 24200
rect 23256 24188 23262 24200
rect 23584 24197 23612 24364
rect 26234 24352 26240 24364
rect 26292 24352 26298 24404
rect 25774 24256 25780 24268
rect 25735 24228 25780 24256
rect 25774 24216 25780 24228
rect 25832 24216 25838 24268
rect 23293 24191 23351 24197
rect 23293 24188 23305 24191
rect 23256 24160 23305 24188
rect 23256 24148 23262 24160
rect 23293 24157 23305 24160
rect 23339 24157 23351 24191
rect 23293 24151 23351 24157
rect 23569 24191 23627 24197
rect 23569 24157 23581 24191
rect 23615 24157 23627 24191
rect 23569 24151 23627 24157
rect 23658 24148 23664 24200
rect 23716 24197 23722 24200
rect 23716 24188 23724 24197
rect 24394 24188 24400 24200
rect 23716 24160 23761 24188
rect 24355 24160 24400 24188
rect 23716 24151 23724 24160
rect 23716 24148 23722 24151
rect 24394 24148 24400 24160
rect 24452 24148 24458 24200
rect 25501 24191 25559 24197
rect 25501 24157 25513 24191
rect 25547 24157 25559 24191
rect 25501 24151 25559 24157
rect 3660 24092 4568 24120
rect 5344 24123 5402 24129
rect 3660 24080 3666 24092
rect 5344 24089 5356 24123
rect 5390 24120 5402 24123
rect 5534 24120 5540 24132
rect 5390 24092 5540 24120
rect 5390 24089 5402 24092
rect 5344 24083 5402 24089
rect 5534 24080 5540 24092
rect 5592 24080 5598 24132
rect 7190 24120 7196 24132
rect 7151 24092 7196 24120
rect 7190 24080 7196 24092
rect 7248 24080 7254 24132
rect 7282 24080 7288 24132
rect 7340 24120 7346 24132
rect 9493 24123 9551 24129
rect 9493 24120 9505 24123
rect 7340 24092 7682 24120
rect 8680 24092 9505 24120
rect 7340 24080 7346 24092
rect 3326 24012 3332 24064
rect 3384 24052 3390 24064
rect 3881 24055 3939 24061
rect 3881 24052 3893 24055
rect 3384 24024 3893 24052
rect 3384 24012 3390 24024
rect 3881 24021 3893 24024
rect 3927 24021 3939 24055
rect 6454 24052 6460 24064
rect 6415 24024 6460 24052
rect 3881 24015 3939 24021
rect 6454 24012 6460 24024
rect 6512 24012 6518 24064
rect 6730 24012 6736 24064
rect 6788 24052 6794 24064
rect 8680 24061 8708 24092
rect 9493 24089 9505 24092
rect 9539 24089 9551 24123
rect 9493 24083 9551 24089
rect 11054 24080 11060 24132
rect 11112 24120 11118 24132
rect 11701 24123 11759 24129
rect 11701 24120 11713 24123
rect 11112 24092 11713 24120
rect 11112 24080 11118 24092
rect 11701 24089 11713 24092
rect 11747 24089 11759 24123
rect 11701 24083 11759 24089
rect 12710 24080 12716 24132
rect 12768 24080 12774 24132
rect 17120 24123 17178 24129
rect 17120 24089 17132 24123
rect 17166 24120 17178 24123
rect 17770 24120 17776 24132
rect 17166 24092 17776 24120
rect 17166 24089 17178 24092
rect 17120 24083 17178 24089
rect 17770 24080 17776 24092
rect 17828 24080 17834 24132
rect 19061 24123 19119 24129
rect 19061 24089 19073 24123
rect 19107 24120 19119 24123
rect 19429 24123 19487 24129
rect 19429 24120 19441 24123
rect 19107 24092 19441 24120
rect 19107 24089 19119 24092
rect 19061 24083 19119 24089
rect 8665 24055 8723 24061
rect 8665 24052 8677 24055
rect 6788 24024 8677 24052
rect 6788 24012 6794 24024
rect 8665 24021 8677 24024
rect 8711 24021 8723 24055
rect 8665 24015 8723 24021
rect 8754 24012 8760 24064
rect 8812 24052 8818 24064
rect 9015 24055 9073 24061
rect 9015 24052 9027 24055
rect 8812 24024 9027 24052
rect 8812 24012 8818 24024
rect 9015 24021 9027 24024
rect 9061 24021 9073 24055
rect 9015 24015 9073 24021
rect 9858 24012 9864 24064
rect 9916 24052 9922 24064
rect 10229 24055 10287 24061
rect 10229 24052 10241 24055
rect 9916 24024 10241 24052
rect 9916 24012 9922 24024
rect 10229 24021 10241 24024
rect 10275 24021 10287 24055
rect 10229 24015 10287 24021
rect 12618 24012 12624 24064
rect 12676 24052 12682 24064
rect 13173 24055 13231 24061
rect 13173 24052 13185 24055
rect 12676 24024 13185 24052
rect 12676 24012 12682 24024
rect 13173 24021 13185 24024
rect 13219 24021 13231 24055
rect 14550 24052 14556 24064
rect 14511 24024 14556 24052
rect 13173 24015 13231 24021
rect 14550 24012 14556 24024
rect 14608 24012 14614 24064
rect 19260 24052 19288 24092
rect 19429 24089 19441 24092
rect 19475 24089 19487 24123
rect 19429 24083 19487 24089
rect 20162 24080 20168 24132
rect 20220 24120 20226 24132
rect 20818 24123 20876 24129
rect 20818 24120 20830 24123
rect 20220 24092 20830 24120
rect 20220 24080 20226 24092
rect 20818 24089 20830 24092
rect 20864 24089 20876 24123
rect 20818 24083 20876 24089
rect 22097 24123 22155 24129
rect 22097 24089 22109 24123
rect 22143 24120 22155 24123
rect 22646 24120 22652 24132
rect 22143 24092 22652 24120
rect 22143 24089 22155 24092
rect 22097 24083 22155 24089
rect 22646 24080 22652 24092
rect 22704 24080 22710 24132
rect 23477 24123 23535 24129
rect 23477 24120 23489 24123
rect 23124 24092 23489 24120
rect 19334 24052 19340 24064
rect 19260 24024 19340 24052
rect 19334 24012 19340 24024
rect 19392 24012 19398 24064
rect 23014 24012 23020 24064
rect 23072 24052 23078 24064
rect 23124 24061 23152 24092
rect 23477 24089 23489 24092
rect 23523 24089 23535 24123
rect 25038 24120 25044 24132
rect 23477 24083 23535 24089
rect 23768 24092 25044 24120
rect 23768 24064 23796 24092
rect 25038 24080 25044 24092
rect 25096 24120 25102 24132
rect 25516 24120 25544 24151
rect 25096 24092 25544 24120
rect 25096 24080 25102 24092
rect 26510 24080 26516 24132
rect 26568 24080 26574 24132
rect 23109 24055 23167 24061
rect 23109 24052 23121 24055
rect 23072 24024 23121 24052
rect 23072 24012 23078 24024
rect 23109 24021 23121 24024
rect 23155 24021 23167 24055
rect 23109 24015 23167 24021
rect 23382 24012 23388 24064
rect 23440 24052 23446 24064
rect 23566 24052 23572 24064
rect 23440 24024 23572 24052
rect 23440 24012 23446 24024
rect 23566 24012 23572 24024
rect 23624 24012 23630 24064
rect 23750 24012 23756 24064
rect 23808 24012 23814 24064
rect 23862 24055 23920 24061
rect 23862 24021 23874 24055
rect 23908 24052 23920 24055
rect 24026 24052 24032 24064
rect 23908 24024 24032 24052
rect 23908 24021 23920 24024
rect 23862 24015 23920 24021
rect 24026 24012 24032 24024
rect 24084 24012 24090 24064
rect 24578 24052 24584 24064
rect 24539 24024 24584 24052
rect 24578 24012 24584 24024
rect 24636 24012 24642 24064
rect 26694 24012 26700 24064
rect 26752 24052 26758 24064
rect 27249 24055 27307 24061
rect 27249 24052 27261 24055
rect 26752 24024 27261 24052
rect 26752 24012 26758 24024
rect 27249 24021 27261 24024
rect 27295 24052 27307 24055
rect 27614 24052 27620 24064
rect 27295 24024 27620 24052
rect 27295 24021 27307 24024
rect 27249 24015 27307 24021
rect 27614 24012 27620 24024
rect 27672 24012 27678 24064
rect 1104 23962 29440 23984
rect 1104 23910 10395 23962
rect 10447 23910 10459 23962
rect 10511 23910 10523 23962
rect 10575 23910 10587 23962
rect 10639 23910 10651 23962
rect 10703 23910 19840 23962
rect 19892 23910 19904 23962
rect 19956 23910 19968 23962
rect 20020 23910 20032 23962
rect 20084 23910 20096 23962
rect 20148 23910 29440 23962
rect 1104 23888 29440 23910
rect 2501 23851 2559 23857
rect 2501 23817 2513 23851
rect 2547 23817 2559 23851
rect 2501 23811 2559 23817
rect 1946 23780 1952 23792
rect 1907 23752 1952 23780
rect 1946 23740 1952 23752
rect 2004 23740 2010 23792
rect 2516 23780 2544 23811
rect 2590 23808 2596 23860
rect 2648 23848 2654 23860
rect 2648 23820 2693 23848
rect 2648 23808 2654 23820
rect 3234 23808 3240 23860
rect 3292 23848 3298 23860
rect 3329 23851 3387 23857
rect 3329 23848 3341 23851
rect 3292 23820 3341 23848
rect 3292 23808 3298 23820
rect 3329 23817 3341 23820
rect 3375 23817 3387 23851
rect 3602 23848 3608 23860
rect 3563 23820 3608 23848
rect 3329 23811 3387 23817
rect 3602 23808 3608 23820
rect 3660 23808 3666 23860
rect 4338 23808 4344 23860
rect 4396 23848 4402 23860
rect 5534 23848 5540 23860
rect 4396 23820 4568 23848
rect 5495 23820 5540 23848
rect 4396 23808 4402 23820
rect 2866 23780 2872 23792
rect 2332 23752 2544 23780
rect 2700 23752 2872 23780
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23681 2191 23715
rect 2133 23675 2191 23681
rect 2148 23508 2176 23675
rect 2332 23576 2360 23752
rect 2389 23715 2447 23721
rect 2389 23681 2401 23715
rect 2435 23712 2447 23715
rect 2700 23712 2728 23752
rect 2866 23740 2872 23752
rect 2924 23780 2930 23792
rect 2961 23783 3019 23789
rect 2961 23780 2973 23783
rect 2924 23752 2973 23780
rect 2924 23740 2930 23752
rect 2961 23749 2973 23752
rect 3007 23749 3019 23783
rect 2961 23743 3019 23749
rect 3142 23740 3148 23792
rect 3200 23780 3206 23792
rect 3200 23752 3740 23780
rect 3200 23740 3206 23752
rect 2435 23684 2728 23712
rect 2435 23681 2447 23684
rect 2389 23675 2447 23681
rect 2774 23672 2780 23724
rect 2832 23712 2838 23724
rect 3712 23721 3740 23752
rect 3421 23715 3479 23721
rect 2832 23684 2877 23712
rect 2832 23672 2838 23684
rect 3421 23681 3433 23715
rect 3467 23681 3479 23715
rect 3421 23675 3479 23681
rect 3697 23715 3755 23721
rect 3697 23681 3709 23715
rect 3743 23712 3755 23715
rect 3786 23712 3792 23724
rect 3743 23684 3792 23712
rect 3743 23681 3755 23684
rect 3697 23675 3755 23681
rect 2685 23647 2743 23653
rect 2685 23613 2697 23647
rect 2731 23644 2743 23647
rect 2731 23616 3004 23644
rect 2731 23613 2743 23616
rect 2685 23607 2743 23613
rect 2774 23576 2780 23588
rect 2332 23548 2780 23576
rect 2774 23536 2780 23548
rect 2832 23536 2838 23588
rect 2976 23576 3004 23616
rect 3050 23604 3056 23656
rect 3108 23644 3114 23656
rect 3145 23647 3203 23653
rect 3145 23644 3157 23647
rect 3108 23616 3157 23644
rect 3108 23604 3114 23616
rect 3145 23613 3157 23616
rect 3191 23644 3203 23647
rect 3436 23644 3464 23675
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 4246 23672 4252 23724
rect 4304 23712 4310 23724
rect 4540 23721 4568 23820
rect 5534 23808 5540 23820
rect 5592 23808 5598 23860
rect 6365 23851 6423 23857
rect 6365 23848 6377 23851
rect 5644 23820 6377 23848
rect 4709 23783 4767 23789
rect 4709 23749 4721 23783
rect 4755 23780 4767 23783
rect 5644 23780 5672 23820
rect 6365 23817 6377 23820
rect 6411 23817 6423 23851
rect 6730 23848 6736 23860
rect 6691 23820 6736 23848
rect 6365 23811 6423 23817
rect 6730 23808 6736 23820
rect 6788 23808 6794 23860
rect 7190 23808 7196 23860
rect 7248 23848 7254 23860
rect 7377 23851 7435 23857
rect 7377 23848 7389 23851
rect 7248 23820 7389 23848
rect 7248 23808 7254 23820
rect 7377 23817 7389 23820
rect 7423 23817 7435 23851
rect 7377 23811 7435 23817
rect 9861 23851 9919 23857
rect 9861 23817 9873 23851
rect 9907 23848 9919 23851
rect 10870 23848 10876 23860
rect 9907 23820 10876 23848
rect 9907 23817 9919 23820
rect 9861 23811 9919 23817
rect 10870 23808 10876 23820
rect 10928 23808 10934 23860
rect 11885 23851 11943 23857
rect 11885 23817 11897 23851
rect 11931 23848 11943 23851
rect 12158 23848 12164 23860
rect 11931 23820 12164 23848
rect 11931 23817 11943 23820
rect 11885 23811 11943 23817
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 12710 23848 12716 23860
rect 12671 23820 12716 23848
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 17497 23851 17555 23857
rect 17497 23848 17509 23851
rect 12820 23820 17509 23848
rect 6454 23780 6460 23792
rect 4755 23752 5672 23780
rect 5736 23752 6460 23780
rect 4755 23749 4767 23752
rect 4709 23743 4767 23749
rect 4341 23715 4399 23721
rect 4341 23712 4353 23715
rect 4304 23684 4353 23712
rect 4304 23672 4310 23684
rect 4341 23681 4353 23684
rect 4387 23681 4399 23715
rect 4341 23675 4399 23681
rect 4525 23715 4583 23721
rect 4525 23681 4537 23715
rect 4571 23681 4583 23715
rect 4798 23712 4804 23724
rect 4759 23684 4804 23712
rect 4525 23675 4583 23681
rect 3878 23644 3884 23656
rect 3191 23616 3884 23644
rect 3191 23613 3203 23616
rect 3145 23607 3203 23613
rect 3878 23604 3884 23616
rect 3936 23604 3942 23656
rect 4540 23644 4568 23675
rect 4798 23672 4804 23684
rect 4856 23672 4862 23724
rect 4982 23721 4988 23724
rect 4945 23715 4988 23721
rect 4945 23681 4957 23715
rect 4945 23675 4988 23681
rect 4982 23672 4988 23675
rect 5040 23672 5046 23724
rect 5736 23721 5764 23752
rect 6454 23740 6460 23752
rect 6512 23780 6518 23792
rect 6825 23783 6883 23789
rect 6825 23780 6837 23783
rect 6512 23752 6837 23780
rect 6512 23740 6518 23752
rect 6825 23749 6837 23752
rect 6871 23749 6883 23783
rect 6825 23743 6883 23749
rect 9953 23783 10011 23789
rect 9953 23749 9965 23783
rect 9999 23780 10011 23783
rect 9999 23752 10548 23780
rect 9999 23749 10011 23752
rect 9953 23743 10011 23749
rect 5721 23715 5779 23721
rect 5721 23681 5733 23715
rect 5767 23681 5779 23715
rect 5721 23675 5779 23681
rect 5813 23715 5871 23721
rect 5813 23681 5825 23715
rect 5859 23681 5871 23715
rect 5813 23675 5871 23681
rect 5828 23644 5856 23675
rect 6546 23672 6552 23724
rect 6604 23712 6610 23724
rect 7466 23712 7472 23724
rect 6604 23684 7472 23712
rect 6604 23672 6610 23684
rect 3988 23616 5856 23644
rect 6089 23647 6147 23653
rect 3988 23576 4016 23616
rect 6089 23613 6101 23647
rect 6135 23644 6147 23647
rect 6822 23644 6828 23656
rect 6135 23616 6828 23644
rect 6135 23613 6147 23616
rect 6089 23607 6147 23613
rect 6822 23604 6828 23616
rect 6880 23604 6886 23656
rect 6932 23653 6960 23684
rect 7466 23672 7472 23684
rect 7524 23672 7530 23724
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23712 7619 23715
rect 8754 23712 8760 23724
rect 7607 23684 8760 23712
rect 7607 23681 7619 23684
rect 7561 23675 7619 23681
rect 8754 23672 8760 23684
rect 8812 23672 8818 23724
rect 9766 23672 9772 23724
rect 9824 23712 9830 23724
rect 10520 23721 10548 23752
rect 10137 23715 10195 23721
rect 10137 23712 10149 23715
rect 9824 23684 10149 23712
rect 9824 23672 9830 23684
rect 10137 23681 10149 23684
rect 10183 23681 10195 23715
rect 10137 23675 10195 23681
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23712 10563 23715
rect 10778 23712 10784 23724
rect 10551 23684 10784 23712
rect 10551 23681 10563 23684
rect 10505 23675 10563 23681
rect 10778 23672 10784 23684
rect 10836 23672 10842 23724
rect 12069 23715 12127 23721
rect 12069 23681 12081 23715
rect 12115 23712 12127 23715
rect 12618 23712 12624 23724
rect 12115 23684 12624 23712
rect 12115 23681 12127 23684
rect 12069 23675 12127 23681
rect 12618 23672 12624 23684
rect 12676 23672 12682 23724
rect 6917 23647 6975 23653
rect 6917 23613 6929 23647
rect 6963 23613 6975 23647
rect 11698 23644 11704 23656
rect 11659 23616 11704 23644
rect 6917 23607 6975 23613
rect 11698 23604 11704 23616
rect 11756 23604 11762 23656
rect 2976 23548 4016 23576
rect 4062 23536 4068 23588
rect 4120 23576 4126 23588
rect 12820 23576 12848 23820
rect 17497 23817 17509 23820
rect 17543 23817 17555 23851
rect 17770 23848 17776 23860
rect 17731 23820 17776 23848
rect 17497 23811 17555 23817
rect 14550 23740 14556 23792
rect 14608 23740 14614 23792
rect 12897 23715 12955 23721
rect 12897 23681 12909 23715
rect 12943 23712 12955 23715
rect 13170 23712 13176 23724
rect 12943 23684 13032 23712
rect 13131 23684 13176 23712
rect 12943 23681 12955 23684
rect 12897 23675 12955 23681
rect 13004 23585 13032 23684
rect 13170 23672 13176 23684
rect 13228 23672 13234 23724
rect 15289 23715 15347 23721
rect 15289 23681 15301 23715
rect 15335 23712 15347 23715
rect 15562 23712 15568 23724
rect 15335 23684 15568 23712
rect 15335 23681 15347 23684
rect 15289 23675 15347 23681
rect 15562 23672 15568 23684
rect 15620 23672 15626 23724
rect 15838 23712 15844 23724
rect 15799 23684 15844 23712
rect 15838 23672 15844 23684
rect 15896 23672 15902 23724
rect 16209 23715 16267 23721
rect 16209 23681 16221 23715
rect 16255 23712 16267 23715
rect 16298 23712 16304 23724
rect 16255 23684 16304 23712
rect 16255 23681 16267 23684
rect 16209 23675 16267 23681
rect 13078 23604 13084 23656
rect 13136 23644 13142 23656
rect 13357 23647 13415 23653
rect 13357 23644 13369 23647
rect 13136 23616 13369 23644
rect 13136 23604 13142 23616
rect 13357 23613 13369 23616
rect 13403 23613 13415 23647
rect 13722 23644 13728 23656
rect 13683 23616 13728 23644
rect 13357 23607 13415 23613
rect 13722 23604 13728 23616
rect 13780 23604 13786 23656
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23644 15255 23647
rect 15746 23644 15752 23656
rect 15243 23616 15752 23644
rect 15243 23613 15255 23616
rect 15197 23607 15255 23613
rect 15746 23604 15752 23616
rect 15804 23604 15810 23656
rect 4120 23548 12848 23576
rect 12989 23579 13047 23585
rect 4120 23536 4126 23548
rect 12989 23545 13001 23579
rect 13035 23545 13047 23579
rect 12989 23539 13047 23545
rect 16025 23579 16083 23585
rect 16025 23545 16037 23579
rect 16071 23576 16083 23579
rect 16224 23576 16252 23675
rect 16298 23672 16304 23684
rect 16356 23672 16362 23724
rect 16853 23715 16911 23721
rect 16853 23712 16865 23715
rect 16408 23684 16865 23712
rect 16408 23585 16436 23684
rect 16853 23681 16865 23684
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 16071 23548 16252 23576
rect 16393 23579 16451 23585
rect 16071 23545 16083 23548
rect 16025 23539 16083 23545
rect 16393 23545 16405 23579
rect 16439 23545 16451 23579
rect 17512 23576 17540 23811
rect 17770 23808 17776 23820
rect 17828 23808 17834 23860
rect 19150 23808 19156 23860
rect 19208 23848 19214 23860
rect 19981 23851 20039 23857
rect 19208 23820 19932 23848
rect 19208 23808 19214 23820
rect 18966 23780 18972 23792
rect 18432 23752 18972 23780
rect 17862 23712 17868 23724
rect 17823 23684 17868 23712
rect 17862 23672 17868 23684
rect 17920 23672 17926 23724
rect 18046 23721 18052 23724
rect 18003 23715 18052 23721
rect 18003 23681 18015 23715
rect 18049 23681 18052 23715
rect 18003 23675 18052 23681
rect 18046 23672 18052 23675
rect 18104 23672 18110 23724
rect 18234 23715 18292 23721
rect 18234 23681 18246 23715
rect 18280 23712 18292 23715
rect 18322 23712 18328 23724
rect 18280 23684 18328 23712
rect 18280 23681 18292 23684
rect 18234 23675 18292 23681
rect 18322 23672 18328 23684
rect 18380 23672 18386 23724
rect 18432 23721 18460 23752
rect 18966 23740 18972 23752
rect 19024 23740 19030 23792
rect 19904 23780 19932 23820
rect 19981 23817 19993 23851
rect 20027 23848 20039 23851
rect 20162 23848 20168 23860
rect 20027 23820 20168 23848
rect 20027 23817 20039 23820
rect 19981 23811 20039 23817
rect 20162 23808 20168 23820
rect 20220 23808 20226 23860
rect 20346 23808 20352 23860
rect 20404 23848 20410 23860
rect 22370 23848 22376 23860
rect 20404 23820 22376 23848
rect 20404 23808 20410 23820
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 22554 23808 22560 23860
rect 22612 23848 22618 23860
rect 23382 23848 23388 23860
rect 22612 23820 23388 23848
rect 22612 23808 22618 23820
rect 23382 23808 23388 23820
rect 23440 23808 23446 23860
rect 23661 23851 23719 23857
rect 23661 23817 23673 23851
rect 23707 23848 23719 23851
rect 24394 23848 24400 23860
rect 23707 23820 24400 23848
rect 23707 23817 23719 23820
rect 23661 23811 23719 23817
rect 24394 23808 24400 23820
rect 24452 23808 24458 23860
rect 25501 23851 25559 23857
rect 25501 23817 25513 23851
rect 25547 23848 25559 23851
rect 26234 23848 26240 23860
rect 25547 23820 26240 23848
rect 25547 23817 25559 23820
rect 25501 23811 25559 23817
rect 26234 23808 26240 23820
rect 26292 23808 26298 23860
rect 24026 23780 24032 23792
rect 19904 23752 23520 23780
rect 23987 23752 24032 23780
rect 18417 23715 18475 23721
rect 18417 23681 18429 23715
rect 18463 23681 18475 23715
rect 18417 23675 18475 23681
rect 18598 23672 18604 23724
rect 18656 23712 18662 23724
rect 18693 23715 18751 23721
rect 18693 23712 18705 23715
rect 18656 23684 18705 23712
rect 18656 23672 18662 23684
rect 18693 23681 18705 23684
rect 18739 23681 18751 23715
rect 18984 23712 19012 23740
rect 19150 23712 19156 23724
rect 18984 23684 19156 23712
rect 18693 23675 18751 23681
rect 19150 23672 19156 23684
rect 19208 23712 19214 23724
rect 19337 23715 19395 23721
rect 19337 23712 19349 23715
rect 19208 23684 19349 23712
rect 19208 23672 19214 23684
rect 19337 23681 19349 23684
rect 19383 23681 19395 23715
rect 19337 23675 19395 23681
rect 19520 23715 19578 23721
rect 19520 23681 19532 23715
rect 19566 23712 19578 23715
rect 19566 23684 19840 23712
rect 19566 23681 19578 23684
rect 19520 23675 19578 23681
rect 18141 23647 18199 23653
rect 18141 23613 18153 23647
rect 18187 23644 18199 23647
rect 18187 23616 18552 23644
rect 18187 23613 18199 23616
rect 18141 23607 18199 23613
rect 18322 23576 18328 23588
rect 17512 23548 18328 23576
rect 16393 23539 16451 23545
rect 18322 23536 18328 23548
rect 18380 23536 18386 23588
rect 4157 23511 4215 23517
rect 4157 23508 4169 23511
rect 2148 23480 4169 23508
rect 4157 23477 4169 23480
rect 4203 23508 4215 23511
rect 4982 23508 4988 23520
rect 4203 23480 4988 23508
rect 4203 23477 4215 23480
rect 4157 23471 4215 23477
rect 4982 23468 4988 23480
rect 5040 23468 5046 23520
rect 5077 23511 5135 23517
rect 5077 23477 5089 23511
rect 5123 23508 5135 23511
rect 5534 23508 5540 23520
rect 5123 23480 5540 23508
rect 5123 23477 5135 23480
rect 5077 23471 5135 23477
rect 5534 23468 5540 23480
rect 5592 23468 5598 23520
rect 5997 23511 6055 23517
rect 5997 23477 6009 23511
rect 6043 23508 6055 23511
rect 6086 23508 6092 23520
rect 6043 23480 6092 23508
rect 6043 23477 6055 23480
rect 5997 23471 6055 23477
rect 6086 23468 6092 23480
rect 6144 23468 6150 23520
rect 10226 23508 10232 23520
rect 10187 23480 10232 23508
rect 10226 23468 10232 23480
rect 10284 23468 10290 23520
rect 10965 23511 11023 23517
rect 10965 23477 10977 23511
rect 11011 23508 11023 23511
rect 11422 23508 11428 23520
rect 11011 23480 11428 23508
rect 11011 23477 11023 23480
rect 10965 23471 11023 23477
rect 11422 23468 11428 23480
rect 11480 23468 11486 23520
rect 11701 23511 11759 23517
rect 11701 23477 11713 23511
rect 11747 23508 11759 23511
rect 11790 23508 11796 23520
rect 11747 23480 11796 23508
rect 11747 23477 11759 23480
rect 11701 23471 11759 23477
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 15470 23508 15476 23520
rect 15431 23480 15476 23508
rect 15470 23468 15476 23480
rect 15528 23468 15534 23520
rect 16666 23508 16672 23520
rect 16627 23480 16672 23508
rect 16666 23468 16672 23480
rect 16724 23468 16730 23520
rect 18524 23517 18552 23616
rect 19058 23604 19064 23656
rect 19116 23644 19122 23656
rect 19613 23647 19671 23653
rect 19613 23644 19625 23647
rect 19116 23616 19625 23644
rect 19116 23604 19122 23616
rect 19613 23613 19625 23616
rect 19659 23613 19671 23647
rect 19613 23607 19671 23613
rect 19705 23647 19763 23653
rect 19705 23613 19717 23647
rect 19751 23613 19763 23647
rect 19705 23607 19763 23613
rect 18966 23536 18972 23588
rect 19024 23576 19030 23588
rect 19720 23576 19748 23607
rect 19024 23548 19748 23576
rect 19812 23576 19840 23684
rect 19886 23672 19892 23724
rect 19944 23712 19950 23724
rect 22002 23712 22008 23724
rect 19944 23684 19989 23712
rect 21963 23684 22008 23712
rect 19944 23672 19950 23684
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 22738 23712 22744 23724
rect 22699 23684 22744 23712
rect 22738 23672 22744 23684
rect 22796 23672 22802 23724
rect 23492 23721 23520 23752
rect 24026 23740 24032 23752
rect 24084 23740 24090 23792
rect 24578 23740 24584 23792
rect 24636 23740 24642 23792
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23681 23535 23715
rect 23477 23675 23535 23681
rect 23750 23644 23756 23656
rect 23711 23616 23756 23644
rect 23750 23604 23756 23616
rect 23808 23604 23814 23656
rect 20257 23579 20315 23585
rect 20257 23576 20269 23579
rect 19812 23548 20269 23576
rect 19024 23536 19030 23548
rect 20257 23545 20269 23548
rect 20303 23576 20315 23579
rect 20303 23548 23888 23576
rect 20303 23545 20315 23548
rect 20257 23539 20315 23545
rect 18509 23511 18567 23517
rect 18509 23477 18521 23511
rect 18555 23508 18567 23511
rect 19058 23508 19064 23520
rect 18555 23480 19064 23508
rect 18555 23477 18567 23480
rect 18509 23471 18567 23477
rect 19058 23468 19064 23480
rect 19116 23468 19122 23520
rect 21818 23508 21824 23520
rect 21779 23480 21824 23508
rect 21818 23468 21824 23480
rect 21876 23468 21882 23520
rect 22557 23511 22615 23517
rect 22557 23477 22569 23511
rect 22603 23508 22615 23511
rect 22922 23508 22928 23520
rect 22603 23480 22928 23508
rect 22603 23477 22615 23480
rect 22557 23471 22615 23477
rect 22922 23468 22928 23480
rect 22980 23468 22986 23520
rect 23860 23508 23888 23548
rect 26326 23508 26332 23520
rect 23860 23480 26332 23508
rect 26326 23468 26332 23480
rect 26384 23468 26390 23520
rect 1104 23418 29440 23440
rect 1104 23366 5672 23418
rect 5724 23366 5736 23418
rect 5788 23366 5800 23418
rect 5852 23366 5864 23418
rect 5916 23366 5928 23418
rect 5980 23366 15118 23418
rect 15170 23366 15182 23418
rect 15234 23366 15246 23418
rect 15298 23366 15310 23418
rect 15362 23366 15374 23418
rect 15426 23366 24563 23418
rect 24615 23366 24627 23418
rect 24679 23366 24691 23418
rect 24743 23366 24755 23418
rect 24807 23366 24819 23418
rect 24871 23366 29440 23418
rect 1104 23344 29440 23366
rect 9677 23307 9735 23313
rect 9677 23273 9689 23307
rect 9723 23304 9735 23307
rect 10042 23304 10048 23316
rect 9723 23276 10048 23304
rect 9723 23273 9735 23276
rect 9677 23267 9735 23273
rect 10042 23264 10048 23276
rect 10100 23264 10106 23316
rect 10134 23264 10140 23316
rect 10192 23304 10198 23316
rect 11238 23304 11244 23316
rect 10192 23276 11244 23304
rect 10192 23264 10198 23276
rect 11238 23264 11244 23276
rect 11296 23264 11302 23316
rect 13541 23307 13599 23313
rect 13541 23273 13553 23307
rect 13587 23304 13599 23307
rect 13722 23304 13728 23316
rect 13587 23276 13728 23304
rect 13587 23273 13599 23276
rect 13541 23267 13599 23273
rect 13722 23264 13728 23276
rect 13780 23264 13786 23316
rect 14366 23304 14372 23316
rect 14327 23276 14372 23304
rect 14366 23264 14372 23276
rect 14424 23264 14430 23316
rect 18506 23264 18512 23316
rect 18564 23304 18570 23316
rect 19245 23307 19303 23313
rect 19245 23304 19257 23307
rect 18564 23276 19257 23304
rect 18564 23264 18570 23276
rect 19245 23273 19257 23276
rect 19291 23273 19303 23307
rect 19245 23267 19303 23273
rect 20806 23264 20812 23316
rect 20864 23304 20870 23316
rect 20993 23307 21051 23313
rect 20993 23304 21005 23307
rect 20864 23276 21005 23304
rect 20864 23264 20870 23276
rect 20993 23273 21005 23276
rect 21039 23304 21051 23307
rect 22094 23304 22100 23316
rect 21039 23276 22100 23304
rect 21039 23273 21051 23276
rect 20993 23267 21051 23273
rect 22094 23264 22100 23276
rect 22152 23264 22158 23316
rect 22738 23264 22744 23316
rect 22796 23304 22802 23316
rect 23293 23307 23351 23313
rect 23293 23304 23305 23307
rect 22796 23276 23305 23304
rect 22796 23264 22802 23276
rect 23293 23273 23305 23276
rect 23339 23273 23351 23307
rect 23293 23267 23351 23273
rect 23842 23264 23848 23316
rect 23900 23304 23906 23316
rect 24394 23304 24400 23316
rect 23900 23276 24400 23304
rect 23900 23264 23906 23276
rect 24394 23264 24400 23276
rect 24452 23304 24458 23316
rect 24581 23307 24639 23313
rect 24581 23304 24593 23307
rect 24452 23276 24593 23304
rect 24452 23264 24458 23276
rect 24581 23273 24593 23276
rect 24627 23273 24639 23307
rect 24581 23267 24639 23273
rect 11422 23236 11428 23248
rect 10152 23208 11428 23236
rect 3970 23128 3976 23180
rect 4028 23168 4034 23180
rect 10152 23177 10180 23208
rect 11422 23196 11428 23208
rect 11480 23196 11486 23248
rect 18046 23196 18052 23248
rect 18104 23236 18110 23248
rect 18601 23239 18659 23245
rect 18601 23236 18613 23239
rect 18104 23208 18613 23236
rect 18104 23196 18110 23208
rect 18601 23205 18613 23208
rect 18647 23236 18659 23239
rect 18966 23236 18972 23248
rect 18647 23208 18972 23236
rect 18647 23205 18659 23208
rect 18601 23199 18659 23205
rect 18966 23196 18972 23208
rect 19024 23196 19030 23248
rect 23109 23239 23167 23245
rect 23109 23205 23121 23239
rect 23155 23236 23167 23239
rect 23658 23236 23664 23248
rect 23155 23208 23664 23236
rect 23155 23205 23167 23208
rect 23109 23199 23167 23205
rect 23658 23196 23664 23208
rect 23716 23236 23722 23248
rect 23716 23208 23888 23236
rect 23716 23196 23722 23208
rect 4065 23171 4123 23177
rect 4065 23168 4077 23171
rect 4028 23140 4077 23168
rect 4028 23128 4034 23140
rect 4065 23137 4077 23140
rect 4111 23137 4123 23171
rect 10045 23171 10103 23177
rect 10045 23168 10057 23171
rect 4065 23131 4123 23137
rect 9324 23140 10057 23168
rect 1949 23103 2007 23109
rect 1949 23069 1961 23103
rect 1995 23100 2007 23103
rect 3326 23100 3332 23112
rect 1995 23072 3332 23100
rect 1995 23069 2007 23072
rect 1949 23063 2007 23069
rect 3326 23060 3332 23072
rect 3384 23060 3390 23112
rect 3786 23100 3792 23112
rect 3747 23072 3792 23100
rect 3786 23060 3792 23072
rect 3844 23060 3850 23112
rect 3878 23060 3884 23112
rect 3936 23100 3942 23112
rect 3936 23072 3981 23100
rect 3936 23060 3942 23072
rect 4706 23060 4712 23112
rect 4764 23100 4770 23112
rect 6089 23103 6147 23109
rect 6089 23100 6101 23103
rect 4764 23072 6101 23100
rect 4764 23060 4770 23072
rect 6089 23069 6101 23072
rect 6135 23069 6147 23103
rect 6089 23063 6147 23069
rect 8205 23103 8263 23109
rect 8205 23069 8217 23103
rect 8251 23069 8263 23103
rect 8205 23063 8263 23069
rect 3234 22992 3240 23044
rect 3292 23032 3298 23044
rect 3292 23004 5488 23032
rect 3292 22992 3298 23004
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 1857 22967 1915 22973
rect 1857 22964 1869 22967
rect 1728 22936 1869 22964
rect 1728 22924 1734 22936
rect 1857 22933 1869 22936
rect 1903 22933 1915 22967
rect 1857 22927 1915 22933
rect 4154 22924 4160 22976
rect 4212 22964 4218 22976
rect 4249 22967 4307 22973
rect 4249 22964 4261 22967
rect 4212 22936 4261 22964
rect 4212 22924 4218 22936
rect 4249 22933 4261 22936
rect 4295 22933 4307 22967
rect 4249 22927 4307 22933
rect 4338 22924 4344 22976
rect 4396 22964 4402 22976
rect 4709 22967 4767 22973
rect 4709 22964 4721 22967
rect 4396 22936 4721 22964
rect 4396 22924 4402 22936
rect 4709 22933 4721 22936
rect 4755 22964 4767 22967
rect 4798 22964 4804 22976
rect 4755 22936 4804 22964
rect 4755 22933 4767 22936
rect 4709 22927 4767 22933
rect 4798 22924 4804 22936
rect 4856 22924 4862 22976
rect 5460 22964 5488 23004
rect 5534 22992 5540 23044
rect 5592 23032 5598 23044
rect 5822 23035 5880 23041
rect 5822 23032 5834 23035
rect 5592 23004 5834 23032
rect 5592 22992 5598 23004
rect 5822 23001 5834 23004
rect 5868 23001 5880 23035
rect 5822 22995 5880 23001
rect 7190 22992 7196 23044
rect 7248 22992 7254 23044
rect 7926 23032 7932 23044
rect 7887 23004 7932 23032
rect 7926 22992 7932 23004
rect 7984 22992 7990 23044
rect 8220 22976 8248 23063
rect 9030 22992 9036 23044
rect 9088 23032 9094 23044
rect 9324 23041 9352 23140
rect 10045 23137 10057 23140
rect 10091 23137 10103 23171
rect 10045 23131 10103 23137
rect 10137 23171 10195 23177
rect 10137 23137 10149 23171
rect 10183 23137 10195 23171
rect 10137 23131 10195 23137
rect 10318 23128 10324 23180
rect 10376 23177 10382 23180
rect 10376 23171 10395 23177
rect 10383 23168 10395 23171
rect 11149 23171 11207 23177
rect 11149 23168 11161 23171
rect 10383 23140 11161 23168
rect 10383 23137 10395 23140
rect 10376 23131 10395 23137
rect 11149 23137 11161 23140
rect 11195 23137 11207 23171
rect 11149 23131 11207 23137
rect 10376 23128 10382 23131
rect 11698 23128 11704 23180
rect 11756 23128 11762 23180
rect 13078 23168 13084 23180
rect 12406 23140 13084 23168
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23069 10011 23103
rect 9953 23063 10011 23069
rect 9309 23035 9367 23041
rect 9309 23032 9321 23035
rect 9088 23004 9321 23032
rect 9088 22992 9094 23004
rect 9309 23001 9321 23004
rect 9355 23001 9367 23035
rect 9309 22995 9367 23001
rect 9723 23035 9781 23041
rect 9723 23001 9735 23035
rect 9769 23032 9781 23035
rect 9858 23032 9864 23044
rect 9769 23004 9864 23032
rect 9769 23001 9781 23004
rect 9723 22995 9781 23001
rect 9858 22992 9864 23004
rect 9916 22992 9922 23044
rect 9968 23032 9996 23063
rect 10226 23060 10232 23112
rect 10284 23100 10290 23112
rect 10873 23103 10931 23109
rect 10873 23100 10885 23103
rect 10284 23072 10885 23100
rect 10284 23060 10290 23072
rect 10873 23069 10885 23072
rect 10919 23069 10931 23103
rect 10873 23063 10931 23069
rect 11057 23103 11115 23109
rect 11057 23069 11069 23103
rect 11103 23100 11115 23103
rect 11238 23100 11244 23112
rect 11103 23072 11244 23100
rect 11103 23069 11115 23072
rect 11057 23063 11115 23069
rect 11238 23060 11244 23072
rect 11296 23060 11302 23112
rect 11517 23103 11575 23109
rect 11517 23069 11529 23103
rect 11563 23100 11575 23103
rect 11716 23100 11744 23128
rect 12406 23100 12434 23140
rect 13078 23128 13084 23140
rect 13136 23128 13142 23180
rect 15470 23128 15476 23180
rect 15528 23168 15534 23180
rect 15657 23171 15715 23177
rect 15657 23168 15669 23171
rect 15528 23140 15669 23168
rect 15528 23128 15534 23140
rect 15657 23137 15669 23140
rect 15703 23137 15715 23171
rect 15657 23131 15715 23137
rect 18782 23128 18788 23180
rect 18840 23168 18846 23180
rect 19797 23171 19855 23177
rect 19797 23168 19809 23171
rect 18840 23140 19809 23168
rect 18840 23128 18846 23140
rect 19797 23137 19809 23140
rect 19843 23137 19855 23171
rect 19797 23131 19855 23137
rect 20990 23128 20996 23180
rect 21048 23168 21054 23180
rect 22741 23171 22799 23177
rect 22741 23168 22753 23171
rect 21048 23140 22753 23168
rect 21048 23128 21054 23140
rect 22741 23137 22753 23140
rect 22787 23168 22799 23171
rect 23750 23168 23756 23180
rect 22787 23140 23756 23168
rect 22787 23137 22799 23140
rect 22741 23131 22799 23137
rect 23750 23128 23756 23140
rect 23808 23128 23814 23180
rect 11563 23072 12434 23100
rect 13265 23103 13323 23109
rect 11563 23069 11575 23072
rect 11517 23063 11575 23069
rect 13265 23069 13277 23103
rect 13311 23100 13323 23103
rect 13357 23103 13415 23109
rect 13357 23100 13369 23103
rect 13311 23072 13369 23100
rect 13311 23069 13323 23072
rect 13265 23063 13323 23069
rect 13357 23069 13369 23072
rect 13403 23069 13415 23103
rect 13357 23063 13415 23069
rect 14185 23103 14243 23109
rect 14185 23069 14197 23103
rect 14231 23069 14243 23103
rect 15102 23100 15108 23112
rect 15063 23072 15108 23100
rect 14185 23063 14243 23069
rect 10597 23035 10655 23041
rect 10597 23032 10609 23035
rect 9968 23004 10609 23032
rect 10597 23001 10609 23004
rect 10643 23001 10655 23035
rect 10597 22995 10655 23001
rect 10781 23035 10839 23041
rect 10781 23001 10793 23035
rect 10827 23032 10839 23035
rect 11330 23032 11336 23044
rect 10827 23004 11192 23032
rect 11291 23004 11336 23032
rect 10827 23001 10839 23004
rect 10781 22995 10839 23001
rect 6457 22967 6515 22973
rect 6457 22964 6469 22967
rect 5460 22936 6469 22964
rect 6457 22933 6469 22936
rect 6503 22964 6515 22967
rect 8110 22964 8116 22976
rect 6503 22936 8116 22964
rect 6503 22933 6515 22936
rect 6457 22927 6515 22933
rect 8110 22924 8116 22936
rect 8168 22924 8174 22976
rect 8202 22924 8208 22976
rect 8260 22964 8266 22976
rect 8297 22967 8355 22973
rect 8297 22964 8309 22967
rect 8260 22936 8309 22964
rect 8260 22924 8266 22936
rect 8297 22933 8309 22936
rect 8343 22933 8355 22967
rect 8297 22927 8355 22933
rect 10226 22924 10232 22976
rect 10284 22964 10290 22976
rect 11164 22964 11192 23004
rect 11330 22992 11336 23004
rect 11388 22992 11394 23044
rect 11701 23035 11759 23041
rect 11701 23001 11713 23035
rect 11747 23032 11759 23035
rect 11790 23032 11796 23044
rect 11747 23004 11796 23032
rect 11747 23001 11759 23004
rect 11701 22995 11759 23001
rect 11790 22992 11796 23004
rect 11848 22992 11854 23044
rect 12894 23032 12900 23044
rect 12855 23004 12900 23032
rect 12894 22992 12900 23004
rect 12952 22992 12958 23044
rect 13081 23035 13139 23041
rect 13081 23001 13093 23035
rect 13127 23001 13139 23035
rect 13081 22995 13139 23001
rect 11514 22964 11520 22976
rect 10284 22936 10329 22964
rect 11164 22936 11520 22964
rect 10284 22924 10290 22936
rect 11514 22924 11520 22936
rect 11572 22964 11578 22976
rect 13096 22964 13124 22995
rect 13170 22992 13176 23044
rect 13228 23032 13234 23044
rect 14200 23032 14228 23063
rect 15102 23060 15108 23072
rect 15160 23060 15166 23112
rect 15286 23100 15292 23112
rect 15247 23072 15292 23100
rect 15286 23060 15292 23072
rect 15344 23060 15350 23112
rect 18414 23100 18420 23112
rect 18375 23072 18420 23100
rect 18414 23060 18420 23072
rect 18472 23060 18478 23112
rect 22925 23103 22983 23109
rect 22925 23069 22937 23103
rect 22971 23100 22983 23103
rect 23201 23103 23259 23109
rect 23201 23100 23213 23103
rect 22971 23072 23213 23100
rect 22971 23069 22983 23072
rect 22925 23063 22983 23069
rect 23201 23069 23213 23072
rect 23247 23069 23259 23103
rect 23201 23063 23259 23069
rect 13228 23004 14228 23032
rect 13228 22992 13234 23004
rect 11572 22936 13124 22964
rect 14200 22964 14228 23004
rect 16672 23044 16724 23050
rect 16758 22992 16764 23044
rect 16816 23032 16822 23044
rect 17126 23032 17132 23044
rect 16816 23004 17132 23032
rect 16816 22992 16822 23004
rect 17126 22992 17132 23004
rect 17184 22992 17190 23044
rect 18690 23032 18696 23044
rect 18651 23004 18696 23032
rect 18690 22992 18696 23004
rect 18748 22992 18754 23044
rect 21818 22992 21824 23044
rect 21876 22992 21882 23044
rect 22462 23032 22468 23044
rect 22423 23004 22468 23032
rect 22462 22992 22468 23004
rect 22520 22992 22526 23044
rect 22554 22992 22560 23044
rect 22612 23032 22618 23044
rect 22940 23032 22968 23063
rect 23290 23060 23296 23112
rect 23348 23100 23354 23112
rect 23860 23109 23888 23208
rect 23477 23103 23535 23109
rect 23477 23100 23489 23103
rect 23348 23072 23489 23100
rect 23348 23060 23354 23072
rect 23477 23069 23489 23072
rect 23523 23069 23535 23103
rect 23477 23063 23535 23069
rect 23850 23103 23908 23109
rect 23850 23069 23862 23103
rect 23896 23069 23908 23103
rect 23850 23063 23908 23069
rect 22612 23004 22968 23032
rect 23661 23035 23719 23041
rect 22612 22992 22618 23004
rect 23661 23001 23673 23035
rect 23707 23001 23719 23035
rect 23661 22995 23719 23001
rect 23753 23035 23811 23041
rect 23753 23001 23765 23035
rect 23799 23032 23811 23035
rect 24489 23035 24547 23041
rect 24489 23032 24501 23035
rect 23799 23004 24501 23032
rect 23799 23001 23811 23004
rect 23753 22995 23811 23001
rect 24489 23001 24501 23004
rect 24535 23032 24547 23035
rect 26234 23032 26240 23044
rect 24535 23004 26240 23032
rect 24535 23001 24547 23004
rect 24489 22995 24547 23001
rect 16672 22986 16724 22992
rect 14921 22967 14979 22973
rect 14921 22964 14933 22967
rect 14200 22936 14933 22964
rect 11572 22924 11578 22936
rect 14921 22933 14933 22936
rect 14967 22933 14979 22967
rect 19610 22964 19616 22976
rect 19571 22936 19616 22964
rect 14921 22927 14979 22933
rect 19610 22924 19616 22936
rect 19668 22924 19674 22976
rect 19702 22924 19708 22976
rect 19760 22964 19766 22976
rect 19760 22936 19805 22964
rect 19760 22924 19766 22936
rect 23014 22924 23020 22976
rect 23072 22964 23078 22976
rect 23198 22964 23204 22976
rect 23072 22936 23204 22964
rect 23072 22924 23078 22936
rect 23198 22924 23204 22936
rect 23256 22924 23262 22976
rect 23676 22964 23704 22995
rect 26234 22992 26240 23004
rect 26292 22992 26298 23044
rect 23842 22964 23848 22976
rect 23676 22936 23848 22964
rect 23842 22924 23848 22936
rect 23900 22924 23906 22976
rect 24046 22967 24104 22973
rect 24046 22933 24058 22967
rect 24092 22964 24104 22967
rect 24210 22964 24216 22976
rect 24092 22936 24216 22964
rect 24092 22933 24104 22936
rect 24046 22927 24104 22933
rect 24210 22924 24216 22936
rect 24268 22924 24274 22976
rect 1104 22874 29440 22896
rect 1104 22822 10395 22874
rect 10447 22822 10459 22874
rect 10511 22822 10523 22874
rect 10575 22822 10587 22874
rect 10639 22822 10651 22874
rect 10703 22822 19840 22874
rect 19892 22822 19904 22874
rect 19956 22822 19968 22874
rect 20020 22822 20032 22874
rect 20084 22822 20096 22874
rect 20148 22822 29440 22874
rect 1104 22800 29440 22822
rect 2777 22763 2835 22769
rect 2777 22729 2789 22763
rect 2823 22760 2835 22763
rect 3050 22760 3056 22772
rect 2823 22732 3056 22760
rect 2823 22729 2835 22732
rect 2777 22723 2835 22729
rect 3050 22720 3056 22732
rect 3108 22720 3114 22772
rect 4338 22760 4344 22772
rect 3160 22732 4344 22760
rect 2866 22692 2872 22704
rect 1412 22664 2872 22692
rect 1412 22633 1440 22664
rect 2866 22652 2872 22664
rect 2924 22652 2930 22704
rect 3160 22701 3188 22732
rect 4338 22720 4344 22732
rect 4396 22720 4402 22772
rect 4430 22720 4436 22772
rect 4488 22760 4494 22772
rect 4525 22763 4583 22769
rect 4525 22760 4537 22763
rect 4488 22732 4537 22760
rect 4488 22720 4494 22732
rect 4525 22729 4537 22732
rect 4571 22729 4583 22763
rect 7190 22760 7196 22772
rect 7151 22732 7196 22760
rect 4525 22723 4583 22729
rect 7190 22720 7196 22732
rect 7248 22720 7254 22772
rect 7926 22720 7932 22772
rect 7984 22760 7990 22772
rect 8832 22763 8890 22769
rect 8832 22760 8844 22763
rect 7984 22732 8844 22760
rect 7984 22720 7990 22732
rect 8832 22729 8844 22732
rect 8878 22729 8890 22763
rect 9766 22760 9772 22772
rect 9727 22732 9772 22760
rect 8832 22723 8890 22729
rect 9766 22720 9772 22732
rect 9824 22720 9830 22772
rect 9858 22720 9864 22772
rect 9916 22760 9922 22772
rect 13265 22763 13323 22769
rect 9916 22732 11100 22760
rect 9916 22720 9922 22732
rect 3145 22695 3203 22701
rect 3145 22661 3157 22695
rect 3191 22661 3203 22695
rect 3145 22655 3203 22661
rect 3329 22695 3387 22701
rect 3329 22661 3341 22695
rect 3375 22692 3387 22695
rect 4246 22692 4252 22704
rect 3375 22664 4252 22692
rect 3375 22661 3387 22664
rect 3329 22655 3387 22661
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 7742 22692 7748 22704
rect 7484 22664 7748 22692
rect 1670 22633 1676 22636
rect 1397 22627 1455 22633
rect 1397 22593 1409 22627
rect 1443 22593 1455 22627
rect 1664 22624 1676 22633
rect 1631 22596 1676 22624
rect 1397 22587 1455 22593
rect 1664 22587 1676 22596
rect 1670 22584 1676 22587
rect 1728 22584 1734 22636
rect 3786 22584 3792 22636
rect 3844 22624 3850 22636
rect 3881 22627 3939 22633
rect 3881 22624 3893 22627
rect 3844 22596 3893 22624
rect 3844 22584 3850 22596
rect 3881 22593 3893 22596
rect 3927 22593 3939 22627
rect 3881 22587 3939 22593
rect 3970 22584 3976 22636
rect 4028 22624 4034 22636
rect 4065 22627 4123 22633
rect 4065 22624 4077 22627
rect 4028 22596 4077 22624
rect 4028 22584 4034 22596
rect 4065 22593 4077 22596
rect 4111 22593 4123 22627
rect 4065 22587 4123 22593
rect 4154 22584 4160 22636
rect 4212 22624 4218 22636
rect 7484 22633 7512 22664
rect 7742 22652 7748 22664
rect 7800 22692 7806 22704
rect 9125 22695 9183 22701
rect 9125 22692 9137 22695
rect 7800 22664 8432 22692
rect 7800 22652 7806 22664
rect 4893 22627 4951 22633
rect 4893 22624 4905 22627
rect 4212 22596 4257 22624
rect 4356 22596 4905 22624
rect 4212 22584 4218 22596
rect 3418 22516 3424 22568
rect 3476 22556 3482 22568
rect 4249 22559 4307 22565
rect 4249 22556 4261 22559
rect 3476 22528 4261 22556
rect 3476 22516 3482 22528
rect 4249 22525 4261 22528
rect 4295 22525 4307 22559
rect 4249 22519 4307 22525
rect 3697 22491 3755 22497
rect 3697 22457 3709 22491
rect 3743 22488 3755 22491
rect 4356 22488 4384 22596
rect 4893 22593 4905 22596
rect 4939 22593 4951 22627
rect 4893 22587 4951 22593
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22593 7435 22627
rect 7377 22587 7435 22593
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22593 7527 22627
rect 7469 22587 7527 22593
rect 7837 22627 7895 22633
rect 7837 22593 7849 22627
rect 7883 22624 7895 22627
rect 7929 22627 7987 22633
rect 7929 22624 7941 22627
rect 7883 22596 7941 22624
rect 7883 22593 7895 22596
rect 7837 22587 7895 22593
rect 7929 22593 7941 22596
rect 7975 22593 7987 22627
rect 7929 22587 7987 22593
rect 7392 22556 7420 22587
rect 8110 22584 8116 22636
rect 8168 22624 8174 22636
rect 8404 22633 8432 22664
rect 8496 22664 9137 22692
rect 8389 22627 8447 22633
rect 8168 22596 8340 22624
rect 8168 22584 8174 22596
rect 8312 22556 8340 22596
rect 8389 22593 8401 22627
rect 8435 22593 8447 22627
rect 8389 22587 8447 22593
rect 8496 22556 8524 22664
rect 9125 22661 9137 22664
rect 9171 22661 9183 22695
rect 9125 22655 9183 22661
rect 9217 22695 9275 22701
rect 9217 22661 9229 22695
rect 9263 22692 9275 22695
rect 9263 22664 9536 22692
rect 9263 22661 9275 22664
rect 9217 22655 9275 22661
rect 9028 22627 9086 22633
rect 9028 22593 9040 22627
rect 9074 22593 9086 22627
rect 9398 22624 9404 22636
rect 9359 22596 9404 22624
rect 9028 22587 9086 22593
rect 7392 22528 8248 22556
rect 8312 22528 8524 22556
rect 9048 22556 9076 22587
rect 9398 22584 9404 22596
rect 9456 22584 9462 22636
rect 9508 22624 9536 22664
rect 9582 22652 9588 22704
rect 9640 22692 9646 22704
rect 9953 22695 10011 22701
rect 9640 22664 9685 22692
rect 9640 22652 9646 22664
rect 9953 22661 9965 22695
rect 9999 22692 10011 22695
rect 10410 22692 10416 22704
rect 9999 22664 10416 22692
rect 9999 22661 10011 22664
rect 9953 22655 10011 22661
rect 10410 22652 10416 22664
rect 10468 22652 10474 22704
rect 10870 22652 10876 22704
rect 10928 22692 10934 22704
rect 11072 22701 11100 22732
rect 13265 22729 13277 22763
rect 13311 22729 13323 22763
rect 13265 22723 13323 22729
rect 11057 22695 11115 22701
rect 10928 22664 11008 22692
rect 10928 22652 10934 22664
rect 10980 22633 11008 22664
rect 11057 22661 11069 22695
rect 11103 22661 11115 22695
rect 11057 22655 11115 22661
rect 11149 22695 11207 22701
rect 11149 22661 11161 22695
rect 11195 22692 11207 22695
rect 12434 22692 12440 22704
rect 11195 22664 12440 22692
rect 11195 22661 11207 22664
rect 11149 22655 11207 22661
rect 10321 22627 10379 22633
rect 10321 22624 10333 22627
rect 9508 22596 10333 22624
rect 10321 22593 10333 22596
rect 10367 22624 10379 22627
rect 10960 22627 11018 22633
rect 10367 22596 10916 22624
rect 10367 22593 10379 22596
rect 10321 22587 10379 22593
rect 10888 22556 10916 22596
rect 10960 22593 10972 22627
rect 11006 22593 11018 22627
rect 11330 22624 11336 22636
rect 11291 22596 11336 22624
rect 10960 22587 11018 22593
rect 11330 22584 11336 22596
rect 11388 22584 11394 22636
rect 11514 22624 11520 22636
rect 11475 22596 11520 22624
rect 11514 22584 11520 22596
rect 11572 22584 11578 22636
rect 11606 22584 11612 22636
rect 11664 22584 11670 22636
rect 11992 22633 12020 22664
rect 12434 22652 12440 22664
rect 12492 22692 12498 22704
rect 12618 22692 12624 22704
rect 12492 22664 12624 22692
rect 12492 22652 12498 22664
rect 12618 22652 12624 22664
rect 12676 22652 12682 22704
rect 11977 22627 12035 22633
rect 11977 22593 11989 22627
rect 12023 22593 12035 22627
rect 11977 22587 12035 22593
rect 13081 22627 13139 22633
rect 13081 22593 13093 22627
rect 13127 22624 13139 22627
rect 13170 22624 13176 22636
rect 13127 22596 13176 22624
rect 13127 22593 13139 22596
rect 13081 22587 13139 22593
rect 13170 22584 13176 22596
rect 13228 22584 13234 22636
rect 13280 22624 13308 22723
rect 15654 22720 15660 22772
rect 15712 22760 15718 22772
rect 19613 22763 19671 22769
rect 15712 22732 19564 22760
rect 15712 22720 15718 22732
rect 15286 22652 15292 22704
rect 15344 22692 15350 22704
rect 16850 22692 16856 22704
rect 15344 22664 16856 22692
rect 15344 22652 15350 22664
rect 16850 22652 16856 22664
rect 16908 22692 16914 22704
rect 16908 22664 17080 22692
rect 16908 22652 16914 22664
rect 13541 22627 13599 22633
rect 13541 22624 13553 22627
rect 13280 22596 13553 22624
rect 13541 22593 13553 22596
rect 13587 22593 13599 22627
rect 13541 22587 13599 22593
rect 14461 22627 14519 22633
rect 14461 22593 14473 22627
rect 14507 22593 14519 22627
rect 14921 22627 14979 22633
rect 14921 22624 14933 22627
rect 14461 22587 14519 22593
rect 14660 22596 14933 22624
rect 11624 22556 11652 22584
rect 9048 22528 10824 22556
rect 10888 22528 11652 22556
rect 3743 22460 4384 22488
rect 3743 22457 3755 22460
rect 3697 22451 3755 22457
rect 4430 22448 4436 22500
rect 4488 22488 4494 22500
rect 8220 22497 8248 22528
rect 4709 22491 4767 22497
rect 4709 22488 4721 22491
rect 4488 22460 4721 22488
rect 4488 22448 4494 22460
rect 4709 22457 4721 22460
rect 4755 22457 4767 22491
rect 4709 22451 4767 22457
rect 7653 22491 7711 22497
rect 7653 22457 7665 22491
rect 7699 22488 7711 22491
rect 7837 22491 7895 22497
rect 7837 22488 7849 22491
rect 7699 22460 7849 22488
rect 7699 22457 7711 22460
rect 7653 22451 7711 22457
rect 7837 22457 7849 22460
rect 7883 22457 7895 22491
rect 7837 22451 7895 22457
rect 8205 22491 8263 22497
rect 8205 22457 8217 22491
rect 8251 22457 8263 22491
rect 8205 22451 8263 22457
rect 9674 22448 9680 22500
rect 9732 22488 9738 22500
rect 10137 22491 10195 22497
rect 10137 22488 10149 22491
rect 9732 22460 10149 22488
rect 9732 22448 9738 22460
rect 10137 22457 10149 22460
rect 10183 22488 10195 22491
rect 10686 22488 10692 22500
rect 10183 22460 10692 22488
rect 10183 22457 10195 22460
rect 10137 22451 10195 22457
rect 10686 22448 10692 22460
rect 10744 22448 10750 22500
rect 10796 22488 10824 22528
rect 11698 22516 11704 22568
rect 11756 22556 11762 22568
rect 12069 22559 12127 22565
rect 12069 22556 12081 22559
rect 11756 22528 12081 22556
rect 11756 22516 11762 22528
rect 12069 22525 12081 22528
rect 12115 22525 12127 22559
rect 12069 22519 12127 22525
rect 12253 22559 12311 22565
rect 12253 22525 12265 22559
rect 12299 22525 12311 22559
rect 13188 22556 13216 22584
rect 14476 22556 14504 22587
rect 13188 22528 14504 22556
rect 12253 22519 12311 22525
rect 11606 22488 11612 22500
rect 10796 22460 11468 22488
rect 11567 22460 11612 22488
rect 3050 22420 3056 22432
rect 3011 22392 3056 22420
rect 3050 22380 3056 22392
rect 3108 22380 3114 22432
rect 3878 22420 3884 22432
rect 3839 22392 3884 22420
rect 3878 22380 3884 22392
rect 3936 22380 3942 22432
rect 4246 22420 4252 22432
rect 4207 22392 4252 22420
rect 4246 22380 4252 22392
rect 4304 22380 4310 22432
rect 7926 22380 7932 22432
rect 7984 22420 7990 22432
rect 8113 22423 8171 22429
rect 8113 22420 8125 22423
rect 7984 22392 8125 22420
rect 7984 22380 7990 22392
rect 8113 22389 8125 22392
rect 8159 22389 8171 22423
rect 8113 22383 8171 22389
rect 10781 22423 10839 22429
rect 10781 22389 10793 22423
rect 10827 22420 10839 22423
rect 11054 22420 11060 22432
rect 10827 22392 11060 22420
rect 10827 22389 10839 22392
rect 10781 22383 10839 22389
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 11440 22420 11468 22460
rect 11606 22448 11612 22460
rect 11664 22448 11670 22500
rect 11790 22448 11796 22500
rect 11848 22488 11854 22500
rect 12268 22488 12296 22519
rect 12526 22488 12532 22500
rect 11848 22460 12296 22488
rect 12406 22460 12532 22488
rect 11848 22448 11854 22460
rect 12406 22420 12434 22460
rect 12526 22448 12532 22460
rect 12584 22448 12590 22500
rect 14660 22497 14688 22596
rect 14921 22593 14933 22596
rect 14967 22593 14979 22627
rect 14921 22587 14979 22593
rect 15102 22584 15108 22636
rect 15160 22624 15166 22636
rect 15470 22624 15476 22636
rect 15160 22596 15476 22624
rect 15160 22584 15166 22596
rect 15470 22584 15476 22596
rect 15528 22624 15534 22636
rect 15565 22627 15623 22633
rect 15565 22624 15577 22627
rect 15528 22596 15577 22624
rect 15528 22584 15534 22596
rect 15565 22593 15577 22596
rect 15611 22624 15623 22627
rect 15838 22624 15844 22636
rect 15611 22596 15844 22624
rect 15611 22593 15623 22596
rect 15565 22587 15623 22593
rect 15838 22584 15844 22596
rect 15896 22584 15902 22636
rect 17052 22633 17080 22664
rect 18690 22652 18696 22704
rect 18748 22692 18754 22704
rect 19536 22692 19564 22732
rect 19613 22729 19625 22763
rect 19659 22760 19671 22763
rect 19702 22760 19708 22772
rect 19659 22732 19708 22760
rect 19659 22729 19671 22732
rect 19613 22723 19671 22729
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 21726 22760 21732 22772
rect 20824 22732 21732 22760
rect 20824 22692 20852 22732
rect 21726 22720 21732 22732
rect 21784 22720 21790 22772
rect 21821 22763 21879 22769
rect 21821 22729 21833 22763
rect 21867 22760 21879 22763
rect 22002 22760 22008 22772
rect 21867 22732 22008 22760
rect 21867 22729 21879 22732
rect 21821 22723 21879 22729
rect 22002 22720 22008 22732
rect 22060 22720 22066 22772
rect 22646 22720 22652 22772
rect 22704 22760 22710 22772
rect 22741 22763 22799 22769
rect 22741 22760 22753 22763
rect 22704 22732 22753 22760
rect 22704 22720 22710 22732
rect 22741 22729 22753 22732
rect 22787 22760 22799 22763
rect 22830 22760 22836 22772
rect 22787 22732 22836 22760
rect 22787 22729 22799 22732
rect 22741 22723 22799 22729
rect 22830 22720 22836 22732
rect 22888 22720 22894 22772
rect 18748 22664 19104 22692
rect 19536 22664 20852 22692
rect 18748 22652 18754 22664
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22593 17095 22627
rect 17037 22587 17095 22593
rect 17304 22627 17362 22633
rect 17304 22593 17316 22627
rect 17350 22624 17362 22627
rect 18601 22627 18659 22633
rect 18601 22624 18613 22627
rect 17350 22596 18613 22624
rect 17350 22593 17362 22596
rect 17304 22587 17362 22593
rect 18601 22593 18613 22596
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 18785 22627 18843 22633
rect 18785 22593 18797 22627
rect 18831 22593 18843 22627
rect 18966 22624 18972 22636
rect 18927 22596 18972 22624
rect 18785 22587 18843 22593
rect 18800 22556 18828 22587
rect 18966 22584 18972 22596
rect 19024 22584 19030 22636
rect 19076 22624 19104 22664
rect 20898 22652 20904 22704
rect 20956 22692 20962 22704
rect 20956 22664 21128 22692
rect 20956 22652 20962 22664
rect 19154 22627 19212 22633
rect 19154 22624 19166 22627
rect 19076 22596 19166 22624
rect 19154 22593 19166 22596
rect 19200 22593 19212 22627
rect 19154 22587 19212 22593
rect 19337 22627 19395 22633
rect 19337 22593 19349 22627
rect 19383 22593 19395 22627
rect 20714 22624 20720 22636
rect 20772 22633 20778 22636
rect 20684 22596 20720 22624
rect 19337 22587 19395 22593
rect 19058 22556 19064 22568
rect 18524 22528 18828 22556
rect 19019 22528 19064 22556
rect 14645 22491 14703 22497
rect 14645 22457 14657 22491
rect 14691 22457 14703 22491
rect 14645 22451 14703 22457
rect 18524 22432 18552 22528
rect 19058 22516 19064 22528
rect 19116 22516 19122 22568
rect 19242 22448 19248 22500
rect 19300 22488 19306 22500
rect 19352 22488 19380 22587
rect 20714 22584 20720 22596
rect 20772 22587 20784 22633
rect 20990 22624 20996 22636
rect 20951 22596 20996 22624
rect 20772 22584 20778 22587
rect 20990 22584 20996 22596
rect 21048 22584 21054 22636
rect 21100 22633 21128 22664
rect 21376 22664 24702 22692
rect 21085 22627 21143 22633
rect 21085 22593 21097 22627
rect 21131 22593 21143 22627
rect 21085 22587 21143 22593
rect 19300 22460 19380 22488
rect 21269 22491 21327 22497
rect 19300 22448 19306 22460
rect 21269 22457 21281 22491
rect 21315 22488 21327 22491
rect 21376 22488 21404 22664
rect 22002 22624 22008 22636
rect 21963 22596 22008 22624
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 22097 22627 22155 22633
rect 22097 22593 22109 22627
rect 22143 22624 22155 22627
rect 22186 22624 22192 22636
rect 22143 22596 22192 22624
rect 22143 22593 22155 22596
rect 22097 22587 22155 22593
rect 22186 22584 22192 22596
rect 22244 22584 22250 22636
rect 22554 22624 22560 22636
rect 22515 22596 22560 22624
rect 22554 22584 22560 22596
rect 22612 22584 22618 22636
rect 22738 22584 22744 22636
rect 22796 22624 22802 22636
rect 23017 22627 23075 22633
rect 23017 22624 23029 22627
rect 22796 22596 23029 22624
rect 22796 22584 22802 22596
rect 23017 22593 23029 22596
rect 23063 22593 23075 22627
rect 23017 22587 23075 22593
rect 23750 22584 23756 22636
rect 23808 22624 23814 22636
rect 23937 22627 23995 22633
rect 23937 22624 23949 22627
rect 23808 22596 23949 22624
rect 23808 22584 23814 22596
rect 23937 22593 23949 22596
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 24210 22556 24216 22568
rect 24171 22528 24216 22556
rect 24210 22516 24216 22528
rect 24268 22516 24274 22568
rect 21315 22460 21404 22488
rect 22833 22491 22891 22497
rect 21315 22457 21327 22460
rect 21269 22451 21327 22457
rect 22833 22457 22845 22491
rect 22879 22488 22891 22491
rect 23290 22488 23296 22500
rect 22879 22460 23296 22488
rect 22879 22457 22891 22460
rect 22833 22451 22891 22457
rect 11440 22392 12434 22420
rect 13354 22380 13360 22432
rect 13412 22420 13418 22432
rect 13412 22392 13457 22420
rect 13412 22380 13418 22392
rect 14734 22380 14740 22432
rect 14792 22420 14798 22432
rect 14792 22392 14837 22420
rect 14792 22380 14798 22392
rect 15654 22380 15660 22432
rect 15712 22420 15718 22432
rect 15749 22423 15807 22429
rect 15749 22420 15761 22423
rect 15712 22392 15761 22420
rect 15712 22380 15718 22392
rect 15749 22389 15761 22392
rect 15795 22389 15807 22423
rect 15749 22383 15807 22389
rect 15838 22380 15844 22432
rect 15896 22420 15902 22432
rect 16025 22423 16083 22429
rect 16025 22420 16037 22423
rect 15896 22392 16037 22420
rect 15896 22380 15902 22392
rect 16025 22389 16037 22392
rect 16071 22389 16083 22423
rect 16025 22383 16083 22389
rect 18417 22423 18475 22429
rect 18417 22389 18429 22423
rect 18463 22420 18475 22423
rect 18506 22420 18512 22432
rect 18463 22392 18512 22420
rect 18463 22389 18475 22392
rect 18417 22383 18475 22389
rect 18506 22380 18512 22392
rect 18564 22380 18570 22432
rect 20622 22380 20628 22432
rect 20680 22420 20686 22432
rect 21284 22420 21312 22451
rect 23290 22448 23296 22460
rect 23348 22448 23354 22500
rect 22278 22420 22284 22432
rect 20680 22392 21312 22420
rect 22239 22392 22284 22420
rect 20680 22380 20686 22392
rect 22278 22380 22284 22392
rect 22336 22380 22342 22432
rect 25685 22423 25743 22429
rect 25685 22389 25697 22423
rect 25731 22420 25743 22423
rect 26234 22420 26240 22432
rect 25731 22392 26240 22420
rect 25731 22389 25743 22392
rect 25685 22383 25743 22389
rect 26234 22380 26240 22392
rect 26292 22380 26298 22432
rect 1104 22330 29440 22352
rect 1104 22278 5672 22330
rect 5724 22278 5736 22330
rect 5788 22278 5800 22330
rect 5852 22278 5864 22330
rect 5916 22278 5928 22330
rect 5980 22278 15118 22330
rect 15170 22278 15182 22330
rect 15234 22278 15246 22330
rect 15298 22278 15310 22330
rect 15362 22278 15374 22330
rect 15426 22278 24563 22330
rect 24615 22278 24627 22330
rect 24679 22278 24691 22330
rect 24743 22278 24755 22330
rect 24807 22278 24819 22330
rect 24871 22278 29440 22330
rect 1104 22256 29440 22278
rect 3418 22176 3424 22228
rect 3476 22216 3482 22228
rect 3789 22219 3847 22225
rect 3789 22216 3801 22219
rect 3476 22188 3801 22216
rect 3476 22176 3482 22188
rect 3789 22185 3801 22188
rect 3835 22185 3847 22219
rect 3789 22179 3847 22185
rect 7180 22219 7238 22225
rect 7180 22185 7192 22219
rect 7226 22216 7238 22219
rect 9033 22219 9091 22225
rect 9033 22216 9045 22219
rect 7226 22188 9045 22216
rect 7226 22185 7238 22188
rect 7180 22179 7238 22185
rect 9033 22185 9045 22188
rect 9079 22185 9091 22219
rect 9033 22179 9091 22185
rect 9398 22176 9404 22228
rect 9456 22216 9462 22228
rect 12802 22216 12808 22228
rect 9456 22188 12808 22216
rect 9456 22176 9462 22188
rect 12802 22176 12808 22188
rect 12860 22176 12866 22228
rect 15010 22176 15016 22228
rect 15068 22216 15074 22228
rect 19334 22216 19340 22228
rect 15068 22188 19340 22216
rect 15068 22176 15074 22188
rect 19334 22176 19340 22188
rect 19392 22176 19398 22228
rect 21256 22219 21314 22225
rect 21256 22185 21268 22219
rect 21302 22216 21314 22219
rect 22370 22216 22376 22228
rect 21302 22188 22376 22216
rect 21302 22185 21314 22188
rect 21256 22179 21314 22185
rect 22370 22176 22376 22188
rect 22428 22176 22434 22228
rect 22462 22176 22468 22228
rect 22520 22216 22526 22228
rect 25590 22216 25596 22228
rect 22520 22188 25596 22216
rect 22520 22176 22526 22188
rect 25590 22176 25596 22188
rect 25648 22176 25654 22228
rect 2866 22108 2872 22160
rect 2924 22108 2930 22160
rect 9950 22108 9956 22160
rect 10008 22148 10014 22160
rect 10226 22148 10232 22160
rect 10008 22120 10232 22148
rect 10008 22108 10014 22120
rect 10226 22108 10232 22120
rect 10284 22108 10290 22160
rect 10594 22148 10600 22160
rect 10352 22120 10600 22148
rect 2884 22080 2912 22108
rect 2884 22052 4752 22080
rect 4724 22024 4752 22052
rect 8202 22040 8208 22092
rect 8260 22080 8266 22092
rect 9766 22080 9772 22092
rect 8260 22052 9772 22080
rect 8260 22040 8266 22052
rect 9766 22040 9772 22052
rect 9824 22040 9830 22092
rect 10352 22080 10380 22120
rect 10594 22108 10600 22120
rect 10652 22148 10658 22160
rect 10652 22120 11100 22148
rect 10652 22108 10658 22120
rect 11072 22089 11100 22120
rect 11514 22108 11520 22160
rect 11572 22148 11578 22160
rect 11701 22151 11759 22157
rect 11701 22148 11713 22151
rect 11572 22120 11713 22148
rect 11572 22108 11578 22120
rect 11701 22117 11713 22120
rect 11747 22117 11759 22151
rect 11701 22111 11759 22117
rect 9951 22052 10380 22080
rect 10781 22083 10839 22089
rect 2774 21972 2780 22024
rect 2832 22012 2838 22024
rect 2869 22015 2927 22021
rect 2869 22012 2881 22015
rect 2832 21984 2881 22012
rect 2832 21972 2838 21984
rect 2869 21981 2881 21984
rect 2915 21981 2927 22015
rect 2869 21975 2927 21981
rect 3878 21972 3884 22024
rect 3936 22012 3942 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3936 21984 3985 22012
rect 3936 21972 3942 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 4065 22015 4123 22021
rect 4065 21981 4077 22015
rect 4111 22012 4123 22015
rect 4154 22012 4160 22024
rect 4111 21984 4160 22012
rect 4111 21981 4123 21984
rect 4065 21975 4123 21981
rect 4154 21972 4160 21984
rect 4212 22012 4218 22024
rect 4430 22012 4436 22024
rect 4212 21984 4436 22012
rect 4212 21972 4218 21984
rect 4430 21972 4436 21984
rect 4488 21972 4494 22024
rect 4706 21972 4712 22024
rect 4764 22012 4770 22024
rect 4893 22015 4951 22021
rect 4893 22012 4905 22015
rect 4764 21984 4905 22012
rect 4764 21972 4770 21984
rect 4893 21981 4905 21984
rect 4939 22012 4951 22015
rect 6914 22012 6920 22024
rect 4939 21984 6920 22012
rect 4939 21981 4951 21984
rect 4893 21975 4951 21981
rect 6914 21972 6920 21984
rect 6972 21972 6978 22024
rect 8938 21972 8944 22024
rect 8996 22012 9002 22024
rect 9171 22015 9229 22021
rect 9171 22012 9183 22015
rect 8996 21984 9183 22012
rect 8996 21972 9002 21984
rect 9171 21981 9183 21984
rect 9217 21981 9229 22015
rect 9171 21975 9229 21981
rect 9306 21972 9312 22024
rect 9364 22012 9370 22024
rect 9582 22012 9588 22024
rect 9364 21984 9409 22012
rect 9543 21984 9588 22012
rect 9364 21972 9370 21984
rect 9582 21972 9588 21984
rect 9640 21972 9646 22024
rect 9951 22021 9979 22052
rect 10781 22049 10793 22083
rect 10827 22080 10839 22083
rect 11057 22083 11115 22089
rect 10827 22052 10916 22080
rect 10827 22049 10839 22052
rect 10781 22043 10839 22049
rect 10888 22024 10916 22052
rect 11057 22049 11069 22083
rect 11103 22080 11115 22083
rect 15028 22080 15056 22176
rect 15105 22151 15163 22157
rect 15105 22117 15117 22151
rect 15151 22148 15163 22151
rect 15470 22148 15476 22160
rect 15151 22120 15476 22148
rect 15151 22117 15163 22120
rect 15105 22111 15163 22117
rect 15470 22108 15476 22120
rect 15528 22108 15534 22160
rect 23485 22151 23543 22157
rect 23485 22117 23497 22151
rect 23531 22117 23543 22151
rect 23485 22111 23543 22117
rect 11103 22052 15056 22080
rect 15565 22083 15623 22089
rect 11103 22049 11115 22052
rect 11057 22043 11115 22049
rect 15565 22049 15577 22083
rect 15611 22080 15623 22083
rect 16482 22080 16488 22092
rect 15611 22052 16488 22080
rect 15611 22049 15623 22052
rect 15565 22043 15623 22049
rect 16482 22040 16488 22052
rect 16540 22040 16546 22092
rect 18506 22080 18512 22092
rect 18467 22052 18512 22080
rect 18506 22040 18512 22052
rect 18564 22040 18570 22092
rect 18601 22083 18659 22089
rect 18601 22049 18613 22083
rect 18647 22080 18659 22083
rect 18782 22080 18788 22092
rect 18647 22052 18788 22080
rect 18647 22049 18659 22052
rect 18601 22043 18659 22049
rect 9951 22015 10011 22021
rect 9951 21984 9965 22015
rect 9953 21981 9965 21984
rect 9999 21981 10011 22015
rect 10413 22015 10471 22021
rect 10413 22012 10425 22015
rect 9953 21975 10011 21981
rect 10060 21984 10425 22012
rect 5160 21947 5218 21953
rect 3068 21916 4384 21944
rect 3068 21885 3096 21916
rect 4356 21888 4384 21916
rect 5160 21913 5172 21947
rect 5206 21944 5218 21947
rect 5350 21944 5356 21956
rect 5206 21916 5356 21944
rect 5206 21913 5218 21916
rect 5160 21907 5218 21913
rect 5350 21904 5356 21916
rect 5408 21904 5414 21956
rect 6454 21944 6460 21956
rect 5460 21916 6460 21944
rect 3053 21879 3111 21885
rect 3053 21845 3065 21879
rect 3099 21845 3111 21879
rect 3053 21839 3111 21845
rect 4157 21879 4215 21885
rect 4157 21845 4169 21879
rect 4203 21876 4215 21879
rect 4246 21876 4252 21888
rect 4203 21848 4252 21876
rect 4203 21845 4215 21848
rect 4157 21839 4215 21845
rect 4246 21836 4252 21848
rect 4304 21836 4310 21888
rect 4338 21836 4344 21888
rect 4396 21876 4402 21888
rect 5460 21876 5488 21916
rect 6454 21904 6460 21916
rect 6512 21904 6518 21956
rect 7926 21904 7932 21956
rect 7984 21904 7990 21956
rect 9677 21947 9735 21953
rect 9677 21944 9689 21947
rect 8680 21916 9689 21944
rect 6270 21876 6276 21888
rect 4396 21848 5488 21876
rect 6231 21848 6276 21876
rect 4396 21836 4402 21848
rect 6270 21836 6276 21848
rect 6328 21836 6334 21888
rect 8680 21885 8708 21916
rect 9677 21913 9689 21916
rect 9723 21944 9735 21947
rect 10060 21944 10088 21984
rect 10413 21981 10425 21984
rect 10459 21981 10471 22015
rect 10413 21975 10471 21981
rect 10686 21972 10692 22024
rect 10744 22012 10750 22024
rect 10744 21984 10789 22012
rect 10744 21972 10750 21984
rect 10870 21972 10876 22024
rect 10928 21972 10934 22024
rect 11514 21972 11520 22024
rect 11572 22012 11578 22024
rect 11885 22015 11943 22021
rect 11885 22012 11897 22015
rect 11572 21984 11897 22012
rect 11572 21972 11578 21984
rect 11885 21981 11897 21984
rect 11931 21981 11943 22015
rect 11885 21975 11943 21981
rect 13262 21972 13268 22024
rect 13320 21972 13326 22024
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 22012 15071 22015
rect 15194 22012 15200 22024
rect 15059 21984 15200 22012
rect 15059 21981 15071 21984
rect 15013 21975 15071 21981
rect 15194 21972 15200 21984
rect 15252 21972 15258 22024
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 21981 15347 22015
rect 18616 22012 18644 22043
rect 18782 22040 18788 22052
rect 18840 22040 18846 22092
rect 19058 22040 19064 22092
rect 19116 22080 19122 22092
rect 19521 22083 19579 22089
rect 19521 22080 19533 22083
rect 19116 22052 19533 22080
rect 19116 22040 19122 22052
rect 19521 22049 19533 22052
rect 19567 22049 19579 22083
rect 19521 22043 19579 22049
rect 19981 22083 20039 22089
rect 19981 22049 19993 22083
rect 20027 22080 20039 22083
rect 20714 22080 20720 22092
rect 20027 22052 20720 22080
rect 20027 22049 20039 22052
rect 19981 22043 20039 22049
rect 20714 22040 20720 22052
rect 20772 22040 20778 22092
rect 20806 22040 20812 22092
rect 20864 22080 20870 22092
rect 20864 22052 22600 22080
rect 20864 22040 20870 22052
rect 15289 21975 15347 21981
rect 17880 21984 18644 22012
rect 9723 21916 10088 21944
rect 10229 21947 10287 21953
rect 9723 21913 9735 21916
rect 9677 21907 9735 21913
rect 10229 21913 10241 21947
rect 10275 21944 10287 21947
rect 10318 21944 10324 21956
rect 10275 21916 10324 21944
rect 10275 21913 10287 21916
rect 10229 21907 10287 21913
rect 10318 21904 10324 21916
rect 10376 21904 10382 21956
rect 10597 21947 10655 21953
rect 10597 21913 10609 21947
rect 10643 21944 10655 21947
rect 11698 21944 11704 21956
rect 10643 21916 11704 21944
rect 10643 21913 10655 21916
rect 10597 21907 10655 21913
rect 11698 21904 11704 21916
rect 11756 21904 11762 21956
rect 12158 21944 12164 21956
rect 12119 21916 12164 21944
rect 12158 21904 12164 21916
rect 12216 21904 12222 21956
rect 14918 21904 14924 21956
rect 14976 21944 14982 21956
rect 15304 21944 15332 21975
rect 14976 21916 15332 21944
rect 15841 21947 15899 21953
rect 14976 21904 14982 21916
rect 15841 21913 15853 21947
rect 15887 21944 15899 21947
rect 15930 21944 15936 21956
rect 15887 21916 15936 21944
rect 15887 21913 15899 21916
rect 15841 21907 15899 21913
rect 15930 21904 15936 21916
rect 15988 21904 15994 21956
rect 16850 21904 16856 21956
rect 16908 21904 16914 21956
rect 17880 21888 17908 21984
rect 19150 21972 19156 22024
rect 19208 22012 19214 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 19208 21984 19257 22012
rect 19208 21972 19214 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 19245 21975 19303 21981
rect 19334 21972 19340 22024
rect 19392 22012 19398 22024
rect 19428 22015 19486 22021
rect 19428 22012 19440 22015
rect 19392 21984 19440 22012
rect 19392 21972 19398 21984
rect 19428 21981 19440 21984
rect 19474 21981 19486 22015
rect 19428 21975 19486 21981
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 18966 21904 18972 21956
rect 19024 21944 19030 21956
rect 19628 21944 19656 21975
rect 19702 21972 19708 22024
rect 19760 22012 19766 22024
rect 19797 22015 19855 22021
rect 19797 22012 19809 22015
rect 19760 21984 19809 22012
rect 19760 21972 19766 21984
rect 19797 21981 19809 21984
rect 19843 21981 19855 22015
rect 19797 21975 19855 21981
rect 20993 22015 21051 22021
rect 20993 21981 21005 22015
rect 21039 21981 21051 22015
rect 20993 21975 21051 21981
rect 19024 21916 19656 21944
rect 19024 21904 19030 21916
rect 8665 21879 8723 21885
rect 8665 21845 8677 21879
rect 8711 21845 8723 21879
rect 8665 21839 8723 21845
rect 8754 21836 8760 21888
rect 8812 21876 8818 21888
rect 9861 21879 9919 21885
rect 9861 21876 9873 21879
rect 8812 21848 9873 21876
rect 8812 21836 8818 21848
rect 9861 21845 9873 21848
rect 9907 21845 9919 21879
rect 9861 21839 9919 21845
rect 12802 21836 12808 21888
rect 12860 21876 12866 21888
rect 12986 21876 12992 21888
rect 12860 21848 12992 21876
rect 12860 21836 12866 21848
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 13538 21836 13544 21888
rect 13596 21876 13602 21888
rect 13633 21879 13691 21885
rect 13633 21876 13645 21879
rect 13596 21848 13645 21876
rect 13596 21836 13602 21848
rect 13633 21845 13645 21848
rect 13679 21845 13691 21879
rect 13633 21839 13691 21845
rect 14829 21879 14887 21885
rect 14829 21845 14841 21879
rect 14875 21876 14887 21879
rect 16022 21876 16028 21888
rect 14875 21848 16028 21876
rect 14875 21845 14887 21848
rect 14829 21839 14887 21845
rect 16022 21836 16028 21848
rect 16080 21836 16086 21888
rect 17313 21879 17371 21885
rect 17313 21845 17325 21879
rect 17359 21876 17371 21879
rect 17862 21876 17868 21888
rect 17359 21848 17868 21876
rect 17359 21845 17371 21848
rect 17313 21839 17371 21845
rect 17862 21836 17868 21848
rect 17920 21836 17926 21888
rect 17954 21836 17960 21888
rect 18012 21876 18018 21888
rect 18049 21879 18107 21885
rect 18049 21876 18061 21879
rect 18012 21848 18061 21876
rect 18012 21836 18018 21848
rect 18049 21845 18061 21848
rect 18095 21845 18107 21879
rect 18049 21839 18107 21845
rect 18322 21836 18328 21888
rect 18380 21876 18386 21888
rect 18417 21879 18475 21885
rect 18417 21876 18429 21879
rect 18380 21848 18429 21876
rect 18380 21836 18386 21848
rect 18417 21845 18429 21848
rect 18463 21845 18475 21879
rect 18417 21839 18475 21845
rect 19334 21836 19340 21888
rect 19392 21876 19398 21888
rect 20073 21879 20131 21885
rect 20073 21876 20085 21879
rect 19392 21848 20085 21876
rect 19392 21836 19398 21848
rect 20073 21845 20085 21848
rect 20119 21845 20131 21879
rect 21008 21876 21036 21975
rect 22278 21904 22284 21956
rect 22336 21904 22342 21956
rect 22572 21944 22600 22052
rect 22646 22040 22652 22092
rect 22704 22080 22710 22092
rect 22704 22052 23060 22080
rect 22704 22040 22710 22052
rect 22830 21972 22836 22024
rect 22888 22012 22894 22024
rect 22925 22015 22983 22021
rect 22925 22012 22937 22015
rect 22888 21984 22937 22012
rect 22888 21972 22894 21984
rect 22925 21981 22937 21984
rect 22971 21981 22983 22015
rect 23032 22012 23060 22052
rect 23106 22040 23112 22092
rect 23164 22080 23170 22092
rect 23492 22080 23520 22111
rect 23566 22080 23572 22092
rect 23164 22052 23428 22080
rect 23492 22052 23572 22080
rect 23164 22040 23170 22052
rect 23298 22015 23356 22021
rect 23298 22012 23310 22015
rect 23032 21984 23310 22012
rect 22925 21975 22983 21981
rect 23298 21981 23310 21984
rect 23344 21981 23356 22015
rect 23400 22012 23428 22052
rect 23566 22040 23572 22052
rect 23624 22040 23630 22092
rect 24118 22080 24124 22092
rect 23676 22052 24124 22080
rect 23676 22012 23704 22052
rect 24118 22040 24124 22052
rect 24176 22040 24182 22092
rect 23842 22012 23848 22024
rect 23400 21984 23704 22012
rect 23803 21984 23848 22012
rect 23298 21975 23356 21981
rect 23842 21972 23848 21984
rect 23900 21972 23906 22024
rect 23106 21944 23112 21956
rect 22572 21916 22968 21944
rect 23067 21916 23112 21944
rect 22094 21876 22100 21888
rect 21008 21848 22100 21876
rect 20073 21839 20131 21845
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 22741 21879 22799 21885
rect 22741 21845 22753 21879
rect 22787 21876 22799 21879
rect 22830 21876 22836 21888
rect 22787 21848 22836 21876
rect 22787 21845 22799 21848
rect 22741 21839 22799 21845
rect 22830 21836 22836 21848
rect 22888 21836 22894 21888
rect 22940 21876 22968 21916
rect 23106 21904 23112 21916
rect 23164 21904 23170 21956
rect 23201 21947 23259 21953
rect 23201 21913 23213 21947
rect 23247 21944 23259 21947
rect 23753 21947 23811 21953
rect 23753 21944 23765 21947
rect 23247 21916 23765 21944
rect 23247 21913 23259 21916
rect 23201 21907 23259 21913
rect 23753 21913 23765 21916
rect 23799 21944 23811 21947
rect 25222 21944 25228 21956
rect 23799 21916 25228 21944
rect 23799 21913 23811 21916
rect 23753 21907 23811 21913
rect 25222 21904 25228 21916
rect 25280 21904 25286 21956
rect 23474 21876 23480 21888
rect 22940 21848 23480 21876
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 24026 21876 24032 21888
rect 23987 21848 24032 21876
rect 24026 21836 24032 21848
rect 24084 21836 24090 21888
rect 1104 21786 29440 21808
rect 1104 21734 10395 21786
rect 10447 21734 10459 21786
rect 10511 21734 10523 21786
rect 10575 21734 10587 21786
rect 10639 21734 10651 21786
rect 10703 21734 19840 21786
rect 19892 21734 19904 21786
rect 19956 21734 19968 21786
rect 20020 21734 20032 21786
rect 20084 21734 20096 21786
rect 20148 21734 29440 21786
rect 1104 21712 29440 21734
rect 4890 21672 4896 21684
rect 4080 21644 4896 21672
rect 3970 21604 3976 21616
rect 3712 21576 3976 21604
rect 3326 21496 3332 21548
rect 3384 21536 3390 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 3384 21508 3433 21536
rect 3384 21496 3390 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3602 21536 3608 21548
rect 3564 21508 3608 21536
rect 3421 21499 3479 21505
rect 3602 21496 3608 21508
rect 3660 21496 3666 21548
rect 3712 21545 3740 21576
rect 3970 21564 3976 21576
rect 4028 21564 4034 21616
rect 4080 21613 4108 21644
rect 4890 21632 4896 21644
rect 4948 21632 4954 21684
rect 6454 21672 6460 21684
rect 6012 21644 6460 21672
rect 4065 21607 4123 21613
rect 4065 21573 4077 21607
rect 4111 21573 4123 21607
rect 4065 21567 4123 21573
rect 3697 21539 3755 21545
rect 3697 21505 3709 21539
rect 3743 21505 3755 21539
rect 3697 21499 3755 21505
rect 3823 21539 3881 21545
rect 3823 21505 3835 21539
rect 3869 21536 3881 21539
rect 4154 21536 4160 21548
rect 3869 21508 4160 21536
rect 3869 21505 3881 21508
rect 3823 21499 3881 21505
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21505 4675 21539
rect 4798 21536 4804 21548
rect 4759 21508 4804 21536
rect 4617 21499 4675 21505
rect 4632 21468 4660 21499
rect 4798 21496 4804 21508
rect 4856 21496 4862 21548
rect 6012 21545 6040 21644
rect 6454 21632 6460 21644
rect 6512 21672 6518 21684
rect 6512 21644 6684 21672
rect 6512 21632 6518 21644
rect 6270 21604 6276 21616
rect 6183 21576 6276 21604
rect 6196 21545 6224 21576
rect 6270 21564 6276 21576
rect 6328 21604 6334 21616
rect 6549 21607 6607 21613
rect 6549 21604 6561 21607
rect 6328 21576 6561 21604
rect 6328 21564 6334 21576
rect 6549 21573 6561 21576
rect 6595 21573 6607 21607
rect 6656 21604 6684 21644
rect 6914 21632 6920 21684
rect 6972 21672 6978 21684
rect 7377 21675 7435 21681
rect 7377 21672 7389 21675
rect 6972 21644 7389 21672
rect 6972 21632 6978 21644
rect 7377 21641 7389 21644
rect 7423 21641 7435 21675
rect 7377 21635 7435 21641
rect 7742 21632 7748 21684
rect 7800 21672 7806 21684
rect 7929 21675 7987 21681
rect 7929 21672 7941 21675
rect 7800 21644 7941 21672
rect 7800 21632 7806 21644
rect 7929 21641 7941 21644
rect 7975 21641 7987 21675
rect 7929 21635 7987 21641
rect 8938 21632 8944 21684
rect 8996 21672 9002 21684
rect 9858 21672 9864 21684
rect 8996 21644 9864 21672
rect 8996 21632 9002 21644
rect 9858 21632 9864 21644
rect 9916 21672 9922 21684
rect 10045 21675 10103 21681
rect 10045 21672 10057 21675
rect 9916 21644 10057 21672
rect 9916 21632 9922 21644
rect 10045 21641 10057 21644
rect 10091 21641 10103 21675
rect 10045 21635 10103 21641
rect 10778 21632 10784 21684
rect 10836 21672 10842 21684
rect 10965 21675 11023 21681
rect 10965 21672 10977 21675
rect 10836 21644 10977 21672
rect 10836 21632 10842 21644
rect 10965 21641 10977 21644
rect 11011 21672 11023 21675
rect 11238 21672 11244 21684
rect 11011 21644 11244 21672
rect 11011 21641 11023 21644
rect 10965 21635 11023 21641
rect 11238 21632 11244 21644
rect 11296 21632 11302 21684
rect 12250 21632 12256 21684
rect 12308 21672 12314 21684
rect 12437 21675 12495 21681
rect 12437 21672 12449 21675
rect 12308 21644 12449 21672
rect 12308 21632 12314 21644
rect 12437 21641 12449 21644
rect 12483 21641 12495 21675
rect 12437 21635 12495 21641
rect 12529 21675 12587 21681
rect 12529 21641 12541 21675
rect 12575 21672 12587 21675
rect 13538 21672 13544 21684
rect 12575 21644 13544 21672
rect 12575 21641 12587 21644
rect 12529 21635 12587 21641
rect 13538 21632 13544 21644
rect 13596 21632 13602 21684
rect 15194 21632 15200 21684
rect 15252 21672 15258 21684
rect 15841 21675 15899 21681
rect 15841 21672 15853 21675
rect 15252 21644 15853 21672
rect 15252 21632 15258 21644
rect 15841 21641 15853 21644
rect 15887 21672 15899 21675
rect 16390 21672 16396 21684
rect 15887 21644 16396 21672
rect 15887 21641 15899 21644
rect 15841 21635 15899 21641
rect 16390 21632 16396 21644
rect 16448 21632 16454 21684
rect 16850 21672 16856 21684
rect 16811 21644 16856 21672
rect 16850 21632 16856 21644
rect 16908 21632 16914 21684
rect 19426 21672 19432 21684
rect 19387 21644 19432 21672
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 22005 21675 22063 21681
rect 22005 21641 22017 21675
rect 22051 21672 22063 21675
rect 22186 21672 22192 21684
rect 22051 21644 22192 21672
rect 22051 21641 22063 21644
rect 22005 21635 22063 21641
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 23201 21675 23259 21681
rect 22388 21644 23060 21672
rect 7469 21607 7527 21613
rect 6656 21576 7144 21604
rect 6549 21567 6607 21573
rect 4893 21539 4951 21545
rect 4893 21505 4905 21539
rect 4939 21505 4951 21539
rect 4893 21499 4951 21505
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21505 6055 21539
rect 5997 21499 6055 21505
rect 6181 21539 6239 21545
rect 6181 21505 6193 21539
rect 6227 21505 6239 21539
rect 6362 21536 6368 21548
rect 6323 21508 6368 21536
rect 6181 21499 6239 21505
rect 4908 21468 4936 21499
rect 6362 21496 6368 21508
rect 6420 21536 6426 21548
rect 6825 21539 6883 21545
rect 6825 21536 6837 21539
rect 6420 21508 6837 21536
rect 6420 21496 6426 21508
rect 6825 21505 6837 21508
rect 6871 21505 6883 21539
rect 6825 21499 6883 21505
rect 7009 21539 7067 21545
rect 7009 21505 7021 21539
rect 7055 21505 7067 21539
rect 7116 21536 7144 21576
rect 7469 21573 7481 21607
rect 7515 21604 7527 21607
rect 8294 21604 8300 21616
rect 7515 21576 8300 21604
rect 7515 21573 7527 21576
rect 7469 21567 7527 21573
rect 8294 21564 8300 21576
rect 8352 21604 8358 21616
rect 8754 21604 8760 21616
rect 8352 21576 8760 21604
rect 8352 21564 8358 21576
rect 8754 21564 8760 21576
rect 8812 21564 8818 21616
rect 9033 21607 9091 21613
rect 9033 21573 9045 21607
rect 9079 21604 9091 21607
rect 9677 21607 9735 21613
rect 9677 21604 9689 21607
rect 9079 21576 9689 21604
rect 9079 21573 9091 21576
rect 9033 21567 9091 21573
rect 9677 21573 9689 21576
rect 9723 21573 9735 21607
rect 9677 21567 9735 21573
rect 10134 21564 10140 21616
rect 10192 21564 10198 21616
rect 10318 21564 10324 21616
rect 10376 21604 10382 21616
rect 12158 21604 12164 21616
rect 10376 21576 11100 21604
rect 12119 21576 12164 21604
rect 10376 21564 10382 21576
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 7116 21508 7665 21536
rect 7009 21499 7067 21505
rect 7653 21505 7665 21508
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 7024 21468 7052 21499
rect 8018 21496 8024 21548
rect 8076 21536 8082 21548
rect 8113 21539 8171 21545
rect 8113 21536 8125 21539
rect 8076 21508 8125 21536
rect 8076 21496 8082 21508
rect 8113 21505 8125 21508
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 9217 21539 9275 21545
rect 9217 21505 9229 21539
rect 9263 21505 9275 21539
rect 9217 21499 9275 21505
rect 9401 21539 9459 21545
rect 9401 21505 9413 21539
rect 9447 21536 9459 21539
rect 9582 21536 9588 21548
rect 9447 21508 9588 21536
rect 9447 21505 9459 21508
rect 9401 21499 9459 21505
rect 7834 21468 7840 21480
rect 4632 21440 6960 21468
rect 7024 21440 7840 21468
rect 4154 21360 4160 21412
rect 4212 21400 4218 21412
rect 5077 21403 5135 21409
rect 5077 21400 5089 21403
rect 4212 21372 5089 21400
rect 4212 21360 4218 21372
rect 5077 21369 5089 21372
rect 5123 21400 5135 21403
rect 5442 21400 5448 21412
rect 5123 21372 5448 21400
rect 5123 21369 5135 21372
rect 5077 21363 5135 21369
rect 5442 21360 5448 21372
rect 5500 21360 5506 21412
rect 6730 21400 6736 21412
rect 6691 21372 6736 21400
rect 6730 21360 6736 21372
rect 6788 21360 6794 21412
rect 6932 21409 6960 21440
rect 7834 21428 7840 21440
rect 7892 21428 7898 21480
rect 9232 21412 9260 21499
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 10152 21536 10180 21564
rect 10229 21539 10287 21545
rect 10229 21536 10241 21539
rect 10152 21508 10241 21536
rect 10229 21505 10241 21508
rect 10275 21505 10287 21539
rect 10778 21536 10784 21548
rect 10739 21508 10784 21536
rect 10229 21499 10287 21505
rect 10778 21496 10784 21508
rect 10836 21496 10842 21548
rect 11072 21545 11100 21576
rect 12158 21564 12164 21576
rect 12216 21564 12222 21616
rect 12345 21607 12403 21613
rect 12345 21573 12357 21607
rect 12391 21604 12403 21607
rect 12716 21607 12774 21613
rect 12391 21576 12664 21604
rect 12391 21573 12403 21576
rect 12345 21567 12403 21573
rect 11057 21539 11115 21545
rect 11057 21505 11069 21539
rect 11103 21536 11115 21539
rect 11149 21539 11207 21545
rect 11149 21536 11161 21539
rect 11103 21508 11161 21536
rect 11103 21505 11115 21508
rect 11057 21499 11115 21505
rect 11149 21505 11161 21508
rect 11195 21505 11207 21539
rect 12636 21536 12664 21576
rect 12716 21573 12728 21607
rect 12762 21604 12774 21607
rect 12986 21604 12992 21616
rect 12762 21576 12992 21604
rect 12762 21573 12774 21576
rect 12716 21567 12774 21573
rect 12986 21564 12992 21576
rect 13044 21564 13050 21616
rect 14734 21564 14740 21616
rect 14792 21564 14798 21616
rect 15470 21564 15476 21616
rect 15528 21604 15534 21616
rect 19444 21604 19472 21632
rect 19797 21607 19855 21613
rect 19797 21604 19809 21607
rect 15528 21576 17632 21604
rect 19444 21576 19809 21604
rect 15528 21564 15534 21576
rect 12802 21536 12808 21548
rect 12636 21508 12808 21536
rect 11149 21499 11207 21505
rect 12802 21496 12808 21508
rect 12860 21496 12866 21548
rect 15381 21539 15439 21545
rect 15381 21536 15393 21539
rect 14936 21508 15393 21536
rect 14936 21480 14964 21508
rect 15381 21505 15393 21508
rect 15427 21536 15439 21539
rect 15657 21539 15715 21545
rect 15657 21536 15669 21539
rect 15427 21508 15669 21536
rect 15427 21505 15439 21508
rect 15381 21499 15439 21505
rect 15657 21505 15669 21508
rect 15703 21505 15715 21539
rect 15657 21499 15715 21505
rect 15838 21496 15844 21548
rect 15896 21536 15902 21548
rect 16117 21539 16175 21545
rect 16117 21536 16129 21539
rect 15896 21508 16129 21536
rect 15896 21496 15902 21508
rect 16117 21505 16129 21508
rect 16163 21505 16175 21539
rect 16117 21499 16175 21505
rect 16485 21539 16543 21545
rect 16485 21505 16497 21539
rect 16531 21536 16543 21539
rect 16669 21539 16727 21545
rect 16669 21536 16681 21539
rect 16531 21508 16681 21536
rect 16531 21505 16543 21508
rect 16485 21499 16543 21505
rect 16669 21505 16681 21508
rect 16715 21505 16727 21539
rect 17604 21536 17632 21576
rect 19797 21573 19809 21576
rect 19843 21573 19855 21607
rect 22388 21604 22416 21644
rect 19797 21567 19855 21573
rect 22066 21576 22416 21604
rect 22465 21607 22523 21613
rect 22066 21548 22094 21576
rect 22465 21573 22477 21607
rect 22511 21604 22523 21607
rect 22830 21604 22836 21616
rect 22511 21576 22836 21604
rect 22511 21573 22523 21576
rect 22465 21567 22523 21573
rect 22830 21564 22836 21576
rect 22888 21564 22894 21616
rect 20898 21536 20904 21548
rect 17604 21508 20904 21536
rect 16669 21499 16727 21505
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21100 21508 21833 21536
rect 9950 21477 9956 21480
rect 9936 21471 9956 21477
rect 9936 21437 9948 21471
rect 9936 21431 9956 21437
rect 9950 21428 9956 21431
rect 10008 21428 10014 21480
rect 10137 21471 10195 21477
rect 10137 21437 10149 21471
rect 10183 21437 10195 21471
rect 10686 21468 10692 21480
rect 10647 21440 10692 21468
rect 10137 21431 10195 21437
rect 6917 21403 6975 21409
rect 6917 21369 6929 21403
rect 6963 21369 6975 21403
rect 9214 21400 9220 21412
rect 6917 21363 6975 21369
rect 7668 21372 9220 21400
rect 3878 21292 3884 21344
rect 3936 21332 3942 21344
rect 4525 21335 4583 21341
rect 4525 21332 4537 21335
rect 3936 21304 4537 21332
rect 3936 21292 3942 21304
rect 4525 21301 4537 21304
rect 4571 21301 4583 21335
rect 6086 21332 6092 21344
rect 6047 21304 6092 21332
rect 4525 21295 4583 21301
rect 6086 21292 6092 21304
rect 6144 21292 6150 21344
rect 6748 21332 6776 21360
rect 7668 21332 7696 21372
rect 9214 21360 9220 21372
rect 9272 21360 9278 21412
rect 9306 21360 9312 21412
rect 9364 21400 9370 21412
rect 10152 21400 10180 21431
rect 10686 21428 10692 21440
rect 10744 21428 10750 21480
rect 11514 21428 11520 21480
rect 11572 21468 11578 21480
rect 13265 21471 13323 21477
rect 13265 21468 13277 21471
rect 11572 21440 13277 21468
rect 11572 21428 11578 21440
rect 13265 21437 13277 21440
rect 13311 21468 13323 21471
rect 13449 21471 13507 21477
rect 13449 21468 13461 21471
rect 13311 21440 13461 21468
rect 13311 21437 13323 21440
rect 13265 21431 13323 21437
rect 13449 21437 13461 21440
rect 13495 21437 13507 21471
rect 13722 21468 13728 21480
rect 13683 21440 13728 21468
rect 13449 21431 13507 21437
rect 13722 21428 13728 21440
rect 13780 21428 13786 21480
rect 14918 21428 14924 21480
rect 14976 21428 14982 21480
rect 15120 21440 21036 21468
rect 10870 21400 10876 21412
rect 9364 21372 9628 21400
rect 10152 21372 10876 21400
rect 9364 21360 9370 21372
rect 7834 21332 7840 21344
rect 6748 21304 7696 21332
rect 7795 21304 7840 21332
rect 7834 21292 7840 21304
rect 7892 21292 7898 21344
rect 9398 21292 9404 21344
rect 9456 21332 9462 21344
rect 9493 21335 9551 21341
rect 9493 21332 9505 21335
rect 9456 21304 9505 21332
rect 9456 21292 9462 21304
rect 9493 21301 9505 21304
rect 9539 21301 9551 21335
rect 9600 21332 9628 21372
rect 10870 21360 10876 21372
rect 10928 21360 10934 21412
rect 11333 21403 11391 21409
rect 11333 21369 11345 21403
rect 11379 21400 11391 21403
rect 11422 21400 11428 21412
rect 11379 21372 11428 21400
rect 11379 21369 11391 21372
rect 11333 21363 11391 21369
rect 11422 21360 11428 21372
rect 11480 21400 11486 21412
rect 12342 21400 12348 21412
rect 11480 21372 12348 21400
rect 11480 21360 11486 21372
rect 12342 21360 12348 21372
rect 12400 21360 12406 21412
rect 10413 21335 10471 21341
rect 10413 21332 10425 21335
rect 9600 21304 10425 21332
rect 9493 21295 9551 21301
rect 10413 21301 10425 21304
rect 10459 21301 10471 21335
rect 10413 21295 10471 21301
rect 10781 21335 10839 21341
rect 10781 21301 10793 21335
rect 10827 21332 10839 21335
rect 11514 21332 11520 21344
rect 10827 21304 11520 21332
rect 10827 21301 10839 21304
rect 10781 21295 10839 21301
rect 11514 21292 11520 21304
rect 11572 21292 11578 21344
rect 14090 21292 14096 21344
rect 14148 21332 14154 21344
rect 15120 21332 15148 21440
rect 15197 21403 15255 21409
rect 15197 21369 15209 21403
rect 15243 21400 15255 21403
rect 16114 21400 16120 21412
rect 15243 21372 16120 21400
rect 15243 21369 15255 21372
rect 15197 21363 15255 21369
rect 16114 21360 16120 21372
rect 16172 21360 16178 21412
rect 16301 21403 16359 21409
rect 16301 21369 16313 21403
rect 16347 21400 16359 21403
rect 16485 21403 16543 21409
rect 16485 21400 16497 21403
rect 16347 21372 16497 21400
rect 16347 21369 16359 21372
rect 16301 21363 16359 21369
rect 16485 21369 16497 21372
rect 16531 21369 16543 21403
rect 16485 21363 16543 21369
rect 18046 21360 18052 21412
rect 18104 21400 18110 21412
rect 19242 21400 19248 21412
rect 18104 21372 19248 21400
rect 18104 21360 18110 21372
rect 19242 21360 19248 21372
rect 19300 21360 19306 21412
rect 19426 21360 19432 21412
rect 19484 21400 19490 21412
rect 19613 21403 19671 21409
rect 19613 21400 19625 21403
rect 19484 21372 19625 21400
rect 19484 21360 19490 21372
rect 19613 21369 19625 21372
rect 19659 21400 19671 21403
rect 20530 21400 20536 21412
rect 19659 21372 20536 21400
rect 19659 21369 19671 21372
rect 19613 21363 19671 21369
rect 20530 21360 20536 21372
rect 20588 21360 20594 21412
rect 14148 21304 15148 21332
rect 14148 21292 14154 21304
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 15565 21335 15623 21341
rect 15565 21332 15577 21335
rect 15528 21304 15577 21332
rect 15528 21292 15534 21304
rect 15565 21301 15577 21304
rect 15611 21301 15623 21335
rect 15565 21295 15623 21301
rect 16206 21292 16212 21344
rect 16264 21332 16270 21344
rect 20898 21332 20904 21344
rect 16264 21304 20904 21332
rect 16264 21292 16270 21304
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 21008 21332 21036 21440
rect 21100 21409 21128 21508
rect 21821 21505 21833 21508
rect 21867 21536 21879 21539
rect 22002 21536 22008 21548
rect 21867 21508 22008 21536
rect 21867 21505 21879 21508
rect 21821 21499 21879 21505
rect 22002 21496 22008 21508
rect 22060 21508 22094 21548
rect 22060 21496 22066 21508
rect 22278 21496 22284 21548
rect 22336 21545 22342 21548
rect 22336 21539 22379 21545
rect 22367 21505 22379 21539
rect 22336 21499 22379 21505
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21505 22615 21539
rect 22738 21536 22744 21548
rect 22699 21508 22744 21536
rect 22557 21499 22615 21505
rect 22336 21496 22342 21499
rect 21085 21403 21143 21409
rect 21085 21369 21097 21403
rect 21131 21369 21143 21403
rect 21085 21363 21143 21369
rect 22189 21403 22247 21409
rect 22189 21369 22201 21403
rect 22235 21400 22247 21403
rect 22370 21400 22376 21412
rect 22235 21372 22376 21400
rect 22235 21369 22247 21372
rect 22189 21363 22247 21369
rect 22370 21360 22376 21372
rect 22428 21360 22434 21412
rect 22462 21360 22468 21412
rect 22520 21400 22526 21412
rect 22572 21400 22600 21499
rect 22738 21496 22744 21508
rect 22796 21496 22802 21548
rect 23032 21545 23060 21644
rect 23201 21641 23213 21675
rect 23247 21672 23259 21675
rect 23842 21672 23848 21684
rect 23247 21644 23848 21672
rect 23247 21641 23259 21644
rect 23201 21635 23259 21641
rect 23842 21632 23848 21644
rect 23900 21632 23906 21684
rect 23566 21604 23572 21616
rect 23527 21576 23572 21604
rect 23566 21564 23572 21576
rect 23624 21564 23630 21616
rect 24026 21564 24032 21616
rect 24084 21564 24090 21616
rect 23017 21539 23075 21545
rect 23017 21505 23029 21539
rect 23063 21505 23075 21539
rect 23017 21499 23075 21505
rect 22646 21428 22652 21480
rect 22704 21468 22710 21480
rect 23293 21471 23351 21477
rect 23293 21468 23305 21471
rect 22704 21440 23305 21468
rect 22704 21428 22710 21440
rect 23293 21437 23305 21440
rect 23339 21437 23351 21471
rect 23293 21431 23351 21437
rect 23106 21400 23112 21412
rect 22520 21372 22600 21400
rect 22664 21372 23112 21400
rect 22520 21360 22526 21372
rect 22664 21332 22692 21372
rect 23106 21360 23112 21372
rect 23164 21360 23170 21412
rect 22830 21332 22836 21344
rect 21008 21304 22692 21332
rect 22791 21304 22836 21332
rect 22830 21292 22836 21304
rect 22888 21292 22894 21344
rect 25041 21335 25099 21341
rect 25041 21301 25053 21335
rect 25087 21332 25099 21335
rect 25222 21332 25228 21344
rect 25087 21304 25228 21332
rect 25087 21301 25099 21304
rect 25041 21295 25099 21301
rect 25222 21292 25228 21304
rect 25280 21292 25286 21344
rect 1104 21242 29440 21264
rect 1104 21190 5672 21242
rect 5724 21190 5736 21242
rect 5788 21190 5800 21242
rect 5852 21190 5864 21242
rect 5916 21190 5928 21242
rect 5980 21190 15118 21242
rect 15170 21190 15182 21242
rect 15234 21190 15246 21242
rect 15298 21190 15310 21242
rect 15362 21190 15374 21242
rect 15426 21190 24563 21242
rect 24615 21190 24627 21242
rect 24679 21190 24691 21242
rect 24743 21190 24755 21242
rect 24807 21190 24819 21242
rect 24871 21190 29440 21242
rect 1104 21168 29440 21190
rect 3602 21128 3608 21140
rect 3436 21100 3608 21128
rect 2866 20992 2872 21004
rect 2827 20964 2872 20992
rect 2866 20952 2872 20964
rect 2924 20952 2930 21004
rect 3436 20992 3464 21100
rect 3602 21088 3608 21100
rect 3660 21128 3666 21140
rect 5350 21128 5356 21140
rect 3660 21100 4936 21128
rect 5311 21100 5356 21128
rect 3660 21088 3666 21100
rect 4062 21020 4068 21072
rect 4120 21060 4126 21072
rect 4908 21060 4936 21100
rect 5350 21088 5356 21100
rect 5408 21088 5414 21140
rect 7377 21131 7435 21137
rect 7377 21097 7389 21131
rect 7423 21128 7435 21131
rect 8938 21128 8944 21140
rect 7423 21100 8944 21128
rect 7423 21097 7435 21100
rect 7377 21091 7435 21097
rect 8938 21088 8944 21100
rect 8996 21088 9002 21140
rect 9030 21088 9036 21140
rect 9088 21128 9094 21140
rect 9493 21131 9551 21137
rect 9493 21128 9505 21131
rect 9088 21100 9505 21128
rect 9088 21088 9094 21100
rect 9493 21097 9505 21100
rect 9539 21097 9551 21131
rect 9493 21091 9551 21097
rect 12434 21088 12440 21140
rect 12492 21128 12498 21140
rect 12621 21131 12679 21137
rect 12621 21128 12633 21131
rect 12492 21100 12633 21128
rect 12492 21088 12498 21100
rect 12621 21097 12633 21100
rect 12667 21097 12679 21131
rect 13814 21128 13820 21140
rect 13775 21100 13820 21128
rect 12621 21091 12679 21097
rect 13814 21088 13820 21100
rect 13872 21088 13878 21140
rect 16942 21088 16948 21140
rect 17000 21128 17006 21140
rect 17313 21131 17371 21137
rect 17313 21128 17325 21131
rect 17000 21100 17325 21128
rect 17000 21088 17006 21100
rect 17313 21097 17325 21100
rect 17359 21097 17371 21131
rect 20806 21128 20812 21140
rect 17313 21091 17371 21097
rect 19260 21100 20812 21128
rect 6086 21060 6092 21072
rect 4120 21032 4844 21060
rect 4908 21032 6092 21060
rect 4120 21020 4126 21032
rect 3160 20964 3464 20992
rect 3160 20933 3188 20964
rect 3145 20927 3203 20933
rect 3145 20893 3157 20927
rect 3191 20893 3203 20927
rect 3326 20924 3332 20936
rect 3287 20896 3332 20924
rect 3145 20887 3203 20893
rect 3326 20884 3332 20896
rect 3384 20884 3390 20936
rect 3436 20933 3464 20964
rect 4709 20995 4767 21001
rect 4709 20961 4721 20995
rect 4755 20961 4767 20995
rect 4816 20992 4844 21032
rect 6086 21020 6092 21032
rect 6144 21020 6150 21072
rect 7834 21020 7840 21072
rect 7892 21060 7898 21072
rect 14918 21060 14924 21072
rect 7892 21032 14924 21060
rect 7892 21020 7898 21032
rect 14918 21020 14924 21032
rect 14976 21020 14982 21072
rect 16485 21063 16543 21069
rect 16485 21029 16497 21063
rect 16531 21060 16543 21063
rect 19260 21060 19288 21100
rect 20806 21088 20812 21100
rect 20864 21088 20870 21140
rect 22002 21088 22008 21140
rect 22060 21128 22066 21140
rect 22060 21100 22416 21128
rect 22060 21088 22066 21100
rect 16531 21032 19288 21060
rect 22388 21060 22416 21100
rect 22462 21088 22468 21140
rect 22520 21128 22526 21140
rect 23017 21131 23075 21137
rect 23017 21128 23029 21131
rect 22520 21100 23029 21128
rect 22520 21088 22526 21100
rect 23017 21097 23029 21100
rect 23063 21097 23075 21131
rect 23017 21091 23075 21097
rect 22388 21032 22784 21060
rect 16531 21029 16543 21032
rect 16485 21023 16543 21029
rect 17221 20995 17279 21001
rect 4816 20964 16896 20992
rect 4709 20955 4767 20961
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20893 3479 20927
rect 3421 20887 3479 20893
rect 3789 20927 3847 20933
rect 3789 20893 3801 20927
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 1854 20816 1860 20868
rect 1912 20856 1918 20868
rect 2602 20859 2660 20865
rect 2602 20856 2614 20859
rect 1912 20828 2614 20856
rect 1912 20816 1918 20828
rect 2602 20825 2614 20828
rect 2648 20825 2660 20859
rect 2958 20856 2964 20868
rect 2919 20828 2964 20856
rect 2602 20819 2660 20825
rect 2958 20816 2964 20828
rect 3016 20816 3022 20868
rect 3234 20816 3240 20868
rect 3292 20856 3298 20868
rect 3804 20856 3832 20887
rect 3970 20884 3976 20936
rect 4028 20924 4034 20936
rect 4085 20927 4143 20933
rect 4085 20924 4097 20927
rect 4028 20896 4097 20924
rect 4028 20884 4034 20896
rect 4085 20893 4097 20896
rect 4131 20893 4143 20927
rect 4338 20924 4344 20936
rect 4299 20896 4344 20924
rect 4085 20887 4143 20893
rect 4338 20884 4344 20896
rect 4396 20884 4402 20936
rect 4614 20884 4620 20936
rect 4672 20924 4678 20936
rect 4724 20924 4752 20955
rect 5442 20924 5448 20936
rect 4672 20896 5120 20924
rect 5403 20896 5448 20924
rect 4672 20884 4678 20896
rect 4525 20859 4583 20865
rect 3292 20828 3832 20856
rect 3896 20828 4292 20856
rect 3292 20816 3298 20828
rect 1394 20748 1400 20800
rect 1452 20788 1458 20800
rect 1489 20791 1547 20797
rect 1489 20788 1501 20791
rect 1452 20760 1501 20788
rect 1452 20748 1458 20760
rect 1489 20757 1501 20760
rect 1535 20757 1547 20791
rect 3510 20788 3516 20800
rect 3471 20760 3516 20788
rect 1489 20751 1547 20757
rect 3510 20748 3516 20760
rect 3568 20788 3574 20800
rect 3896 20797 3924 20828
rect 3881 20791 3939 20797
rect 3881 20788 3893 20791
rect 3568 20760 3893 20788
rect 3568 20748 3574 20760
rect 3881 20757 3893 20760
rect 3927 20757 3939 20791
rect 3881 20751 3939 20757
rect 3973 20791 4031 20797
rect 3973 20757 3985 20791
rect 4019 20788 4031 20791
rect 4154 20788 4160 20800
rect 4019 20760 4160 20788
rect 4019 20757 4031 20760
rect 3973 20751 4031 20757
rect 4154 20748 4160 20760
rect 4212 20748 4218 20800
rect 4264 20788 4292 20828
rect 4525 20825 4537 20859
rect 4571 20856 4583 20859
rect 4985 20859 5043 20865
rect 4985 20856 4997 20859
rect 4571 20828 4997 20856
rect 4571 20825 4583 20828
rect 4525 20819 4583 20825
rect 4985 20825 4997 20828
rect 5031 20825 5043 20859
rect 5092 20856 5120 20896
rect 5442 20884 5448 20896
rect 5500 20884 5506 20936
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20924 5779 20927
rect 6086 20924 6092 20936
rect 5767 20896 6092 20924
rect 5767 20893 5779 20896
rect 5721 20887 5779 20893
rect 6086 20884 6092 20896
rect 6144 20884 6150 20936
rect 6914 20884 6920 20936
rect 6972 20924 6978 20936
rect 7193 20927 7251 20933
rect 7193 20924 7205 20927
rect 6972 20896 7205 20924
rect 6972 20884 6978 20896
rect 7193 20893 7205 20896
rect 7239 20893 7251 20927
rect 7193 20887 7251 20893
rect 7745 20927 7803 20933
rect 7745 20893 7757 20927
rect 7791 20893 7803 20927
rect 7926 20924 7932 20936
rect 7887 20896 7932 20924
rect 7745 20887 7803 20893
rect 7760 20856 7788 20887
rect 7926 20884 7932 20896
rect 7984 20884 7990 20936
rect 9306 20884 9312 20936
rect 9364 20924 9370 20936
rect 9401 20927 9459 20933
rect 9401 20924 9413 20927
rect 9364 20896 9413 20924
rect 9364 20884 9370 20896
rect 9401 20893 9413 20896
rect 9447 20893 9459 20927
rect 12618 20924 12624 20936
rect 12579 20896 12624 20924
rect 9401 20887 9459 20893
rect 12618 20884 12624 20896
rect 12676 20884 12682 20936
rect 12805 20927 12863 20933
rect 12805 20893 12817 20927
rect 12851 20924 12863 20927
rect 13538 20924 13544 20936
rect 12851 20896 13544 20924
rect 12851 20893 12863 20896
rect 12805 20887 12863 20893
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 13633 20927 13691 20933
rect 13633 20893 13645 20927
rect 13679 20893 13691 20927
rect 14550 20924 14556 20936
rect 14511 20896 14556 20924
rect 13633 20887 13691 20893
rect 9122 20856 9128 20868
rect 5092 20828 5580 20856
rect 7760 20828 9128 20856
rect 4985 20819 5043 20825
rect 4798 20788 4804 20800
rect 4264 20760 4804 20788
rect 4798 20748 4804 20760
rect 4856 20788 4862 20800
rect 5552 20797 5580 20828
rect 9122 20816 9128 20828
rect 9180 20816 9186 20868
rect 9217 20859 9275 20865
rect 9217 20825 9229 20859
rect 9263 20825 9275 20859
rect 13648 20856 13676 20887
rect 14550 20884 14556 20896
rect 14608 20884 14614 20936
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20924 14887 20927
rect 15194 20924 15200 20936
rect 14875 20896 15200 20924
rect 14875 20893 14887 20896
rect 14829 20887 14887 20893
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 15654 20884 15660 20936
rect 15712 20924 15718 20936
rect 16301 20927 16359 20933
rect 16301 20924 16313 20927
rect 15712 20896 16313 20924
rect 15712 20884 15718 20896
rect 16301 20893 16313 20896
rect 16347 20893 16359 20927
rect 16301 20887 16359 20893
rect 16761 20927 16819 20933
rect 16761 20893 16773 20927
rect 16807 20893 16819 20927
rect 16868 20924 16896 20964
rect 17221 20961 17233 20995
rect 17267 20992 17279 20995
rect 17865 20995 17923 21001
rect 17865 20992 17877 20995
rect 17267 20964 17877 20992
rect 17267 20961 17279 20964
rect 17221 20955 17279 20961
rect 17865 20961 17877 20964
rect 17911 20992 17923 20995
rect 17954 20992 17960 21004
rect 17911 20964 17960 20992
rect 17911 20961 17923 20964
rect 17865 20955 17923 20961
rect 17954 20952 17960 20964
rect 18012 20952 18018 21004
rect 18601 20995 18659 21001
rect 18156 20964 18460 20992
rect 18156 20933 18184 20964
rect 18141 20927 18199 20933
rect 18141 20924 18153 20927
rect 16868 20896 18153 20924
rect 16761 20887 16819 20893
rect 18141 20893 18153 20896
rect 18187 20893 18199 20927
rect 18325 20927 18383 20933
rect 18325 20924 18337 20927
rect 18141 20887 18199 20893
rect 18248 20896 18337 20924
rect 9217 20819 9275 20825
rect 13004 20828 13676 20856
rect 4893 20791 4951 20797
rect 4893 20788 4905 20791
rect 4856 20760 4905 20788
rect 4856 20748 4862 20760
rect 4893 20757 4905 20760
rect 4939 20757 4951 20791
rect 4893 20751 4951 20757
rect 5537 20791 5595 20797
rect 5537 20757 5549 20791
rect 5583 20757 5595 20791
rect 5537 20751 5595 20757
rect 7466 20748 7472 20800
rect 7524 20788 7530 20800
rect 7561 20791 7619 20797
rect 7561 20788 7573 20791
rect 7524 20760 7573 20788
rect 7524 20748 7530 20760
rect 7561 20757 7573 20760
rect 7607 20757 7619 20791
rect 8110 20788 8116 20800
rect 8071 20760 8116 20788
rect 7561 20751 7619 20757
rect 8110 20748 8116 20760
rect 8168 20748 8174 20800
rect 9232 20788 9260 20819
rect 13004 20800 13032 20828
rect 14090 20816 14096 20868
rect 14148 20856 14154 20868
rect 14461 20859 14519 20865
rect 14461 20856 14473 20859
rect 14148 20828 14473 20856
rect 14148 20816 14154 20828
rect 14461 20825 14473 20828
rect 14507 20825 14519 20859
rect 16114 20856 16120 20868
rect 16075 20828 16120 20856
rect 14461 20819 14519 20825
rect 16114 20816 16120 20828
rect 16172 20816 16178 20868
rect 16776 20856 16804 20887
rect 17221 20859 17279 20865
rect 17221 20856 17233 20859
rect 16776 20828 17233 20856
rect 17221 20825 17233 20828
rect 17267 20825 17279 20859
rect 17221 20819 17279 20825
rect 18046 20816 18052 20868
rect 18104 20856 18110 20868
rect 18248 20856 18276 20896
rect 18325 20893 18337 20896
rect 18371 20893 18383 20927
rect 18432 20924 18460 20964
rect 18601 20961 18613 20995
rect 18647 20992 18659 20995
rect 19058 20992 19064 21004
rect 18647 20964 19064 20992
rect 18647 20961 18659 20964
rect 18601 20955 18659 20961
rect 19058 20952 19064 20964
rect 19116 20952 19122 21004
rect 22646 20992 22652 21004
rect 22296 20964 22652 20992
rect 18490 20927 18548 20933
rect 18490 20924 18502 20927
rect 18432 20896 18502 20924
rect 18325 20887 18383 20893
rect 18490 20893 18502 20896
rect 18536 20893 18548 20927
rect 18490 20887 18548 20893
rect 18693 20927 18751 20933
rect 18693 20893 18705 20927
rect 18739 20924 18751 20927
rect 18782 20924 18788 20936
rect 18739 20896 18788 20924
rect 18739 20893 18751 20896
rect 18693 20887 18751 20893
rect 18782 20884 18788 20896
rect 18840 20884 18846 20936
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 18892 20856 18920 20887
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19610 20924 19616 20936
rect 19392 20896 19616 20924
rect 19392 20884 19398 20896
rect 19610 20884 19616 20896
rect 19668 20884 19674 20936
rect 20714 20924 20720 20936
rect 20675 20896 20720 20924
rect 20714 20884 20720 20896
rect 20772 20884 20778 20936
rect 20898 20884 20904 20936
rect 20956 20924 20962 20936
rect 20956 20896 22140 20924
rect 20956 20884 20962 20896
rect 18104 20828 18276 20856
rect 18432 20828 18920 20856
rect 18104 20816 18110 20828
rect 9769 20791 9827 20797
rect 9769 20788 9781 20791
rect 9232 20760 9781 20788
rect 9769 20757 9781 20760
rect 9815 20788 9827 20791
rect 11514 20788 11520 20800
rect 9815 20760 11520 20788
rect 9815 20757 9827 20760
rect 9769 20751 9827 20757
rect 11514 20748 11520 20760
rect 11572 20748 11578 20800
rect 12986 20788 12992 20800
rect 12947 20760 12992 20788
rect 12986 20748 12992 20760
rect 13044 20748 13050 20800
rect 13449 20791 13507 20797
rect 13449 20757 13461 20791
rect 13495 20788 13507 20791
rect 13630 20788 13636 20800
rect 13495 20760 13636 20788
rect 13495 20757 13507 20760
rect 13449 20751 13507 20757
rect 13630 20748 13636 20760
rect 13688 20748 13694 20800
rect 15470 20748 15476 20800
rect 15528 20788 15534 20800
rect 15746 20788 15752 20800
rect 15528 20760 15752 20788
rect 15528 20748 15534 20760
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 16666 20788 16672 20800
rect 16627 20760 16672 20788
rect 16666 20748 16672 20760
rect 16724 20748 16730 20800
rect 17402 20748 17408 20800
rect 17460 20788 17466 20800
rect 17681 20791 17739 20797
rect 17681 20788 17693 20791
rect 17460 20760 17693 20788
rect 17460 20748 17466 20760
rect 17681 20757 17693 20760
rect 17727 20757 17739 20791
rect 17681 20751 17739 20757
rect 17773 20791 17831 20797
rect 17773 20757 17785 20791
rect 17819 20788 17831 20791
rect 18432 20788 18460 20828
rect 17819 20760 18460 20788
rect 18892 20788 18920 20828
rect 19061 20859 19119 20865
rect 19061 20825 19073 20859
rect 19107 20856 19119 20859
rect 20450 20859 20508 20865
rect 20450 20856 20462 20859
rect 19107 20828 20462 20856
rect 19107 20825 19119 20828
rect 19061 20819 19119 20825
rect 20450 20825 20462 20828
rect 20496 20825 20508 20859
rect 20450 20819 20508 20825
rect 20806 20816 20812 20868
rect 20864 20856 20870 20868
rect 22014 20859 22072 20865
rect 22014 20856 22026 20859
rect 20864 20828 22026 20856
rect 20864 20816 20870 20828
rect 22014 20825 22026 20828
rect 22060 20825 22072 20859
rect 22112 20856 22140 20896
rect 22186 20884 22192 20936
rect 22244 20924 22250 20936
rect 22296 20933 22324 20964
rect 22646 20952 22652 20964
rect 22704 20952 22710 21004
rect 22281 20927 22339 20933
rect 22281 20924 22293 20927
rect 22244 20896 22293 20924
rect 22244 20884 22250 20896
rect 22281 20893 22293 20896
rect 22327 20893 22339 20927
rect 22281 20887 22339 20893
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20924 22615 20927
rect 22756 20924 22784 21032
rect 23382 21020 23388 21072
rect 23440 21020 23446 21072
rect 23937 21063 23995 21069
rect 23937 21029 23949 21063
rect 23983 21060 23995 21063
rect 24118 21060 24124 21072
rect 23983 21032 24124 21060
rect 23983 21029 23995 21032
rect 23937 21023 23995 21029
rect 24118 21020 24124 21032
rect 24176 21020 24182 21072
rect 23106 20952 23112 21004
rect 23164 20992 23170 21004
rect 23400 20992 23428 21020
rect 23164 20964 23612 20992
rect 23164 20952 23170 20964
rect 22603 20896 22784 20924
rect 22603 20893 22615 20896
rect 22557 20887 22615 20893
rect 23198 20884 23204 20936
rect 23256 20924 23262 20936
rect 23584 20933 23612 20964
rect 23385 20927 23443 20933
rect 23385 20924 23397 20927
rect 23256 20896 23397 20924
rect 23256 20884 23262 20896
rect 23385 20893 23397 20896
rect 23431 20893 23443 20927
rect 23385 20887 23443 20893
rect 23569 20927 23627 20933
rect 23569 20893 23581 20927
rect 23615 20893 23627 20927
rect 23569 20887 23627 20893
rect 23805 20927 23863 20933
rect 23805 20893 23817 20927
rect 23851 20924 23863 20927
rect 23934 20924 23940 20936
rect 23851 20896 23940 20924
rect 23851 20893 23863 20896
rect 23805 20887 23863 20893
rect 23934 20884 23940 20896
rect 23992 20884 23998 20936
rect 23661 20859 23719 20865
rect 23661 20856 23673 20859
rect 22112 20828 23673 20856
rect 22014 20819 22072 20825
rect 23661 20825 23673 20828
rect 23707 20856 23719 20859
rect 24121 20859 24179 20865
rect 24121 20856 24133 20859
rect 23707 20828 24133 20856
rect 23707 20825 23719 20828
rect 23661 20819 23719 20825
rect 24121 20825 24133 20828
rect 24167 20856 24179 20859
rect 25590 20856 25596 20868
rect 24167 20828 25596 20856
rect 24167 20825 24179 20828
rect 24121 20819 24179 20825
rect 25590 20816 25596 20828
rect 25648 20816 25654 20868
rect 19337 20791 19395 20797
rect 19337 20788 19349 20791
rect 18892 20760 19349 20788
rect 17819 20757 17831 20760
rect 17773 20751 17831 20757
rect 19337 20757 19349 20760
rect 19383 20757 19395 20791
rect 19337 20751 19395 20757
rect 20346 20748 20352 20800
rect 20404 20788 20410 20800
rect 20901 20791 20959 20797
rect 20901 20788 20913 20791
rect 20404 20760 20913 20788
rect 20404 20748 20410 20760
rect 20901 20757 20913 20760
rect 20947 20757 20959 20791
rect 20901 20751 20959 20757
rect 22186 20748 22192 20800
rect 22244 20788 22250 20800
rect 22373 20791 22431 20797
rect 22373 20788 22385 20791
rect 22244 20760 22385 20788
rect 22244 20748 22250 20760
rect 22373 20757 22385 20760
rect 22419 20757 22431 20791
rect 22373 20751 22431 20757
rect 23106 20748 23112 20800
rect 23164 20788 23170 20800
rect 23201 20791 23259 20797
rect 23201 20788 23213 20791
rect 23164 20760 23213 20788
rect 23164 20748 23170 20760
rect 23201 20757 23213 20760
rect 23247 20757 23259 20791
rect 23201 20751 23259 20757
rect 1104 20698 29440 20720
rect 1104 20646 10395 20698
rect 10447 20646 10459 20698
rect 10511 20646 10523 20698
rect 10575 20646 10587 20698
rect 10639 20646 10651 20698
rect 10703 20646 19840 20698
rect 19892 20646 19904 20698
rect 19956 20646 19968 20698
rect 20020 20646 20032 20698
rect 20084 20646 20096 20698
rect 20148 20646 29440 20698
rect 1104 20624 29440 20646
rect 2406 20584 2412 20596
rect 2367 20556 2412 20584
rect 2406 20544 2412 20556
rect 2464 20544 2470 20596
rect 2501 20587 2559 20593
rect 2501 20553 2513 20587
rect 2547 20584 2559 20587
rect 3050 20584 3056 20596
rect 2547 20556 3056 20584
rect 2547 20553 2559 20556
rect 2501 20547 2559 20553
rect 3050 20544 3056 20556
rect 3108 20544 3114 20596
rect 3970 20584 3976 20596
rect 3931 20556 3976 20584
rect 3970 20544 3976 20556
rect 4028 20544 4034 20596
rect 6089 20587 6147 20593
rect 6089 20553 6101 20587
rect 6135 20584 6147 20587
rect 6362 20584 6368 20596
rect 6135 20556 6368 20584
rect 6135 20553 6147 20556
rect 6089 20547 6147 20553
rect 6362 20544 6368 20556
rect 6420 20544 6426 20596
rect 6454 20544 6460 20596
rect 6512 20584 6518 20596
rect 6914 20584 6920 20596
rect 6512 20556 6557 20584
rect 6875 20556 6920 20584
rect 6512 20544 6518 20556
rect 6914 20544 6920 20556
rect 6972 20544 6978 20596
rect 9585 20587 9643 20593
rect 9585 20553 9597 20587
rect 9631 20584 9643 20587
rect 9861 20587 9919 20593
rect 9861 20584 9873 20587
rect 9631 20556 9873 20584
rect 9631 20553 9643 20556
rect 9585 20547 9643 20553
rect 9861 20553 9873 20556
rect 9907 20553 9919 20587
rect 9861 20547 9919 20553
rect 10229 20587 10287 20593
rect 10229 20553 10241 20587
rect 10275 20584 10287 20587
rect 13817 20587 13875 20593
rect 13817 20584 13829 20587
rect 10275 20556 13829 20584
rect 10275 20553 10287 20556
rect 10229 20547 10287 20553
rect 13817 20553 13829 20556
rect 13863 20553 13875 20587
rect 17310 20584 17316 20596
rect 17271 20556 17316 20584
rect 13817 20547 13875 20553
rect 17310 20544 17316 20556
rect 17368 20544 17374 20596
rect 17773 20587 17831 20593
rect 17773 20553 17785 20587
rect 17819 20584 17831 20587
rect 20346 20584 20352 20596
rect 17819 20556 20352 20584
rect 17819 20553 17831 20556
rect 17773 20547 17831 20553
rect 20346 20544 20352 20556
rect 20404 20544 20410 20596
rect 20441 20587 20499 20593
rect 20441 20553 20453 20587
rect 20487 20584 20499 20587
rect 20806 20584 20812 20596
rect 20487 20556 20812 20584
rect 20487 20553 20499 20556
rect 20441 20547 20499 20553
rect 20806 20544 20812 20556
rect 20864 20544 20870 20596
rect 21542 20544 21548 20596
rect 21600 20584 21606 20596
rect 21913 20587 21971 20593
rect 21913 20584 21925 20587
rect 21600 20556 21925 20584
rect 21600 20544 21606 20556
rect 21913 20553 21925 20556
rect 21959 20553 21971 20587
rect 23382 20584 23388 20596
rect 21913 20547 21971 20553
rect 22112 20556 23388 20584
rect 1854 20516 1860 20528
rect 1815 20488 1860 20516
rect 1854 20476 1860 20488
rect 1912 20476 1918 20528
rect 2041 20519 2099 20525
rect 2041 20485 2053 20519
rect 2087 20516 2099 20519
rect 2958 20516 2964 20528
rect 2087 20488 2964 20516
rect 2087 20485 2099 20488
rect 2041 20479 2099 20485
rect 2958 20476 2964 20488
rect 3016 20476 3022 20528
rect 3326 20476 3332 20528
rect 3384 20476 3390 20528
rect 4246 20516 4252 20528
rect 3620 20488 4252 20516
rect 2593 20451 2651 20457
rect 2593 20417 2605 20451
rect 2639 20448 2651 20451
rect 2866 20448 2872 20460
rect 2639 20420 2872 20448
rect 2639 20417 2651 20420
rect 2593 20411 2651 20417
rect 2866 20408 2872 20420
rect 2924 20448 2930 20460
rect 3344 20448 3372 20476
rect 3620 20460 3648 20488
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 7377 20519 7435 20525
rect 7377 20485 7389 20519
rect 7423 20516 7435 20519
rect 7466 20516 7472 20528
rect 7423 20488 7472 20516
rect 7423 20485 7435 20488
rect 7377 20479 7435 20485
rect 7466 20476 7472 20488
rect 7524 20476 7530 20528
rect 8110 20476 8116 20528
rect 8168 20476 8174 20528
rect 10321 20519 10379 20525
rect 10321 20485 10333 20519
rect 10367 20516 10379 20519
rect 13906 20516 13912 20528
rect 10367 20488 12204 20516
rect 10367 20485 10379 20488
rect 10321 20479 10379 20485
rect 12176 20460 12204 20488
rect 12636 20488 13912 20516
rect 3602 20448 3608 20460
rect 2924 20420 3372 20448
rect 3563 20420 3608 20448
rect 2924 20408 2930 20420
rect 3602 20408 3608 20420
rect 3660 20408 3666 20460
rect 4154 20408 4160 20460
rect 4212 20448 4218 20460
rect 4433 20451 4491 20457
rect 4433 20448 4445 20451
rect 4212 20420 4445 20448
rect 4212 20408 4218 20420
rect 4433 20417 4445 20420
rect 4479 20417 4491 20451
rect 4433 20411 4491 20417
rect 4976 20451 5034 20457
rect 4976 20417 4988 20451
rect 5022 20448 5034 20451
rect 5258 20448 5264 20460
rect 5022 20420 5264 20448
rect 5022 20417 5034 20420
rect 4976 20411 5034 20417
rect 5258 20408 5264 20420
rect 5316 20408 5322 20460
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20448 6607 20451
rect 6638 20448 6644 20460
rect 6595 20420 6644 20448
rect 6595 20417 6607 20420
rect 6549 20411 6607 20417
rect 6638 20408 6644 20420
rect 6696 20408 6702 20460
rect 6730 20408 6736 20460
rect 6788 20448 6794 20460
rect 6825 20451 6883 20457
rect 6825 20448 6837 20451
rect 6788 20420 6837 20448
rect 6788 20408 6794 20420
rect 6825 20417 6837 20420
rect 6871 20417 6883 20451
rect 6825 20411 6883 20417
rect 10042 20408 10048 20460
rect 10100 20448 10106 20460
rect 10686 20448 10692 20460
rect 10100 20420 10692 20448
rect 10100 20408 10106 20420
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 10962 20408 10968 20460
rect 11020 20448 11026 20460
rect 11149 20451 11207 20457
rect 11149 20448 11161 20451
rect 11020 20420 11161 20448
rect 11020 20408 11026 20420
rect 11149 20417 11161 20420
rect 11195 20417 11207 20451
rect 11149 20411 11207 20417
rect 11238 20408 11244 20460
rect 11296 20448 11302 20460
rect 11517 20451 11575 20457
rect 11296 20420 11341 20448
rect 11296 20408 11302 20420
rect 11517 20417 11529 20451
rect 11563 20448 11575 20451
rect 11606 20448 11612 20460
rect 11563 20420 11612 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 11606 20408 11612 20420
rect 11664 20408 11670 20460
rect 11793 20451 11851 20457
rect 11793 20417 11805 20451
rect 11839 20417 11851 20451
rect 11974 20448 11980 20460
rect 11935 20420 11980 20448
rect 11793 20411 11851 20417
rect 2297 20383 2355 20389
rect 2297 20380 2309 20383
rect 1688 20352 2309 20380
rect 1394 20204 1400 20256
rect 1452 20244 1458 20256
rect 1688 20253 1716 20352
rect 2297 20349 2309 20352
rect 2343 20349 2355 20383
rect 2297 20343 2355 20349
rect 3050 20340 3056 20392
rect 3108 20380 3114 20392
rect 3234 20380 3240 20392
rect 3108 20352 3240 20380
rect 3108 20340 3114 20352
rect 3234 20340 3240 20352
rect 3292 20380 3298 20392
rect 3329 20383 3387 20389
rect 3329 20380 3341 20383
rect 3292 20352 3341 20380
rect 3292 20340 3298 20352
rect 3329 20349 3341 20352
rect 3375 20349 3387 20383
rect 3510 20380 3516 20392
rect 3471 20352 3516 20380
rect 3329 20343 3387 20349
rect 3510 20340 3516 20352
rect 3568 20340 3574 20392
rect 4706 20380 4712 20392
rect 4667 20352 4712 20380
rect 4706 20340 4712 20352
rect 4764 20340 4770 20392
rect 7101 20383 7159 20389
rect 7101 20349 7113 20383
rect 7147 20380 7159 20383
rect 7466 20380 7472 20392
rect 7147 20352 7472 20380
rect 7147 20349 7159 20352
rect 7101 20343 7159 20349
rect 7466 20340 7472 20352
rect 7524 20380 7530 20392
rect 8110 20380 8116 20392
rect 7524 20352 8116 20380
rect 7524 20340 7530 20352
rect 8110 20340 8116 20352
rect 8168 20340 8174 20392
rect 9493 20383 9551 20389
rect 9493 20349 9505 20383
rect 9539 20349 9551 20383
rect 9674 20380 9680 20392
rect 9635 20352 9680 20380
rect 9493 20343 9551 20349
rect 9122 20312 9128 20324
rect 9083 20284 9128 20312
rect 9122 20272 9128 20284
rect 9180 20272 9186 20324
rect 1673 20247 1731 20253
rect 1673 20244 1685 20247
rect 1452 20216 1685 20244
rect 1452 20204 1458 20216
rect 1673 20213 1685 20216
rect 1719 20213 1731 20247
rect 4338 20244 4344 20256
rect 4299 20216 4344 20244
rect 1673 20207 1731 20213
rect 4338 20204 4344 20216
rect 4396 20204 4402 20256
rect 6638 20244 6644 20256
rect 6599 20216 6644 20244
rect 6638 20204 6644 20216
rect 6696 20204 6702 20256
rect 8386 20204 8392 20256
rect 8444 20244 8450 20256
rect 8849 20247 8907 20253
rect 8849 20244 8861 20247
rect 8444 20216 8861 20244
rect 8444 20204 8450 20216
rect 8849 20213 8861 20216
rect 8895 20244 8907 20247
rect 9508 20244 9536 20343
rect 9674 20340 9680 20352
rect 9732 20340 9738 20392
rect 10505 20383 10563 20389
rect 10505 20349 10517 20383
rect 10551 20380 10563 20383
rect 10980 20380 11008 20408
rect 10551 20352 11008 20380
rect 11808 20380 11836 20411
rect 11974 20408 11980 20420
rect 12032 20408 12038 20460
rect 12158 20408 12164 20460
rect 12216 20448 12222 20460
rect 12636 20457 12664 20488
rect 13906 20476 13912 20488
rect 13964 20476 13970 20528
rect 14369 20519 14427 20525
rect 14369 20485 14381 20519
rect 14415 20516 14427 20519
rect 14826 20516 14832 20528
rect 14415 20488 14832 20516
rect 14415 20485 14427 20488
rect 14369 20479 14427 20485
rect 14826 20476 14832 20488
rect 14884 20476 14890 20528
rect 15304 20488 16804 20516
rect 12529 20451 12587 20457
rect 12216 20420 12309 20448
rect 12216 20408 12222 20420
rect 12529 20417 12541 20451
rect 12575 20417 12587 20451
rect 12529 20411 12587 20417
rect 12621 20451 12679 20457
rect 12621 20417 12633 20451
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20448 12955 20451
rect 13078 20448 13084 20460
rect 12943 20420 13084 20448
rect 12943 20417 12955 20420
rect 12897 20411 12955 20417
rect 12544 20380 12572 20411
rect 13078 20408 13084 20420
rect 13136 20408 13142 20460
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20448 13231 20451
rect 13354 20448 13360 20460
rect 13219 20420 13360 20448
rect 13219 20417 13231 20420
rect 13173 20411 13231 20417
rect 13354 20408 13360 20420
rect 13412 20408 13418 20460
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20448 13507 20451
rect 14090 20448 14096 20460
rect 13495 20420 14096 20448
rect 13495 20417 13507 20420
rect 13449 20411 13507 20417
rect 14090 20408 14096 20420
rect 14148 20408 14154 20460
rect 14182 20408 14188 20460
rect 14240 20448 14246 20460
rect 14553 20451 14611 20457
rect 14553 20448 14565 20451
rect 14240 20420 14565 20448
rect 14240 20408 14246 20420
rect 14553 20417 14565 20420
rect 14599 20417 14611 20451
rect 14553 20411 14611 20417
rect 14737 20451 14795 20457
rect 14737 20417 14749 20451
rect 14783 20417 14795 20451
rect 14737 20411 14795 20417
rect 13981 20383 14039 20389
rect 11808 20352 12434 20380
rect 12544 20352 12756 20380
rect 10551 20349 10563 20352
rect 10505 20343 10563 20349
rect 10778 20312 10784 20324
rect 10691 20284 10784 20312
rect 10778 20272 10784 20284
rect 10836 20312 10842 20324
rect 10836 20284 11100 20312
rect 10836 20272 10842 20284
rect 8895 20216 9536 20244
rect 11072 20244 11100 20284
rect 11146 20272 11152 20324
rect 11204 20312 11210 20324
rect 11609 20315 11667 20321
rect 11609 20312 11621 20315
rect 11204 20284 11621 20312
rect 11204 20272 11210 20284
rect 11609 20281 11621 20284
rect 11655 20281 11667 20315
rect 12406 20312 12434 20352
rect 12621 20315 12679 20321
rect 12621 20312 12633 20315
rect 12406 20284 12633 20312
rect 11609 20275 11667 20281
rect 12621 20281 12633 20284
rect 12667 20281 12679 20315
rect 12621 20275 12679 20281
rect 12728 20244 12756 20352
rect 13981 20349 13993 20383
rect 14027 20380 14039 20383
rect 14366 20380 14372 20392
rect 14027 20352 14372 20380
rect 14027 20349 14039 20352
rect 13981 20343 14039 20349
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 14461 20383 14519 20389
rect 14461 20349 14473 20383
rect 14507 20380 14519 20383
rect 14642 20380 14648 20392
rect 14507 20352 14648 20380
rect 14507 20349 14519 20352
rect 14461 20343 14519 20349
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 13630 20272 13636 20324
rect 13688 20312 13694 20324
rect 14752 20312 14780 20411
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 15304 20457 15332 20488
rect 16776 20460 16804 20488
rect 15289 20451 15347 20457
rect 15289 20448 15301 20451
rect 15252 20420 15301 20448
rect 15252 20408 15258 20420
rect 15289 20417 15301 20420
rect 15335 20417 15347 20451
rect 15289 20411 15347 20417
rect 15381 20451 15439 20457
rect 15381 20417 15393 20451
rect 15427 20448 15439 20451
rect 15654 20448 15660 20460
rect 15427 20420 15660 20448
rect 15427 20417 15439 20420
rect 15381 20411 15439 20417
rect 15105 20383 15163 20389
rect 15105 20349 15117 20383
rect 15151 20380 15163 20383
rect 15396 20380 15424 20411
rect 15654 20408 15660 20420
rect 15712 20408 15718 20460
rect 15746 20408 15752 20460
rect 15804 20448 15810 20460
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 15804 20420 15853 20448
rect 15804 20408 15810 20420
rect 15841 20417 15853 20420
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 16022 20408 16028 20460
rect 16080 20448 16086 20460
rect 16117 20451 16175 20457
rect 16117 20448 16129 20451
rect 16080 20420 16129 20448
rect 16080 20408 16086 20420
rect 16117 20417 16129 20420
rect 16163 20417 16175 20451
rect 16298 20448 16304 20460
rect 16259 20420 16304 20448
rect 16117 20411 16175 20417
rect 16298 20408 16304 20420
rect 16356 20408 16362 20460
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 15930 20380 15936 20392
rect 15151 20352 15424 20380
rect 15891 20352 15936 20380
rect 15151 20349 15163 20352
rect 15105 20343 15163 20349
rect 15930 20340 15936 20352
rect 15988 20340 15994 20392
rect 16684 20380 16712 20411
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 16816 20420 16909 20448
rect 16816 20408 16822 20420
rect 17494 20408 17500 20460
rect 17552 20448 17558 20460
rect 17681 20451 17739 20457
rect 17681 20448 17693 20451
rect 17552 20420 17693 20448
rect 17552 20408 17558 20420
rect 17681 20417 17693 20420
rect 17727 20417 17739 20451
rect 17681 20411 17739 20417
rect 18414 20408 18420 20460
rect 18472 20448 18478 20460
rect 18601 20451 18659 20457
rect 18601 20448 18613 20451
rect 18472 20420 18613 20448
rect 18472 20408 18478 20420
rect 18601 20417 18613 20420
rect 18647 20417 18659 20451
rect 18601 20411 18659 20417
rect 18690 20408 18696 20460
rect 18748 20448 18754 20460
rect 18877 20451 18935 20457
rect 18877 20448 18889 20451
rect 18748 20420 18889 20448
rect 18748 20408 18754 20420
rect 18877 20417 18889 20420
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 19242 20408 19248 20460
rect 19300 20448 19306 20460
rect 20364 20457 20392 20544
rect 22112 20528 22140 20556
rect 23382 20544 23388 20556
rect 23440 20584 23446 20596
rect 25590 20584 25596 20596
rect 23440 20556 23704 20584
rect 25551 20556 25596 20584
rect 23440 20544 23446 20556
rect 20530 20476 20536 20528
rect 20588 20516 20594 20528
rect 21453 20519 21511 20525
rect 21453 20516 21465 20519
rect 20588 20488 21465 20516
rect 20588 20476 20594 20488
rect 21453 20485 21465 20488
rect 21499 20485 21511 20519
rect 21453 20479 21511 20485
rect 21637 20519 21695 20525
rect 21637 20485 21649 20519
rect 21683 20516 21695 20519
rect 22094 20516 22100 20528
rect 21683 20488 22100 20516
rect 21683 20485 21695 20488
rect 21637 20479 21695 20485
rect 22094 20476 22100 20488
rect 22152 20476 22158 20528
rect 22370 20476 22376 20528
rect 22428 20476 22434 20528
rect 19797 20451 19855 20457
rect 19797 20448 19809 20451
rect 19300 20420 19809 20448
rect 19300 20408 19306 20420
rect 19797 20417 19809 20420
rect 19843 20417 19855 20451
rect 19797 20411 19855 20417
rect 19980 20451 20038 20457
rect 19980 20417 19992 20451
rect 20026 20448 20038 20451
rect 20349 20451 20407 20457
rect 20026 20420 20300 20448
rect 20026 20417 20038 20420
rect 19980 20411 20038 20417
rect 16132 20352 16712 20380
rect 17865 20383 17923 20389
rect 16132 20324 16160 20352
rect 17865 20349 17877 20383
rect 17911 20380 17923 20383
rect 17954 20380 17960 20392
rect 17911 20352 17960 20380
rect 17911 20349 17923 20352
rect 17865 20343 17923 20349
rect 17954 20340 17960 20352
rect 18012 20380 18018 20392
rect 18966 20380 18972 20392
rect 18012 20352 18972 20380
rect 18012 20340 18018 20352
rect 18966 20340 18972 20352
rect 19024 20340 19030 20392
rect 20073 20383 20131 20389
rect 20073 20349 20085 20383
rect 20119 20349 20131 20383
rect 20073 20343 20131 20349
rect 20165 20383 20223 20389
rect 20165 20349 20177 20383
rect 20211 20349 20223 20383
rect 20272 20380 20300 20420
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 20438 20408 20444 20460
rect 20496 20448 20502 20460
rect 23676 20457 23704 20556
rect 25590 20544 25596 20556
rect 25648 20544 25654 20596
rect 24118 20516 24124 20528
rect 24079 20488 24124 20516
rect 24118 20476 24124 20488
rect 24176 20476 24182 20528
rect 25130 20476 25136 20528
rect 25188 20476 25194 20528
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 20496 20420 20637 20448
rect 20496 20408 20502 20420
rect 20625 20417 20637 20420
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 23661 20451 23719 20457
rect 23661 20417 23673 20451
rect 23707 20448 23719 20451
rect 23845 20451 23903 20457
rect 23845 20448 23857 20451
rect 23707 20420 23857 20448
rect 23707 20417 23719 20420
rect 23661 20411 23719 20417
rect 23845 20417 23857 20420
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 20456 20380 20484 20408
rect 20272 20352 20484 20380
rect 20165 20343 20223 20349
rect 13688 20284 14780 20312
rect 15013 20315 15071 20321
rect 13688 20272 13694 20284
rect 15013 20281 15025 20315
rect 15059 20281 15071 20315
rect 15013 20275 15071 20281
rect 13446 20244 13452 20256
rect 11072 20216 13452 20244
rect 8895 20213 8907 20216
rect 8849 20207 8907 20213
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 14550 20204 14556 20256
rect 14608 20244 14614 20256
rect 15028 20244 15056 20275
rect 15286 20272 15292 20324
rect 15344 20312 15350 20324
rect 15654 20312 15660 20324
rect 15344 20284 15660 20312
rect 15344 20272 15350 20284
rect 15654 20272 15660 20284
rect 15712 20272 15718 20324
rect 16114 20272 16120 20324
rect 16172 20272 16178 20324
rect 19058 20312 19064 20324
rect 19019 20284 19064 20312
rect 19058 20272 19064 20284
rect 19116 20312 19122 20324
rect 19610 20312 19616 20324
rect 19116 20284 19616 20312
rect 19116 20272 19122 20284
rect 19610 20272 19616 20284
rect 19668 20312 19674 20324
rect 20088 20312 20116 20343
rect 19668 20284 20116 20312
rect 20180 20312 20208 20343
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 23385 20383 23443 20389
rect 23385 20380 23397 20383
rect 23348 20352 23397 20380
rect 23348 20340 23354 20352
rect 23385 20349 23397 20352
rect 23431 20349 23443 20383
rect 23385 20343 23443 20349
rect 20438 20312 20444 20324
rect 20180 20284 20444 20312
rect 19668 20272 19674 20284
rect 14608 20216 15056 20244
rect 14608 20204 14614 20216
rect 16298 20204 16304 20256
rect 16356 20244 16362 20256
rect 16666 20244 16672 20256
rect 16356 20216 16672 20244
rect 16356 20204 16362 20216
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 17034 20244 17040 20256
rect 16995 20216 17040 20244
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 18782 20244 18788 20256
rect 18695 20216 18788 20244
rect 18782 20204 18788 20216
rect 18840 20244 18846 20256
rect 20180 20244 20208 20284
rect 20438 20272 20444 20284
rect 20496 20272 20502 20324
rect 18840 20216 20208 20244
rect 18840 20204 18846 20216
rect 1104 20154 29440 20176
rect 1104 20102 5672 20154
rect 5724 20102 5736 20154
rect 5788 20102 5800 20154
rect 5852 20102 5864 20154
rect 5916 20102 5928 20154
rect 5980 20102 15118 20154
rect 15170 20102 15182 20154
rect 15234 20102 15246 20154
rect 15298 20102 15310 20154
rect 15362 20102 15374 20154
rect 15426 20102 24563 20154
rect 24615 20102 24627 20154
rect 24679 20102 24691 20154
rect 24743 20102 24755 20154
rect 24807 20102 24819 20154
rect 24871 20102 29440 20154
rect 1104 20080 29440 20102
rect 2498 20040 2504 20052
rect 2459 20012 2504 20040
rect 2498 20000 2504 20012
rect 2556 20000 2562 20052
rect 2866 20040 2872 20052
rect 2827 20012 2872 20040
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 5258 20040 5264 20052
rect 5219 20012 5264 20040
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 7926 20040 7932 20052
rect 7887 20012 7932 20040
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 8202 20040 8208 20052
rect 8163 20012 8208 20040
rect 8202 20000 8208 20012
rect 8260 20040 8266 20052
rect 9033 20043 9091 20049
rect 9033 20040 9045 20043
rect 8260 20012 9045 20040
rect 8260 20000 8266 20012
rect 9033 20009 9045 20012
rect 9079 20009 9091 20043
rect 9033 20003 9091 20009
rect 10965 20043 11023 20049
rect 10965 20009 10977 20043
rect 11011 20040 11023 20043
rect 11146 20040 11152 20052
rect 11011 20012 11152 20040
rect 11011 20009 11023 20012
rect 10965 20003 11023 20009
rect 11146 20000 11152 20012
rect 11204 20040 11210 20052
rect 11974 20040 11980 20052
rect 11204 20012 11980 20040
rect 11204 20000 11210 20012
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 14553 20043 14611 20049
rect 14553 20040 14565 20043
rect 13872 20012 14565 20040
rect 13872 20000 13878 20012
rect 14553 20009 14565 20012
rect 14599 20009 14611 20043
rect 14553 20003 14611 20009
rect 14921 20043 14979 20049
rect 14921 20009 14933 20043
rect 14967 20040 14979 20043
rect 15562 20040 15568 20052
rect 14967 20012 15568 20040
rect 14967 20009 14979 20012
rect 14921 20003 14979 20009
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 15746 20040 15752 20052
rect 15707 20012 15752 20040
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 16574 20040 16580 20052
rect 16535 20012 16580 20040
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 18141 20043 18199 20049
rect 18141 20009 18153 20043
rect 18187 20040 18199 20043
rect 18414 20040 18420 20052
rect 18187 20012 18420 20040
rect 18187 20009 18199 20012
rect 18141 20003 18199 20009
rect 18414 20000 18420 20012
rect 18472 20000 18478 20052
rect 22370 20040 22376 20052
rect 22331 20012 22376 20040
rect 22370 20000 22376 20012
rect 22428 20000 22434 20052
rect 23201 20043 23259 20049
rect 23201 20009 23213 20043
rect 23247 20040 23259 20043
rect 23290 20040 23296 20052
rect 23247 20012 23296 20040
rect 23247 20009 23259 20012
rect 23201 20003 23259 20009
rect 23290 20000 23296 20012
rect 23348 20000 23354 20052
rect 24394 20040 24400 20052
rect 24355 20012 24400 20040
rect 24394 20000 24400 20012
rect 24452 20000 24458 20052
rect 25130 20040 25136 20052
rect 25091 20012 25136 20040
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 3421 19975 3479 19981
rect 3421 19941 3433 19975
rect 3467 19972 3479 19975
rect 4338 19972 4344 19984
rect 3467 19944 4344 19972
rect 3467 19941 3479 19944
rect 3421 19935 3479 19941
rect 4338 19932 4344 19944
rect 4396 19972 4402 19984
rect 4396 19944 4844 19972
rect 4396 19932 4402 19944
rect 3881 19907 3939 19913
rect 3881 19904 3893 19907
rect 3252 19876 3893 19904
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19836 2743 19839
rect 3051 19839 3109 19845
rect 3051 19836 3063 19839
rect 2731 19808 3063 19836
rect 2731 19805 2743 19808
rect 2685 19799 2743 19805
rect 3051 19805 3063 19808
rect 3097 19836 3109 19839
rect 3252 19836 3280 19876
rect 3881 19873 3893 19876
rect 3927 19873 3939 19907
rect 4614 19904 4620 19916
rect 4575 19876 4620 19904
rect 3881 19867 3939 19873
rect 4614 19864 4620 19876
rect 4672 19864 4678 19916
rect 4816 19913 4844 19944
rect 11072 19944 13308 19972
rect 4801 19907 4859 19913
rect 4801 19873 4813 19907
rect 4847 19873 4859 19907
rect 4801 19867 4859 19873
rect 3097 19808 3280 19836
rect 3513 19839 3571 19845
rect 3097 19805 3109 19808
rect 3051 19799 3109 19805
rect 3513 19805 3525 19839
rect 3559 19805 3571 19839
rect 3970 19836 3976 19848
rect 3931 19808 3976 19836
rect 3513 19799 3571 19805
rect 3234 19728 3240 19780
rect 3292 19768 3298 19780
rect 3528 19768 3556 19799
rect 3970 19796 3976 19808
rect 4028 19796 4034 19848
rect 6825 19839 6883 19845
rect 6825 19805 6837 19839
rect 6871 19836 6883 19839
rect 6914 19836 6920 19848
rect 6871 19808 6920 19836
rect 6871 19805 6883 19808
rect 6825 19799 6883 19805
rect 6914 19796 6920 19808
rect 6972 19796 6978 19848
rect 7742 19836 7748 19848
rect 7703 19808 7748 19836
rect 7742 19796 7748 19808
rect 7800 19796 7806 19848
rect 8294 19836 8300 19848
rect 8255 19808 8300 19836
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 10686 19796 10692 19848
rect 10744 19836 10750 19848
rect 11072 19845 11100 19944
rect 11238 19904 11244 19916
rect 11151 19876 11244 19904
rect 11238 19864 11244 19876
rect 11296 19904 11302 19916
rect 12621 19907 12679 19913
rect 12621 19904 12633 19907
rect 11296 19876 12633 19904
rect 11296 19864 11302 19876
rect 12621 19873 12633 19876
rect 12667 19873 12679 19907
rect 12621 19867 12679 19873
rect 11057 19839 11115 19845
rect 11057 19836 11069 19839
rect 10744 19808 11069 19836
rect 10744 19796 10750 19808
rect 11057 19805 11069 19808
rect 11103 19805 11115 19839
rect 11330 19836 11336 19848
rect 11291 19808 11336 19836
rect 11057 19799 11115 19805
rect 11330 19796 11336 19808
rect 11388 19796 11394 19848
rect 11422 19796 11428 19848
rect 11480 19836 11486 19848
rect 11609 19839 11667 19845
rect 11480 19808 11525 19836
rect 11480 19796 11486 19808
rect 11609 19805 11621 19839
rect 11655 19836 11667 19839
rect 11882 19836 11888 19848
rect 11655 19808 11888 19836
rect 11655 19805 11667 19808
rect 11609 19799 11667 19805
rect 11882 19796 11888 19808
rect 11940 19796 11946 19848
rect 12986 19836 12992 19848
rect 12947 19808 12992 19836
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 5350 19768 5356 19780
rect 3292 19740 5356 19768
rect 3292 19728 3298 19740
rect 5350 19728 5356 19740
rect 5408 19728 5414 19780
rect 6362 19728 6368 19780
rect 6420 19768 6426 19780
rect 6457 19771 6515 19777
rect 6457 19768 6469 19771
rect 6420 19740 6469 19768
rect 6420 19728 6426 19740
rect 6457 19737 6469 19740
rect 6503 19737 6515 19771
rect 6457 19731 6515 19737
rect 6638 19728 6644 19780
rect 6696 19768 6702 19780
rect 7282 19768 7288 19780
rect 6696 19740 7288 19768
rect 6696 19728 6702 19740
rect 7282 19728 7288 19740
rect 7340 19728 7346 19780
rect 12710 19728 12716 19780
rect 12768 19768 12774 19780
rect 12805 19771 12863 19777
rect 12805 19768 12817 19771
rect 12768 19740 12817 19768
rect 12768 19728 12774 19740
rect 12805 19737 12817 19740
rect 12851 19737 12863 19771
rect 13170 19768 13176 19780
rect 13131 19740 13176 19768
rect 12805 19731 12863 19737
rect 13170 19728 13176 19740
rect 13228 19728 13234 19780
rect 13280 19768 13308 19944
rect 17034 19932 17040 19984
rect 17092 19972 17098 19984
rect 22554 19972 22560 19984
rect 17092 19944 22560 19972
rect 17092 19932 17098 19944
rect 22554 19932 22560 19944
rect 22612 19932 22618 19984
rect 24121 19975 24179 19981
rect 24121 19941 24133 19975
rect 24167 19972 24179 19975
rect 25038 19972 25044 19984
rect 24167 19944 25044 19972
rect 24167 19941 24179 19944
rect 24121 19935 24179 19941
rect 25038 19932 25044 19944
rect 25096 19932 25102 19984
rect 13538 19864 13544 19916
rect 13596 19864 13602 19916
rect 14366 19864 14372 19916
rect 14424 19904 14430 19916
rect 15381 19907 15439 19913
rect 15381 19904 15393 19907
rect 14424 19876 15393 19904
rect 14424 19864 14430 19876
rect 15381 19873 15393 19876
rect 15427 19873 15439 19907
rect 17862 19904 17868 19916
rect 15381 19867 15439 19873
rect 16868 19876 17868 19904
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19836 13415 19839
rect 13556 19836 13584 19864
rect 14550 19836 14556 19848
rect 13403 19808 13584 19836
rect 14511 19808 14556 19836
rect 13403 19805 13415 19808
rect 13357 19799 13415 19805
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 14737 19839 14795 19845
rect 14737 19805 14749 19839
rect 14783 19805 14795 19839
rect 15562 19836 15568 19848
rect 15523 19808 15568 19836
rect 14737 19799 14795 19805
rect 13541 19771 13599 19777
rect 13541 19768 13553 19771
rect 13280 19740 13553 19768
rect 13541 19737 13553 19740
rect 13587 19768 13599 19771
rect 14752 19768 14780 19799
rect 15562 19796 15568 19808
rect 15620 19836 15626 19848
rect 16114 19836 16120 19848
rect 15620 19808 16120 19836
rect 15620 19796 15626 19808
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19836 16727 19839
rect 16758 19836 16764 19848
rect 16715 19808 16764 19836
rect 16715 19805 16727 19808
rect 16669 19799 16727 19805
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 16868 19845 16896 19876
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 23198 19904 23204 19916
rect 22664 19876 23204 19904
rect 16853 19839 16911 19845
rect 16853 19805 16865 19839
rect 16899 19805 16911 19839
rect 17954 19836 17960 19848
rect 17915 19808 17960 19836
rect 16853 19799 16911 19805
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19805 18291 19839
rect 22186 19836 22192 19848
rect 22147 19808 22192 19836
rect 18233 19799 18291 19805
rect 15470 19768 15476 19780
rect 13587 19740 15476 19768
rect 13587 19737 13599 19740
rect 13541 19731 13599 19737
rect 15470 19728 15476 19740
rect 15528 19728 15534 19780
rect 17770 19728 17776 19780
rect 17828 19768 17834 19780
rect 18248 19768 18276 19799
rect 22186 19796 22192 19808
rect 22244 19796 22250 19848
rect 22554 19796 22560 19848
rect 22612 19836 22618 19848
rect 22664 19845 22692 19876
rect 23198 19864 23204 19876
rect 23256 19864 23262 19916
rect 23492 19876 23980 19904
rect 22649 19839 22707 19845
rect 22649 19836 22661 19839
rect 22612 19808 22661 19836
rect 22612 19796 22618 19808
rect 22649 19805 22661 19808
rect 22695 19805 22707 19839
rect 22925 19839 22983 19845
rect 22925 19836 22937 19839
rect 22649 19799 22707 19805
rect 22756 19808 22937 19836
rect 17828 19740 18276 19768
rect 17828 19728 17834 19740
rect 21542 19728 21548 19780
rect 21600 19768 21606 19780
rect 22756 19768 22784 19808
rect 22925 19805 22937 19808
rect 22971 19805 22983 19839
rect 22925 19799 22983 19805
rect 23069 19839 23127 19845
rect 23069 19805 23081 19839
rect 23115 19836 23127 19839
rect 23492 19836 23520 19876
rect 23952 19848 23980 19876
rect 23115 19808 23520 19836
rect 23569 19839 23627 19845
rect 23115 19805 23127 19808
rect 23069 19799 23127 19805
rect 23569 19805 23581 19839
rect 23615 19805 23627 19839
rect 23569 19799 23627 19805
rect 21600 19740 22784 19768
rect 22833 19771 22891 19777
rect 21600 19728 21606 19740
rect 22833 19737 22845 19771
rect 22879 19737 22891 19771
rect 22833 19731 22891 19737
rect 3050 19700 3056 19712
rect 3011 19672 3056 19700
rect 3050 19660 3056 19672
rect 3108 19660 3114 19712
rect 4890 19660 4896 19712
rect 4948 19700 4954 19712
rect 6270 19700 6276 19712
rect 4948 19672 4993 19700
rect 6183 19672 6276 19700
rect 4948 19660 4954 19672
rect 6270 19660 6276 19672
rect 6328 19700 6334 19712
rect 6656 19700 6684 19728
rect 6328 19672 6684 19700
rect 6328 19660 6334 19672
rect 11238 19660 11244 19712
rect 11296 19700 11302 19712
rect 13630 19700 13636 19712
rect 11296 19672 13636 19700
rect 11296 19660 11302 19672
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 18417 19703 18475 19709
rect 18417 19669 18429 19703
rect 18463 19700 18475 19703
rect 18598 19700 18604 19712
rect 18463 19672 18604 19700
rect 18463 19669 18475 19672
rect 18417 19663 18475 19669
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 19702 19660 19708 19712
rect 19760 19700 19766 19712
rect 20254 19700 20260 19712
rect 19760 19672 20260 19700
rect 19760 19660 19766 19672
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 22557 19703 22615 19709
rect 22557 19669 22569 19703
rect 22603 19700 22615 19703
rect 22848 19700 22876 19731
rect 23198 19728 23204 19780
rect 23256 19768 23262 19780
rect 23584 19768 23612 19799
rect 23934 19796 23940 19848
rect 23992 19845 23998 19848
rect 23992 19836 24000 19845
rect 23992 19808 24037 19836
rect 23992 19799 24000 19808
rect 23992 19796 23998 19799
rect 24670 19796 24676 19848
rect 24728 19836 24734 19848
rect 24949 19839 25007 19845
rect 24949 19836 24961 19839
rect 24728 19808 24961 19836
rect 24728 19796 24734 19808
rect 24949 19805 24961 19808
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 23256 19740 23612 19768
rect 23753 19771 23811 19777
rect 23256 19728 23262 19740
rect 23753 19737 23765 19771
rect 23799 19737 23811 19771
rect 23753 19731 23811 19737
rect 23845 19771 23903 19777
rect 23845 19737 23857 19771
rect 23891 19768 23903 19771
rect 26510 19768 26516 19780
rect 23891 19740 26516 19768
rect 23891 19737 23903 19740
rect 23845 19731 23903 19737
rect 23014 19700 23020 19712
rect 22603 19672 23020 19700
rect 22603 19669 22615 19672
rect 22557 19663 22615 19669
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 23768 19700 23796 19731
rect 26510 19728 26516 19740
rect 26568 19768 26574 19780
rect 27522 19768 27528 19780
rect 26568 19740 27528 19768
rect 26568 19728 26574 19740
rect 27522 19728 27528 19740
rect 27580 19728 27586 19780
rect 24026 19700 24032 19712
rect 23768 19672 24032 19700
rect 24026 19660 24032 19672
rect 24084 19700 24090 19712
rect 24394 19700 24400 19712
rect 24084 19672 24400 19700
rect 24084 19660 24090 19672
rect 24394 19660 24400 19672
rect 24452 19660 24458 19712
rect 1104 19610 29440 19632
rect 1104 19558 10395 19610
rect 10447 19558 10459 19610
rect 10511 19558 10523 19610
rect 10575 19558 10587 19610
rect 10639 19558 10651 19610
rect 10703 19558 19840 19610
rect 19892 19558 19904 19610
rect 19956 19558 19968 19610
rect 20020 19558 20032 19610
rect 20084 19558 20096 19610
rect 20148 19558 29440 19610
rect 1104 19536 29440 19558
rect 2777 19499 2835 19505
rect 2777 19465 2789 19499
rect 2823 19496 2835 19499
rect 3602 19496 3608 19508
rect 2823 19468 3608 19496
rect 2823 19465 2835 19468
rect 2777 19459 2835 19465
rect 3602 19456 3608 19468
rect 3660 19456 3666 19508
rect 4338 19496 4344 19508
rect 4299 19468 4344 19496
rect 4338 19456 4344 19468
rect 4396 19456 4402 19508
rect 4801 19499 4859 19505
rect 4801 19465 4813 19499
rect 4847 19496 4859 19499
rect 8297 19499 8355 19505
rect 4847 19468 5304 19496
rect 4847 19465 4859 19468
rect 4801 19459 4859 19465
rect 4246 19388 4252 19440
rect 4304 19428 4310 19440
rect 5276 19437 5304 19468
rect 8297 19465 8309 19499
rect 8343 19465 8355 19499
rect 8297 19459 8355 19465
rect 5261 19431 5319 19437
rect 4304 19400 5120 19428
rect 4304 19388 4310 19400
rect 4430 19360 4436 19372
rect 4391 19332 4436 19360
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 4890 19320 4896 19372
rect 4948 19360 4954 19372
rect 5092 19369 5120 19400
rect 5261 19397 5273 19431
rect 5307 19397 5319 19431
rect 5261 19391 5319 19397
rect 5092 19363 5175 19369
rect 4948 19332 5028 19360
rect 5092 19332 5129 19363
rect 4948 19320 4954 19332
rect 2590 19252 2596 19304
rect 2648 19292 2654 19304
rect 2869 19295 2927 19301
rect 2869 19292 2881 19295
rect 2648 19264 2881 19292
rect 2648 19252 2654 19264
rect 2869 19261 2881 19264
rect 2915 19261 2927 19295
rect 3050 19292 3056 19304
rect 3011 19264 3056 19292
rect 2869 19255 2927 19261
rect 3050 19252 3056 19264
rect 3108 19292 3114 19304
rect 4157 19295 4215 19301
rect 4157 19292 4169 19295
rect 3108 19264 4169 19292
rect 3108 19252 3114 19264
rect 4157 19261 4169 19264
rect 4203 19292 4215 19295
rect 4522 19292 4528 19304
rect 4203 19264 4528 19292
rect 4203 19261 4215 19264
rect 4157 19255 4215 19261
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 5000 19233 5028 19332
rect 5117 19329 5129 19332
rect 5163 19329 5175 19363
rect 5350 19360 5356 19372
rect 5311 19332 5356 19360
rect 5117 19323 5175 19329
rect 5350 19320 5356 19332
rect 5408 19320 5414 19372
rect 5534 19360 5540 19372
rect 5495 19332 5540 19360
rect 5534 19320 5540 19332
rect 5592 19320 5598 19372
rect 6362 19360 6368 19372
rect 6323 19332 6368 19360
rect 6362 19320 6368 19332
rect 6420 19320 6426 19372
rect 7742 19320 7748 19372
rect 7800 19360 7806 19372
rect 8113 19363 8171 19369
rect 8113 19360 8125 19363
rect 7800 19332 8125 19360
rect 7800 19320 7806 19332
rect 8113 19329 8125 19332
rect 8159 19329 8171 19363
rect 8312 19360 8340 19459
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 10689 19499 10747 19505
rect 10689 19496 10701 19499
rect 9732 19468 10701 19496
rect 9732 19456 9738 19468
rect 10689 19465 10701 19468
rect 10735 19465 10747 19499
rect 11330 19496 11336 19508
rect 10689 19459 10747 19465
rect 10796 19468 11336 19496
rect 10413 19431 10471 19437
rect 10413 19397 10425 19431
rect 10459 19428 10471 19431
rect 10594 19428 10600 19440
rect 10459 19400 10600 19428
rect 10459 19397 10471 19400
rect 10413 19391 10471 19397
rect 10594 19388 10600 19400
rect 10652 19388 10658 19440
rect 8573 19363 8631 19369
rect 8573 19360 8585 19363
rect 8312 19332 8585 19360
rect 8113 19323 8171 19329
rect 8573 19329 8585 19332
rect 8619 19329 8631 19363
rect 8573 19323 8631 19329
rect 10505 19363 10563 19369
rect 10505 19329 10517 19363
rect 10551 19360 10563 19363
rect 10796 19360 10824 19468
rect 11330 19456 11336 19468
rect 11388 19456 11394 19508
rect 11974 19496 11980 19508
rect 11935 19468 11980 19496
rect 11974 19456 11980 19468
rect 12032 19496 12038 19508
rect 13173 19499 13231 19505
rect 12032 19468 12434 19496
rect 12032 19456 12038 19468
rect 11238 19428 11244 19440
rect 10888 19400 11244 19428
rect 10888 19369 10916 19400
rect 11238 19388 11244 19400
rect 11296 19388 11302 19440
rect 11606 19428 11612 19440
rect 11348 19400 11612 19428
rect 10551 19332 10824 19360
rect 10873 19363 10931 19369
rect 10551 19329 10563 19332
rect 10505 19323 10563 19329
rect 10873 19329 10885 19363
rect 10919 19329 10931 19363
rect 11054 19360 11060 19372
rect 11015 19332 11060 19360
rect 10873 19323 10931 19329
rect 11054 19320 11060 19332
rect 11112 19320 11118 19372
rect 11146 19320 11152 19372
rect 11204 19360 11210 19372
rect 11348 19369 11376 19400
rect 11606 19388 11612 19400
rect 11664 19388 11670 19440
rect 11698 19388 11704 19440
rect 11756 19428 11762 19440
rect 12250 19428 12256 19440
rect 11756 19400 12256 19428
rect 11756 19388 11762 19400
rect 12250 19388 12256 19400
rect 12308 19388 12314 19440
rect 12406 19428 12434 19468
rect 13173 19465 13185 19499
rect 13219 19496 13231 19499
rect 13722 19496 13728 19508
rect 13219 19468 13728 19496
rect 13219 19465 13231 19468
rect 13173 19459 13231 19465
rect 13722 19456 13728 19468
rect 13780 19456 13786 19508
rect 13998 19456 14004 19508
rect 14056 19496 14062 19508
rect 14366 19496 14372 19508
rect 14056 19468 14372 19496
rect 14056 19456 14062 19468
rect 14366 19456 14372 19468
rect 14424 19496 14430 19508
rect 14645 19499 14703 19505
rect 14645 19496 14657 19499
rect 14424 19468 14657 19496
rect 14424 19456 14430 19468
rect 14645 19465 14657 19468
rect 14691 19465 14703 19499
rect 14645 19459 14703 19465
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 12406 19400 14688 19428
rect 11333 19363 11391 19369
rect 11204 19332 11249 19360
rect 11204 19320 11210 19332
rect 11333 19329 11345 19363
rect 11379 19329 11391 19363
rect 11333 19323 11391 19329
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19360 11575 19363
rect 11716 19360 11744 19388
rect 14660 19372 14688 19400
rect 11563 19332 11744 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 12066 19320 12072 19372
rect 12124 19360 12130 19372
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 12124 19332 12173 19360
rect 12124 19320 12130 19332
rect 12161 19329 12173 19332
rect 12207 19329 12219 19363
rect 12161 19323 12219 19329
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19360 12587 19363
rect 12710 19360 12716 19372
rect 12575 19332 12716 19360
rect 12575 19329 12587 19332
rect 12529 19323 12587 19329
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 12802 19320 12808 19372
rect 12860 19360 12866 19372
rect 13078 19369 13084 19372
rect 12897 19363 12955 19369
rect 12897 19360 12909 19363
rect 12860 19332 12909 19360
rect 12860 19320 12866 19332
rect 12897 19329 12909 19332
rect 12943 19329 12955 19363
rect 12897 19323 12955 19329
rect 13035 19363 13084 19369
rect 13035 19329 13047 19363
rect 13081 19329 13084 19363
rect 13035 19323 13084 19329
rect 13078 19320 13084 19323
rect 13136 19320 13142 19372
rect 14642 19320 14648 19372
rect 14700 19320 14706 19372
rect 14826 19360 14832 19372
rect 14787 19332 14832 19360
rect 14826 19320 14832 19332
rect 14884 19320 14890 19372
rect 15838 19320 15844 19372
rect 15896 19360 15902 19372
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 15896 19332 16681 19360
rect 15896 19320 15902 19332
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 16868 19360 16896 19459
rect 18230 19456 18236 19508
rect 18288 19496 18294 19508
rect 18325 19499 18383 19505
rect 18325 19496 18337 19499
rect 18288 19468 18337 19496
rect 18288 19456 18294 19468
rect 18325 19465 18337 19468
rect 18371 19465 18383 19499
rect 19702 19496 19708 19508
rect 18325 19459 18383 19465
rect 19536 19468 19708 19496
rect 19536 19372 19564 19468
rect 19702 19456 19708 19468
rect 19760 19456 19766 19508
rect 19981 19499 20039 19505
rect 19981 19465 19993 19499
rect 20027 19496 20039 19499
rect 20254 19496 20260 19508
rect 20027 19468 20260 19496
rect 20027 19465 20039 19468
rect 19981 19459 20039 19465
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 20346 19456 20352 19508
rect 20404 19496 20410 19508
rect 21545 19499 21603 19505
rect 21545 19496 21557 19499
rect 20404 19468 21557 19496
rect 20404 19456 20410 19468
rect 21545 19465 21557 19468
rect 21591 19465 21603 19499
rect 24670 19496 24676 19508
rect 24631 19468 24676 19496
rect 21545 19459 21603 19465
rect 24670 19456 24676 19468
rect 24728 19456 24734 19508
rect 26510 19496 26516 19508
rect 26471 19468 26516 19496
rect 26510 19456 26516 19468
rect 26568 19456 26574 19508
rect 20070 19428 20076 19440
rect 19720 19400 20076 19428
rect 17129 19363 17187 19369
rect 17129 19360 17141 19363
rect 16868 19332 17141 19360
rect 16669 19323 16727 19329
rect 17129 19329 17141 19332
rect 17175 19329 17187 19363
rect 17129 19323 17187 19329
rect 17218 19320 17224 19372
rect 17276 19360 17282 19372
rect 17770 19360 17776 19372
rect 17276 19332 17776 19360
rect 17276 19320 17282 19332
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 17865 19363 17923 19369
rect 17865 19329 17877 19363
rect 17911 19360 17923 19363
rect 17954 19360 17960 19372
rect 17911 19332 17960 19360
rect 17911 19329 17923 19332
rect 17865 19323 17923 19329
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 18690 19360 18696 19372
rect 18651 19332 18696 19360
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 19242 19320 19248 19372
rect 19300 19360 19306 19372
rect 19337 19363 19395 19369
rect 19337 19360 19349 19363
rect 19300 19332 19349 19360
rect 19300 19320 19306 19332
rect 19337 19329 19349 19332
rect 19383 19329 19395 19363
rect 19337 19323 19395 19329
rect 19520 19366 19578 19372
rect 19520 19332 19532 19366
rect 19566 19332 19578 19366
rect 19520 19326 19578 19332
rect 12621 19295 12679 19301
rect 12621 19261 12633 19295
rect 12667 19261 12679 19295
rect 12728 19292 12756 19320
rect 13354 19292 13360 19304
rect 12728 19264 13360 19292
rect 12621 19255 12679 19261
rect 4985 19227 5043 19233
rect 4985 19193 4997 19227
rect 5031 19193 5043 19227
rect 4985 19187 5043 19193
rect 10965 19227 11023 19233
rect 10965 19193 10977 19227
rect 11011 19224 11023 19227
rect 12636 19224 12664 19255
rect 13354 19252 13360 19264
rect 13412 19292 13418 19304
rect 16206 19292 16212 19304
rect 13412 19264 16212 19292
rect 13412 19252 13418 19264
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 18782 19292 18788 19304
rect 18743 19264 18788 19292
rect 18782 19252 18788 19264
rect 18840 19252 18846 19304
rect 18966 19292 18972 19304
rect 18927 19264 18972 19292
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19610 19292 19616 19304
rect 19571 19264 19616 19292
rect 19610 19252 19616 19264
rect 19668 19252 19674 19304
rect 19720 19301 19748 19400
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 20714 19428 20720 19440
rect 20180 19400 20720 19428
rect 19886 19360 19892 19372
rect 19847 19332 19892 19360
rect 19886 19320 19892 19332
rect 19944 19320 19950 19372
rect 20180 19369 20208 19400
rect 20714 19388 20720 19400
rect 20772 19388 20778 19440
rect 23382 19388 23388 19440
rect 23440 19428 23446 19440
rect 25038 19428 25044 19440
rect 23440 19400 24808 19428
rect 24999 19400 25044 19428
rect 23440 19388 23446 19400
rect 20165 19363 20223 19369
rect 20165 19329 20177 19363
rect 20211 19329 20223 19363
rect 20165 19323 20223 19329
rect 19705 19295 19763 19301
rect 19705 19261 19717 19295
rect 19751 19261 19763 19295
rect 20180 19292 20208 19323
rect 20254 19320 20260 19372
rect 20312 19360 20318 19372
rect 20421 19363 20479 19369
rect 20421 19360 20433 19363
rect 20312 19332 20433 19360
rect 20312 19320 20318 19332
rect 20421 19329 20433 19332
rect 20467 19329 20479 19363
rect 24486 19360 24492 19372
rect 24447 19332 24492 19360
rect 20421 19323 20479 19329
rect 24486 19320 24492 19332
rect 24544 19320 24550 19372
rect 24780 19369 24808 19400
rect 25038 19388 25044 19400
rect 25096 19388 25102 19440
rect 26050 19388 26056 19440
rect 26108 19388 26114 19440
rect 24765 19363 24823 19369
rect 24765 19329 24777 19363
rect 24811 19329 24823 19363
rect 24765 19323 24823 19329
rect 19705 19255 19763 19261
rect 19812 19264 20208 19292
rect 11011 19196 11744 19224
rect 12636 19196 13032 19224
rect 11011 19193 11023 19196
rect 10965 19187 11023 19193
rect 2406 19156 2412 19168
rect 2367 19128 2412 19156
rect 2406 19116 2412 19128
rect 2464 19116 2470 19168
rect 5534 19116 5540 19168
rect 5592 19156 5598 19168
rect 5629 19159 5687 19165
rect 5629 19156 5641 19159
rect 5592 19128 5641 19156
rect 5592 19116 5598 19128
rect 5629 19125 5641 19128
rect 5675 19156 5687 19159
rect 6549 19159 6607 19165
rect 6549 19156 6561 19159
rect 5675 19128 6561 19156
rect 5675 19125 5687 19128
rect 5629 19119 5687 19125
rect 6549 19125 6561 19128
rect 6595 19125 6607 19159
rect 8754 19156 8760 19168
rect 8715 19128 8760 19156
rect 6549 19119 6607 19125
rect 8754 19116 8760 19128
rect 8812 19116 8818 19168
rect 11716 19165 11744 19196
rect 13004 19168 13032 19196
rect 18230 19184 18236 19236
rect 18288 19224 18294 19236
rect 19812 19224 19840 19264
rect 18288 19196 19840 19224
rect 18288 19184 18294 19196
rect 11701 19159 11759 19165
rect 11701 19125 11713 19159
rect 11747 19156 11759 19159
rect 12066 19156 12072 19168
rect 11747 19128 12072 19156
rect 11747 19125 11759 19128
rect 11701 19119 11759 19125
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 12986 19116 12992 19168
rect 13044 19116 13050 19168
rect 17310 19156 17316 19168
rect 17271 19128 17316 19156
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 19886 19116 19892 19168
rect 19944 19156 19950 19168
rect 20346 19156 20352 19168
rect 19944 19128 20352 19156
rect 19944 19116 19950 19128
rect 20346 19116 20352 19128
rect 20404 19116 20410 19168
rect 1104 19066 29440 19088
rect 1104 19014 5672 19066
rect 5724 19014 5736 19066
rect 5788 19014 5800 19066
rect 5852 19014 5864 19066
rect 5916 19014 5928 19066
rect 5980 19014 15118 19066
rect 15170 19014 15182 19066
rect 15234 19014 15246 19066
rect 15298 19014 15310 19066
rect 15362 19014 15374 19066
rect 15426 19014 24563 19066
rect 24615 19014 24627 19066
rect 24679 19014 24691 19066
rect 24743 19014 24755 19066
rect 24807 19014 24819 19066
rect 24871 19014 29440 19066
rect 1104 18992 29440 19014
rect 7469 18955 7527 18961
rect 7469 18952 7481 18955
rect 5644 18924 7481 18952
rect 2300 18819 2358 18825
rect 2300 18785 2312 18819
rect 2346 18816 2358 18819
rect 2406 18816 2412 18828
rect 2346 18788 2412 18816
rect 2346 18785 2358 18788
rect 2300 18779 2358 18785
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 2590 18816 2596 18828
rect 2551 18788 2596 18816
rect 2590 18776 2596 18788
rect 2648 18776 2654 18828
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18748 2099 18751
rect 2498 18748 2504 18760
rect 2087 18720 2504 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 2498 18708 2504 18720
rect 2556 18708 2562 18760
rect 4798 18748 4804 18760
rect 2746 18720 4804 18748
rect 1854 18680 1860 18692
rect 1815 18652 1860 18680
rect 1854 18640 1860 18652
rect 1912 18640 1918 18692
rect 2746 18680 2774 18720
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 5644 18757 5672 18924
rect 7469 18921 7481 18924
rect 7515 18921 7527 18955
rect 13078 18952 13084 18964
rect 7469 18915 7527 18921
rect 7760 18924 8524 18952
rect 7760 18828 7788 18924
rect 7742 18816 7748 18828
rect 7655 18788 7748 18816
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18816 7895 18819
rect 8202 18816 8208 18828
rect 7883 18788 8208 18816
rect 7883 18785 7895 18788
rect 7837 18779 7895 18785
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 5077 18751 5135 18757
rect 5077 18717 5089 18751
rect 5123 18748 5135 18751
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 5123 18720 5365 18748
rect 5123 18717 5135 18720
rect 5077 18711 5135 18717
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 5629 18751 5687 18757
rect 5629 18717 5641 18751
rect 5675 18717 5687 18751
rect 5629 18711 5687 18717
rect 5813 18751 5871 18757
rect 5813 18717 5825 18751
rect 5859 18748 5871 18751
rect 7466 18748 7472 18760
rect 5859 18720 7472 18748
rect 5859 18717 5871 18720
rect 5813 18711 5871 18717
rect 7466 18708 7472 18720
rect 7524 18708 7530 18760
rect 7653 18751 7711 18757
rect 7653 18717 7665 18751
rect 7699 18717 7711 18751
rect 7653 18711 7711 18717
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18748 7987 18751
rect 8018 18748 8024 18760
rect 7975 18720 8024 18748
rect 7975 18717 7987 18720
rect 7929 18711 7987 18717
rect 5534 18680 5540 18692
rect 2424 18652 2774 18680
rect 3804 18652 5540 18680
rect 2424 18621 2452 18652
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18581 2467 18615
rect 2409 18575 2467 18581
rect 2501 18615 2559 18621
rect 2501 18581 2513 18615
rect 2547 18612 2559 18615
rect 2682 18612 2688 18624
rect 2547 18584 2688 18612
rect 2547 18581 2559 18584
rect 2501 18575 2559 18581
rect 2682 18572 2688 18584
rect 2740 18612 2746 18624
rect 3804 18621 3832 18652
rect 5534 18640 5540 18652
rect 5592 18640 5598 18692
rect 5721 18683 5779 18689
rect 5721 18649 5733 18683
rect 5767 18680 5779 18683
rect 6058 18683 6116 18689
rect 6058 18680 6070 18683
rect 5767 18652 6070 18680
rect 5767 18649 5779 18652
rect 5721 18643 5779 18649
rect 6058 18649 6070 18652
rect 6104 18649 6116 18683
rect 6058 18643 6116 18649
rect 7558 18640 7564 18692
rect 7616 18680 7622 18692
rect 7668 18680 7696 18711
rect 8018 18708 8024 18720
rect 8076 18708 8082 18760
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18748 8171 18751
rect 8297 18751 8355 18757
rect 8297 18748 8309 18751
rect 8159 18720 8309 18748
rect 8159 18717 8171 18720
rect 8113 18711 8171 18717
rect 8297 18717 8309 18720
rect 8343 18717 8355 18751
rect 8297 18711 8355 18717
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8496 18748 8524 18924
rect 11716 18924 13084 18952
rect 8662 18844 8668 18896
rect 8720 18884 8726 18896
rect 10870 18884 10876 18896
rect 8720 18856 10876 18884
rect 8720 18844 8726 18856
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 11422 18884 11428 18896
rect 11256 18856 11428 18884
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 9861 18819 9919 18825
rect 9861 18816 9873 18819
rect 8628 18788 9873 18816
rect 8628 18776 8634 18788
rect 9861 18785 9873 18788
rect 9907 18785 9919 18819
rect 9861 18779 9919 18785
rect 9950 18776 9956 18828
rect 10008 18816 10014 18828
rect 11256 18816 11284 18856
rect 11422 18844 11428 18856
rect 11480 18844 11486 18896
rect 10008 18788 11284 18816
rect 11333 18819 11391 18825
rect 10008 18776 10014 18788
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 8496 18720 9597 18748
rect 8389 18711 8447 18717
rect 9585 18717 9597 18720
rect 9631 18748 9643 18751
rect 9769 18751 9827 18757
rect 9631 18720 9720 18748
rect 9631 18717 9643 18720
rect 9585 18711 9643 18717
rect 8404 18680 8432 18711
rect 8662 18680 8668 18692
rect 7616 18652 8668 18680
rect 7616 18640 7622 18652
rect 8662 18640 8668 18652
rect 8720 18640 8726 18692
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 2740 18584 3801 18612
rect 2740 18572 2746 18584
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 5077 18615 5135 18621
rect 5077 18581 5089 18615
rect 5123 18612 5135 18615
rect 5261 18615 5319 18621
rect 5261 18612 5273 18615
rect 5123 18584 5273 18612
rect 5123 18581 5135 18584
rect 5077 18575 5135 18581
rect 5261 18581 5273 18584
rect 5307 18612 5319 18615
rect 6270 18612 6276 18624
rect 5307 18584 6276 18612
rect 5307 18581 5319 18584
rect 5261 18575 5319 18581
rect 6270 18572 6276 18584
rect 6328 18572 6334 18624
rect 7193 18615 7251 18621
rect 7193 18581 7205 18615
rect 7239 18612 7251 18615
rect 7576 18612 7604 18640
rect 7239 18584 7604 18612
rect 9692 18612 9720 18720
rect 9769 18717 9781 18751
rect 9815 18717 9827 18751
rect 10042 18748 10048 18760
rect 10003 18720 10048 18748
rect 9769 18711 9827 18717
rect 9784 18680 9812 18711
rect 10042 18708 10048 18720
rect 10100 18708 10106 18760
rect 10244 18757 10272 18788
rect 11333 18785 11345 18819
rect 11379 18816 11391 18819
rect 11609 18819 11667 18825
rect 11609 18816 11621 18819
rect 11379 18788 11621 18816
rect 11379 18785 11391 18788
rect 11333 18779 11391 18785
rect 11609 18785 11621 18788
rect 11655 18785 11667 18819
rect 11609 18779 11667 18785
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18717 10287 18751
rect 10229 18711 10287 18717
rect 10318 18708 10324 18760
rect 10376 18748 10382 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 10376 18720 10425 18748
rect 10376 18708 10382 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 11149 18751 11207 18757
rect 11149 18717 11161 18751
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18748 11483 18751
rect 11716 18748 11744 18924
rect 13078 18912 13084 18924
rect 13136 18952 13142 18964
rect 13909 18955 13967 18961
rect 13909 18952 13921 18955
rect 13136 18924 13921 18952
rect 13136 18912 13142 18924
rect 13909 18921 13921 18924
rect 13955 18921 13967 18955
rect 13909 18915 13967 18921
rect 19061 18955 19119 18961
rect 19061 18921 19073 18955
rect 19107 18952 19119 18955
rect 19242 18952 19248 18964
rect 19107 18924 19248 18952
rect 19107 18921 19119 18924
rect 19061 18915 19119 18921
rect 11977 18887 12035 18893
rect 11977 18853 11989 18887
rect 12023 18884 12035 18887
rect 12066 18884 12072 18896
rect 12023 18856 12072 18884
rect 12023 18853 12035 18856
rect 11977 18847 12035 18853
rect 12066 18844 12072 18856
rect 12124 18844 12130 18896
rect 12526 18844 12532 18896
rect 12584 18844 12590 18896
rect 12894 18884 12900 18896
rect 12855 18856 12900 18884
rect 12894 18844 12900 18856
rect 12952 18844 12958 18896
rect 11793 18819 11851 18825
rect 11793 18785 11805 18819
rect 11839 18816 11851 18819
rect 12434 18816 12440 18828
rect 11839 18788 12440 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 12434 18776 12440 18788
rect 12492 18776 12498 18828
rect 12544 18816 12572 18844
rect 13538 18816 13544 18828
rect 12544 18788 12848 18816
rect 11471 18720 11744 18748
rect 12069 18751 12127 18757
rect 11471 18717 11483 18720
rect 11425 18711 11483 18717
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 12161 18751 12219 18757
rect 12161 18748 12173 18751
rect 12115 18720 12173 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 12161 18717 12173 18720
rect 12207 18717 12219 18751
rect 12526 18748 12532 18760
rect 12487 18720 12532 18748
rect 12161 18711 12219 18717
rect 10965 18683 11023 18689
rect 10965 18680 10977 18683
rect 9784 18652 10977 18680
rect 10965 18649 10977 18652
rect 11011 18649 11023 18683
rect 11164 18680 11192 18711
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 12710 18748 12716 18760
rect 12671 18720 12716 18748
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 11698 18680 11704 18692
rect 11164 18652 11704 18680
rect 10965 18643 11023 18649
rect 11698 18640 11704 18652
rect 11756 18640 11762 18692
rect 12437 18683 12495 18689
rect 12437 18649 12449 18683
rect 12483 18680 12495 18683
rect 12820 18680 12848 18788
rect 13372 18788 13544 18816
rect 12986 18748 12992 18760
rect 12947 18720 12992 18748
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 13372 18757 13400 18788
rect 13538 18776 13544 18788
rect 13596 18776 13602 18828
rect 13924 18816 13952 18915
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 19518 18912 19524 18964
rect 19576 18952 19582 18964
rect 19981 18955 20039 18961
rect 19981 18952 19993 18955
rect 19576 18924 19993 18952
rect 19576 18912 19582 18924
rect 19981 18921 19993 18924
rect 20027 18921 20039 18955
rect 19981 18915 20039 18921
rect 20070 18912 20076 18964
rect 20128 18952 20134 18964
rect 20438 18952 20444 18964
rect 20128 18924 20444 18952
rect 20128 18912 20134 18924
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 22281 18955 22339 18961
rect 22281 18952 22293 18955
rect 20640 18924 22293 18952
rect 18782 18844 18788 18896
rect 18840 18884 18846 18896
rect 20640 18884 20668 18924
rect 22281 18921 22293 18924
rect 22327 18921 22339 18955
rect 22554 18952 22560 18964
rect 22515 18924 22560 18952
rect 22281 18915 22339 18921
rect 22554 18912 22560 18924
rect 22612 18912 22618 18964
rect 22922 18912 22928 18964
rect 22980 18952 22986 18964
rect 22980 18924 23612 18952
rect 22980 18912 22986 18924
rect 18840 18856 20668 18884
rect 18840 18844 18846 18856
rect 14461 18819 14519 18825
rect 13924 18788 14320 18816
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13372 18680 13400 18711
rect 13446 18708 13452 18760
rect 13504 18748 13510 18760
rect 13504 18720 13549 18748
rect 13504 18708 13510 18720
rect 13630 18708 13636 18760
rect 13688 18748 13694 18760
rect 13725 18751 13783 18757
rect 13725 18748 13737 18751
rect 13688 18720 13737 18748
rect 13688 18708 13694 18720
rect 13725 18717 13737 18720
rect 13771 18717 13783 18751
rect 14182 18748 14188 18760
rect 14143 18720 14188 18748
rect 13725 18711 13783 18717
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 14292 18748 14320 18788
rect 14461 18785 14473 18819
rect 14507 18816 14519 18819
rect 14642 18816 14648 18828
rect 14507 18788 14648 18816
rect 14507 18785 14519 18788
rect 14461 18779 14519 18785
rect 14642 18776 14648 18788
rect 14700 18776 14706 18828
rect 14921 18819 14979 18825
rect 14921 18785 14933 18819
rect 14967 18816 14979 18819
rect 16025 18819 16083 18825
rect 14967 18788 15884 18816
rect 14967 18785 14979 18788
rect 14921 18779 14979 18785
rect 14366 18757 14372 18760
rect 14350 18751 14372 18757
rect 14350 18748 14362 18751
rect 14279 18720 14362 18748
rect 14350 18717 14362 18720
rect 14350 18711 14372 18717
rect 14366 18708 14372 18711
rect 14424 18708 14430 18760
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 14737 18751 14795 18757
rect 14608 18720 14653 18748
rect 14608 18708 14614 18720
rect 14737 18717 14749 18751
rect 14783 18717 14795 18751
rect 14737 18711 14795 18717
rect 15197 18751 15255 18757
rect 15197 18717 15209 18751
rect 15243 18717 15255 18751
rect 15470 18748 15476 18760
rect 15431 18720 15476 18748
rect 15197 18711 15255 18717
rect 14752 18680 14780 18711
rect 14826 18680 14832 18692
rect 12483 18652 13400 18680
rect 14660 18652 14832 18680
rect 12483 18649 12495 18652
rect 12437 18643 12495 18649
rect 10505 18615 10563 18621
rect 10505 18612 10517 18615
rect 9692 18584 10517 18612
rect 7239 18581 7251 18584
rect 7193 18575 7251 18581
rect 10505 18581 10517 18584
rect 10551 18581 10563 18615
rect 10505 18575 10563 18581
rect 10870 18572 10876 18624
rect 10928 18612 10934 18624
rect 12161 18615 12219 18621
rect 12161 18612 12173 18615
rect 10928 18584 12173 18612
rect 10928 18572 10934 18584
rect 12161 18581 12173 18584
rect 12207 18581 12219 18615
rect 12161 18575 12219 18581
rect 12710 18572 12716 18624
rect 12768 18612 12774 18624
rect 13078 18612 13084 18624
rect 12768 18584 13084 18612
rect 12768 18572 12774 18584
rect 13078 18572 13084 18584
rect 13136 18612 13142 18624
rect 14660 18612 14688 18652
rect 14826 18640 14832 18652
rect 14884 18680 14890 18692
rect 15105 18683 15163 18689
rect 15105 18680 15117 18683
rect 14884 18652 15117 18680
rect 14884 18640 14890 18652
rect 15105 18649 15117 18652
rect 15151 18649 15163 18683
rect 15212 18680 15240 18711
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 15654 18748 15660 18760
rect 15615 18720 15660 18748
rect 15654 18708 15660 18720
rect 15712 18708 15718 18760
rect 15856 18757 15884 18788
rect 16025 18785 16037 18819
rect 16071 18785 16083 18819
rect 16482 18816 16488 18828
rect 16443 18788 16488 18816
rect 16025 18779 16083 18785
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18748 15899 18751
rect 15930 18748 15936 18760
rect 15887 18720 15936 18748
rect 15887 18717 15899 18720
rect 15841 18711 15899 18717
rect 15930 18708 15936 18720
rect 15988 18708 15994 18760
rect 16040 18680 16068 18779
rect 16482 18776 16488 18788
rect 16540 18816 16546 18828
rect 18230 18816 18236 18828
rect 16540 18788 18236 18816
rect 16540 18776 16546 18788
rect 18230 18776 18236 18788
rect 18288 18816 18294 18828
rect 18509 18819 18567 18825
rect 18509 18816 18521 18819
rect 18288 18788 18521 18816
rect 18288 18776 18294 18788
rect 18509 18785 18521 18788
rect 18555 18785 18567 18819
rect 18509 18779 18567 18785
rect 18966 18776 18972 18828
rect 19024 18816 19030 18828
rect 19337 18819 19395 18825
rect 19337 18816 19349 18819
rect 19024 18788 19349 18816
rect 19024 18776 19030 18788
rect 19337 18785 19349 18788
rect 19383 18785 19395 18819
rect 19337 18779 19395 18785
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 20349 18819 20407 18825
rect 20349 18816 20361 18819
rect 19760 18788 20361 18816
rect 19760 18776 19766 18788
rect 20349 18785 20361 18788
rect 20395 18785 20407 18819
rect 20349 18779 20407 18785
rect 20438 18776 20444 18828
rect 20496 18816 20502 18828
rect 20496 18788 20541 18816
rect 20496 18776 20502 18788
rect 16114 18708 16120 18760
rect 16172 18748 16178 18760
rect 16298 18748 16304 18760
rect 16172 18720 16217 18748
rect 16259 18720 16304 18748
rect 16172 18708 16178 18720
rect 16298 18708 16304 18720
rect 16356 18708 16362 18760
rect 18782 18708 18788 18760
rect 18840 18748 18846 18760
rect 18877 18751 18935 18757
rect 18877 18748 18889 18751
rect 18840 18720 18889 18748
rect 18840 18708 18846 18720
rect 18877 18717 18889 18720
rect 18923 18717 18935 18751
rect 18877 18711 18935 18717
rect 19518 18708 19524 18760
rect 19576 18748 19582 18760
rect 20640 18757 20668 18856
rect 20714 18776 20720 18828
rect 20772 18816 20778 18828
rect 20901 18819 20959 18825
rect 20901 18816 20913 18819
rect 20772 18788 20913 18816
rect 20772 18776 20778 18788
rect 20901 18785 20913 18788
rect 20947 18785 20959 18819
rect 22572 18816 22600 18912
rect 23385 18887 23443 18893
rect 23385 18853 23397 18887
rect 23431 18884 23443 18887
rect 23474 18884 23480 18896
rect 23431 18856 23480 18884
rect 23431 18853 23443 18856
rect 23385 18847 23443 18853
rect 23474 18844 23480 18856
rect 23532 18844 23538 18896
rect 23584 18884 23612 18924
rect 23750 18912 23756 18964
rect 23808 18952 23814 18964
rect 23934 18952 23940 18964
rect 23808 18924 23940 18952
rect 23808 18912 23814 18924
rect 23934 18912 23940 18924
rect 23992 18912 23998 18964
rect 25961 18955 26019 18961
rect 25961 18921 25973 18955
rect 26007 18952 26019 18955
rect 26050 18952 26056 18964
rect 26007 18924 26056 18952
rect 26007 18921 26019 18924
rect 25961 18915 26019 18921
rect 26050 18912 26056 18924
rect 26108 18912 26114 18964
rect 24029 18887 24087 18893
rect 24029 18884 24041 18887
rect 23584 18856 24041 18884
rect 24029 18853 24041 18856
rect 24075 18853 24087 18887
rect 24029 18847 24087 18853
rect 24857 18887 24915 18893
rect 24857 18853 24869 18887
rect 24903 18853 24915 18887
rect 24857 18847 24915 18853
rect 25501 18887 25559 18893
rect 25501 18853 25513 18887
rect 25547 18853 25559 18887
rect 25501 18847 25559 18853
rect 23750 18816 23756 18828
rect 22572 18788 22876 18816
rect 20901 18779 20959 18785
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19576 18720 19625 18748
rect 19576 18708 19582 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 20073 18751 20131 18757
rect 20073 18717 20085 18751
rect 20119 18717 20131 18751
rect 20073 18711 20131 18717
rect 20256 18751 20314 18757
rect 20256 18717 20268 18751
rect 20302 18748 20314 18751
rect 20625 18751 20683 18757
rect 20302 18720 20576 18748
rect 20302 18717 20314 18720
rect 20256 18711 20314 18717
rect 16761 18683 16819 18689
rect 16761 18680 16773 18683
rect 15212 18652 15700 18680
rect 16040 18652 16773 18680
rect 15105 18643 15163 18649
rect 15286 18612 15292 18624
rect 13136 18584 14688 18612
rect 15247 18584 15292 18612
rect 13136 18572 13142 18584
rect 15286 18572 15292 18584
rect 15344 18612 15350 18624
rect 15562 18612 15568 18624
rect 15344 18584 15568 18612
rect 15344 18572 15350 18584
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 15672 18612 15700 18652
rect 16761 18649 16773 18652
rect 16807 18649 16819 18683
rect 16761 18643 16819 18649
rect 17310 18640 17316 18692
rect 17368 18640 17374 18692
rect 18693 18683 18751 18689
rect 18693 18649 18705 18683
rect 18739 18680 18751 18683
rect 19426 18680 19432 18692
rect 18739 18652 19432 18680
rect 18739 18649 18751 18652
rect 18693 18643 18751 18649
rect 19426 18640 19432 18652
rect 19484 18640 19490 18692
rect 19886 18680 19892 18692
rect 19536 18652 19892 18680
rect 16206 18612 16212 18624
rect 15672 18584 16212 18612
rect 16206 18572 16212 18584
rect 16264 18572 16270 18624
rect 18233 18615 18291 18621
rect 18233 18581 18245 18615
rect 18279 18612 18291 18615
rect 18414 18612 18420 18624
rect 18279 18584 18420 18612
rect 18279 18581 18291 18584
rect 18233 18575 18291 18581
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 19536 18621 19564 18652
rect 19886 18640 19892 18652
rect 19944 18640 19950 18692
rect 20088 18680 20116 18711
rect 20548 18680 20576 18720
rect 20625 18717 20637 18751
rect 20671 18717 20683 18751
rect 22738 18748 22744 18760
rect 22699 18720 22744 18748
rect 20625 18711 20683 18717
rect 22738 18708 22744 18720
rect 22796 18708 22802 18760
rect 22848 18757 22876 18788
rect 23492 18788 23756 18816
rect 22833 18751 22891 18757
rect 22833 18717 22845 18751
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 22922 18708 22928 18760
rect 22980 18748 22986 18760
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 22980 18720 23029 18748
rect 22980 18708 22986 18720
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 23253 18751 23311 18757
rect 23253 18717 23265 18751
rect 23299 18748 23311 18751
rect 23492 18748 23520 18788
rect 23750 18776 23756 18788
rect 23808 18776 23814 18828
rect 23299 18720 23520 18748
rect 23569 18751 23627 18757
rect 23299 18717 23311 18720
rect 23253 18711 23311 18717
rect 23569 18717 23581 18751
rect 23615 18748 23627 18751
rect 23615 18720 23980 18748
rect 23615 18717 23627 18720
rect 23569 18711 23627 18717
rect 20714 18680 20720 18692
rect 20088 18652 20300 18680
rect 20548 18652 20720 18680
rect 20272 18624 20300 18652
rect 20714 18640 20720 18652
rect 20772 18640 20778 18692
rect 20809 18683 20867 18689
rect 20809 18649 20821 18683
rect 20855 18680 20867 18683
rect 21146 18683 21204 18689
rect 21146 18680 21158 18683
rect 20855 18652 21158 18680
rect 20855 18649 20867 18652
rect 20809 18643 20867 18649
rect 21146 18649 21158 18652
rect 21192 18649 21204 18683
rect 21146 18643 21204 18649
rect 22370 18640 22376 18692
rect 22428 18680 22434 18692
rect 22940 18680 22968 18708
rect 22428 18652 22968 18680
rect 22428 18640 22434 18652
rect 23106 18640 23112 18692
rect 23164 18680 23170 18692
rect 23845 18683 23903 18689
rect 23845 18680 23857 18683
rect 23164 18652 23857 18680
rect 23164 18640 23170 18652
rect 23845 18649 23857 18652
rect 23891 18649 23903 18683
rect 23845 18643 23903 18649
rect 19521 18615 19579 18621
rect 19521 18581 19533 18615
rect 19567 18581 19579 18615
rect 19521 18575 19579 18581
rect 20254 18572 20260 18624
rect 20312 18572 20318 18624
rect 22646 18572 22652 18624
rect 22704 18612 22710 18624
rect 23952 18612 23980 18720
rect 24486 18708 24492 18760
rect 24544 18748 24550 18760
rect 24673 18751 24731 18757
rect 24673 18748 24685 18751
rect 24544 18720 24685 18748
rect 24544 18708 24550 18720
rect 24673 18717 24685 18720
rect 24719 18717 24731 18751
rect 24872 18748 24900 18847
rect 25133 18751 25191 18757
rect 25133 18748 25145 18751
rect 24872 18720 25145 18748
rect 24673 18711 24731 18717
rect 25133 18717 25145 18720
rect 25179 18717 25191 18751
rect 25133 18711 25191 18717
rect 25317 18751 25375 18757
rect 25317 18717 25329 18751
rect 25363 18717 25375 18751
rect 25516 18748 25544 18847
rect 25777 18751 25835 18757
rect 25777 18748 25789 18751
rect 25516 18720 25789 18748
rect 25317 18711 25375 18717
rect 25777 18717 25789 18720
rect 25823 18717 25835 18751
rect 25777 18711 25835 18717
rect 24688 18680 24716 18711
rect 25332 18680 25360 18711
rect 24688 18652 25360 18680
rect 24946 18612 24952 18624
rect 22704 18584 23980 18612
rect 24907 18584 24952 18612
rect 22704 18572 22710 18584
rect 24946 18572 24952 18584
rect 25004 18572 25010 18624
rect 1104 18522 29440 18544
rect 1104 18470 10395 18522
rect 10447 18470 10459 18522
rect 10511 18470 10523 18522
rect 10575 18470 10587 18522
rect 10639 18470 10651 18522
rect 10703 18470 19840 18522
rect 19892 18470 19904 18522
rect 19956 18470 19968 18522
rect 20020 18470 20032 18522
rect 20084 18470 20096 18522
rect 20148 18470 29440 18522
rect 1104 18448 29440 18470
rect 1854 18408 1860 18420
rect 1815 18380 1860 18408
rect 1854 18368 1860 18380
rect 1912 18368 1918 18420
rect 1949 18411 2007 18417
rect 1949 18377 1961 18411
rect 1995 18408 2007 18411
rect 2222 18408 2228 18420
rect 1995 18380 2228 18408
rect 1995 18377 2007 18380
rect 1949 18371 2007 18377
rect 2222 18368 2228 18380
rect 2280 18408 2286 18420
rect 2590 18408 2596 18420
rect 2280 18380 2596 18408
rect 2280 18368 2286 18380
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 2682 18368 2688 18420
rect 2740 18408 2746 18420
rect 3605 18411 3663 18417
rect 2740 18380 3096 18408
rect 2740 18368 2746 18380
rect 3068 18349 3096 18380
rect 3605 18377 3617 18411
rect 3651 18377 3663 18411
rect 3605 18371 3663 18377
rect 3973 18411 4031 18417
rect 3973 18377 3985 18411
rect 4019 18408 4031 18411
rect 4430 18408 4436 18420
rect 4019 18380 4436 18408
rect 4019 18377 4031 18380
rect 3973 18371 4031 18377
rect 2409 18343 2467 18349
rect 2409 18309 2421 18343
rect 2455 18340 2467 18343
rect 3053 18343 3111 18349
rect 2455 18312 2912 18340
rect 2455 18309 2467 18312
rect 2409 18303 2467 18309
rect 2884 18281 2912 18312
rect 3053 18309 3065 18343
rect 3099 18309 3111 18343
rect 3053 18303 3111 18309
rect 3145 18343 3203 18349
rect 3145 18309 3157 18343
rect 3191 18340 3203 18343
rect 3620 18340 3648 18371
rect 4430 18368 4436 18380
rect 4488 18368 4494 18420
rect 7466 18408 7472 18420
rect 7427 18380 7472 18408
rect 7466 18368 7472 18380
rect 7524 18408 7530 18420
rect 8202 18408 8208 18420
rect 7524 18380 8208 18408
rect 7524 18368 7530 18380
rect 3191 18312 3648 18340
rect 3988 18312 4384 18340
rect 3191 18309 3203 18312
rect 3145 18303 3203 18309
rect 2593 18275 2651 18281
rect 2593 18241 2605 18275
rect 2639 18241 2651 18275
rect 2593 18235 2651 18241
rect 2777 18275 2835 18281
rect 2777 18241 2789 18275
rect 2823 18241 2835 18275
rect 2777 18235 2835 18241
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18241 2927 18275
rect 2869 18235 2927 18241
rect 3289 18275 3347 18281
rect 3289 18241 3301 18275
rect 3335 18272 3347 18275
rect 3988 18272 4016 18312
rect 4356 18284 4384 18312
rect 3335 18244 4016 18272
rect 3335 18241 3347 18244
rect 3289 18235 3347 18241
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18204 2191 18207
rect 2498 18204 2504 18216
rect 2179 18176 2504 18204
rect 2179 18173 2191 18176
rect 2133 18167 2191 18173
rect 2498 18164 2504 18176
rect 2556 18164 2562 18216
rect 2608 18136 2636 18235
rect 2792 18204 2820 18235
rect 4338 18232 4344 18284
rect 4396 18232 4402 18284
rect 4614 18272 4620 18284
rect 4575 18244 4620 18272
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 6362 18272 6368 18284
rect 6043 18244 6368 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 7558 18272 7564 18284
rect 7519 18244 7564 18272
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 7742 18272 7748 18284
rect 7703 18244 7748 18272
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 8036 18281 8064 18380
rect 8202 18368 8208 18380
rect 8260 18408 8266 18420
rect 9214 18408 9220 18420
rect 8260 18380 9220 18408
rect 8260 18368 8266 18380
rect 9214 18368 9220 18380
rect 9272 18408 9278 18420
rect 9953 18411 10011 18417
rect 9953 18408 9965 18411
rect 9272 18380 9965 18408
rect 9272 18368 9278 18380
rect 9953 18377 9965 18380
rect 9999 18377 10011 18411
rect 9953 18371 10011 18377
rect 12342 18368 12348 18420
rect 12400 18408 12406 18420
rect 12989 18411 13047 18417
rect 12400 18380 12848 18408
rect 12400 18368 12406 18380
rect 8297 18343 8355 18349
rect 8297 18309 8309 18343
rect 8343 18340 8355 18343
rect 8570 18340 8576 18352
rect 8343 18312 8576 18340
rect 8343 18309 8355 18312
rect 8297 18303 8355 18309
rect 8570 18300 8576 18312
rect 8628 18300 8634 18352
rect 8754 18300 8760 18352
rect 8812 18300 8818 18352
rect 11149 18343 11207 18349
rect 11149 18309 11161 18343
rect 11195 18340 11207 18343
rect 11238 18340 11244 18352
rect 11195 18312 11244 18340
rect 11195 18309 11207 18312
rect 11149 18303 11207 18309
rect 11238 18300 11244 18312
rect 11296 18300 11302 18352
rect 11698 18300 11704 18352
rect 11756 18340 11762 18352
rect 11756 18312 12572 18340
rect 11756 18300 11762 18312
rect 8021 18275 8079 18281
rect 8021 18241 8033 18275
rect 8067 18241 8079 18275
rect 8021 18235 8079 18241
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18241 11391 18275
rect 11333 18235 11391 18241
rect 4062 18204 4068 18216
rect 2792 18176 4068 18204
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18173 4215 18207
rect 4157 18167 4215 18173
rect 9769 18207 9827 18213
rect 9769 18173 9781 18207
rect 9815 18204 9827 18207
rect 10318 18204 10324 18216
rect 9815 18176 10324 18204
rect 9815 18173 9827 18176
rect 9769 18167 9827 18173
rect 3234 18136 3240 18148
rect 2608 18108 3240 18136
rect 3234 18096 3240 18108
rect 3292 18096 3298 18148
rect 3510 18136 3516 18148
rect 3344 18108 3516 18136
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 2498 18028 2504 18080
rect 2556 18068 2562 18080
rect 3344 18068 3372 18108
rect 3510 18096 3516 18108
rect 3568 18096 3574 18148
rect 4172 18136 4200 18167
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 11238 18164 11244 18216
rect 11296 18204 11302 18216
rect 11348 18204 11376 18235
rect 11422 18232 11428 18284
rect 11480 18272 11486 18284
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 11480 18244 11529 18272
rect 11480 18232 11486 18244
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 12342 18272 12348 18284
rect 12303 18244 12348 18272
rect 11517 18235 11575 18241
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 12544 18272 12572 18312
rect 12618 18300 12624 18352
rect 12676 18340 12682 18352
rect 12820 18340 12848 18380
rect 12989 18377 13001 18411
rect 13035 18408 13047 18411
rect 14182 18408 14188 18420
rect 13035 18380 14188 18408
rect 13035 18377 13047 18380
rect 12989 18371 13047 18377
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 16298 18408 16304 18420
rect 15396 18380 16304 18408
rect 15396 18349 15424 18380
rect 16298 18368 16304 18380
rect 16356 18368 16362 18420
rect 17037 18411 17095 18417
rect 17037 18377 17049 18411
rect 17083 18408 17095 18411
rect 17083 18380 22094 18408
rect 17083 18377 17095 18380
rect 17037 18371 17095 18377
rect 13817 18343 13875 18349
rect 13817 18340 13829 18343
rect 12676 18312 12756 18340
rect 12820 18312 13829 18340
rect 12676 18300 12682 18312
rect 12728 18281 12756 18312
rect 13817 18309 13829 18312
rect 13863 18340 13875 18343
rect 15381 18343 15439 18349
rect 13863 18312 14872 18340
rect 13863 18309 13875 18312
rect 13817 18303 13875 18309
rect 12713 18275 12771 18281
rect 12544 18244 12664 18272
rect 11296 18176 11560 18204
rect 11296 18164 11302 18176
rect 4433 18139 4491 18145
rect 4433 18136 4445 18139
rect 4172 18108 4445 18136
rect 4433 18105 4445 18108
rect 4479 18136 4491 18139
rect 4522 18136 4528 18148
rect 4479 18108 4528 18136
rect 4479 18105 4491 18108
rect 4433 18099 4491 18105
rect 4522 18096 4528 18108
rect 4580 18096 4586 18148
rect 7834 18136 7840 18148
rect 7795 18108 7840 18136
rect 7834 18096 7840 18108
rect 7892 18096 7898 18148
rect 10042 18096 10048 18148
rect 10100 18136 10106 18148
rect 11532 18136 11560 18176
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 12636 18213 12664 18244
rect 12713 18241 12725 18275
rect 12759 18241 12771 18275
rect 12713 18235 12771 18241
rect 13170 18232 13176 18284
rect 13228 18272 13234 18284
rect 13725 18275 13783 18281
rect 13725 18272 13737 18275
rect 13228 18244 13737 18272
rect 13228 18232 13234 18244
rect 13725 18241 13737 18244
rect 13771 18241 13783 18275
rect 13998 18272 14004 18284
rect 13959 18244 14004 18272
rect 13725 18235 13783 18241
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 14277 18275 14335 18281
rect 14277 18241 14289 18275
rect 14323 18272 14335 18275
rect 14366 18272 14372 18284
rect 14323 18244 14372 18272
rect 14323 18241 14335 18244
rect 14277 18235 14335 18241
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 14737 18275 14795 18281
rect 14737 18241 14749 18275
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 12529 18207 12587 18213
rect 12529 18204 12541 18207
rect 12124 18176 12541 18204
rect 12124 18164 12130 18176
rect 12529 18173 12541 18176
rect 12575 18173 12587 18207
rect 12529 18167 12587 18173
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18173 12679 18207
rect 12621 18167 12679 18173
rect 12805 18207 12863 18213
rect 12805 18173 12817 18207
rect 12851 18204 12863 18207
rect 13354 18204 13360 18216
rect 12851 18176 13360 18204
rect 12851 18173 12863 18176
rect 12805 18167 12863 18173
rect 12636 18136 12664 18167
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 14016 18204 14044 18232
rect 14752 18204 14780 18235
rect 14016 18176 14780 18204
rect 14844 18204 14872 18312
rect 15381 18309 15393 18343
rect 15427 18309 15439 18343
rect 15381 18303 15439 18309
rect 15470 18300 15476 18352
rect 15528 18340 15534 18352
rect 15749 18343 15807 18349
rect 15749 18340 15761 18343
rect 15528 18312 15761 18340
rect 15528 18300 15534 18312
rect 15749 18309 15761 18312
rect 15795 18340 15807 18343
rect 15795 18312 16712 18340
rect 15795 18309 15807 18312
rect 15749 18303 15807 18309
rect 15013 18275 15071 18281
rect 15013 18241 15025 18275
rect 15059 18272 15071 18275
rect 15286 18272 15292 18284
rect 15059 18244 15292 18272
rect 15059 18241 15071 18244
rect 15013 18235 15071 18241
rect 15286 18232 15292 18244
rect 15344 18232 15350 18284
rect 16684 18281 16712 18312
rect 18414 18300 18420 18352
rect 18472 18340 18478 18352
rect 19426 18340 19432 18352
rect 18472 18312 19432 18340
rect 18472 18300 18478 18312
rect 19426 18300 19432 18312
rect 19484 18340 19490 18352
rect 22066 18340 22094 18380
rect 22922 18368 22928 18420
rect 22980 18408 22986 18420
rect 23106 18408 23112 18420
rect 22980 18380 23112 18408
rect 22980 18368 22986 18380
rect 23106 18368 23112 18380
rect 23164 18408 23170 18420
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 23164 18380 24869 18408
rect 23164 18368 23170 18380
rect 24857 18377 24869 18380
rect 24903 18377 24915 18411
rect 24857 18371 24915 18377
rect 23382 18340 23388 18352
rect 19484 18312 19932 18340
rect 22066 18312 22692 18340
rect 19484 18300 19490 18312
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 16669 18275 16727 18281
rect 16669 18241 16681 18275
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 18693 18275 18751 18281
rect 18693 18241 18705 18275
rect 18739 18272 18751 18275
rect 18782 18272 18788 18284
rect 18739 18244 18788 18272
rect 18739 18241 18751 18244
rect 18693 18235 18751 18241
rect 15580 18204 15608 18235
rect 18782 18232 18788 18244
rect 18840 18232 18846 18284
rect 19610 18232 19616 18284
rect 19668 18272 19674 18284
rect 19705 18275 19763 18281
rect 19705 18272 19717 18275
rect 19668 18244 19717 18272
rect 19668 18232 19674 18244
rect 19705 18241 19717 18244
rect 19751 18241 19763 18275
rect 19705 18235 19763 18241
rect 16758 18204 16764 18216
rect 14844 18176 15608 18204
rect 16719 18176 16764 18204
rect 16758 18164 16764 18176
rect 16816 18164 16822 18216
rect 19904 18213 19932 18312
rect 22664 18284 22692 18312
rect 23124 18312 23388 18340
rect 22646 18272 22652 18284
rect 22559 18244 22652 18272
rect 22646 18232 22652 18244
rect 22704 18232 22710 18284
rect 23124 18281 23152 18312
rect 23382 18300 23388 18312
rect 23440 18300 23446 18352
rect 24946 18340 24952 18352
rect 24610 18312 24952 18340
rect 24946 18300 24952 18312
rect 25004 18300 25010 18352
rect 23109 18275 23167 18281
rect 23109 18241 23121 18275
rect 23155 18241 23167 18275
rect 23109 18235 23167 18241
rect 19797 18207 19855 18213
rect 19797 18173 19809 18207
rect 19843 18173 19855 18207
rect 19797 18167 19855 18173
rect 19889 18207 19947 18213
rect 19889 18173 19901 18207
rect 19935 18173 19947 18207
rect 19889 18167 19947 18173
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18204 23443 18207
rect 23474 18204 23480 18216
rect 23431 18176 23480 18204
rect 23431 18173 23443 18176
rect 23385 18167 23443 18173
rect 13170 18136 13176 18148
rect 10100 18108 11468 18136
rect 11532 18108 12434 18136
rect 12636 18108 13176 18136
rect 10100 18096 10106 18108
rect 11440 18080 11468 18108
rect 2556 18040 3372 18068
rect 3421 18071 3479 18077
rect 2556 18028 2562 18040
rect 3421 18037 3433 18071
rect 3467 18068 3479 18071
rect 4154 18068 4160 18080
rect 3467 18040 4160 18068
rect 3467 18037 3479 18040
rect 3421 18031 3479 18037
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 5905 18071 5963 18077
rect 5905 18037 5917 18071
rect 5951 18068 5963 18071
rect 6086 18068 6092 18080
rect 5951 18040 6092 18068
rect 5951 18037 5963 18040
rect 5905 18031 5963 18037
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 11057 18071 11115 18077
rect 11057 18037 11069 18071
rect 11103 18068 11115 18071
rect 11330 18068 11336 18080
rect 11103 18040 11336 18068
rect 11103 18037 11115 18040
rect 11057 18031 11115 18037
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 11422 18028 11428 18080
rect 11480 18068 11486 18080
rect 11701 18071 11759 18077
rect 11701 18068 11713 18071
rect 11480 18040 11713 18068
rect 11480 18028 11486 18040
rect 11701 18037 11713 18040
rect 11747 18037 11759 18071
rect 12406 18068 12434 18108
rect 13170 18096 13176 18108
rect 13228 18096 13234 18148
rect 13814 18136 13820 18148
rect 13280 18108 13820 18136
rect 13280 18068 13308 18108
rect 13814 18096 13820 18108
rect 13872 18096 13878 18148
rect 14093 18139 14151 18145
rect 14093 18105 14105 18139
rect 14139 18136 14151 18139
rect 14642 18136 14648 18148
rect 14139 18108 14648 18136
rect 14139 18105 14151 18108
rect 14093 18099 14151 18105
rect 14642 18096 14648 18108
rect 14700 18096 14706 18148
rect 14826 18136 14832 18148
rect 14787 18108 14832 18136
rect 14826 18096 14832 18108
rect 14884 18096 14890 18148
rect 19334 18136 19340 18148
rect 19295 18108 19340 18136
rect 19334 18096 19340 18108
rect 19392 18096 19398 18148
rect 19702 18096 19708 18148
rect 19760 18136 19766 18148
rect 19812 18136 19840 18167
rect 23474 18164 23480 18176
rect 23532 18164 23538 18216
rect 19760 18108 19840 18136
rect 19760 18096 19766 18108
rect 12406 18040 13308 18068
rect 11701 18031 11759 18037
rect 13354 18028 13360 18080
rect 13412 18068 13418 18080
rect 13541 18071 13599 18077
rect 13541 18068 13553 18071
rect 13412 18040 13553 18068
rect 13412 18028 13418 18040
rect 13541 18037 13553 18040
rect 13587 18037 13599 18071
rect 13541 18031 13599 18037
rect 14918 18028 14924 18080
rect 14976 18068 14982 18080
rect 15197 18071 15255 18077
rect 15197 18068 15209 18071
rect 14976 18040 15209 18068
rect 14976 18028 14982 18040
rect 15197 18037 15209 18040
rect 15243 18037 15255 18071
rect 15197 18031 15255 18037
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 16669 18071 16727 18077
rect 16669 18068 16681 18071
rect 16632 18040 16681 18068
rect 16632 18028 16638 18040
rect 16669 18037 16681 18040
rect 16715 18037 16727 18071
rect 16669 18031 16727 18037
rect 18877 18071 18935 18077
rect 18877 18037 18889 18071
rect 18923 18068 18935 18071
rect 20254 18068 20260 18080
rect 18923 18040 20260 18068
rect 18923 18037 18935 18040
rect 18877 18031 18935 18037
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20901 18071 20959 18077
rect 20901 18068 20913 18071
rect 20772 18040 20913 18068
rect 20772 18028 20778 18040
rect 20901 18037 20913 18040
rect 20947 18037 20959 18071
rect 22738 18068 22744 18080
rect 22651 18040 22744 18068
rect 20901 18031 20959 18037
rect 22738 18028 22744 18040
rect 22796 18068 22802 18080
rect 23198 18068 23204 18080
rect 22796 18040 23204 18068
rect 22796 18028 22802 18040
rect 23198 18028 23204 18040
rect 23256 18028 23262 18080
rect 1104 17978 29440 18000
rect 1104 17926 5672 17978
rect 5724 17926 5736 17978
rect 5788 17926 5800 17978
rect 5852 17926 5864 17978
rect 5916 17926 5928 17978
rect 5980 17926 15118 17978
rect 15170 17926 15182 17978
rect 15234 17926 15246 17978
rect 15298 17926 15310 17978
rect 15362 17926 15374 17978
rect 15426 17926 24563 17978
rect 24615 17926 24627 17978
rect 24679 17926 24691 17978
rect 24743 17926 24755 17978
rect 24807 17926 24819 17978
rect 24871 17926 29440 17978
rect 1104 17904 29440 17926
rect 14 17824 20 17876
rect 72 17864 78 17876
rect 7190 17864 7196 17876
rect 72 17836 7196 17864
rect 72 17824 78 17836
rect 7190 17824 7196 17836
rect 7248 17824 7254 17876
rect 9214 17864 9220 17876
rect 9175 17836 9220 17864
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 11698 17864 11704 17876
rect 9324 17836 11704 17864
rect 6638 17796 6644 17808
rect 6599 17768 6644 17796
rect 6638 17756 6644 17768
rect 6696 17756 6702 17808
rect 7101 17799 7159 17805
rect 7101 17765 7113 17799
rect 7147 17796 7159 17799
rect 9324 17796 9352 17836
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 11974 17864 11980 17876
rect 11935 17836 11980 17864
rect 11974 17824 11980 17836
rect 12032 17824 12038 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 12802 17864 12808 17876
rect 12492 17836 12537 17864
rect 12636 17836 12808 17864
rect 12492 17824 12498 17836
rect 7147 17768 9352 17796
rect 10965 17799 11023 17805
rect 7147 17765 7159 17768
rect 7101 17759 7159 17765
rect 10965 17765 10977 17799
rect 11011 17796 11023 17799
rect 11054 17796 11060 17808
rect 11011 17768 11060 17796
rect 11011 17765 11023 17768
rect 10965 17759 11023 17765
rect 7116 17728 7144 17759
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 12161 17799 12219 17805
rect 12161 17765 12173 17799
rect 12207 17796 12219 17799
rect 12636 17796 12664 17836
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 13357 17867 13415 17873
rect 13357 17833 13369 17867
rect 13403 17864 13415 17867
rect 13446 17864 13452 17876
rect 13403 17836 13452 17864
rect 13403 17833 13415 17836
rect 13357 17827 13415 17833
rect 13446 17824 13452 17836
rect 13504 17864 13510 17876
rect 14826 17864 14832 17876
rect 13504 17836 14832 17864
rect 13504 17824 13510 17836
rect 14826 17824 14832 17836
rect 14884 17824 14890 17876
rect 15105 17867 15163 17873
rect 15105 17833 15117 17867
rect 15151 17864 15163 17867
rect 16298 17864 16304 17876
rect 15151 17836 16304 17864
rect 15151 17833 15163 17836
rect 15105 17827 15163 17833
rect 16298 17824 16304 17836
rect 16356 17824 16362 17876
rect 17586 17824 17592 17876
rect 17644 17864 17650 17876
rect 17865 17867 17923 17873
rect 17865 17864 17877 17867
rect 17644 17836 17877 17864
rect 17644 17824 17650 17836
rect 17865 17833 17877 17836
rect 17911 17833 17923 17867
rect 17865 17827 17923 17833
rect 14182 17796 14188 17808
rect 12207 17768 12664 17796
rect 14143 17768 14188 17796
rect 12207 17765 12219 17768
rect 12161 17759 12219 17765
rect 14182 17756 14188 17768
rect 14240 17796 14246 17808
rect 16669 17799 16727 17805
rect 16669 17796 16681 17799
rect 14240 17768 15516 17796
rect 14240 17756 14246 17768
rect 6748 17700 7144 17728
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17660 1455 17663
rect 3881 17663 3939 17669
rect 1443 17632 3096 17660
rect 1443 17629 1455 17632
rect 1397 17623 1455 17629
rect 1486 17552 1492 17604
rect 1544 17592 1550 17604
rect 1642 17595 1700 17601
rect 1642 17592 1654 17595
rect 1544 17564 1654 17592
rect 1544 17552 1550 17564
rect 1642 17561 1654 17564
rect 1688 17561 1700 17595
rect 1642 17555 1700 17561
rect 3068 17536 3096 17632
rect 3881 17629 3893 17663
rect 3927 17660 3939 17663
rect 4706 17660 4712 17672
rect 3927 17632 4712 17660
rect 3927 17629 3939 17632
rect 3881 17623 3939 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 6457 17663 6515 17669
rect 6457 17629 6469 17663
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 3786 17552 3792 17604
rect 3844 17592 3850 17604
rect 4126 17595 4184 17601
rect 4126 17592 4138 17595
rect 3844 17564 4138 17592
rect 3844 17552 3850 17564
rect 4126 17561 4138 17564
rect 4172 17561 4184 17595
rect 6472 17592 6500 17623
rect 6546 17620 6552 17672
rect 6604 17660 6610 17672
rect 6748 17669 6776 17700
rect 7374 17688 7380 17740
rect 7432 17728 7438 17740
rect 13538 17728 13544 17740
rect 7432 17700 13544 17728
rect 7432 17688 7438 17700
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 15488 17737 15516 17768
rect 15672 17768 16681 17796
rect 15672 17740 15700 17768
rect 16669 17765 16681 17768
rect 16715 17796 16727 17799
rect 16758 17796 16764 17808
rect 16715 17768 16764 17796
rect 16715 17765 16727 17768
rect 16669 17759 16727 17765
rect 16758 17756 16764 17768
rect 16816 17756 16822 17808
rect 17405 17799 17463 17805
rect 17405 17765 17417 17799
rect 17451 17796 17463 17799
rect 17678 17796 17684 17808
rect 17451 17768 17684 17796
rect 17451 17765 17463 17768
rect 17405 17759 17463 17765
rect 17678 17756 17684 17768
rect 17736 17756 17742 17808
rect 15105 17731 15163 17737
rect 15105 17728 15117 17731
rect 13872 17700 15117 17728
rect 13872 17688 13878 17700
rect 6733 17663 6791 17669
rect 6604 17632 6649 17660
rect 6604 17620 6610 17632
rect 6733 17629 6745 17663
rect 6779 17629 6791 17663
rect 6733 17623 6791 17629
rect 6822 17620 6828 17672
rect 6880 17660 6886 17672
rect 6917 17663 6975 17669
rect 6917 17660 6929 17663
rect 6880 17632 6929 17660
rect 6880 17620 6886 17632
rect 6917 17629 6929 17632
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 7837 17663 7895 17669
rect 7837 17660 7849 17663
rect 7800 17632 7849 17660
rect 7800 17620 7806 17632
rect 7837 17629 7849 17632
rect 7883 17629 7895 17663
rect 7837 17623 7895 17629
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17660 8171 17663
rect 8159 17632 8800 17660
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 7006 17592 7012 17604
rect 4126 17555 4184 17561
rect 5092 17564 6408 17592
rect 6472 17564 7012 17592
rect 2774 17524 2780 17536
rect 2735 17496 2780 17524
rect 2774 17484 2780 17496
rect 2832 17484 2838 17536
rect 3050 17524 3056 17536
rect 3011 17496 3056 17524
rect 3050 17484 3056 17496
rect 3108 17484 3114 17536
rect 3510 17484 3516 17536
rect 3568 17524 3574 17536
rect 5092 17524 5120 17564
rect 5258 17524 5264 17536
rect 3568 17496 5120 17524
rect 5219 17496 5264 17524
rect 3568 17484 3574 17496
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 6273 17527 6331 17533
rect 6273 17524 6285 17527
rect 6052 17496 6285 17524
rect 6052 17484 6058 17496
rect 6273 17493 6285 17496
rect 6319 17493 6331 17527
rect 6380 17524 6408 17564
rect 7006 17552 7012 17564
rect 7064 17552 7070 17604
rect 8772 17592 8800 17632
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 8904 17632 9781 17660
rect 8904 17620 8910 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 10778 17660 10784 17672
rect 10739 17632 10784 17660
rect 9769 17623 9827 17629
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 10870 17620 10876 17672
rect 10928 17660 10934 17672
rect 11149 17663 11207 17669
rect 10928 17632 10973 17660
rect 10928 17620 10934 17632
rect 11149 17629 11161 17663
rect 11195 17629 11207 17663
rect 11149 17623 11207 17629
rect 9490 17592 9496 17604
rect 7300 17564 8248 17592
rect 8772 17564 9496 17592
rect 7300 17524 7328 17564
rect 8110 17524 8116 17536
rect 6380 17496 7328 17524
rect 8071 17496 8116 17524
rect 6273 17487 6331 17493
rect 8110 17484 8116 17496
rect 8168 17484 8174 17536
rect 8220 17524 8248 17564
rect 9490 17552 9496 17564
rect 9548 17592 9554 17604
rect 9585 17595 9643 17601
rect 9585 17592 9597 17595
rect 9548 17564 9597 17592
rect 9548 17552 9554 17564
rect 9585 17561 9597 17564
rect 9631 17561 9643 17595
rect 9585 17555 9643 17561
rect 9953 17595 10011 17601
rect 9953 17561 9965 17595
rect 9999 17592 10011 17595
rect 10318 17592 10324 17604
rect 9999 17564 10324 17592
rect 9999 17561 10011 17564
rect 9953 17555 10011 17561
rect 10318 17552 10324 17564
rect 10376 17552 10382 17604
rect 10796 17592 10824 17620
rect 11164 17592 11192 17623
rect 11238 17620 11244 17672
rect 11296 17660 11302 17672
rect 11517 17663 11575 17669
rect 11517 17660 11529 17663
rect 11296 17632 11529 17660
rect 11296 17620 11302 17632
rect 11517 17629 11529 17632
rect 11563 17629 11575 17663
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11517 17623 11575 17629
rect 11716 17632 11805 17660
rect 11716 17592 11744 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11974 17660 11980 17672
rect 11935 17632 11980 17660
rect 11793 17623 11851 17629
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 12066 17620 12072 17672
rect 12124 17660 12130 17672
rect 12529 17663 12587 17669
rect 12529 17660 12541 17663
rect 12124 17632 12541 17660
rect 12124 17620 12130 17632
rect 12529 17629 12541 17632
rect 12575 17629 12587 17663
rect 12529 17623 12587 17629
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17660 12771 17663
rect 12802 17660 12808 17672
rect 12759 17632 12808 17660
rect 12759 17629 12771 17632
rect 12713 17623 12771 17629
rect 12728 17592 12756 17623
rect 12802 17620 12808 17632
rect 12860 17620 12866 17672
rect 13078 17620 13084 17672
rect 13136 17660 13142 17672
rect 13265 17663 13323 17669
rect 13265 17660 13277 17663
rect 13136 17632 13277 17660
rect 13136 17620 13142 17632
rect 13265 17629 13277 17632
rect 13311 17629 13323 17663
rect 13265 17623 13323 17629
rect 13357 17663 13415 17669
rect 13357 17629 13369 17663
rect 13403 17660 13415 17663
rect 13449 17663 13507 17669
rect 13449 17660 13461 17663
rect 13403 17632 13461 17660
rect 13403 17629 13415 17632
rect 13357 17623 13415 17629
rect 13449 17629 13461 17632
rect 13495 17660 13507 17663
rect 13998 17660 14004 17672
rect 13495 17632 14004 17660
rect 13495 17629 13507 17632
rect 13449 17623 13507 17629
rect 13998 17620 14004 17632
rect 14056 17620 14062 17672
rect 14108 17669 14136 17700
rect 15105 17697 15117 17700
rect 15151 17697 15163 17731
rect 15105 17691 15163 17697
rect 15473 17731 15531 17737
rect 15473 17697 15485 17731
rect 15519 17697 15531 17731
rect 15654 17728 15660 17740
rect 15615 17700 15660 17728
rect 15473 17691 15531 17697
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 15933 17731 15991 17737
rect 15933 17697 15945 17731
rect 15979 17728 15991 17731
rect 16574 17728 16580 17740
rect 15979 17700 16580 17728
rect 15979 17697 15991 17700
rect 15933 17691 15991 17697
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 14826 17620 14832 17672
rect 14884 17660 14890 17672
rect 15565 17663 15623 17669
rect 15565 17660 15577 17663
rect 14884 17632 15577 17660
rect 14884 17620 14890 17632
rect 15565 17629 15577 17632
rect 15611 17629 15623 17663
rect 16022 17660 16028 17672
rect 15983 17632 16028 17660
rect 15565 17623 15623 17629
rect 16022 17620 16028 17632
rect 16080 17620 16086 17672
rect 16761 17663 16819 17669
rect 16761 17629 16773 17663
rect 16807 17660 16819 17663
rect 16850 17660 16856 17672
rect 16807 17632 16856 17660
rect 16807 17629 16819 17632
rect 16761 17623 16819 17629
rect 16850 17620 16856 17632
rect 16908 17620 16914 17672
rect 17218 17660 17224 17672
rect 17131 17632 17224 17660
rect 10796 17564 11192 17592
rect 11256 17564 11744 17592
rect 11808 17564 12756 17592
rect 9766 17524 9772 17536
rect 8220 17496 9772 17524
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 10870 17484 10876 17536
rect 10928 17524 10934 17536
rect 11256 17533 11284 17564
rect 11241 17527 11299 17533
rect 11241 17524 11253 17527
rect 10928 17496 11253 17524
rect 10928 17484 10934 17496
rect 11241 17493 11253 17496
rect 11287 17493 11299 17527
rect 11241 17487 11299 17493
rect 11701 17527 11759 17533
rect 11701 17493 11713 17527
rect 11747 17524 11759 17527
rect 11808 17524 11836 17564
rect 13170 17552 13176 17604
rect 13228 17592 13234 17604
rect 15197 17595 15255 17601
rect 15197 17592 15209 17595
rect 13228 17564 15209 17592
rect 13228 17552 13234 17564
rect 15197 17561 15209 17564
rect 15243 17561 15255 17595
rect 15197 17555 15255 17561
rect 16040 17564 16344 17592
rect 11747 17496 11836 17524
rect 11747 17493 11759 17496
rect 11701 17487 11759 17493
rect 11882 17484 11888 17536
rect 11940 17524 11946 17536
rect 12989 17527 13047 17533
rect 12989 17524 13001 17527
rect 11940 17496 13001 17524
rect 11940 17484 11946 17496
rect 12989 17493 13001 17496
rect 13035 17493 13047 17527
rect 12989 17487 13047 17493
rect 13262 17484 13268 17536
rect 13320 17524 13326 17536
rect 13449 17527 13507 17533
rect 13449 17524 13461 17527
rect 13320 17496 13461 17524
rect 13320 17484 13326 17496
rect 13449 17493 13461 17496
rect 13495 17493 13507 17527
rect 13449 17487 13507 17493
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 16040 17524 16068 17564
rect 14700 17496 16068 17524
rect 14700 17484 14706 17496
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 16209 17527 16267 17533
rect 16209 17524 16221 17527
rect 16172 17496 16221 17524
rect 16172 17484 16178 17496
rect 16209 17493 16221 17496
rect 16255 17493 16267 17527
rect 16316 17524 16344 17564
rect 16390 17552 16396 17604
rect 16448 17592 16454 17604
rect 17144 17592 17172 17632
rect 17218 17620 17224 17632
rect 17276 17620 17282 17672
rect 16448 17564 17172 17592
rect 17880 17592 17908 17827
rect 18506 17824 18512 17876
rect 18564 17864 18570 17876
rect 20073 17867 20131 17873
rect 18564 17836 19840 17864
rect 18564 17824 18570 17836
rect 19702 17796 19708 17808
rect 18248 17768 19708 17796
rect 18248 17669 18276 17768
rect 19702 17756 19708 17768
rect 19760 17756 19766 17808
rect 19150 17688 19156 17740
rect 19208 17728 19214 17740
rect 19426 17728 19432 17740
rect 19208 17700 19432 17728
rect 19208 17688 19214 17700
rect 19426 17688 19432 17700
rect 19484 17688 19490 17740
rect 19812 17728 19840 17836
rect 20073 17833 20085 17867
rect 20119 17864 20131 17867
rect 20162 17864 20168 17876
rect 20119 17836 20168 17864
rect 20119 17833 20131 17836
rect 20073 17827 20131 17833
rect 20162 17824 20168 17836
rect 20220 17824 20226 17876
rect 20441 17731 20499 17737
rect 20441 17728 20453 17731
rect 19812 17700 20453 17728
rect 20441 17697 20453 17700
rect 20487 17697 20499 17731
rect 20441 17691 20499 17697
rect 22462 17688 22468 17740
rect 22520 17728 22526 17740
rect 23382 17728 23388 17740
rect 22520 17700 23388 17728
rect 22520 17688 22526 17700
rect 23382 17688 23388 17700
rect 23440 17728 23446 17740
rect 24394 17728 24400 17740
rect 23440 17700 24400 17728
rect 23440 17688 23446 17700
rect 24394 17688 24400 17700
rect 24452 17728 24458 17740
rect 24581 17731 24639 17737
rect 24581 17728 24593 17731
rect 24452 17700 24593 17728
rect 24452 17688 24458 17700
rect 24581 17697 24593 17700
rect 24627 17697 24639 17731
rect 24581 17691 24639 17697
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17629 18291 17663
rect 18414 17660 18420 17672
rect 18375 17632 18420 17660
rect 18233 17623 18291 17629
rect 18414 17620 18420 17632
rect 18472 17620 18478 17672
rect 18506 17620 18512 17672
rect 18564 17660 18570 17672
rect 18637 17660 18695 17666
rect 18564 17632 18609 17660
rect 18564 17620 18570 17632
rect 18637 17626 18649 17660
rect 18683 17626 18695 17660
rect 18637 17620 18695 17626
rect 18785 17663 18843 17669
rect 18785 17629 18797 17663
rect 18831 17660 18843 17663
rect 20162 17660 20168 17672
rect 18831 17632 20168 17660
rect 18831 17629 18843 17632
rect 18785 17623 18843 17629
rect 20162 17620 20168 17632
rect 20220 17620 20226 17672
rect 20346 17660 20352 17672
rect 20307 17632 20352 17660
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20530 17660 20536 17672
rect 20491 17632 20536 17660
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 20717 17663 20775 17669
rect 20717 17629 20729 17663
rect 20763 17629 20775 17663
rect 20717 17623 20775 17629
rect 18652 17592 18680 17620
rect 17880 17564 18680 17592
rect 19613 17595 19671 17601
rect 16448 17552 16454 17564
rect 19613 17561 19625 17595
rect 19659 17592 19671 17595
rect 20732 17592 20760 17623
rect 22646 17620 22652 17672
rect 22704 17660 22710 17672
rect 22925 17663 22983 17669
rect 22925 17660 22937 17663
rect 22704 17632 22937 17660
rect 22704 17620 22710 17632
rect 22925 17629 22937 17632
rect 22971 17629 22983 17663
rect 23198 17660 23204 17672
rect 23159 17632 23204 17660
rect 22925 17623 22983 17629
rect 23198 17620 23204 17632
rect 23256 17620 23262 17672
rect 19659 17564 20760 17592
rect 19659 17561 19671 17564
rect 19613 17555 19671 17561
rect 17310 17524 17316 17536
rect 16316 17496 17316 17524
rect 16209 17487 16267 17493
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 18138 17524 18144 17536
rect 18099 17496 18144 17524
rect 18138 17484 18144 17496
rect 18196 17484 18202 17536
rect 19334 17484 19340 17536
rect 19392 17524 19398 17536
rect 19705 17527 19763 17533
rect 19705 17524 19717 17527
rect 19392 17496 19717 17524
rect 19392 17484 19398 17496
rect 19705 17493 19717 17496
rect 19751 17493 19763 17527
rect 20732 17524 20760 17564
rect 20901 17595 20959 17601
rect 20901 17561 20913 17595
rect 20947 17592 20959 17595
rect 22198 17595 22256 17601
rect 22198 17592 22210 17595
rect 20947 17564 22210 17592
rect 20947 17561 20959 17564
rect 20901 17555 20959 17561
rect 22198 17561 22210 17564
rect 22244 17561 22256 17595
rect 24854 17592 24860 17604
rect 24815 17564 24860 17592
rect 22198 17555 22256 17561
rect 24854 17552 24860 17564
rect 24912 17552 24918 17604
rect 25498 17552 25504 17604
rect 25556 17552 25562 17604
rect 21085 17527 21143 17533
rect 21085 17524 21097 17527
rect 20732 17496 21097 17524
rect 19705 17487 19763 17493
rect 21085 17493 21097 17496
rect 21131 17493 21143 17527
rect 21085 17487 21143 17493
rect 23109 17527 23167 17533
rect 23109 17493 23121 17527
rect 23155 17524 23167 17527
rect 23198 17524 23204 17536
rect 23155 17496 23204 17524
rect 23155 17493 23167 17496
rect 23109 17487 23167 17493
rect 23198 17484 23204 17496
rect 23256 17484 23262 17536
rect 23385 17527 23443 17533
rect 23385 17493 23397 17527
rect 23431 17524 23443 17527
rect 24210 17524 24216 17536
rect 23431 17496 24216 17524
rect 23431 17493 23443 17496
rect 23385 17487 23443 17493
rect 24210 17484 24216 17496
rect 24268 17484 24274 17536
rect 24762 17484 24768 17536
rect 24820 17524 24826 17536
rect 26329 17527 26387 17533
rect 26329 17524 26341 17527
rect 24820 17496 26341 17524
rect 24820 17484 24826 17496
rect 26329 17493 26341 17496
rect 26375 17493 26387 17527
rect 26329 17487 26387 17493
rect 1104 17434 29440 17456
rect 1104 17382 10395 17434
rect 10447 17382 10459 17434
rect 10511 17382 10523 17434
rect 10575 17382 10587 17434
rect 10639 17382 10651 17434
rect 10703 17382 19840 17434
rect 19892 17382 19904 17434
rect 19956 17382 19968 17434
rect 20020 17382 20032 17434
rect 20084 17382 20096 17434
rect 20148 17382 29440 17434
rect 1104 17360 29440 17382
rect 2222 17320 2228 17332
rect 2183 17292 2228 17320
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 2593 17323 2651 17329
rect 2593 17289 2605 17323
rect 2639 17320 2651 17323
rect 2774 17320 2780 17332
rect 2639 17292 2780 17320
rect 2639 17289 2651 17292
rect 2593 17283 2651 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 4154 17320 4160 17332
rect 4115 17292 4160 17320
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 7006 17280 7012 17332
rect 7064 17320 7070 17332
rect 7190 17320 7196 17332
rect 7064 17292 7196 17320
rect 7064 17280 7070 17292
rect 7190 17280 7196 17292
rect 7248 17280 7254 17332
rect 7558 17320 7564 17332
rect 7519 17292 7564 17320
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 7650 17280 7656 17332
rect 7708 17320 7714 17332
rect 8846 17320 8852 17332
rect 7708 17292 8156 17320
rect 8807 17292 8852 17320
rect 7708 17280 7714 17292
rect 2792 17252 2820 17280
rect 4985 17255 5043 17261
rect 2792 17224 3648 17252
rect 3053 17187 3111 17193
rect 3053 17184 3065 17187
rect 2792 17156 3065 17184
rect 2685 17119 2743 17125
rect 2685 17085 2697 17119
rect 2731 17116 2743 17119
rect 2792 17116 2820 17156
rect 3053 17153 3065 17156
rect 3099 17153 3111 17187
rect 3053 17147 3111 17153
rect 3142 17144 3148 17196
rect 3200 17184 3206 17196
rect 3620 17193 3648 17224
rect 4985 17221 4997 17255
rect 5031 17252 5043 17255
rect 5258 17252 5264 17264
rect 5031 17224 5264 17252
rect 5031 17221 5043 17224
rect 4985 17215 5043 17221
rect 5258 17212 5264 17224
rect 5316 17212 5322 17264
rect 6822 17252 6828 17264
rect 6783 17224 6828 17252
rect 6822 17212 6828 17224
rect 6880 17212 6886 17264
rect 6917 17255 6975 17261
rect 6917 17221 6929 17255
rect 6963 17252 6975 17255
rect 6963 17224 8064 17252
rect 6963 17221 6975 17224
rect 6917 17215 6975 17221
rect 3238 17187 3296 17193
rect 3238 17184 3250 17187
rect 3200 17156 3250 17184
rect 3200 17144 3206 17156
rect 3238 17153 3250 17156
rect 3284 17153 3296 17187
rect 3238 17147 3296 17153
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17153 3663 17187
rect 3605 17147 3663 17153
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17184 3755 17187
rect 4890 17184 4896 17196
rect 3743 17156 4896 17184
rect 3743 17153 3755 17156
rect 3697 17147 3755 17153
rect 4890 17144 4896 17156
rect 4948 17144 4954 17196
rect 5169 17187 5227 17193
rect 5169 17153 5181 17187
rect 5215 17184 5227 17187
rect 5534 17184 5540 17196
rect 5215 17156 5540 17184
rect 5215 17153 5227 17156
rect 5169 17147 5227 17153
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 6546 17184 6552 17196
rect 6507 17156 6552 17184
rect 6546 17144 6552 17156
rect 6604 17184 6610 17196
rect 7098 17184 7104 17196
rect 6604 17156 7104 17184
rect 6604 17144 6610 17156
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 7190 17144 7196 17196
rect 7248 17184 7254 17196
rect 7466 17193 7472 17196
rect 7449 17187 7472 17193
rect 7248 17156 7293 17184
rect 7248 17144 7254 17156
rect 7449 17153 7461 17187
rect 7449 17147 7472 17153
rect 7466 17144 7472 17147
rect 7524 17144 7530 17196
rect 7834 17184 7840 17196
rect 7567 17156 7840 17184
rect 2731 17088 2820 17116
rect 2869 17119 2927 17125
rect 2731 17085 2743 17088
rect 2685 17079 2743 17085
rect 2869 17085 2881 17119
rect 2915 17085 2927 17119
rect 4246 17116 4252 17128
rect 4207 17088 4252 17116
rect 2869 17079 2927 17085
rect 2884 17048 2912 17079
rect 4246 17076 4252 17088
rect 4304 17076 4310 17128
rect 4430 17116 4436 17128
rect 4391 17088 4436 17116
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 6733 17119 6791 17125
rect 6733 17085 6745 17119
rect 6779 17116 6791 17119
rect 6914 17116 6920 17128
rect 6779 17088 6920 17116
rect 6779 17085 6791 17088
rect 6733 17079 6791 17085
rect 6914 17076 6920 17088
rect 6972 17116 6978 17128
rect 7567 17116 7595 17156
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 8036 17128 8064 17224
rect 8128 17184 8156 17292
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 9214 17280 9220 17332
rect 9272 17280 9278 17332
rect 10778 17320 10784 17332
rect 10739 17292 10784 17320
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 11238 17280 11244 17332
rect 11296 17320 11302 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11296 17292 11621 17320
rect 11296 17280 11302 17292
rect 11609 17289 11621 17292
rect 11655 17320 11667 17323
rect 12066 17320 12072 17332
rect 11655 17292 12072 17320
rect 11655 17289 11667 17292
rect 11609 17283 11667 17289
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 12342 17280 12348 17332
rect 12400 17320 12406 17332
rect 12621 17323 12679 17329
rect 12621 17320 12633 17323
rect 12400 17292 12633 17320
rect 12400 17280 12406 17292
rect 12621 17289 12633 17292
rect 12667 17289 12679 17323
rect 12621 17283 12679 17289
rect 13538 17280 13544 17332
rect 13596 17320 13602 17332
rect 13596 17292 13768 17320
rect 13596 17280 13602 17292
rect 9232 17252 9260 17280
rect 9232 17224 9444 17252
rect 8205 17187 8263 17193
rect 8205 17184 8217 17187
rect 8128 17156 8217 17184
rect 8205 17153 8217 17156
rect 8251 17153 8263 17187
rect 8665 17187 8723 17193
rect 8665 17184 8677 17187
rect 8205 17147 8263 17153
rect 8312 17156 8677 17184
rect 6972 17088 7595 17116
rect 7653 17119 7711 17125
rect 6972 17076 6978 17088
rect 7653 17085 7665 17119
rect 7699 17085 7711 17119
rect 7653 17079 7711 17085
rect 2958 17048 2964 17060
rect 2884 17020 2964 17048
rect 2958 17008 2964 17020
rect 3016 17008 3022 17060
rect 7374 17048 7380 17060
rect 3620 17020 7380 17048
rect 1302 16940 1308 16992
rect 1360 16980 1366 16992
rect 3620 16980 3648 17020
rect 7374 17008 7380 17020
rect 7432 17008 7438 17060
rect 3786 16980 3792 16992
rect 1360 16952 3648 16980
rect 3747 16952 3792 16980
rect 1360 16940 1366 16952
rect 3786 16940 3792 16952
rect 3844 16940 3850 16992
rect 4890 16980 4896 16992
rect 4851 16952 4896 16980
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 6638 16940 6644 16992
rect 6696 16980 6702 16992
rect 7193 16983 7251 16989
rect 7193 16980 7205 16983
rect 6696 16952 7205 16980
rect 6696 16940 6702 16952
rect 7193 16949 7205 16952
rect 7239 16980 7251 16983
rect 7466 16980 7472 16992
rect 7239 16952 7472 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 7668 16980 7696 17079
rect 7742 17076 7748 17128
rect 7800 17116 7806 17128
rect 7800 17088 7893 17116
rect 7800 17076 7806 17088
rect 8018 17076 8024 17128
rect 8076 17116 8082 17128
rect 8312 17116 8340 17156
rect 8665 17153 8677 17156
rect 8711 17153 8723 17187
rect 8665 17147 8723 17153
rect 9214 17144 9220 17196
rect 9272 17184 9278 17196
rect 9416 17193 9444 17224
rect 10318 17212 10324 17264
rect 10376 17252 10382 17264
rect 13740 17261 13768 17292
rect 13998 17280 14004 17332
rect 14056 17280 14062 17332
rect 15010 17320 15016 17332
rect 14971 17292 15016 17320
rect 15010 17280 15016 17292
rect 15068 17280 15074 17332
rect 17037 17323 17095 17329
rect 17037 17320 17049 17323
rect 15120 17292 17049 17320
rect 13725 17255 13783 17261
rect 10376 17224 13676 17252
rect 10376 17212 10382 17224
rect 9309 17187 9367 17193
rect 9309 17184 9321 17187
rect 9272 17156 9321 17184
rect 9272 17144 9278 17156
rect 9309 17153 9321 17156
rect 9355 17153 9367 17187
rect 9309 17147 9367 17153
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17153 9459 17187
rect 9401 17147 9459 17153
rect 9668 17187 9726 17193
rect 9668 17153 9680 17187
rect 9714 17184 9726 17187
rect 9950 17184 9956 17196
rect 9714 17156 9956 17184
rect 9714 17153 9726 17156
rect 9668 17147 9726 17153
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 10962 17144 10968 17196
rect 11020 17184 11026 17196
rect 11514 17184 11520 17196
rect 11020 17156 11520 17184
rect 11020 17144 11026 17156
rect 11514 17144 11520 17156
rect 11572 17144 11578 17196
rect 12618 17144 12624 17196
rect 12676 17184 12682 17196
rect 12713 17187 12771 17193
rect 12713 17184 12725 17187
rect 12676 17156 12725 17184
rect 12676 17144 12682 17156
rect 12713 17153 12725 17156
rect 12759 17153 12771 17187
rect 12713 17147 12771 17153
rect 12897 17187 12955 17193
rect 12897 17153 12909 17187
rect 12943 17153 12955 17187
rect 13078 17184 13084 17196
rect 13039 17156 13084 17184
rect 12897 17147 12955 17153
rect 8076 17088 8340 17116
rect 8389 17119 8447 17125
rect 8076 17076 8082 17088
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 8478 17116 8484 17128
rect 8435 17088 8484 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 8478 17076 8484 17088
rect 8536 17076 8542 17128
rect 9033 17119 9091 17125
rect 9033 17085 9045 17119
rect 9079 17085 9091 17119
rect 12912 17116 12940 17147
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 13354 17184 13360 17196
rect 13315 17156 13360 17184
rect 13354 17144 13360 17156
rect 13412 17144 13418 17196
rect 13538 17184 13544 17196
rect 13499 17156 13544 17184
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 13648 17184 13676 17224
rect 13725 17221 13737 17255
rect 13771 17221 13783 17255
rect 14016 17252 14044 17280
rect 15120 17252 15148 17292
rect 17037 17289 17049 17292
rect 17083 17289 17095 17323
rect 17037 17283 17095 17289
rect 17681 17323 17739 17329
rect 17681 17289 17693 17323
rect 17727 17320 17739 17323
rect 18046 17320 18052 17332
rect 17727 17292 18052 17320
rect 17727 17289 17739 17292
rect 17681 17283 17739 17289
rect 18046 17280 18052 17292
rect 18104 17320 18110 17332
rect 18782 17320 18788 17332
rect 18104 17292 18788 17320
rect 18104 17280 18110 17292
rect 18782 17280 18788 17292
rect 18840 17280 18846 17332
rect 19613 17323 19671 17329
rect 19613 17289 19625 17323
rect 19659 17320 19671 17323
rect 19702 17320 19708 17332
rect 19659 17292 19708 17320
rect 19659 17289 19671 17292
rect 19613 17283 19671 17289
rect 19702 17280 19708 17292
rect 19760 17280 19766 17332
rect 20346 17280 20352 17332
rect 20404 17320 20410 17332
rect 21085 17323 21143 17329
rect 21085 17320 21097 17323
rect 20404 17292 21097 17320
rect 20404 17280 20410 17292
rect 21085 17289 21097 17292
rect 21131 17320 21143 17323
rect 21174 17320 21180 17332
rect 21131 17292 21180 17320
rect 21131 17289 21143 17292
rect 21085 17283 21143 17289
rect 21174 17280 21180 17292
rect 21232 17280 21238 17332
rect 25498 17320 25504 17332
rect 25459 17292 25504 17320
rect 25498 17280 25504 17292
rect 25556 17280 25562 17332
rect 25682 17280 25688 17332
rect 25740 17320 25746 17332
rect 25777 17323 25835 17329
rect 25777 17320 25789 17323
rect 25740 17292 25789 17320
rect 25740 17280 25746 17292
rect 25777 17289 25789 17292
rect 25823 17289 25835 17323
rect 25777 17283 25835 17289
rect 14016 17224 15148 17252
rect 13725 17215 13783 17221
rect 15930 17212 15936 17264
rect 15988 17212 15994 17264
rect 16758 17252 16764 17264
rect 16316 17224 16764 17252
rect 14642 17184 14648 17196
rect 13648 17156 14648 17184
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 15565 17187 15623 17193
rect 15565 17184 15577 17187
rect 14844 17156 15577 17184
rect 13265 17119 13323 17125
rect 12912 17088 13216 17116
rect 9033 17079 9091 17085
rect 7760 17048 7788 17076
rect 7929 17051 7987 17057
rect 7929 17048 7941 17051
rect 7760 17020 7941 17048
rect 7929 17017 7941 17020
rect 7975 17048 7987 17051
rect 9048 17048 9076 17079
rect 7975 17020 9076 17048
rect 13188 17048 13216 17088
rect 13265 17085 13277 17119
rect 13311 17116 13323 17119
rect 14734 17116 14740 17128
rect 13311 17088 14740 17116
rect 13311 17085 13323 17088
rect 13265 17079 13323 17085
rect 14734 17076 14740 17088
rect 14792 17076 14798 17128
rect 14642 17048 14648 17060
rect 13188 17020 14648 17048
rect 7975 17017 7987 17020
rect 7929 17011 7987 17017
rect 14642 17008 14648 17020
rect 14700 17048 14706 17060
rect 14844 17048 14872 17156
rect 15565 17153 15577 17156
rect 15611 17153 15623 17187
rect 15565 17147 15623 17153
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17184 15899 17187
rect 15948 17184 15976 17212
rect 15887 17156 15976 17184
rect 16117 17187 16175 17193
rect 15887 17153 15899 17156
rect 15841 17147 15899 17153
rect 16117 17153 16129 17187
rect 16163 17184 16175 17187
rect 16206 17184 16212 17196
rect 16163 17156 16212 17184
rect 16163 17153 16175 17156
rect 16117 17147 16175 17153
rect 16206 17144 16212 17156
rect 16264 17144 16270 17196
rect 16316 17193 16344 17224
rect 16758 17212 16764 17224
rect 16816 17212 16822 17264
rect 18138 17212 18144 17264
rect 18196 17252 18202 17264
rect 18478 17255 18536 17261
rect 18478 17252 18490 17255
rect 18196 17224 18490 17252
rect 18196 17212 18202 17224
rect 18478 17221 18490 17224
rect 18524 17221 18536 17255
rect 18478 17215 18536 17221
rect 19150 17212 19156 17264
rect 19208 17212 19214 17264
rect 23842 17252 23848 17264
rect 23690 17224 23848 17252
rect 23842 17212 23848 17224
rect 23900 17212 23906 17264
rect 24210 17212 24216 17264
rect 24268 17252 24274 17264
rect 24762 17252 24768 17264
rect 24268 17224 24624 17252
rect 24723 17224 24768 17252
rect 24268 17212 24274 17224
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 16632 17156 16681 17184
rect 16632 17144 16638 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 17218 17144 17224 17196
rect 17276 17184 17282 17196
rect 17405 17187 17463 17193
rect 17405 17184 17417 17187
rect 17276 17156 17417 17184
rect 17276 17144 17282 17156
rect 17405 17153 17417 17156
rect 17451 17184 17463 17187
rect 17497 17187 17555 17193
rect 17497 17184 17509 17187
rect 17451 17156 17509 17184
rect 17451 17153 17463 17156
rect 17405 17147 17463 17153
rect 17497 17153 17509 17156
rect 17543 17153 17555 17187
rect 17954 17184 17960 17196
rect 17915 17156 17960 17184
rect 17497 17147 17555 17153
rect 17954 17144 17960 17156
rect 18012 17144 18018 17196
rect 18230 17184 18236 17196
rect 18191 17156 18236 17184
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 19168 17184 19196 17212
rect 18340 17156 19196 17184
rect 24489 17187 24547 17193
rect 15654 17076 15660 17128
rect 15712 17116 15718 17128
rect 15933 17119 15991 17125
rect 15933 17116 15945 17119
rect 15712 17088 15945 17116
rect 15712 17076 15718 17088
rect 15933 17085 15945 17088
rect 15979 17085 15991 17119
rect 15933 17079 15991 17085
rect 16761 17119 16819 17125
rect 16761 17085 16773 17119
rect 16807 17116 16819 17119
rect 16850 17116 16856 17128
rect 16807 17088 16856 17116
rect 16807 17085 16819 17088
rect 16761 17079 16819 17085
rect 16850 17076 16856 17088
rect 16908 17116 16914 17128
rect 18340 17116 18368 17156
rect 24489 17153 24501 17187
rect 24535 17184 24547 17187
rect 24596 17184 24624 17224
rect 24762 17212 24768 17224
rect 24820 17252 24826 17264
rect 25593 17255 25651 17261
rect 25593 17252 25605 17255
rect 24820 17224 25605 17252
rect 24820 17212 24826 17224
rect 25593 17221 25605 17224
rect 25639 17221 25651 17255
rect 25593 17215 25651 17221
rect 24946 17193 24952 17196
rect 24535 17156 24624 17184
rect 24673 17187 24731 17193
rect 24535 17153 24547 17156
rect 24489 17147 24547 17153
rect 24673 17153 24685 17187
rect 24719 17153 24731 17187
rect 24673 17147 24731 17153
rect 24909 17187 24952 17193
rect 24909 17153 24921 17187
rect 24909 17147 24952 17153
rect 22646 17116 22652 17128
rect 16908 17088 18368 17116
rect 22607 17088 22652 17116
rect 16908 17076 16914 17088
rect 22646 17076 22652 17088
rect 22704 17076 22710 17128
rect 23474 17076 23480 17128
rect 23532 17116 23538 17128
rect 24121 17119 24179 17125
rect 24121 17116 24133 17119
rect 23532 17088 24133 17116
rect 23532 17076 23538 17088
rect 24121 17085 24133 17088
rect 24167 17085 24179 17119
rect 24394 17116 24400 17128
rect 24355 17088 24400 17116
rect 24121 17079 24179 17085
rect 24394 17076 24400 17088
rect 24452 17076 24458 17128
rect 24688 17116 24716 17147
rect 24946 17144 24952 17147
rect 25004 17144 25010 17196
rect 25314 17184 25320 17196
rect 25275 17156 25320 17184
rect 25314 17144 25320 17156
rect 25372 17144 25378 17196
rect 25682 17116 25688 17128
rect 24688 17088 25688 17116
rect 25682 17076 25688 17088
rect 25740 17076 25746 17128
rect 14700 17020 14872 17048
rect 14700 17008 14706 17020
rect 16574 17008 16580 17060
rect 16632 17048 16638 17060
rect 17221 17051 17279 17057
rect 17221 17048 17233 17051
rect 16632 17020 17233 17048
rect 16632 17008 16638 17020
rect 17221 17017 17233 17020
rect 17267 17048 17279 17051
rect 17267 17020 17908 17048
rect 17267 17017 17279 17020
rect 17221 17011 17279 17017
rect 8481 16983 8539 16989
rect 8481 16980 8493 16983
rect 7668 16952 8493 16980
rect 8481 16949 8493 16952
rect 8527 16980 8539 16983
rect 8570 16980 8576 16992
rect 8527 16952 8576 16980
rect 8527 16949 8539 16952
rect 8481 16943 8539 16949
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 9217 16983 9275 16989
rect 9217 16949 9229 16983
rect 9263 16980 9275 16983
rect 9306 16980 9312 16992
rect 9263 16952 9312 16980
rect 9263 16949 9275 16952
rect 9217 16943 9275 16949
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 11790 16980 11796 16992
rect 9824 16952 11796 16980
rect 9824 16940 9830 16952
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 16666 16980 16672 16992
rect 16627 16952 16672 16980
rect 16666 16940 16672 16952
rect 16724 16940 16730 16992
rect 17770 16980 17776 16992
rect 17731 16952 17776 16980
rect 17770 16940 17776 16952
rect 17828 16940 17834 16992
rect 17880 16980 17908 17020
rect 24854 17008 24860 17060
rect 24912 17048 24918 17060
rect 25041 17051 25099 17057
rect 25041 17048 25053 17051
rect 24912 17020 25053 17048
rect 24912 17008 24918 17020
rect 25041 17017 25053 17020
rect 25087 17017 25099 17051
rect 25041 17011 25099 17017
rect 24302 16980 24308 16992
rect 17880 16952 24308 16980
rect 24302 16940 24308 16952
rect 24360 16940 24366 16992
rect 1104 16890 29440 16912
rect 1104 16838 5672 16890
rect 5724 16838 5736 16890
rect 5788 16838 5800 16890
rect 5852 16838 5864 16890
rect 5916 16838 5928 16890
rect 5980 16838 15118 16890
rect 15170 16838 15182 16890
rect 15234 16838 15246 16890
rect 15298 16838 15310 16890
rect 15362 16838 15374 16890
rect 15426 16838 24563 16890
rect 24615 16838 24627 16890
rect 24679 16838 24691 16890
rect 24743 16838 24755 16890
rect 24807 16838 24819 16890
rect 24871 16838 29440 16890
rect 1104 16816 29440 16838
rect 2685 16779 2743 16785
rect 2685 16745 2697 16779
rect 2731 16776 2743 16779
rect 2731 16748 2912 16776
rect 2731 16745 2743 16748
rect 2685 16739 2743 16745
rect 2884 16720 2912 16748
rect 3050 16736 3056 16788
rect 3108 16776 3114 16788
rect 7561 16779 7619 16785
rect 7561 16776 7573 16779
rect 3108 16748 7573 16776
rect 3108 16736 3114 16748
rect 2866 16668 2872 16720
rect 2924 16708 2930 16720
rect 3142 16708 3148 16720
rect 2924 16680 3148 16708
rect 2924 16668 2930 16680
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 2958 16600 2964 16652
rect 3016 16640 3022 16652
rect 4706 16640 4712 16652
rect 3016 16612 4712 16640
rect 3016 16600 3022 16612
rect 4706 16600 4712 16612
rect 4764 16640 4770 16652
rect 5368 16649 5396 16748
rect 7561 16745 7573 16748
rect 7607 16776 7619 16779
rect 8202 16776 8208 16788
rect 7607 16748 8208 16776
rect 7607 16745 7619 16748
rect 7561 16739 7619 16745
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 8570 16776 8576 16788
rect 8531 16748 8576 16776
rect 8570 16736 8576 16748
rect 8628 16736 8634 16788
rect 12986 16776 12992 16788
rect 12947 16748 12992 16776
rect 12986 16736 12992 16748
rect 13044 16736 13050 16788
rect 13262 16776 13268 16788
rect 13223 16748 13268 16776
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 13538 16776 13544 16788
rect 13372 16748 13544 16776
rect 7006 16708 7012 16720
rect 6967 16680 7012 16708
rect 7006 16668 7012 16680
rect 7064 16668 7070 16720
rect 7285 16711 7343 16717
rect 7285 16677 7297 16711
rect 7331 16708 7343 16711
rect 8018 16708 8024 16720
rect 7331 16680 8024 16708
rect 7331 16677 7343 16680
rect 7285 16671 7343 16677
rect 8018 16668 8024 16680
rect 8076 16668 8082 16720
rect 8389 16711 8447 16717
rect 8389 16677 8401 16711
rect 8435 16708 8447 16711
rect 9214 16708 9220 16720
rect 8435 16680 9220 16708
rect 8435 16677 8447 16680
rect 8389 16671 8447 16677
rect 9214 16668 9220 16680
rect 9272 16708 9278 16720
rect 9950 16708 9956 16720
rect 9272 16680 9536 16708
rect 9911 16680 9956 16708
rect 9272 16668 9278 16680
rect 4801 16643 4859 16649
rect 4801 16640 4813 16643
rect 4764 16612 4813 16640
rect 4764 16600 4770 16612
rect 4801 16609 4813 16612
rect 4847 16609 4859 16643
rect 4801 16603 4859 16609
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16609 5411 16643
rect 7024 16640 7052 16668
rect 7653 16643 7711 16649
rect 7653 16640 7665 16643
rect 7024 16612 7665 16640
rect 5353 16603 5411 16609
rect 7653 16609 7665 16612
rect 7699 16640 7711 16643
rect 7834 16640 7840 16652
rect 7699 16612 7840 16640
rect 7699 16609 7711 16612
rect 7653 16603 7711 16609
rect 7834 16600 7840 16612
rect 7892 16640 7898 16652
rect 8478 16640 8484 16652
rect 7892 16612 8484 16640
rect 7892 16600 7898 16612
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 9306 16640 9312 16652
rect 9267 16612 9312 16640
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 9508 16649 9536 16680
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16609 9551 16643
rect 9493 16603 9551 16609
rect 9674 16600 9680 16652
rect 9732 16640 9738 16652
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 9732 16612 10057 16640
rect 9732 16600 9738 16612
rect 10045 16609 10057 16612
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16609 11575 16643
rect 13170 16640 13176 16652
rect 11517 16603 11575 16609
rect 12544 16612 13176 16640
rect 2774 16572 2780 16584
rect 2735 16544 2780 16572
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 4430 16572 4436 16584
rect 2884 16544 4436 16572
rect 2498 16464 2504 16516
rect 2556 16504 2562 16516
rect 2884 16504 2912 16544
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16572 4675 16575
rect 5258 16572 5264 16584
rect 4663 16544 5264 16572
rect 4663 16541 4675 16544
rect 4617 16535 4675 16541
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 5620 16575 5678 16581
rect 5620 16541 5632 16575
rect 5666 16572 5678 16575
rect 5994 16572 6000 16584
rect 5666 16544 6000 16572
rect 5666 16541 5678 16544
rect 5620 16535 5678 16541
rect 5994 16532 6000 16544
rect 6052 16532 6058 16584
rect 7377 16575 7435 16581
rect 7377 16541 7389 16575
rect 7423 16572 7435 16575
rect 7558 16572 7564 16584
rect 7423 16544 7564 16572
rect 7423 16541 7435 16544
rect 7377 16535 7435 16541
rect 2556 16476 2912 16504
rect 2961 16507 3019 16513
rect 2556 16464 2562 16476
rect 2961 16473 2973 16507
rect 3007 16504 3019 16507
rect 4890 16504 4896 16516
rect 3007 16476 4896 16504
rect 3007 16473 3019 16476
rect 2961 16467 3019 16473
rect 4890 16464 4896 16476
rect 4948 16464 4954 16516
rect 7392 16504 7420 16535
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16572 7987 16575
rect 8570 16572 8576 16584
rect 7975 16544 8576 16572
rect 7975 16541 7987 16544
rect 7929 16535 7987 16541
rect 8570 16532 8576 16544
rect 8628 16572 8634 16584
rect 8665 16575 8723 16581
rect 8665 16572 8677 16575
rect 8628 16544 8677 16572
rect 8628 16532 8634 16544
rect 8665 16541 8677 16544
rect 8711 16541 8723 16575
rect 8665 16535 8723 16541
rect 8846 16532 8852 16584
rect 8904 16572 8910 16584
rect 9217 16575 9275 16581
rect 9217 16572 9229 16575
rect 8904 16544 9229 16572
rect 8904 16532 8910 16544
rect 9217 16541 9229 16544
rect 9263 16541 9275 16575
rect 9217 16535 9275 16541
rect 9585 16575 9643 16581
rect 9585 16541 9597 16575
rect 9631 16572 9643 16575
rect 10870 16572 10876 16584
rect 9631 16544 10876 16572
rect 9631 16541 9643 16544
rect 9585 16535 9643 16541
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 11238 16572 11244 16584
rect 11199 16544 11244 16572
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 11422 16572 11428 16584
rect 11383 16544 11428 16572
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 6748 16476 7420 16504
rect 4246 16436 4252 16448
rect 4207 16408 4252 16436
rect 4246 16396 4252 16408
rect 4304 16396 4310 16448
rect 4706 16396 4712 16448
rect 4764 16436 4770 16448
rect 6748 16445 6776 16476
rect 7466 16464 7472 16516
rect 7524 16504 7530 16516
rect 8021 16507 8079 16513
rect 8021 16504 8033 16507
rect 7524 16476 8033 16504
rect 7524 16464 7530 16476
rect 8021 16473 8033 16476
rect 8067 16473 8079 16507
rect 8021 16467 8079 16473
rect 8205 16507 8263 16513
rect 8205 16473 8217 16507
rect 8251 16504 8263 16507
rect 8294 16504 8300 16516
rect 8251 16476 8300 16504
rect 8251 16473 8263 16476
rect 8205 16467 8263 16473
rect 6733 16439 6791 16445
rect 4764 16408 4809 16436
rect 4764 16396 4770 16408
rect 6733 16405 6745 16439
rect 6779 16405 6791 16439
rect 6733 16399 6791 16405
rect 7374 16396 7380 16448
rect 7432 16436 7438 16448
rect 8220 16436 8248 16467
rect 8294 16464 8300 16476
rect 8352 16464 8358 16516
rect 11330 16464 11336 16516
rect 11388 16504 11394 16516
rect 11532 16504 11560 16603
rect 11701 16575 11759 16581
rect 11701 16541 11713 16575
rect 11747 16541 11759 16575
rect 11701 16535 11759 16541
rect 11977 16575 12035 16581
rect 11977 16541 11989 16575
rect 12023 16572 12035 16575
rect 12250 16572 12256 16584
rect 12023 16544 12256 16572
rect 12023 16541 12035 16544
rect 11977 16535 12035 16541
rect 11388 16476 11560 16504
rect 11716 16504 11744 16535
rect 12250 16532 12256 16544
rect 12308 16532 12314 16584
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16572 12403 16575
rect 12544 16572 12572 16612
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16640 13323 16643
rect 13372 16640 13400 16748
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 14642 16736 14648 16788
rect 14700 16776 14706 16788
rect 14737 16779 14795 16785
rect 14737 16776 14749 16779
rect 14700 16748 14749 16776
rect 14700 16736 14706 16748
rect 14737 16745 14749 16748
rect 14783 16745 14795 16779
rect 14737 16739 14795 16745
rect 15010 16736 15016 16788
rect 15068 16776 15074 16788
rect 19702 16776 19708 16788
rect 15068 16748 19708 16776
rect 15068 16736 15074 16748
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 20346 16776 20352 16788
rect 19904 16748 20352 16776
rect 18506 16708 18512 16720
rect 18467 16680 18512 16708
rect 18506 16668 18512 16680
rect 18564 16708 18570 16720
rect 19904 16708 19932 16748
rect 20162 16708 20168 16720
rect 18564 16680 19932 16708
rect 19996 16680 20168 16708
rect 18564 16668 18570 16680
rect 15105 16643 15163 16649
rect 13311 16612 13400 16640
rect 13740 16612 14412 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 12391 16544 12572 16572
rect 12621 16575 12679 16581
rect 12391 16541 12403 16544
rect 12345 16535 12403 16541
rect 12621 16541 12633 16575
rect 12667 16572 12679 16575
rect 12802 16572 12808 16584
rect 12667 16544 12808 16572
rect 12667 16541 12679 16544
rect 12621 16535 12679 16541
rect 12360 16504 12388 16535
rect 12802 16532 12808 16544
rect 12860 16532 12866 16584
rect 13354 16572 13360 16584
rect 13315 16544 13360 16572
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 13449 16575 13507 16581
rect 13449 16541 13461 16575
rect 13495 16541 13507 16575
rect 13449 16535 13507 16541
rect 11716 16476 12388 16504
rect 11388 16464 11394 16476
rect 12434 16464 12440 16516
rect 12492 16504 12498 16516
rect 12713 16507 12771 16513
rect 12713 16504 12725 16507
rect 12492 16476 12725 16504
rect 12492 16464 12498 16476
rect 12713 16473 12725 16476
rect 12759 16473 12771 16507
rect 12713 16467 12771 16473
rect 13262 16464 13268 16516
rect 13320 16504 13326 16516
rect 13464 16504 13492 16535
rect 13538 16532 13544 16584
rect 13596 16572 13602 16584
rect 13740 16572 13768 16612
rect 14384 16581 14412 16612
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 15470 16640 15476 16652
rect 15151 16612 15476 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 15470 16600 15476 16612
rect 15528 16640 15534 16652
rect 18230 16640 18236 16652
rect 15528 16612 18236 16640
rect 15528 16600 15534 16612
rect 18230 16600 18236 16612
rect 18288 16600 18294 16652
rect 13596 16544 13768 16572
rect 14369 16575 14427 16581
rect 13596 16532 13602 16544
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 14826 16572 14832 16584
rect 14787 16544 14832 16572
rect 14369 16535 14427 16541
rect 14826 16532 14832 16544
rect 14884 16532 14890 16584
rect 17310 16532 17316 16584
rect 17368 16572 17374 16584
rect 17589 16575 17647 16581
rect 17589 16572 17601 16575
rect 17368 16544 17601 16572
rect 17368 16532 17374 16544
rect 17589 16541 17601 16544
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 17770 16532 17776 16584
rect 17828 16572 17834 16584
rect 19996 16581 20024 16680
rect 20162 16668 20168 16680
rect 20220 16668 20226 16720
rect 20272 16649 20300 16748
rect 20346 16736 20352 16748
rect 20404 16736 20410 16788
rect 22646 16776 22652 16788
rect 22607 16748 22652 16776
rect 22646 16736 22652 16748
rect 22704 16736 22710 16788
rect 23385 16779 23443 16785
rect 23385 16745 23397 16779
rect 23431 16776 23443 16779
rect 23474 16776 23480 16788
rect 23431 16748 23480 16776
rect 23431 16745 23443 16748
rect 23385 16739 23443 16745
rect 23474 16736 23480 16748
rect 23532 16736 23538 16788
rect 23842 16776 23848 16788
rect 23803 16748 23848 16776
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 25133 16779 25191 16785
rect 25133 16745 25145 16779
rect 25179 16776 25191 16779
rect 25314 16776 25320 16788
rect 25179 16748 25320 16776
rect 25179 16745 25191 16748
rect 25133 16739 25191 16745
rect 25314 16736 25320 16748
rect 25372 16736 25378 16788
rect 20530 16668 20536 16720
rect 20588 16668 20594 16720
rect 20257 16643 20315 16649
rect 20257 16609 20269 16643
rect 20303 16609 20315 16643
rect 20257 16603 20315 16609
rect 20349 16643 20407 16649
rect 20349 16609 20361 16643
rect 20395 16640 20407 16643
rect 20548 16640 20576 16668
rect 20395 16612 20576 16640
rect 22281 16643 22339 16649
rect 20395 16609 20407 16612
rect 20349 16603 20407 16609
rect 22281 16609 22293 16643
rect 22327 16640 22339 16643
rect 22462 16640 22468 16652
rect 22327 16612 22468 16640
rect 22327 16609 22339 16612
rect 22281 16603 22339 16609
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17828 16544 18061 16572
rect 17828 16532 17834 16544
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 18325 16575 18383 16581
rect 18325 16541 18337 16575
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16541 20039 16575
rect 20162 16572 20168 16584
rect 20123 16544 20168 16572
rect 19981 16535 20039 16541
rect 13320 16476 13492 16504
rect 13320 16464 13326 16476
rect 14458 16436 14464 16448
rect 7432 16408 8248 16436
rect 14419 16408 14464 16436
rect 7432 16396 7438 16408
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 14844 16436 14872 16532
rect 15381 16507 15439 16513
rect 15381 16473 15393 16507
rect 15427 16504 15439 16507
rect 15654 16504 15660 16516
rect 15427 16476 15660 16504
rect 15427 16473 15439 16476
rect 15381 16467 15439 16473
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 16114 16464 16120 16516
rect 16172 16464 16178 16516
rect 18340 16504 18368 16535
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 20364 16504 20392 16603
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 22664 16640 22692 16736
rect 23584 16680 24992 16708
rect 22664 16612 23152 16640
rect 23124 16581 23152 16612
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16541 20591 16575
rect 20533 16535 20591 16541
rect 22833 16575 22891 16581
rect 22833 16541 22845 16575
rect 22879 16541 22891 16575
rect 22833 16535 22891 16541
rect 23109 16575 23167 16581
rect 23109 16541 23121 16575
rect 23155 16574 23167 16575
rect 23253 16575 23311 16581
rect 23155 16546 23189 16574
rect 23155 16541 23167 16546
rect 23109 16535 23167 16541
rect 23253 16541 23265 16575
rect 23299 16572 23311 16575
rect 23382 16572 23388 16584
rect 23299 16544 23388 16572
rect 23299 16541 23311 16544
rect 23253 16535 23311 16541
rect 20438 16504 20444 16516
rect 17420 16476 18368 16504
rect 18432 16476 20444 16504
rect 16666 16436 16672 16448
rect 14844 16408 16672 16436
rect 16666 16396 16672 16408
rect 16724 16436 16730 16448
rect 16853 16439 16911 16445
rect 16853 16436 16865 16439
rect 16724 16408 16865 16436
rect 16724 16396 16730 16408
rect 16853 16405 16865 16408
rect 16899 16405 16911 16439
rect 16853 16399 16911 16405
rect 17218 16396 17224 16448
rect 17276 16436 17282 16448
rect 17420 16445 17448 16476
rect 18432 16448 18460 16476
rect 20438 16464 20444 16476
rect 20496 16464 20502 16516
rect 17405 16439 17463 16445
rect 17405 16436 17417 16439
rect 17276 16408 17417 16436
rect 17276 16396 17282 16408
rect 17405 16405 17417 16408
rect 17451 16405 17463 16439
rect 17405 16399 17463 16405
rect 18233 16439 18291 16445
rect 18233 16405 18245 16439
rect 18279 16436 18291 16439
rect 18414 16436 18420 16448
rect 18279 16408 18420 16436
rect 18279 16405 18291 16408
rect 18233 16399 18291 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 19426 16396 19432 16448
rect 19484 16436 19490 16448
rect 20548 16436 20576 16535
rect 20717 16507 20775 16513
rect 20717 16473 20729 16507
rect 20763 16504 20775 16507
rect 22014 16507 22072 16513
rect 22014 16504 22026 16507
rect 20763 16476 22026 16504
rect 20763 16473 20775 16476
rect 20717 16467 20775 16473
rect 22014 16473 22026 16476
rect 22060 16473 22072 16507
rect 22014 16467 22072 16473
rect 20901 16439 20959 16445
rect 20901 16436 20913 16439
rect 19484 16408 20913 16436
rect 19484 16396 19490 16408
rect 20901 16405 20913 16408
rect 20947 16405 20959 16439
rect 22848 16436 22876 16535
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 23584 16581 23612 16680
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16541 23627 16575
rect 24029 16575 24087 16581
rect 24029 16574 24041 16575
rect 23952 16572 24041 16574
rect 23569 16535 23627 16541
rect 23768 16546 24041 16572
rect 23768 16544 23980 16546
rect 23017 16507 23075 16513
rect 23017 16473 23029 16507
rect 23063 16504 23075 16507
rect 23474 16504 23480 16516
rect 23063 16476 23480 16504
rect 23063 16473 23075 16476
rect 23017 16467 23075 16473
rect 23474 16464 23480 16476
rect 23532 16464 23538 16516
rect 23566 16436 23572 16448
rect 22848 16408 23572 16436
rect 20901 16399 20959 16405
rect 23566 16396 23572 16408
rect 23624 16396 23630 16448
rect 23768 16445 23796 16544
rect 24029 16541 24041 16546
rect 24075 16541 24087 16575
rect 24029 16535 24087 16541
rect 24302 16532 24308 16584
rect 24360 16572 24366 16584
rect 24964 16581 24992 16680
rect 24397 16575 24455 16581
rect 24397 16572 24409 16575
rect 24360 16544 24409 16572
rect 24360 16532 24366 16544
rect 24397 16541 24409 16544
rect 24443 16541 24455 16575
rect 24397 16535 24455 16541
rect 24949 16575 25007 16581
rect 24949 16541 24961 16575
rect 24995 16541 25007 16575
rect 24949 16535 25007 16541
rect 25685 16575 25743 16581
rect 25685 16541 25697 16575
rect 25731 16541 25743 16575
rect 25685 16535 25743 16541
rect 26053 16575 26111 16581
rect 26053 16541 26065 16575
rect 26099 16541 26111 16575
rect 26053 16535 26111 16541
rect 24486 16464 24492 16516
rect 24544 16504 24550 16516
rect 24964 16504 24992 16535
rect 24544 16476 24992 16504
rect 24544 16464 24550 16476
rect 23753 16439 23811 16445
rect 23753 16405 23765 16439
rect 23799 16405 23811 16439
rect 23753 16399 23811 16405
rect 24118 16396 24124 16448
rect 24176 16436 24182 16448
rect 24578 16436 24584 16448
rect 24176 16408 24221 16436
rect 24491 16408 24584 16436
rect 24176 16396 24182 16408
rect 24578 16396 24584 16408
rect 24636 16436 24642 16448
rect 25700 16436 25728 16535
rect 24636 16408 25728 16436
rect 25869 16439 25927 16445
rect 24636 16396 24642 16408
rect 25869 16405 25881 16439
rect 25915 16436 25927 16439
rect 26068 16436 26096 16535
rect 25915 16408 26096 16436
rect 25915 16405 25927 16408
rect 25869 16399 25927 16405
rect 26142 16396 26148 16448
rect 26200 16436 26206 16448
rect 26237 16439 26295 16445
rect 26237 16436 26249 16439
rect 26200 16408 26249 16436
rect 26200 16396 26206 16408
rect 26237 16405 26249 16408
rect 26283 16405 26295 16439
rect 26237 16399 26295 16405
rect 1104 16346 29440 16368
rect 1104 16294 10395 16346
rect 10447 16294 10459 16346
rect 10511 16294 10523 16346
rect 10575 16294 10587 16346
rect 10639 16294 10651 16346
rect 10703 16294 19840 16346
rect 19892 16294 19904 16346
rect 19956 16294 19968 16346
rect 20020 16294 20032 16346
rect 20084 16294 20096 16346
rect 20148 16294 29440 16346
rect 1104 16272 29440 16294
rect 3881 16235 3939 16241
rect 3881 16201 3893 16235
rect 3927 16232 3939 16235
rect 4522 16232 4528 16244
rect 3927 16204 4528 16232
rect 3927 16201 3939 16204
rect 3881 16195 3939 16201
rect 4522 16192 4528 16204
rect 4580 16192 4586 16244
rect 4617 16235 4675 16241
rect 4617 16201 4629 16235
rect 4663 16232 4675 16235
rect 4706 16232 4712 16244
rect 4663 16204 4712 16232
rect 4663 16201 4675 16204
rect 4617 16195 4675 16201
rect 4706 16192 4712 16204
rect 4764 16192 4770 16244
rect 5350 16192 5356 16244
rect 5408 16232 5414 16244
rect 5408 16204 5856 16232
rect 5408 16192 5414 16204
rect 2222 16124 2228 16176
rect 2280 16164 2286 16176
rect 3145 16167 3203 16173
rect 2280 16136 3096 16164
rect 2280 16124 2286 16136
rect 2130 16096 2136 16108
rect 2091 16068 2136 16096
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 2225 16031 2283 16037
rect 2225 15997 2237 16031
rect 2271 15997 2283 16031
rect 2225 15991 2283 15997
rect 2409 16031 2467 16037
rect 2409 15997 2421 16031
rect 2455 16028 2467 16031
rect 2498 16028 2504 16040
rect 2455 16000 2504 16028
rect 2455 15997 2467 16000
rect 2409 15991 2467 15997
rect 2240 15960 2268 15991
rect 2498 15988 2504 16000
rect 2556 15988 2562 16040
rect 2869 15963 2927 15969
rect 2869 15960 2881 15963
rect 2240 15932 2881 15960
rect 2869 15929 2881 15932
rect 2915 15960 2927 15963
rect 2958 15960 2964 15972
rect 2915 15932 2964 15960
rect 2915 15929 2927 15932
rect 2869 15923 2927 15929
rect 2958 15920 2964 15932
rect 3016 15920 3022 15972
rect 3068 15960 3096 16136
rect 3145 16133 3157 16167
rect 3191 16164 3203 16167
rect 3786 16164 3792 16176
rect 3191 16136 3792 16164
rect 3191 16133 3203 16136
rect 3145 16127 3203 16133
rect 3786 16124 3792 16136
rect 3844 16124 3850 16176
rect 3970 16124 3976 16176
rect 4028 16164 4034 16176
rect 4028 16136 5580 16164
rect 4028 16124 4034 16136
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16096 3479 16099
rect 3602 16096 3608 16108
rect 3467 16068 3608 16096
rect 3467 16065 3479 16068
rect 3421 16059 3479 16065
rect 3602 16056 3608 16068
rect 3660 16056 3666 16108
rect 3697 16099 3755 16105
rect 3697 16065 3709 16099
rect 3743 16096 3755 16099
rect 4154 16096 4160 16108
rect 3743 16068 4160 16096
rect 3743 16065 3755 16068
rect 3697 16059 3755 16065
rect 4154 16056 4160 16068
rect 4212 16056 4218 16108
rect 4767 16099 4825 16105
rect 4767 16065 4779 16099
rect 4813 16096 4825 16099
rect 4890 16096 4896 16108
rect 4813 16068 4896 16096
rect 4813 16065 4825 16068
rect 4767 16059 4825 16065
rect 4890 16056 4896 16068
rect 4948 16056 4954 16108
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16096 5135 16099
rect 5258 16096 5264 16108
rect 5123 16068 5264 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 5552 16105 5580 16136
rect 5828 16105 5856 16204
rect 7098 16192 7104 16244
rect 7156 16232 7162 16244
rect 7193 16235 7251 16241
rect 7193 16232 7205 16235
rect 7156 16204 7205 16232
rect 7156 16192 7162 16204
rect 7193 16201 7205 16204
rect 7239 16201 7251 16235
rect 8389 16235 8447 16241
rect 7193 16195 7251 16201
rect 7300 16204 8156 16232
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16065 5595 16099
rect 5537 16059 5595 16065
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 7300 16096 7328 16204
rect 7834 16164 7840 16176
rect 7795 16136 7840 16164
rect 7834 16124 7840 16136
rect 7892 16164 7898 16176
rect 8128 16164 8156 16204
rect 8389 16201 8401 16235
rect 8435 16232 8447 16235
rect 8435 16204 8616 16232
rect 8435 16201 8447 16204
rect 8389 16195 8447 16201
rect 8588 16173 8616 16204
rect 8662 16192 8668 16244
rect 8720 16232 8726 16244
rect 9401 16235 9459 16241
rect 9401 16232 9413 16235
rect 8720 16204 9413 16232
rect 8720 16192 8726 16204
rect 9401 16201 9413 16204
rect 9447 16232 9459 16235
rect 9490 16232 9496 16244
rect 9447 16204 9496 16232
rect 9447 16201 9459 16204
rect 9401 16195 9459 16201
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 16022 16192 16028 16244
rect 16080 16232 16086 16244
rect 16117 16235 16175 16241
rect 16117 16232 16129 16235
rect 16080 16204 16129 16232
rect 16080 16192 16086 16204
rect 16117 16201 16129 16204
rect 16163 16201 16175 16235
rect 16117 16195 16175 16201
rect 18141 16235 18199 16241
rect 18141 16201 18153 16235
rect 18187 16232 18199 16235
rect 18322 16232 18328 16244
rect 18187 16204 18328 16232
rect 18187 16201 18199 16204
rect 18141 16195 18199 16201
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 18874 16192 18880 16244
rect 18932 16232 18938 16244
rect 18969 16235 19027 16241
rect 18969 16232 18981 16235
rect 18932 16204 18981 16232
rect 18932 16192 18938 16204
rect 18969 16201 18981 16204
rect 19015 16201 19027 16235
rect 19426 16232 19432 16244
rect 19387 16204 19432 16232
rect 18969 16195 19027 16201
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 20530 16232 20536 16244
rect 20088 16204 20536 16232
rect 8573 16167 8631 16173
rect 7892 16136 8064 16164
rect 8128 16136 8524 16164
rect 7892 16124 7898 16136
rect 5859 16068 7328 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 7374 16056 7380 16108
rect 7432 16096 7438 16108
rect 8036 16105 8064 16136
rect 8021 16099 8079 16105
rect 7432 16068 7477 16096
rect 7432 16056 7438 16068
rect 8021 16065 8033 16099
rect 8067 16065 8079 16099
rect 8021 16059 8079 16065
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16096 8263 16099
rect 8386 16096 8392 16108
rect 8251 16068 8392 16096
rect 8251 16065 8263 16068
rect 8205 16059 8263 16065
rect 8386 16056 8392 16068
rect 8444 16056 8450 16108
rect 8496 16096 8524 16136
rect 8573 16133 8585 16167
rect 8619 16133 8631 16167
rect 14642 16164 14648 16176
rect 14306 16136 14648 16164
rect 8573 16127 8631 16133
rect 14642 16124 14648 16136
rect 14700 16124 14706 16176
rect 14734 16124 14740 16176
rect 14792 16164 14798 16176
rect 14792 16136 14837 16164
rect 14792 16124 14798 16136
rect 17586 16124 17592 16176
rect 17644 16164 17650 16176
rect 18509 16167 18567 16173
rect 18509 16164 18521 16167
rect 17644 16136 18521 16164
rect 17644 16124 17650 16136
rect 18509 16133 18521 16136
rect 18555 16133 18567 16167
rect 18509 16127 18567 16133
rect 18601 16167 18659 16173
rect 18601 16133 18613 16167
rect 18647 16164 18659 16167
rect 20088 16164 20116 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 21085 16235 21143 16241
rect 21085 16201 21097 16235
rect 21131 16232 21143 16235
rect 21174 16232 21180 16244
rect 21131 16204 21180 16232
rect 21131 16201 21143 16204
rect 21085 16195 21143 16201
rect 21100 16164 21128 16195
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 23198 16192 23204 16244
rect 23256 16232 23262 16244
rect 23382 16232 23388 16244
rect 23256 16204 23388 16232
rect 23256 16192 23262 16204
rect 23382 16192 23388 16204
rect 23440 16192 23446 16244
rect 23566 16192 23572 16244
rect 23624 16232 23630 16244
rect 24210 16232 24216 16244
rect 23624 16204 24216 16232
rect 23624 16192 23630 16204
rect 24210 16192 24216 16204
rect 24268 16192 24274 16244
rect 26142 16192 26148 16244
rect 26200 16192 26206 16244
rect 18647 16136 20116 16164
rect 20272 16136 21128 16164
rect 18647 16133 18659 16136
rect 18601 16127 18659 16133
rect 20272 16122 20300 16136
rect 23658 16124 23664 16176
rect 23716 16164 23722 16176
rect 24118 16164 24124 16176
rect 23716 16136 24124 16164
rect 23716 16124 23722 16136
rect 24118 16124 24124 16136
rect 24176 16124 24182 16176
rect 26160 16150 26188 16192
rect 8754 16096 8760 16108
rect 8496 16068 8760 16096
rect 8754 16056 8760 16068
rect 8812 16056 8818 16108
rect 8849 16099 8907 16105
rect 8849 16065 8861 16099
rect 8895 16065 8907 16099
rect 9490 16096 9496 16108
rect 9451 16068 9496 16096
rect 8849 16059 8907 16065
rect 3510 16028 3516 16040
rect 3471 16000 3516 16028
rect 3510 15988 3516 16000
rect 3568 15988 3574 16040
rect 5169 16031 5227 16037
rect 5169 15997 5181 16031
rect 5215 16028 5227 16031
rect 5442 16028 5448 16040
rect 5215 16000 5448 16028
rect 5215 15997 5227 16000
rect 5169 15991 5227 15997
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 5721 16031 5779 16037
rect 5721 15997 5733 16031
rect 5767 16028 5779 16031
rect 6086 16028 6092 16040
rect 5767 16000 6092 16028
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 6086 15988 6092 16000
rect 6144 15988 6150 16040
rect 6730 15988 6736 16040
rect 6788 16028 6794 16040
rect 8665 16031 8723 16037
rect 8665 16028 8677 16031
rect 6788 16000 8677 16028
rect 6788 15988 6794 16000
rect 8665 15997 8677 16000
rect 8711 15997 8723 16031
rect 8665 15991 8723 15997
rect 8864 15960 8892 16059
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16096 15439 16099
rect 15838 16096 15844 16108
rect 15427 16068 15844 16096
rect 15427 16065 15439 16068
rect 15381 16059 15439 16065
rect 15838 16056 15844 16068
rect 15896 16096 15902 16108
rect 15933 16099 15991 16105
rect 15933 16096 15945 16099
rect 15896 16068 15945 16096
rect 15896 16056 15902 16068
rect 15933 16065 15945 16068
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 17957 16099 18015 16105
rect 17957 16065 17969 16099
rect 18003 16096 18015 16099
rect 18046 16096 18052 16108
rect 18003 16068 18052 16096
rect 18003 16065 18015 16068
rect 17957 16059 18015 16065
rect 18046 16056 18052 16068
rect 18104 16096 18110 16108
rect 18414 16096 18420 16108
rect 18104 16068 18420 16096
rect 18104 16056 18110 16068
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 19242 16056 19248 16108
rect 19300 16096 19306 16108
rect 19337 16099 19395 16105
rect 19337 16096 19349 16099
rect 19300 16068 19349 16096
rect 19300 16056 19306 16068
rect 19337 16065 19349 16068
rect 19383 16065 19395 16099
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 19337 16059 19395 16065
rect 19444 16068 19993 16096
rect 10134 15988 10140 16040
rect 10192 16028 10198 16040
rect 14366 16028 14372 16040
rect 10192 16000 14372 16028
rect 10192 15988 10198 16000
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 16028 15071 16031
rect 15470 16028 15476 16040
rect 15059 16000 15476 16028
rect 15059 15997 15071 16000
rect 15013 15991 15071 15997
rect 15470 15988 15476 16000
rect 15528 15988 15534 16040
rect 18782 16028 18788 16040
rect 18743 16000 18788 16028
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 18874 15988 18880 16040
rect 18932 16028 18938 16040
rect 19444 16028 19472 16068
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 20164 16102 20222 16108
rect 20164 16068 20176 16102
rect 20210 16099 20222 16102
rect 20271 16099 20300 16122
rect 20438 16105 20444 16108
rect 20210 16094 20300 16099
rect 20395 16099 20444 16105
rect 20210 16071 20299 16094
rect 20210 16068 20222 16071
rect 20164 16062 20222 16068
rect 20395 16065 20407 16099
rect 20441 16065 20444 16099
rect 20395 16059 20444 16065
rect 20438 16056 20444 16059
rect 20496 16056 20502 16108
rect 20530 16056 20536 16108
rect 20588 16096 20594 16108
rect 20588 16068 20633 16096
rect 20588 16056 20594 16068
rect 24394 16056 24400 16108
rect 24452 16096 24458 16108
rect 24949 16099 25007 16105
rect 24949 16096 24961 16099
rect 24452 16068 24961 16096
rect 24452 16056 24458 16068
rect 24949 16065 24961 16068
rect 24995 16065 25007 16099
rect 24949 16059 25007 16065
rect 18932 16000 19472 16028
rect 19613 16031 19671 16037
rect 18932 15988 18938 16000
rect 19613 15997 19625 16031
rect 19659 15997 19671 16031
rect 19613 15991 19671 15997
rect 20257 16031 20315 16037
rect 20257 15997 20269 16031
rect 20303 15997 20315 16031
rect 25222 16028 25228 16040
rect 25183 16000 25228 16028
rect 20257 15991 20315 15997
rect 3068 15932 3464 15960
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 2314 15852 2320 15904
rect 2372 15892 2378 15904
rect 3436 15901 3464 15932
rect 7668 15932 8892 15960
rect 9033 15963 9091 15969
rect 7668 15904 7696 15932
rect 9033 15929 9045 15963
rect 9079 15960 9091 15963
rect 13354 15960 13360 15972
rect 9079 15932 13360 15960
rect 9079 15929 9091 15932
rect 9033 15923 9091 15929
rect 13354 15920 13360 15932
rect 13412 15920 13418 15972
rect 2685 15895 2743 15901
rect 2685 15892 2697 15895
rect 2372 15864 2697 15892
rect 2372 15852 2378 15864
rect 2685 15861 2697 15864
rect 2731 15861 2743 15895
rect 2685 15855 2743 15861
rect 3421 15895 3479 15901
rect 3421 15861 3433 15895
rect 3467 15861 3479 15895
rect 3421 15855 3479 15861
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 5353 15895 5411 15901
rect 5353 15892 5365 15895
rect 3936 15864 5365 15892
rect 3936 15852 3942 15864
rect 5353 15861 5365 15864
rect 5399 15861 5411 15895
rect 5353 15855 5411 15861
rect 6546 15852 6552 15904
rect 6604 15892 6610 15904
rect 6641 15895 6699 15901
rect 6641 15892 6653 15895
rect 6604 15864 6653 15892
rect 6604 15852 6610 15864
rect 6641 15861 6653 15864
rect 6687 15861 6699 15895
rect 7650 15892 7656 15904
rect 7611 15864 7656 15892
rect 6641 15855 6699 15861
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 7742 15852 7748 15904
rect 7800 15892 7806 15904
rect 8018 15892 8024 15904
rect 7800 15864 8024 15892
rect 7800 15852 7806 15864
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 8205 15895 8263 15901
rect 8205 15861 8217 15895
rect 8251 15892 8263 15895
rect 8478 15892 8484 15904
rect 8251 15864 8484 15892
rect 8251 15861 8263 15864
rect 8205 15855 8263 15861
rect 8478 15852 8484 15864
rect 8536 15852 8542 15904
rect 8754 15892 8760 15904
rect 8715 15864 8760 15892
rect 8754 15852 8760 15864
rect 8812 15852 8818 15904
rect 9674 15892 9680 15904
rect 9635 15864 9680 15892
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 13262 15892 13268 15904
rect 13223 15864 13268 15892
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 14918 15852 14924 15904
rect 14976 15892 14982 15904
rect 15197 15895 15255 15901
rect 15197 15892 15209 15895
rect 14976 15864 15209 15892
rect 14976 15852 14982 15864
rect 15197 15861 15209 15864
rect 15243 15861 15255 15895
rect 15197 15855 15255 15861
rect 17773 15895 17831 15901
rect 17773 15861 17785 15895
rect 17819 15892 17831 15895
rect 17954 15892 17960 15904
rect 17819 15864 17960 15892
rect 17819 15861 17831 15864
rect 17773 15855 17831 15861
rect 17954 15852 17960 15864
rect 18012 15852 18018 15904
rect 18782 15852 18788 15904
rect 18840 15892 18846 15904
rect 19150 15892 19156 15904
rect 18840 15864 19156 15892
rect 18840 15852 18846 15864
rect 19150 15852 19156 15864
rect 19208 15892 19214 15904
rect 19628 15892 19656 15991
rect 19208 15864 19656 15892
rect 20271 15892 20299 15991
rect 25222 15988 25228 16000
rect 25280 15988 25286 16040
rect 20438 15920 20444 15972
rect 20496 15960 20502 15972
rect 20809 15963 20867 15969
rect 20809 15960 20821 15963
rect 20496 15932 20821 15960
rect 20496 15920 20502 15932
rect 20809 15929 20821 15932
rect 20855 15929 20867 15963
rect 20809 15923 20867 15929
rect 20346 15892 20352 15904
rect 20271 15864 20352 15892
rect 19208 15852 19214 15864
rect 20346 15852 20352 15864
rect 20404 15852 20410 15904
rect 20622 15892 20628 15904
rect 20583 15864 20628 15892
rect 20622 15852 20628 15864
rect 20680 15852 20686 15904
rect 26697 15895 26755 15901
rect 26697 15861 26709 15895
rect 26743 15892 26755 15895
rect 26786 15892 26792 15904
rect 26743 15864 26792 15892
rect 26743 15861 26755 15864
rect 26697 15855 26755 15861
rect 26786 15852 26792 15864
rect 26844 15852 26850 15904
rect 1104 15802 29440 15824
rect 1104 15750 5672 15802
rect 5724 15750 5736 15802
rect 5788 15750 5800 15802
rect 5852 15750 5864 15802
rect 5916 15750 5928 15802
rect 5980 15750 15118 15802
rect 15170 15750 15182 15802
rect 15234 15750 15246 15802
rect 15298 15750 15310 15802
rect 15362 15750 15374 15802
rect 15426 15750 24563 15802
rect 24615 15750 24627 15802
rect 24679 15750 24691 15802
rect 24743 15750 24755 15802
rect 24807 15750 24819 15802
rect 24871 15750 29440 15802
rect 1104 15728 29440 15750
rect 2130 15688 2136 15700
rect 2091 15660 2136 15688
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 2958 15688 2964 15700
rect 2919 15660 2964 15688
rect 2958 15648 2964 15660
rect 3016 15648 3022 15700
rect 3145 15691 3203 15697
rect 3145 15657 3157 15691
rect 3191 15688 3203 15691
rect 3510 15688 3516 15700
rect 3191 15660 3516 15688
rect 3191 15657 3203 15660
rect 3145 15651 3203 15657
rect 3510 15648 3516 15660
rect 3568 15648 3574 15700
rect 5353 15691 5411 15697
rect 5353 15688 5365 15691
rect 3988 15660 5365 15688
rect 1578 15580 1584 15632
rect 1636 15620 1642 15632
rect 3988 15620 4016 15660
rect 5353 15657 5365 15660
rect 5399 15688 5411 15691
rect 6546 15688 6552 15700
rect 5399 15660 6552 15688
rect 5399 15657 5411 15660
rect 5353 15651 5411 15657
rect 6546 15648 6552 15660
rect 6604 15688 6610 15700
rect 8294 15688 8300 15700
rect 6604 15660 6868 15688
rect 6604 15648 6610 15660
rect 4154 15620 4160 15632
rect 1636 15592 4016 15620
rect 4115 15592 4160 15620
rect 1636 15580 1642 15592
rect 4154 15580 4160 15592
rect 4212 15580 4218 15632
rect 3878 15552 3884 15564
rect 3839 15524 3884 15552
rect 3878 15512 3884 15524
rect 3936 15512 3942 15564
rect 2314 15484 2320 15496
rect 2275 15456 2320 15484
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 2774 15444 2780 15496
rect 2832 15484 2838 15496
rect 2961 15487 3019 15493
rect 2832 15456 2877 15484
rect 2832 15444 2838 15456
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 4246 15484 4252 15496
rect 3007 15456 4252 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 6730 15484 6736 15496
rect 6691 15456 6736 15484
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 6840 15484 6868 15660
rect 7852 15660 8300 15688
rect 7098 15580 7104 15632
rect 7156 15580 7162 15632
rect 7116 15552 7144 15580
rect 7282 15552 7288 15564
rect 7116 15524 7288 15552
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 7009 15487 7067 15493
rect 7009 15484 7021 15487
rect 6840 15456 7021 15484
rect 7009 15453 7021 15456
rect 7055 15453 7067 15487
rect 7009 15447 7067 15453
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 7193 15487 7251 15493
rect 7193 15484 7205 15487
rect 7156 15456 7205 15484
rect 7156 15444 7162 15456
rect 7193 15453 7205 15456
rect 7239 15453 7251 15487
rect 7193 15447 7251 15453
rect 7374 15444 7380 15496
rect 7432 15484 7438 15496
rect 7561 15487 7619 15493
rect 7432 15456 7477 15484
rect 7432 15444 7438 15456
rect 7561 15453 7573 15487
rect 7607 15453 7619 15487
rect 7742 15484 7748 15496
rect 7703 15456 7748 15484
rect 7561 15447 7619 15453
rect 6488 15419 6546 15425
rect 6488 15385 6500 15419
rect 6534 15416 6546 15419
rect 6825 15419 6883 15425
rect 6825 15416 6837 15419
rect 6534 15388 6837 15416
rect 6534 15385 6546 15388
rect 6488 15379 6546 15385
rect 6825 15385 6837 15388
rect 6871 15385 6883 15419
rect 6825 15379 6883 15385
rect 7466 15376 7472 15428
rect 7524 15416 7530 15428
rect 7576 15416 7604 15447
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 7852 15484 7880 15660
rect 8294 15648 8300 15660
rect 8352 15688 8358 15700
rect 8389 15691 8447 15697
rect 8389 15688 8401 15691
rect 8352 15660 8401 15688
rect 8352 15648 8358 15660
rect 8389 15657 8401 15660
rect 8435 15657 8447 15691
rect 8389 15651 8447 15657
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 10781 15691 10839 15697
rect 10781 15688 10793 15691
rect 10100 15660 10793 15688
rect 10100 15648 10106 15660
rect 10781 15657 10793 15660
rect 10827 15688 10839 15691
rect 10962 15688 10968 15700
rect 10827 15660 10968 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 11606 15688 11612 15700
rect 11112 15660 11612 15688
rect 11112 15648 11118 15660
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 12618 15648 12624 15700
rect 12676 15688 12682 15700
rect 12713 15691 12771 15697
rect 12713 15688 12725 15691
rect 12676 15660 12725 15688
rect 12676 15648 12682 15660
rect 12713 15657 12725 15660
rect 12759 15657 12771 15691
rect 14642 15688 14648 15700
rect 14603 15660 14648 15688
rect 12713 15651 12771 15657
rect 14642 15648 14648 15660
rect 14700 15648 14706 15700
rect 17497 15691 17555 15697
rect 17497 15657 17509 15691
rect 17543 15688 17555 15691
rect 17586 15688 17592 15700
rect 17543 15660 17592 15688
rect 17543 15657 17555 15660
rect 17497 15651 17555 15657
rect 17586 15648 17592 15660
rect 17644 15648 17650 15700
rect 17862 15648 17868 15700
rect 17920 15688 17926 15700
rect 18509 15691 18567 15697
rect 18509 15688 18521 15691
rect 17920 15660 18521 15688
rect 17920 15648 17926 15660
rect 18509 15657 18521 15660
rect 18555 15688 18567 15691
rect 18874 15688 18880 15700
rect 18555 15660 18880 15688
rect 18555 15657 18567 15660
rect 18509 15651 18567 15657
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 20257 15691 20315 15697
rect 20257 15657 20269 15691
rect 20303 15688 20315 15691
rect 20530 15688 20536 15700
rect 20303 15660 20536 15688
rect 20303 15657 20315 15660
rect 20257 15651 20315 15657
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 24486 15648 24492 15700
rect 24544 15688 24550 15700
rect 24581 15691 24639 15697
rect 24581 15688 24593 15691
rect 24544 15660 24593 15688
rect 24544 15648 24550 15660
rect 24581 15657 24593 15660
rect 24627 15657 24639 15691
rect 24581 15651 24639 15657
rect 25222 15648 25228 15700
rect 25280 15688 25286 15700
rect 25317 15691 25375 15697
rect 25317 15688 25329 15691
rect 25280 15660 25329 15688
rect 25280 15648 25286 15660
rect 25317 15657 25329 15660
rect 25363 15657 25375 15691
rect 25317 15651 25375 15657
rect 8018 15580 8024 15632
rect 8076 15620 8082 15632
rect 8941 15623 8999 15629
rect 8941 15620 8953 15623
rect 8076 15592 8953 15620
rect 8076 15580 8082 15592
rect 8941 15589 8953 15592
rect 8987 15589 8999 15623
rect 24026 15620 24032 15632
rect 8941 15583 8999 15589
rect 23768 15592 24032 15620
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 9033 15555 9091 15561
rect 8168 15524 8248 15552
rect 8168 15512 8174 15524
rect 7920 15487 7978 15493
rect 7920 15484 7932 15487
rect 7852 15456 7932 15484
rect 7920 15453 7932 15456
rect 7966 15453 7978 15487
rect 7920 15447 7978 15453
rect 8018 15444 8024 15496
rect 8076 15484 8082 15496
rect 8220 15493 8248 15524
rect 9033 15521 9045 15555
rect 9079 15552 9091 15555
rect 10962 15552 10968 15564
rect 9079 15524 10968 15552
rect 9079 15521 9091 15524
rect 9033 15515 9091 15521
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 11241 15555 11299 15561
rect 11241 15521 11253 15555
rect 11287 15552 11299 15555
rect 11330 15552 11336 15564
rect 11287 15524 11336 15552
rect 11287 15521 11299 15524
rect 11241 15515 11299 15521
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 17126 15512 17132 15564
rect 17184 15552 17190 15564
rect 17957 15555 18015 15561
rect 17184 15524 17816 15552
rect 17184 15512 17190 15524
rect 8205 15487 8263 15493
rect 8076 15456 8121 15484
rect 8076 15444 8082 15456
rect 8205 15453 8217 15487
rect 8251 15453 8263 15487
rect 8205 15447 8263 15453
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 8573 15487 8631 15493
rect 8352 15456 8397 15484
rect 8352 15444 8358 15456
rect 8573 15453 8585 15487
rect 8619 15484 8631 15487
rect 8662 15484 8668 15496
rect 8619 15456 8668 15484
rect 8619 15453 8631 15456
rect 8573 15447 8631 15453
rect 8662 15444 8668 15456
rect 8720 15444 8726 15496
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15484 14887 15487
rect 14918 15484 14924 15496
rect 14875 15456 14924 15484
rect 14875 15453 14887 15456
rect 14829 15447 14887 15453
rect 14918 15444 14924 15456
rect 14976 15444 14982 15496
rect 16114 15484 16120 15496
rect 16075 15456 16120 15484
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 17681 15487 17739 15493
rect 17681 15453 17693 15487
rect 17727 15453 17739 15487
rect 17788 15484 17816 15524
rect 17957 15521 17969 15555
rect 18003 15552 18015 15555
rect 18138 15552 18144 15564
rect 18003 15524 18144 15552
rect 18003 15521 18015 15524
rect 17957 15515 18015 15521
rect 18138 15512 18144 15524
rect 18196 15512 18202 15564
rect 19242 15552 19248 15564
rect 18248 15524 19248 15552
rect 18248 15493 18276 15524
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 17846 15487 17904 15493
rect 17846 15484 17858 15487
rect 17788 15456 17858 15484
rect 17681 15447 17739 15453
rect 17846 15453 17858 15456
rect 17892 15453 17904 15487
rect 17846 15447 17904 15453
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15453 18107 15487
rect 18049 15447 18107 15453
rect 18233 15487 18291 15493
rect 18233 15453 18245 15487
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 7524 15388 7604 15416
rect 9309 15419 9367 15425
rect 7524 15376 7530 15388
rect 9309 15385 9321 15419
rect 9355 15416 9367 15419
rect 9398 15416 9404 15428
rect 9355 15388 9404 15416
rect 9355 15385 9367 15388
rect 9309 15379 9367 15385
rect 9398 15376 9404 15388
rect 9456 15376 9462 15428
rect 10318 15376 10324 15428
rect 10376 15376 10382 15428
rect 11698 15376 11704 15428
rect 11756 15376 11762 15428
rect 12526 15376 12532 15428
rect 12584 15416 12590 15428
rect 13357 15419 13415 15425
rect 13357 15416 13369 15419
rect 12584 15388 13369 15416
rect 12584 15376 12590 15388
rect 13357 15385 13369 15388
rect 13403 15385 13415 15419
rect 13357 15379 13415 15385
rect 16384 15419 16442 15425
rect 16384 15385 16396 15419
rect 16430 15416 16442 15419
rect 17310 15416 17316 15428
rect 16430 15388 17316 15416
rect 16430 15385 16442 15388
rect 16384 15379 16442 15385
rect 17310 15376 17316 15388
rect 17368 15376 17374 15428
rect 17696 15416 17724 15447
rect 17954 15416 17960 15428
rect 17696 15388 17960 15416
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 18064 15416 18092 15447
rect 18414 15444 18420 15496
rect 18472 15484 18478 15496
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18472 15456 18705 15484
rect 18472 15444 18478 15456
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 18693 15447 18751 15453
rect 20622 15444 20628 15496
rect 20680 15484 20686 15496
rect 21370 15487 21428 15493
rect 21370 15484 21382 15487
rect 20680 15456 21382 15484
rect 20680 15444 20686 15456
rect 21370 15453 21382 15456
rect 21416 15453 21428 15487
rect 21634 15484 21640 15496
rect 21595 15456 21640 15484
rect 21370 15447 21428 15453
rect 21634 15444 21640 15456
rect 21692 15484 21698 15496
rect 21729 15487 21787 15493
rect 21729 15484 21741 15487
rect 21692 15456 21741 15484
rect 21692 15444 21698 15456
rect 21729 15453 21741 15456
rect 21775 15453 21787 15487
rect 23566 15484 23572 15496
rect 23527 15456 23572 15484
rect 21729 15447 21787 15453
rect 23566 15444 23572 15456
rect 23624 15444 23630 15496
rect 23768 15493 23796 15592
rect 24026 15580 24032 15592
rect 24084 15580 24090 15632
rect 24121 15623 24179 15629
rect 24121 15589 24133 15623
rect 24167 15620 24179 15623
rect 25038 15620 25044 15632
rect 24167 15592 25044 15620
rect 24167 15589 24179 15592
rect 24121 15583 24179 15589
rect 25038 15580 25044 15592
rect 25096 15580 25102 15632
rect 26510 15552 26516 15564
rect 23860 15524 26516 15552
rect 23860 15493 23888 15524
rect 26510 15512 26516 15524
rect 26568 15512 26574 15564
rect 23753 15487 23811 15493
rect 23753 15453 23765 15487
rect 23799 15453 23811 15487
rect 23753 15447 23811 15453
rect 23845 15487 23903 15493
rect 23845 15453 23857 15487
rect 23891 15453 23903 15487
rect 23845 15447 23903 15453
rect 23989 15487 24047 15493
rect 23989 15453 24001 15487
rect 24035 15484 24047 15487
rect 24035 15456 24164 15484
rect 24035 15453 24047 15456
rect 23989 15447 24047 15453
rect 18598 15416 18604 15428
rect 18064 15388 18604 15416
rect 18598 15376 18604 15388
rect 18656 15376 18662 15428
rect 22002 15425 22008 15428
rect 21996 15416 22008 15425
rect 21963 15388 22008 15416
rect 21996 15379 22008 15388
rect 22002 15376 22008 15379
rect 22060 15376 22066 15428
rect 23198 15376 23204 15428
rect 23256 15416 23262 15428
rect 24136 15416 24164 15456
rect 24302 15444 24308 15496
rect 24360 15484 24366 15496
rect 24397 15487 24455 15493
rect 24397 15484 24409 15487
rect 24360 15456 24409 15484
rect 24360 15444 24366 15456
rect 24397 15453 24409 15456
rect 24443 15453 24455 15487
rect 24397 15447 24455 15453
rect 24673 15487 24731 15493
rect 24673 15453 24685 15487
rect 24719 15484 24731 15487
rect 24765 15487 24823 15493
rect 24765 15484 24777 15487
rect 24719 15456 24777 15484
rect 24719 15453 24731 15456
rect 24673 15447 24731 15453
rect 24765 15453 24777 15456
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 24854 15444 24860 15496
rect 24912 15484 24918 15496
rect 25138 15487 25196 15493
rect 25138 15484 25150 15487
rect 24912 15456 25150 15484
rect 24912 15444 24918 15456
rect 25138 15453 25150 15456
rect 25184 15453 25196 15487
rect 26786 15484 26792 15496
rect 25138 15447 25196 15453
rect 25516 15456 26792 15484
rect 24872 15416 24900 15444
rect 23256 15388 24900 15416
rect 24949 15419 25007 15425
rect 23256 15376 23262 15388
rect 24949 15385 24961 15419
rect 24995 15385 25007 15419
rect 24949 15379 25007 15385
rect 25041 15419 25099 15425
rect 25041 15385 25053 15419
rect 25087 15416 25099 15419
rect 25516 15416 25544 15456
rect 26786 15444 26792 15456
rect 26844 15444 26850 15496
rect 25087 15388 25544 15416
rect 25087 15385 25099 15388
rect 25041 15379 25099 15385
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15348 4399 15351
rect 4982 15348 4988 15360
rect 4387 15320 4988 15348
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 4982 15308 4988 15320
rect 5040 15308 5046 15360
rect 8570 15308 8576 15360
rect 8628 15348 8634 15360
rect 8665 15351 8723 15357
rect 8665 15348 8677 15351
rect 8628 15320 8677 15348
rect 8628 15308 8634 15320
rect 8665 15317 8677 15320
rect 8711 15317 8723 15351
rect 8665 15311 8723 15317
rect 8941 15351 8999 15357
rect 8941 15317 8953 15351
rect 8987 15348 8999 15351
rect 17126 15348 17132 15360
rect 8987 15320 17132 15348
rect 8987 15317 8999 15320
rect 8941 15311 8999 15317
rect 17126 15308 17132 15320
rect 17184 15308 17190 15360
rect 18322 15348 18328 15360
rect 18283 15320 18328 15348
rect 18322 15308 18328 15320
rect 18380 15308 18386 15360
rect 22278 15308 22284 15360
rect 22336 15348 22342 15360
rect 23109 15351 23167 15357
rect 23109 15348 23121 15351
rect 22336 15320 23121 15348
rect 22336 15308 22342 15320
rect 23109 15317 23121 15320
rect 23155 15317 23167 15351
rect 23109 15311 23167 15317
rect 24210 15308 24216 15360
rect 24268 15348 24274 15360
rect 24673 15351 24731 15357
rect 24673 15348 24685 15351
rect 24268 15320 24685 15348
rect 24268 15308 24274 15320
rect 24673 15317 24685 15320
rect 24719 15317 24731 15351
rect 24964 15348 24992 15379
rect 25130 15348 25136 15360
rect 24964 15320 25136 15348
rect 24673 15311 24731 15317
rect 25130 15308 25136 15320
rect 25188 15348 25194 15360
rect 25406 15348 25412 15360
rect 25188 15320 25412 15348
rect 25188 15308 25194 15320
rect 25406 15308 25412 15320
rect 25464 15348 25470 15360
rect 25501 15351 25559 15357
rect 25501 15348 25513 15351
rect 25464 15320 25513 15348
rect 25464 15308 25470 15320
rect 25501 15317 25513 15320
rect 25547 15317 25559 15351
rect 25501 15311 25559 15317
rect 1104 15258 29440 15280
rect 1104 15206 10395 15258
rect 10447 15206 10459 15258
rect 10511 15206 10523 15258
rect 10575 15206 10587 15258
rect 10639 15206 10651 15258
rect 10703 15206 19840 15258
rect 19892 15206 19904 15258
rect 19956 15206 19968 15258
rect 20020 15206 20032 15258
rect 20084 15206 20096 15258
rect 20148 15206 29440 15258
rect 1104 15184 29440 15206
rect 2777 15147 2835 15153
rect 2777 15113 2789 15147
rect 2823 15144 2835 15147
rect 3234 15144 3240 15156
rect 2823 15116 3240 15144
rect 2823 15113 2835 15116
rect 2777 15107 2835 15113
rect 3234 15104 3240 15116
rect 3292 15144 3298 15156
rect 3329 15147 3387 15153
rect 3329 15144 3341 15147
rect 3292 15116 3341 15144
rect 3292 15104 3298 15116
rect 3329 15113 3341 15116
rect 3375 15113 3387 15147
rect 3329 15107 3387 15113
rect 4341 15147 4399 15153
rect 4341 15113 4353 15147
rect 4387 15144 4399 15147
rect 4801 15147 4859 15153
rect 4801 15144 4813 15147
rect 4387 15116 4813 15144
rect 4387 15113 4399 15116
rect 4341 15107 4399 15113
rect 4801 15113 4813 15116
rect 4847 15113 4859 15147
rect 4801 15107 4859 15113
rect 6457 15147 6515 15153
rect 6457 15113 6469 15147
rect 6503 15144 6515 15147
rect 7374 15144 7380 15156
rect 6503 15116 7380 15144
rect 6503 15113 6515 15116
rect 6457 15107 6515 15113
rect 7374 15104 7380 15116
rect 7432 15104 7438 15156
rect 7745 15147 7803 15153
rect 7745 15113 7757 15147
rect 7791 15144 7803 15147
rect 7834 15144 7840 15156
rect 7791 15116 7840 15144
rect 7791 15113 7803 15116
rect 7745 15107 7803 15113
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 8018 15104 8024 15156
rect 8076 15104 8082 15156
rect 8205 15147 8263 15153
rect 8205 15113 8217 15147
rect 8251 15144 8263 15147
rect 8294 15144 8300 15156
rect 8251 15116 8300 15144
rect 8251 15113 8263 15116
rect 8205 15107 8263 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 10597 15147 10655 15153
rect 10597 15144 10609 15147
rect 10376 15116 10609 15144
rect 10376 15104 10382 15116
rect 10597 15113 10609 15116
rect 10643 15113 10655 15147
rect 11698 15144 11704 15156
rect 11659 15116 11704 15144
rect 10597 15107 10655 15113
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 16393 15147 16451 15153
rect 16393 15144 16405 15147
rect 12676 15116 16405 15144
rect 12676 15104 12682 15116
rect 1664 15079 1722 15085
rect 1664 15045 1676 15079
rect 1710 15076 1722 15079
rect 1762 15076 1768 15088
rect 1710 15048 1768 15076
rect 1710 15045 1722 15048
rect 1664 15039 1722 15045
rect 1762 15036 1768 15048
rect 1820 15036 1826 15088
rect 4154 15036 4160 15088
rect 4212 15076 4218 15088
rect 4433 15079 4491 15085
rect 4433 15076 4445 15079
rect 4212 15048 4445 15076
rect 4212 15036 4218 15048
rect 4433 15045 4445 15048
rect 4479 15045 4491 15079
rect 4433 15039 4491 15045
rect 6914 15036 6920 15088
rect 6972 15076 6978 15088
rect 7101 15079 7159 15085
rect 7101 15076 7113 15079
rect 6972 15048 7113 15076
rect 6972 15036 6978 15048
rect 7101 15045 7113 15048
rect 7147 15045 7159 15079
rect 7101 15039 7159 15045
rect 7193 15079 7251 15085
rect 7193 15045 7205 15079
rect 7239 15076 7251 15079
rect 8036 15076 8064 15104
rect 8312 15076 8340 15104
rect 13262 15076 13268 15088
rect 7239 15048 8248 15076
rect 8312 15048 8800 15076
rect 7239 15045 7251 15048
rect 7193 15039 7251 15045
rect 4982 15008 4988 15020
rect 4943 14980 4988 15008
rect 4982 14968 4988 14980
rect 5040 14968 5046 15020
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 15008 6607 15011
rect 7834 15008 7840 15020
rect 6595 14980 6776 15008
rect 7795 14980 7840 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 1394 14940 1400 14952
rect 1355 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14900 1458 14952
rect 3418 14940 3424 14952
rect 3379 14912 3424 14940
rect 3418 14900 3424 14912
rect 3476 14900 3482 14952
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 2958 14872 2964 14884
rect 2919 14844 2964 14872
rect 2958 14832 2964 14844
rect 3016 14832 3022 14884
rect 3620 14872 3648 14903
rect 4430 14900 4436 14952
rect 4488 14940 4494 14952
rect 4525 14943 4583 14949
rect 4525 14940 4537 14943
rect 4488 14912 4537 14940
rect 4488 14900 4494 14912
rect 4525 14909 4537 14912
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 4614 14872 4620 14884
rect 3620 14844 4620 14872
rect 4614 14832 4620 14844
rect 4672 14832 4678 14884
rect 3970 14804 3976 14816
rect 3931 14776 3976 14804
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 6748 14813 6776 14980
rect 7834 14968 7840 14980
rect 7892 14968 7898 15020
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 14977 8079 15011
rect 8220 15008 8248 15048
rect 8772 15017 8800 15048
rect 9692 15048 13268 15076
rect 8665 15011 8723 15017
rect 8665 15008 8677 15011
rect 8220 14980 8677 15008
rect 8021 14971 8079 14977
rect 8665 14977 8677 14980
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 14977 8815 15011
rect 8757 14971 8815 14977
rect 9033 15011 9091 15017
rect 9033 14977 9045 15011
rect 9079 15008 9091 15011
rect 9306 15008 9312 15020
rect 9079 14980 9312 15008
rect 9079 14977 9091 14980
rect 9033 14971 9091 14977
rect 7282 14900 7288 14952
rect 7340 14940 7346 14952
rect 7340 14912 7385 14940
rect 7340 14900 7346 14912
rect 8036 14872 8064 14971
rect 8680 14940 8708 14971
rect 9306 14968 9312 14980
rect 9364 15008 9370 15020
rect 9692 15017 9720 15048
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 9364 14980 9505 15008
rect 9364 14968 9370 14980
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 14977 9735 15011
rect 10042 15008 10048 15020
rect 10003 14980 10048 15008
rect 9677 14971 9735 14977
rect 10042 14968 10048 14980
rect 10100 14968 10106 15020
rect 10778 15008 10784 15020
rect 10739 14980 10784 15008
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 11057 15011 11115 15017
rect 11057 15008 11069 15011
rect 10928 14980 11069 15008
rect 10928 14968 10934 14980
rect 11057 14977 11069 14980
rect 11103 14977 11115 15011
rect 11517 15011 11575 15017
rect 11517 15008 11529 15011
rect 11057 14971 11115 14977
rect 11256 14980 11529 15008
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 8680 14912 9229 14940
rect 9217 14909 9229 14912
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 8662 14872 8668 14884
rect 8036 14844 8668 14872
rect 8662 14832 8668 14844
rect 8720 14832 8726 14884
rect 8941 14875 8999 14881
rect 8941 14841 8953 14875
rect 8987 14872 8999 14875
rect 9490 14872 9496 14884
rect 8987 14844 9496 14872
rect 8987 14841 8999 14844
rect 8941 14835 8999 14841
rect 9490 14832 9496 14844
rect 9548 14872 9554 14884
rect 11256 14881 11284 14980
rect 11517 14977 11529 14980
rect 11563 14977 11575 15011
rect 11517 14971 11575 14977
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12437 15011 12495 15017
rect 12437 15008 12449 15011
rect 12032 14980 12449 15008
rect 12032 14968 12038 14980
rect 12437 14977 12449 14980
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12526 14968 12532 15020
rect 12584 15008 12590 15020
rect 12621 15011 12679 15017
rect 12621 15008 12633 15011
rect 12584 14980 12633 15008
rect 12584 14968 12590 14980
rect 12621 14977 12633 14980
rect 12667 14977 12679 15011
rect 12621 14971 12679 14977
rect 12713 15011 12771 15017
rect 12713 14977 12725 15011
rect 12759 14977 12771 15011
rect 12713 14971 12771 14977
rect 12728 14940 12756 14971
rect 12802 14968 12808 15020
rect 12860 15017 12866 15020
rect 12860 15008 12868 15017
rect 12860 14980 12905 15008
rect 12860 14971 12868 14980
rect 12860 14968 12866 14971
rect 12406 14912 12756 14940
rect 9677 14875 9735 14881
rect 9677 14872 9689 14875
rect 9548 14844 9689 14872
rect 9548 14832 9554 14844
rect 9677 14841 9689 14844
rect 9723 14841 9735 14875
rect 9677 14835 9735 14841
rect 11241 14875 11299 14881
rect 11241 14841 11253 14875
rect 11287 14841 11299 14875
rect 12406 14872 12434 14912
rect 11241 14835 11299 14841
rect 11348 14844 12434 14872
rect 6733 14807 6791 14813
rect 6733 14773 6745 14807
rect 6779 14804 6791 14807
rect 7098 14804 7104 14816
rect 6779 14776 7104 14804
rect 6779 14773 6791 14776
rect 6733 14767 6791 14773
rect 7098 14764 7104 14776
rect 7156 14764 7162 14816
rect 8294 14764 8300 14816
rect 8352 14804 8358 14816
rect 8481 14807 8539 14813
rect 8481 14804 8493 14807
rect 8352 14776 8493 14804
rect 8352 14764 8358 14776
rect 8481 14773 8493 14776
rect 8527 14773 8539 14807
rect 8481 14767 8539 14773
rect 9030 14764 9036 14816
rect 9088 14804 9094 14816
rect 11348 14804 11376 14844
rect 9088 14776 11376 14804
rect 9088 14764 9094 14776
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 12618 14804 12624 14816
rect 11480 14776 12624 14804
rect 11480 14764 11486 14776
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 12728 14804 12756 14912
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 13357 14943 13415 14949
rect 13357 14940 13369 14943
rect 13320 14912 13369 14940
rect 13320 14900 13326 14912
rect 13357 14909 13369 14912
rect 13403 14909 13415 14943
rect 13633 14943 13691 14949
rect 13633 14940 13645 14943
rect 13357 14903 13415 14909
rect 13464 14912 13645 14940
rect 12989 14875 13047 14881
rect 12989 14841 13001 14875
rect 13035 14872 13047 14875
rect 13464 14872 13492 14912
rect 13633 14909 13645 14912
rect 13679 14909 13691 14943
rect 13633 14903 13691 14909
rect 13035 14844 13492 14872
rect 14752 14872 14780 14994
rect 14918 14968 14924 15020
rect 14976 15008 14982 15020
rect 15473 15011 15531 15017
rect 14976 14980 15424 15008
rect 14976 14968 14982 14980
rect 15289 14875 15347 14881
rect 15289 14872 15301 14875
rect 14752 14844 15301 14872
rect 13035 14841 13047 14844
rect 12989 14835 13047 14841
rect 15289 14841 15301 14844
rect 15335 14841 15347 14875
rect 15289 14835 15347 14841
rect 13265 14807 13323 14813
rect 13265 14804 13277 14807
rect 12728 14776 13277 14804
rect 13265 14773 13277 14776
rect 13311 14804 13323 14807
rect 15105 14807 15163 14813
rect 15105 14804 15117 14807
rect 13311 14776 15117 14804
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 15105 14773 15117 14776
rect 15151 14773 15163 14807
rect 15396 14804 15424 14980
rect 15473 14977 15485 15011
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 15488 14872 15516 14971
rect 15562 14968 15568 15020
rect 15620 15008 15626 15020
rect 15620 14980 15665 15008
rect 15620 14968 15626 14980
rect 16040 14940 16068 15116
rect 16393 15113 16405 15116
rect 16439 15113 16451 15147
rect 17310 15144 17316 15156
rect 17271 15116 17316 15144
rect 16393 15107 16451 15113
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 18598 15144 18604 15156
rect 17727 15116 18604 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 19242 15144 19248 15156
rect 19203 15116 19248 15144
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 19334 15104 19340 15156
rect 19392 15144 19398 15156
rect 19797 15147 19855 15153
rect 19797 15144 19809 15147
rect 19392 15116 19809 15144
rect 19392 15104 19398 15116
rect 19797 15113 19809 15116
rect 19843 15113 19855 15147
rect 19797 15107 19855 15113
rect 22370 15104 22376 15156
rect 22428 15144 22434 15156
rect 23845 15147 23903 15153
rect 23845 15144 23857 15147
rect 22428 15116 23857 15144
rect 22428 15104 22434 15116
rect 23845 15113 23857 15116
rect 23891 15144 23903 15147
rect 23934 15144 23940 15156
rect 23891 15116 23940 15144
rect 23891 15113 23903 15116
rect 23845 15107 23903 15113
rect 23934 15104 23940 15116
rect 23992 15104 23998 15156
rect 24026 15104 24032 15156
rect 24084 15144 24090 15156
rect 24305 15147 24363 15153
rect 24305 15144 24317 15147
rect 24084 15116 24317 15144
rect 24084 15104 24090 15116
rect 24305 15113 24317 15116
rect 24351 15113 24363 15147
rect 24305 15107 24363 15113
rect 16114 15036 16120 15088
rect 16172 15076 16178 15088
rect 18132 15079 18190 15085
rect 16172 15048 17908 15076
rect 16172 15036 16178 15048
rect 16666 15008 16672 15020
rect 16627 14980 16672 15008
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 16834 15011 16892 15017
rect 16834 15008 16846 15011
rect 16776 14980 16846 15008
rect 16776 14940 16804 14980
rect 16834 14977 16846 14980
rect 16880 14977 16892 15011
rect 17034 15008 17040 15020
rect 16947 14980 17040 15008
rect 16834 14971 16892 14977
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17586 15008 17592 15020
rect 17267 14980 17592 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 17586 14968 17592 14980
rect 17644 14968 17650 15020
rect 17880 15017 17908 15048
rect 18132 15045 18144 15079
rect 18178 15076 18190 15079
rect 18322 15076 18328 15088
rect 18178 15048 18328 15076
rect 18178 15045 18190 15048
rect 18132 15039 18190 15045
rect 18322 15036 18328 15048
rect 18380 15036 18386 15088
rect 25038 15076 25044 15088
rect 22480 15048 24808 15076
rect 24999 15048 25044 15076
rect 17865 15011 17923 15017
rect 17865 14977 17877 15011
rect 17911 15008 17923 15011
rect 17954 15008 17960 15020
rect 17911 14980 17960 15008
rect 17911 14977 17923 14980
rect 17865 14971 17923 14977
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 18966 14968 18972 15020
rect 19024 15008 19030 15020
rect 20910 15011 20968 15017
rect 20910 15008 20922 15011
rect 19024 14980 20922 15008
rect 19024 14968 19030 14980
rect 20910 14977 20922 14980
rect 20956 14977 20968 15011
rect 20910 14971 20968 14977
rect 16942 14940 16948 14952
rect 16040 14912 16804 14940
rect 16903 14912 16948 14940
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 17052 14940 17080 14968
rect 17681 14943 17739 14949
rect 17681 14940 17693 14943
rect 17052 14912 17693 14940
rect 17681 14909 17693 14912
rect 17727 14909 17739 14943
rect 21174 14940 21180 14952
rect 21135 14912 21180 14940
rect 17681 14903 17739 14909
rect 21174 14900 21180 14912
rect 21232 14940 21238 14952
rect 21634 14940 21640 14952
rect 21232 14912 21640 14940
rect 21232 14900 21238 14912
rect 21634 14900 21640 14912
rect 21692 14940 21698 14952
rect 22480 14949 22508 15048
rect 22554 14968 22560 15020
rect 22612 15008 22618 15020
rect 22721 15011 22779 15017
rect 22721 15008 22733 15011
rect 22612 14980 22733 15008
rect 22612 14968 22618 14980
rect 22721 14977 22733 14980
rect 22767 14977 22779 15011
rect 22721 14971 22779 14977
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 15008 24271 15011
rect 24486 15008 24492 15020
rect 24259 14980 24492 15008
rect 24259 14977 24271 14980
rect 24213 14971 24271 14977
rect 24486 14968 24492 14980
rect 24544 14968 24550 15020
rect 24780 15017 24808 15048
rect 25038 15036 25044 15048
rect 25096 15036 25102 15088
rect 25590 15036 25596 15088
rect 25648 15036 25654 15088
rect 24765 15011 24823 15017
rect 24765 14977 24777 15011
rect 24811 14977 24823 15011
rect 24765 14971 24823 14977
rect 22465 14943 22523 14949
rect 22465 14940 22477 14943
rect 21692 14912 22477 14940
rect 21692 14900 21698 14912
rect 22465 14909 22477 14912
rect 22511 14909 22523 14943
rect 22465 14903 22523 14909
rect 24029 14875 24087 14881
rect 24029 14872 24041 14875
rect 15488 14844 17908 14872
rect 15749 14807 15807 14813
rect 15749 14804 15761 14807
rect 15396 14776 15761 14804
rect 15105 14767 15163 14773
rect 15749 14773 15761 14776
rect 15795 14804 15807 14807
rect 16666 14804 16672 14816
rect 15795 14776 16672 14804
rect 15795 14773 15807 14776
rect 15749 14767 15807 14773
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 17126 14764 17132 14816
rect 17184 14804 17190 14816
rect 17497 14807 17555 14813
rect 17497 14804 17509 14807
rect 17184 14776 17509 14804
rect 17184 14764 17190 14776
rect 17497 14773 17509 14776
rect 17543 14773 17555 14807
rect 17880 14804 17908 14844
rect 23400 14844 24041 14872
rect 23400 14804 23428 14844
rect 24029 14841 24041 14844
rect 24075 14841 24087 14875
rect 24029 14835 24087 14841
rect 17880 14776 23428 14804
rect 24673 14807 24731 14813
rect 17497 14767 17555 14773
rect 24673 14773 24685 14807
rect 24719 14804 24731 14807
rect 25406 14804 25412 14816
rect 24719 14776 25412 14804
rect 24719 14773 24731 14776
rect 24673 14767 24731 14773
rect 25406 14764 25412 14776
rect 25464 14764 25470 14816
rect 26510 14804 26516 14816
rect 26471 14776 26516 14804
rect 26510 14764 26516 14776
rect 26568 14764 26574 14816
rect 1104 14714 29440 14736
rect 1104 14662 5672 14714
rect 5724 14662 5736 14714
rect 5788 14662 5800 14714
rect 5852 14662 5864 14714
rect 5916 14662 5928 14714
rect 5980 14662 15118 14714
rect 15170 14662 15182 14714
rect 15234 14662 15246 14714
rect 15298 14662 15310 14714
rect 15362 14662 15374 14714
rect 15426 14662 24563 14714
rect 24615 14662 24627 14714
rect 24679 14662 24691 14714
rect 24743 14662 24755 14714
rect 24807 14662 24819 14714
rect 24871 14662 29440 14714
rect 1104 14640 29440 14662
rect 3053 14603 3111 14609
rect 3053 14569 3065 14603
rect 3099 14600 3111 14603
rect 3418 14600 3424 14612
rect 3099 14572 3424 14600
rect 3099 14569 3111 14572
rect 3053 14563 3111 14569
rect 3418 14560 3424 14572
rect 3476 14560 3482 14612
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4525 14603 4583 14609
rect 4525 14600 4537 14603
rect 4212 14572 4537 14600
rect 4212 14560 4218 14572
rect 4525 14569 4537 14572
rect 4571 14569 4583 14603
rect 4525 14563 4583 14569
rect 5534 14560 5540 14612
rect 5592 14600 5598 14612
rect 5629 14603 5687 14609
rect 5629 14600 5641 14603
rect 5592 14572 5641 14600
rect 5592 14560 5598 14572
rect 5629 14569 5641 14572
rect 5675 14569 5687 14603
rect 10778 14600 10784 14612
rect 5629 14563 5687 14569
rect 5736 14572 9904 14600
rect 10739 14572 10784 14600
rect 4062 14492 4068 14544
rect 4120 14532 4126 14544
rect 5736 14532 5764 14572
rect 4120 14504 5764 14532
rect 4120 14492 4126 14504
rect 6178 14492 6184 14544
rect 6236 14532 6242 14544
rect 6236 14504 9812 14532
rect 6236 14492 6242 14504
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 4672 14436 5089 14464
rect 4672 14424 4678 14436
rect 5077 14433 5089 14436
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 2498 14396 2504 14408
rect 2459 14368 2504 14396
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 2921 14399 2979 14405
rect 2921 14365 2933 14399
rect 2967 14396 2979 14399
rect 3142 14396 3148 14408
rect 2967 14368 3148 14396
rect 2967 14365 2979 14368
rect 2921 14359 2979 14365
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 3292 14368 3337 14396
rect 3292 14356 3298 14368
rect 5258 14356 5264 14408
rect 5316 14396 5322 14408
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 5316 14368 5549 14396
rect 5316 14356 5322 14368
rect 5537 14365 5549 14368
rect 5583 14365 5595 14399
rect 5537 14359 5595 14365
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 7101 14399 7159 14405
rect 7101 14396 7113 14399
rect 6972 14368 7113 14396
rect 6972 14356 6978 14368
rect 7101 14365 7113 14368
rect 7147 14396 7159 14399
rect 7742 14396 7748 14408
rect 7147 14368 7748 14396
rect 7147 14365 7159 14368
rect 7101 14359 7159 14365
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 8294 14396 8300 14408
rect 8255 14368 8300 14396
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14396 8447 14399
rect 9674 14396 9680 14408
rect 8435 14368 9680 14396
rect 8435 14365 8447 14368
rect 8389 14359 8447 14365
rect 2685 14331 2743 14337
rect 2685 14297 2697 14331
rect 2731 14297 2743 14331
rect 2685 14291 2743 14297
rect 2777 14331 2835 14337
rect 2777 14297 2789 14331
rect 2823 14328 2835 14331
rect 3252 14328 3280 14356
rect 2823 14300 3280 14328
rect 4893 14331 4951 14337
rect 2823 14297 2835 14300
rect 2777 14291 2835 14297
rect 4893 14297 4905 14331
rect 4939 14328 4951 14331
rect 5074 14328 5080 14340
rect 4939 14300 5080 14328
rect 4939 14297 4951 14300
rect 4893 14291 4951 14297
rect 2700 14260 2728 14291
rect 5074 14288 5080 14300
rect 5132 14328 5138 14340
rect 5353 14331 5411 14337
rect 5353 14328 5365 14331
rect 5132 14300 5365 14328
rect 5132 14288 5138 14300
rect 5353 14297 5365 14300
rect 5399 14297 5411 14331
rect 8404 14328 8432 14359
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 5353 14291 5411 14297
rect 7944 14300 8432 14328
rect 9784 14328 9812 14504
rect 9876 14464 9904 14572
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 11149 14603 11207 14609
rect 11149 14569 11161 14603
rect 11195 14600 11207 14603
rect 16485 14603 16543 14609
rect 11195 14572 14228 14600
rect 11195 14569 11207 14572
rect 11149 14563 11207 14569
rect 10689 14535 10747 14541
rect 10689 14501 10701 14535
rect 10735 14532 10747 14535
rect 11164 14532 11192 14563
rect 10735 14504 11192 14532
rect 10735 14501 10747 14504
rect 10689 14495 10747 14501
rect 11606 14492 11612 14544
rect 11664 14532 11670 14544
rect 11664 14504 12020 14532
rect 11664 14492 11670 14504
rect 11992 14464 12020 14504
rect 13170 14464 13176 14476
rect 9876 14436 11928 14464
rect 11992 14436 13176 14464
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14396 10471 14399
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 10459 14368 10701 14396
rect 10459 14365 10471 14368
rect 10413 14359 10471 14365
rect 10689 14365 10701 14368
rect 10735 14396 10747 14399
rect 10778 14396 10784 14408
rect 10735 14368 10784 14396
rect 10735 14365 10747 14368
rect 10689 14359 10747 14365
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11606 14396 11612 14408
rect 11011 14368 11612 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 11422 14328 11428 14340
rect 9784 14300 11428 14328
rect 3329 14263 3387 14269
rect 3329 14260 3341 14263
rect 2700 14232 3341 14260
rect 3329 14229 3341 14232
rect 3375 14229 3387 14263
rect 3329 14223 3387 14229
rect 4985 14263 5043 14269
rect 4985 14229 4997 14263
rect 5031 14260 5043 14263
rect 5626 14260 5632 14272
rect 5031 14232 5632 14260
rect 5031 14229 5043 14232
rect 4985 14223 5043 14229
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 7006 14260 7012 14272
rect 6967 14232 7012 14260
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7190 14220 7196 14272
rect 7248 14260 7254 14272
rect 7742 14260 7748 14272
rect 7248 14232 7748 14260
rect 7248 14220 7254 14232
rect 7742 14220 7748 14232
rect 7800 14260 7806 14272
rect 7944 14269 7972 14300
rect 11422 14288 11428 14300
rect 11480 14288 11486 14340
rect 7929 14263 7987 14269
rect 7929 14260 7941 14263
rect 7800 14232 7941 14260
rect 7800 14220 7806 14232
rect 7929 14229 7941 14232
rect 7975 14229 7987 14263
rect 8202 14260 8208 14272
rect 8163 14232 8208 14260
rect 7929 14223 7987 14229
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 10597 14263 10655 14269
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 10870 14260 10876 14272
rect 10643 14232 10876 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 11790 14260 11796 14272
rect 11751 14232 11796 14260
rect 11790 14220 11796 14232
rect 11848 14220 11854 14272
rect 11900 14260 11928 14436
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 13262 14424 13268 14476
rect 13320 14464 13326 14476
rect 13541 14467 13599 14473
rect 13541 14464 13553 14467
rect 13320 14436 13553 14464
rect 13320 14424 13326 14436
rect 13541 14433 13553 14436
rect 13587 14433 13599 14467
rect 14200 14464 14228 14572
rect 16485 14569 16497 14603
rect 16531 14600 16543 14603
rect 17034 14600 17040 14612
rect 16531 14572 17040 14600
rect 16531 14569 16543 14572
rect 16485 14563 16543 14569
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 18966 14600 18972 14612
rect 18927 14572 18972 14600
rect 18966 14560 18972 14572
rect 19024 14560 19030 14612
rect 19610 14560 19616 14612
rect 19668 14600 19674 14612
rect 22002 14600 22008 14612
rect 19668 14572 19840 14600
rect 21963 14572 22008 14600
rect 19668 14560 19674 14572
rect 14274 14492 14280 14544
rect 14332 14532 14338 14544
rect 16574 14532 16580 14544
rect 14332 14504 16580 14532
rect 14332 14492 14338 14504
rect 16574 14492 16580 14504
rect 16632 14492 16638 14544
rect 16761 14535 16819 14541
rect 16761 14501 16773 14535
rect 16807 14532 16819 14535
rect 16942 14532 16948 14544
rect 16807 14504 16948 14532
rect 16807 14501 16819 14504
rect 16761 14495 16819 14501
rect 16942 14492 16948 14504
rect 17000 14532 17006 14544
rect 18138 14532 18144 14544
rect 17000 14504 18144 14532
rect 17000 14492 17006 14504
rect 18138 14492 18144 14504
rect 18196 14532 18202 14544
rect 18196 14504 19563 14532
rect 18196 14492 18202 14504
rect 17678 14464 17684 14476
rect 14200 14436 17684 14464
rect 13541 14427 13599 14433
rect 17678 14424 17684 14436
rect 17736 14424 17742 14476
rect 18616 14473 18644 14504
rect 19535 14473 19563 14504
rect 18601 14467 18659 14473
rect 18601 14433 18613 14467
rect 18647 14433 18659 14467
rect 18601 14427 18659 14433
rect 19521 14467 19579 14473
rect 19521 14433 19533 14467
rect 19567 14433 19579 14467
rect 19521 14427 19579 14433
rect 13814 14396 13820 14408
rect 13775 14368 13820 14396
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14396 15163 14399
rect 15562 14396 15568 14408
rect 15151 14368 15568 14396
rect 15151 14365 15163 14368
rect 15105 14359 15163 14365
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14365 16359 14399
rect 16574 14396 16580 14408
rect 16535 14368 16580 14396
rect 16301 14359 16359 14365
rect 12526 14260 12532 14272
rect 11900 14232 12532 14260
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 12820 14260 12848 14314
rect 12986 14288 12992 14340
rect 13044 14328 13050 14340
rect 13265 14331 13323 14337
rect 13265 14328 13277 14331
rect 13044 14300 13277 14328
rect 13044 14288 13050 14300
rect 13265 14297 13277 14300
rect 13311 14297 13323 14331
rect 13265 14291 13323 14297
rect 13722 14288 13728 14340
rect 13780 14328 13786 14340
rect 16206 14328 16212 14340
rect 13780 14300 16212 14328
rect 13780 14288 13786 14300
rect 16206 14288 16212 14300
rect 16264 14288 16270 14340
rect 16316 14328 16344 14359
rect 16574 14356 16580 14368
rect 16632 14396 16638 14408
rect 17218 14396 17224 14408
rect 16632 14368 17224 14396
rect 16632 14356 16638 14368
rect 17218 14356 17224 14368
rect 17276 14396 17282 14408
rect 17405 14399 17463 14405
rect 17405 14396 17417 14399
rect 17276 14368 17417 14396
rect 17276 14356 17282 14368
rect 17405 14365 17417 14368
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 17770 14356 17776 14408
rect 17828 14396 17834 14408
rect 17865 14399 17923 14405
rect 17865 14396 17877 14399
rect 17828 14368 17877 14396
rect 17828 14356 17834 14368
rect 17865 14365 17877 14368
rect 17911 14365 17923 14399
rect 17865 14359 17923 14365
rect 18046 14356 18052 14408
rect 18104 14396 18110 14408
rect 18322 14396 18328 14408
rect 18104 14368 18328 14396
rect 18104 14356 18110 14368
rect 18322 14356 18328 14368
rect 18380 14356 18386 14408
rect 18490 14399 18548 14405
rect 18490 14396 18502 14399
rect 18432 14368 18502 14396
rect 16850 14328 16856 14340
rect 16316 14300 16856 14328
rect 16850 14288 16856 14300
rect 16908 14328 16914 14340
rect 17788 14328 17816 14356
rect 18432 14328 18460 14368
rect 18490 14365 18502 14368
rect 18536 14365 18548 14399
rect 18490 14359 18548 14365
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 18877 14399 18935 14405
rect 18877 14365 18889 14399
rect 18923 14396 18935 14399
rect 19058 14396 19064 14408
rect 18923 14368 19064 14396
rect 18923 14365 18935 14368
rect 18877 14359 18935 14365
rect 16908 14300 17816 14328
rect 18156 14300 18460 14328
rect 16908 14288 16914 14300
rect 18156 14272 18184 14300
rect 18598 14288 18604 14340
rect 18656 14328 18662 14340
rect 18708 14328 18736 14359
rect 19058 14356 19064 14368
rect 19116 14356 19122 14408
rect 19150 14356 19156 14408
rect 19208 14396 19214 14408
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 19208 14368 19257 14396
rect 19208 14356 19214 14368
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 19812 14405 19840 14572
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 25590 14600 25596 14612
rect 25551 14572 25596 14600
rect 25590 14560 25596 14572
rect 25648 14560 25654 14612
rect 21634 14492 21640 14544
rect 21692 14532 21698 14544
rect 22370 14532 22376 14544
rect 21692 14504 22376 14532
rect 21692 14492 21698 14504
rect 22370 14492 22376 14504
rect 22428 14492 22434 14544
rect 20162 14464 20168 14476
rect 20075 14436 20168 14464
rect 20162 14424 20168 14436
rect 20220 14464 20226 14476
rect 26694 14464 26700 14476
rect 20220 14436 26700 14464
rect 20220 14424 20226 14436
rect 26694 14424 26700 14436
rect 26752 14424 26758 14476
rect 19428 14399 19486 14405
rect 19428 14396 19440 14399
rect 19392 14368 19440 14396
rect 19392 14356 19398 14368
rect 19428 14365 19440 14368
rect 19474 14365 19486 14399
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 19428 14359 19486 14365
rect 19535 14368 19625 14396
rect 19535 14328 19563 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 19797 14399 19855 14405
rect 19797 14365 19809 14399
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 21453 14399 21511 14405
rect 21453 14365 21465 14399
rect 21499 14396 21511 14399
rect 21542 14396 21548 14408
rect 21499 14368 21548 14396
rect 21499 14365 21511 14368
rect 21453 14359 21511 14365
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 21818 14356 21824 14408
rect 21876 14405 21882 14408
rect 21876 14396 21884 14405
rect 25406 14396 25412 14408
rect 21876 14368 21921 14396
rect 25367 14368 25412 14396
rect 21876 14359 21884 14368
rect 21876 14356 21882 14359
rect 25406 14356 25412 14368
rect 25464 14356 25470 14408
rect 18656 14300 19288 14328
rect 18656 14288 18662 14300
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 12820 14232 13645 14260
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 14918 14260 14924 14272
rect 14879 14232 14924 14260
rect 13633 14223 13691 14229
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 17586 14260 17592 14272
rect 17547 14232 17592 14260
rect 17586 14220 17592 14232
rect 17644 14220 17650 14272
rect 17678 14220 17684 14272
rect 17736 14260 17742 14272
rect 18138 14260 18144 14272
rect 17736 14232 17781 14260
rect 18099 14232 18144 14260
rect 17736 14220 17742 14232
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 18322 14220 18328 14272
rect 18380 14260 18386 14272
rect 19150 14260 19156 14272
rect 18380 14232 19156 14260
rect 18380 14220 18386 14232
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 19260 14260 19288 14300
rect 19505 14300 19563 14328
rect 19981 14331 20039 14337
rect 19505 14260 19533 14300
rect 19981 14297 19993 14331
rect 20027 14328 20039 14331
rect 20898 14328 20904 14340
rect 20027 14300 20904 14328
rect 20027 14297 20039 14300
rect 19981 14291 20039 14297
rect 20898 14288 20904 14300
rect 20956 14288 20962 14340
rect 21634 14328 21640 14340
rect 21595 14300 21640 14328
rect 21634 14288 21640 14300
rect 21692 14288 21698 14340
rect 21729 14331 21787 14337
rect 21729 14297 21741 14331
rect 21775 14328 21787 14331
rect 21775 14300 22094 14328
rect 21775 14297 21787 14300
rect 21729 14291 21787 14297
rect 19260 14232 19533 14260
rect 22066 14260 22094 14300
rect 22278 14260 22284 14272
rect 22066 14232 22284 14260
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 1104 14170 29440 14192
rect 1104 14118 10395 14170
rect 10447 14118 10459 14170
rect 10511 14118 10523 14170
rect 10575 14118 10587 14170
rect 10639 14118 10651 14170
rect 10703 14118 19840 14170
rect 19892 14118 19904 14170
rect 19956 14118 19968 14170
rect 20020 14118 20032 14170
rect 20084 14118 20096 14170
rect 20148 14118 29440 14170
rect 1104 14096 29440 14118
rect 2498 14056 2504 14068
rect 2411 14028 2504 14056
rect 2498 14016 2504 14028
rect 2556 14056 2562 14068
rect 3421 14059 3479 14065
rect 3421 14056 3433 14059
rect 2556 14028 3433 14056
rect 2556 14016 2562 14028
rect 3421 14025 3433 14028
rect 3467 14025 3479 14059
rect 3421 14019 3479 14025
rect 4985 14059 5043 14065
rect 4985 14025 4997 14059
rect 5031 14056 5043 14059
rect 5074 14056 5080 14068
rect 5031 14028 5080 14056
rect 5031 14025 5043 14028
rect 4985 14019 5043 14025
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 5684 14028 5733 14056
rect 5684 14016 5690 14028
rect 5721 14025 5733 14028
rect 5767 14025 5779 14059
rect 5721 14019 5779 14025
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 7190 14056 7196 14068
rect 6687 14028 7196 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 7650 14056 7656 14068
rect 7392 14028 7656 14056
rect 2516 13929 2544 14016
rect 3053 13991 3111 13997
rect 3053 13988 3065 13991
rect 2700 13960 3065 13988
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13889 2559 13923
rect 2501 13883 2559 13889
rect 2590 13880 2596 13932
rect 2648 13920 2654 13932
rect 2700 13929 2728 13960
rect 3053 13957 3065 13960
rect 3099 13957 3111 13991
rect 3053 13951 3111 13957
rect 3142 13948 3148 14000
rect 3200 13988 3206 14000
rect 3237 13991 3295 13997
rect 3237 13988 3249 13991
rect 3200 13960 3249 13988
rect 3200 13948 3206 13960
rect 3237 13957 3249 13960
rect 3283 13957 3295 13991
rect 3237 13951 3295 13957
rect 3872 13991 3930 13997
rect 3872 13957 3884 13991
rect 3918 13988 3930 13991
rect 3970 13988 3976 14000
rect 3918 13960 3976 13988
rect 3918 13957 3930 13960
rect 3872 13951 3930 13957
rect 2685 13923 2743 13929
rect 2685 13920 2697 13923
rect 2648 13892 2697 13920
rect 2648 13880 2654 13892
rect 2685 13889 2697 13892
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13920 2835 13923
rect 2866 13920 2872 13932
rect 2823 13892 2872 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 3252 13920 3280 13951
rect 3970 13948 3976 13960
rect 4028 13948 4034 14000
rect 3329 13923 3387 13929
rect 3329 13920 3341 13923
rect 3252 13892 3341 13920
rect 3329 13889 3341 13892
rect 3375 13889 3387 13923
rect 5092 13920 5120 14016
rect 7392 13997 7420 14028
rect 7650 14016 7656 14028
rect 7708 14056 7714 14068
rect 8294 14056 8300 14068
rect 7708 14028 8300 14056
rect 7708 14016 7714 14028
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 9306 14056 9312 14068
rect 9267 14028 9312 14056
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 10045 14059 10103 14065
rect 10045 14025 10057 14059
rect 10091 14025 10103 14059
rect 10045 14019 10103 14025
rect 8202 13997 8208 14000
rect 7377 13991 7435 13997
rect 7377 13988 7389 13991
rect 6748 13960 7389 13988
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 5092 13892 5181 13920
rect 3329 13883 3387 13889
rect 5169 13889 5181 13892
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 5534 13880 5540 13932
rect 5592 13929 5598 13932
rect 5592 13923 5629 13929
rect 5617 13889 5629 13923
rect 5592 13883 5629 13889
rect 5592 13880 5598 13883
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 6748 13929 6776 13960
rect 7377 13957 7389 13960
rect 7423 13957 7435 13991
rect 8196 13988 8208 13997
rect 8163 13960 8208 13988
rect 7377 13951 7435 13957
rect 8196 13951 8208 13960
rect 8202 13948 8208 13951
rect 8260 13948 8266 14000
rect 10060 13988 10088 14019
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10778 14056 10784 14068
rect 10192 14028 10237 14056
rect 10739 14028 10784 14056
rect 10192 14016 10198 14028
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11790 14016 11796 14068
rect 11848 14056 11854 14068
rect 12066 14056 12072 14068
rect 11848 14028 12072 14056
rect 11848 14016 11854 14028
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 12362 14059 12420 14065
rect 12362 14025 12374 14059
rect 12408 14056 12420 14059
rect 12986 14056 12992 14068
rect 12408 14028 12992 14056
rect 12408 14025 12420 14028
rect 12362 14019 12420 14025
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 13814 14056 13820 14068
rect 13587 14028 13820 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14025 14151 14059
rect 14093 14019 14151 14025
rect 10060 13960 10640 13988
rect 6733 13923 6791 13929
rect 6733 13920 6745 13923
rect 6328 13892 6745 13920
rect 6328 13880 6334 13892
rect 6733 13889 6745 13892
rect 6779 13889 6791 13923
rect 7006 13920 7012 13932
rect 6967 13892 7012 13920
rect 6733 13883 6791 13889
rect 7006 13880 7012 13892
rect 7064 13880 7070 13932
rect 7098 13880 7104 13932
rect 7156 13920 7162 13932
rect 7285 13923 7343 13929
rect 7156 13892 7201 13920
rect 7156 13880 7162 13892
rect 7285 13889 7297 13923
rect 7331 13920 7343 13923
rect 7466 13920 7472 13932
rect 7331 13892 7472 13920
rect 7331 13889 7343 13892
rect 7285 13883 7343 13889
rect 7466 13880 7472 13892
rect 7524 13920 7530 13932
rect 9861 13923 9919 13929
rect 7524 13892 8984 13920
rect 7524 13880 7530 13892
rect 1394 13812 1400 13864
rect 1452 13852 1458 13864
rect 3605 13855 3663 13861
rect 3605 13852 3617 13855
rect 1452 13824 3617 13852
rect 1452 13812 1458 13824
rect 3605 13821 3617 13824
rect 3651 13821 3663 13855
rect 5258 13852 5264 13864
rect 5219 13824 5264 13852
rect 3605 13815 3663 13821
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 6914 13852 6920 13864
rect 6875 13824 6920 13852
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 7929 13855 7987 13861
rect 7929 13821 7941 13855
rect 7975 13821 7987 13855
rect 8956 13852 8984 13892
rect 9861 13889 9873 13923
rect 9907 13920 9919 13923
rect 10134 13920 10140 13932
rect 9907 13892 10140 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 10612 13929 10640 13960
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13889 10379 13923
rect 10321 13883 10379 13889
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 10336 13852 10364 13883
rect 10796 13852 10824 14016
rect 12621 13991 12679 13997
rect 12621 13988 12633 13991
rect 11992 13960 12633 13988
rect 11793 13923 11851 13929
rect 11793 13889 11805 13923
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 11808 13852 11836 13883
rect 11882 13880 11888 13932
rect 11940 13920 11946 13932
rect 11992 13929 12020 13960
rect 12621 13957 12633 13960
rect 12667 13988 12679 13991
rect 12710 13988 12716 14000
rect 12667 13960 12716 13988
rect 12667 13957 12679 13960
rect 12621 13951 12679 13957
rect 12710 13948 12716 13960
rect 12768 13948 12774 14000
rect 13170 13948 13176 14000
rect 13228 13988 13234 14000
rect 14108 13988 14136 14019
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 16393 14059 16451 14065
rect 16393 14056 16405 14059
rect 15528 14028 16405 14056
rect 15528 14016 15534 14028
rect 16393 14025 16405 14028
rect 16439 14056 16451 14059
rect 18690 14056 18696 14068
rect 16439 14028 18368 14056
rect 18651 14028 18696 14056
rect 16439 14025 16451 14028
rect 16393 14019 16451 14025
rect 18340 13988 18368 14028
rect 18690 14016 18696 14028
rect 18748 14016 18754 14068
rect 19610 14016 19616 14068
rect 19668 14056 19674 14068
rect 19797 14059 19855 14065
rect 19797 14056 19809 14059
rect 19668 14028 19809 14056
rect 19668 14016 19674 14028
rect 19797 14025 19809 14028
rect 19843 14025 19855 14059
rect 19797 14019 19855 14025
rect 22002 14016 22008 14068
rect 22060 14056 22066 14068
rect 23014 14056 23020 14068
rect 22060 14028 23020 14056
rect 22060 14016 22066 14028
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 19061 13991 19119 13997
rect 19061 13988 19073 13991
rect 13228 13960 14136 13988
rect 15028 13960 17172 13988
rect 18340 13960 19073 13988
rect 13228 13948 13234 13960
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 11940 13892 11989 13920
rect 11940 13880 11946 13892
rect 11977 13889 11989 13892
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12066 13880 12072 13932
rect 12124 13920 12130 13932
rect 12213 13923 12271 13929
rect 12124 13892 12169 13920
rect 12124 13880 12130 13892
rect 12213 13889 12225 13923
rect 12259 13920 12271 13923
rect 12802 13920 12808 13932
rect 12259 13892 12808 13920
rect 12259 13889 12271 13892
rect 12213 13883 12271 13889
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 13814 13920 13820 13932
rect 13403 13892 13820 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13920 14059 13923
rect 14274 13920 14280 13932
rect 14047 13892 14280 13920
rect 14047 13889 14059 13892
rect 14001 13883 14059 13889
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 15028 13929 15056 13960
rect 17144 13932 17172 13960
rect 19061 13957 19073 13960
rect 19107 13957 19119 13991
rect 19061 13951 19119 13957
rect 20898 13948 20904 14000
rect 20956 13997 20962 14000
rect 20956 13988 20968 13997
rect 20956 13960 21001 13988
rect 21836 13960 24992 13988
rect 20956 13951 20968 13960
rect 20956 13948 20962 13951
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 15280 13923 15338 13929
rect 15280 13889 15292 13923
rect 15326 13920 15338 13923
rect 15562 13920 15568 13932
rect 15326 13892 15568 13920
rect 15326 13889 15338 13892
rect 15280 13883 15338 13889
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 16850 13920 16856 13932
rect 16811 13892 16856 13920
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17126 13920 17132 13932
rect 17087 13892 17132 13920
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 17218 13880 17224 13932
rect 17276 13924 17282 13932
rect 17276 13920 17356 13924
rect 17396 13923 17454 13929
rect 17396 13920 17408 13923
rect 17276 13896 17408 13920
rect 17276 13880 17282 13896
rect 17328 13892 17408 13896
rect 17396 13889 17408 13892
rect 17442 13889 17454 13923
rect 21634 13920 21640 13932
rect 17396 13883 17454 13889
rect 18156 13892 21640 13920
rect 14918 13852 14924 13864
rect 8956 13824 10272 13852
rect 10336 13824 10824 13852
rect 10888 13824 11744 13852
rect 11808 13824 12020 13852
rect 7929 13815 7987 13821
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 7944 13784 7972 13815
rect 6788 13756 7972 13784
rect 10244 13784 10272 13824
rect 10888 13784 10916 13824
rect 10244 13756 10916 13784
rect 6788 13744 6794 13756
rect 2314 13716 2320 13728
rect 2275 13688 2320 13716
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 10410 13716 10416 13728
rect 10371 13688 10416 13716
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 11716 13716 11744 13824
rect 11992 13796 12020 13824
rect 12084 13824 14924 13852
rect 11974 13744 11980 13796
rect 12032 13744 12038 13796
rect 12084 13716 12112 13824
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 16206 13812 16212 13864
rect 16264 13852 16270 13864
rect 16264 13824 17172 13852
rect 16264 13812 16270 13824
rect 13814 13784 13820 13796
rect 13775 13756 13820 13784
rect 13814 13744 13820 13756
rect 13872 13784 13878 13796
rect 14274 13784 14280 13796
rect 13872 13756 14280 13784
rect 13872 13744 13878 13756
rect 14274 13744 14280 13756
rect 14332 13744 14338 13796
rect 16666 13716 16672 13728
rect 11716 13688 12112 13716
rect 16627 13688 16672 13716
rect 16666 13676 16672 13688
rect 16724 13676 16730 13728
rect 17144 13716 17172 13824
rect 18156 13716 18184 13892
rect 21634 13880 21640 13892
rect 21692 13880 21698 13932
rect 19153 13855 19211 13861
rect 19153 13852 19165 13855
rect 18524 13824 19165 13852
rect 18524 13728 18552 13824
rect 19153 13821 19165 13824
rect 19199 13821 19211 13855
rect 19153 13815 19211 13821
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13821 19303 13855
rect 21174 13852 21180 13864
rect 21135 13824 21180 13852
rect 19245 13815 19303 13821
rect 18598 13744 18604 13796
rect 18656 13784 18662 13796
rect 18782 13784 18788 13796
rect 18656 13756 18788 13784
rect 18656 13744 18662 13756
rect 18782 13744 18788 13756
rect 18840 13784 18846 13796
rect 19260 13784 19288 13815
rect 21174 13812 21180 13824
rect 21232 13852 21238 13864
rect 21836 13861 21864 13960
rect 22094 13929 22100 13932
rect 22088 13920 22100 13929
rect 22055 13892 22100 13920
rect 22088 13883 22100 13892
rect 22094 13880 22100 13883
rect 22152 13880 22158 13932
rect 23400 13864 23428 13960
rect 23658 13929 23664 13932
rect 23652 13920 23664 13929
rect 23619 13892 23664 13920
rect 23652 13883 23664 13892
rect 23658 13880 23664 13883
rect 23716 13880 23722 13932
rect 24964 13929 24992 13960
rect 24949 13923 25007 13929
rect 24949 13889 24961 13923
rect 24995 13889 25007 13923
rect 24949 13883 25007 13889
rect 25038 13880 25044 13932
rect 25096 13920 25102 13932
rect 25205 13923 25263 13929
rect 25205 13920 25217 13923
rect 25096 13892 25217 13920
rect 25096 13880 25102 13892
rect 25205 13889 25217 13892
rect 25251 13889 25263 13923
rect 25205 13883 25263 13889
rect 21821 13855 21879 13861
rect 21821 13852 21833 13855
rect 21232 13824 21833 13852
rect 21232 13812 21238 13824
rect 21821 13821 21833 13824
rect 21867 13821 21879 13855
rect 23382 13852 23388 13864
rect 23343 13824 23388 13852
rect 21821 13815 21879 13821
rect 23382 13812 23388 13824
rect 23440 13812 23446 13864
rect 18840 13756 19288 13784
rect 18840 13744 18846 13756
rect 18506 13716 18512 13728
rect 17144 13688 18184 13716
rect 18467 13688 18512 13716
rect 18506 13676 18512 13688
rect 18564 13676 18570 13728
rect 22738 13676 22744 13728
rect 22796 13716 22802 13728
rect 23201 13719 23259 13725
rect 23201 13716 23213 13719
rect 22796 13688 23213 13716
rect 22796 13676 22802 13688
rect 23201 13685 23213 13688
rect 23247 13716 23259 13719
rect 23290 13716 23296 13728
rect 23247 13688 23296 13716
rect 23247 13685 23259 13688
rect 23201 13679 23259 13685
rect 23290 13676 23296 13688
rect 23348 13676 23354 13728
rect 24118 13676 24124 13728
rect 24176 13716 24182 13728
rect 24765 13719 24823 13725
rect 24765 13716 24777 13719
rect 24176 13688 24777 13716
rect 24176 13676 24182 13688
rect 24765 13685 24777 13688
rect 24811 13685 24823 13719
rect 24765 13679 24823 13685
rect 25130 13676 25136 13728
rect 25188 13716 25194 13728
rect 26329 13719 26387 13725
rect 26329 13716 26341 13719
rect 25188 13688 26341 13716
rect 25188 13676 25194 13688
rect 26329 13685 26341 13688
rect 26375 13685 26387 13719
rect 26329 13679 26387 13685
rect 1104 13626 29440 13648
rect 1104 13574 5672 13626
rect 5724 13574 5736 13626
rect 5788 13574 5800 13626
rect 5852 13574 5864 13626
rect 5916 13574 5928 13626
rect 5980 13574 15118 13626
rect 15170 13574 15182 13626
rect 15234 13574 15246 13626
rect 15298 13574 15310 13626
rect 15362 13574 15374 13626
rect 15426 13574 24563 13626
rect 24615 13574 24627 13626
rect 24679 13574 24691 13626
rect 24743 13574 24755 13626
rect 24807 13574 24819 13626
rect 24871 13574 29440 13626
rect 1104 13552 29440 13574
rect 2225 13515 2283 13521
rect 2225 13481 2237 13515
rect 2271 13512 2283 13515
rect 2774 13512 2780 13524
rect 2271 13484 2780 13512
rect 2271 13481 2283 13484
rect 2225 13475 2283 13481
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 5350 13472 5356 13524
rect 5408 13512 5414 13524
rect 8294 13512 8300 13524
rect 5408 13484 7880 13512
rect 8255 13484 8300 13512
rect 5408 13472 5414 13484
rect 7852 13444 7880 13484
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 10983 13515 11041 13521
rect 10983 13481 10995 13515
rect 11029 13512 11041 13515
rect 11425 13515 11483 13521
rect 11425 13512 11437 13515
rect 11029 13484 11437 13512
rect 11029 13481 11041 13484
rect 10983 13475 11041 13481
rect 11425 13481 11437 13484
rect 11471 13481 11483 13515
rect 11425 13475 11483 13481
rect 14366 13472 14372 13524
rect 14424 13512 14430 13524
rect 17129 13515 17187 13521
rect 17129 13512 17141 13515
rect 14424 13484 17141 13512
rect 14424 13472 14430 13484
rect 17129 13481 17141 13484
rect 17175 13481 17187 13515
rect 17129 13475 17187 13481
rect 9493 13447 9551 13453
rect 9493 13444 9505 13447
rect 7852 13416 9505 13444
rect 9493 13413 9505 13416
rect 9539 13444 9551 13447
rect 9539 13416 9674 13444
rect 9539 13413 9551 13416
rect 9493 13407 9551 13413
rect 2314 13336 2320 13388
rect 2372 13376 2378 13388
rect 2685 13379 2743 13385
rect 2685 13376 2697 13379
rect 2372 13348 2697 13376
rect 2372 13336 2378 13348
rect 2685 13345 2697 13348
rect 2731 13345 2743 13379
rect 2685 13339 2743 13345
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13376 2927 13379
rect 4614 13376 4620 13388
rect 2915 13348 4620 13376
rect 2915 13345 2927 13348
rect 2869 13339 2927 13345
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 6917 13379 6975 13385
rect 6917 13376 6929 13379
rect 6788 13348 6929 13376
rect 6788 13336 6794 13348
rect 6917 13345 6929 13348
rect 6963 13345 6975 13379
rect 6917 13339 6975 13345
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 5442 13308 5448 13320
rect 5399 13280 5448 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 5620 13311 5678 13317
rect 5620 13277 5632 13311
rect 5666 13308 5678 13311
rect 6086 13308 6092 13320
rect 5666 13280 6092 13308
rect 5666 13277 5678 13280
rect 5620 13271 5678 13277
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 7190 13317 7196 13320
rect 7184 13308 7196 13317
rect 7151 13280 7196 13308
rect 7184 13271 7196 13280
rect 7190 13268 7196 13271
rect 7248 13268 7254 13320
rect 2590 13172 2596 13184
rect 2551 13144 2596 13172
rect 2590 13132 2596 13144
rect 2648 13132 2654 13184
rect 6638 13132 6644 13184
rect 6696 13172 6702 13184
rect 6733 13175 6791 13181
rect 6733 13172 6745 13175
rect 6696 13144 6745 13172
rect 6696 13132 6702 13144
rect 6733 13141 6745 13144
rect 6779 13141 6791 13175
rect 9646 13172 9674 13416
rect 11974 13404 11980 13456
rect 12032 13404 12038 13456
rect 12526 13404 12532 13456
rect 12584 13404 12590 13456
rect 12713 13447 12771 13453
rect 12713 13413 12725 13447
rect 12759 13444 12771 13447
rect 12986 13444 12992 13456
rect 12759 13416 12992 13444
rect 12759 13413 12771 13416
rect 12713 13407 12771 13413
rect 12986 13404 12992 13416
rect 13044 13404 13050 13456
rect 15562 13444 15568 13456
rect 15523 13416 15568 13444
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 10962 13336 10968 13388
rect 11020 13376 11026 13388
rect 11241 13379 11299 13385
rect 11241 13376 11253 13379
rect 11020 13348 11253 13376
rect 11020 13336 11026 13348
rect 11241 13345 11253 13348
rect 11287 13345 11299 13379
rect 11241 13339 11299 13345
rect 11790 13336 11796 13388
rect 11848 13336 11854 13388
rect 11992 13376 12020 13404
rect 12544 13376 12572 13404
rect 13538 13376 13544 13388
rect 11992 13348 12204 13376
rect 11604 13311 11662 13317
rect 11604 13277 11616 13311
rect 11650 13308 11662 13311
rect 11808 13308 11836 13336
rect 11650 13280 11836 13308
rect 11977 13311 12035 13317
rect 11650 13277 11662 13280
rect 11604 13271 11662 13277
rect 11977 13277 11989 13311
rect 12023 13308 12035 13311
rect 12066 13308 12072 13320
rect 12023 13280 12072 13308
rect 12023 13277 12035 13280
rect 11977 13271 12035 13277
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12176 13317 12204 13348
rect 12452 13348 13544 13376
rect 12452 13317 12480 13348
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 15197 13379 15255 13385
rect 15197 13345 15209 13379
rect 15243 13376 15255 13379
rect 16666 13376 16672 13388
rect 15243 13348 16672 13376
rect 15243 13345 15255 13348
rect 15197 13339 15255 13345
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 12161 13311 12219 13317
rect 12161 13277 12173 13311
rect 12207 13277 12219 13311
rect 12161 13271 12219 13277
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 12581 13311 12639 13317
rect 12581 13277 12593 13311
rect 12627 13308 12639 13311
rect 12802 13308 12808 13320
rect 12627 13280 12808 13308
rect 12627 13277 12639 13280
rect 12581 13271 12639 13277
rect 12802 13268 12808 13280
rect 12860 13268 12866 13320
rect 14826 13308 14832 13320
rect 14787 13280 14832 13308
rect 14826 13268 14832 13280
rect 14884 13268 14890 13320
rect 14994 13308 15052 13314
rect 14994 13274 15006 13308
rect 15040 13274 15052 13308
rect 14994 13268 15052 13274
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13277 15163 13311
rect 15105 13271 15163 13277
rect 15381 13311 15439 13317
rect 15381 13277 15393 13311
rect 15427 13308 15439 13311
rect 15470 13308 15476 13320
rect 15427 13280 15476 13308
rect 15427 13277 15439 13280
rect 15381 13271 15439 13277
rect 10410 13200 10416 13252
rect 10468 13200 10474 13252
rect 11701 13243 11759 13249
rect 11701 13209 11713 13243
rect 11747 13209 11759 13243
rect 11701 13203 11759 13209
rect 11793 13243 11851 13249
rect 11793 13209 11805 13243
rect 11839 13240 11851 13243
rect 11882 13240 11888 13252
rect 11839 13212 11888 13240
rect 11839 13209 11851 13212
rect 11793 13203 11851 13209
rect 11716 13172 11744 13203
rect 11882 13200 11888 13212
rect 11940 13240 11946 13252
rect 12250 13240 12256 13252
rect 11940 13212 12256 13240
rect 11940 13200 11946 13212
rect 12250 13200 12256 13212
rect 12308 13200 12314 13252
rect 12345 13243 12403 13249
rect 12345 13209 12357 13243
rect 12391 13240 12403 13243
rect 15009 13240 15037 13268
rect 12391 13212 13032 13240
rect 12391 13209 12403 13212
rect 12345 13203 12403 13209
rect 12544 13184 12572 13212
rect 9646 13144 11744 13172
rect 6733 13135 6791 13141
rect 12526 13132 12532 13184
rect 12584 13132 12590 13184
rect 13004 13181 13032 13212
rect 14660 13212 15037 13240
rect 15120 13240 15148 13271
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13308 15899 13311
rect 16574 13308 16580 13320
rect 15887 13280 16580 13308
rect 15887 13277 15899 13280
rect 15841 13271 15899 13277
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 17144 13240 17172 13475
rect 19702 13472 19708 13524
rect 19760 13512 19766 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 19760 13484 19901 13512
rect 19760 13472 19766 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 19889 13475 19947 13481
rect 20901 13515 20959 13521
rect 20901 13481 20913 13515
rect 20947 13512 20959 13515
rect 21174 13512 21180 13524
rect 20947 13484 21180 13512
rect 20947 13481 20959 13484
rect 20901 13475 20959 13481
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 21637 13515 21695 13521
rect 21637 13481 21649 13515
rect 21683 13512 21695 13515
rect 22094 13512 22100 13524
rect 21683 13484 22100 13512
rect 21683 13481 21695 13484
rect 21637 13475 21695 13481
rect 22094 13472 22100 13484
rect 22152 13472 22158 13524
rect 22373 13515 22431 13521
rect 22373 13481 22385 13515
rect 22419 13512 22431 13515
rect 22554 13512 22560 13524
rect 22419 13484 22560 13512
rect 22419 13481 22431 13484
rect 22373 13475 22431 13481
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 23658 13472 23664 13524
rect 23716 13512 23722 13524
rect 23845 13515 23903 13521
rect 23845 13512 23857 13515
rect 23716 13484 23857 13512
rect 23716 13472 23722 13484
rect 23845 13481 23857 13484
rect 23891 13481 23903 13515
rect 24121 13515 24179 13521
rect 24121 13512 24133 13515
rect 23845 13475 23903 13481
rect 23952 13484 24133 13512
rect 17218 13404 17224 13456
rect 17276 13444 17282 13456
rect 17313 13447 17371 13453
rect 17313 13444 17325 13447
rect 17276 13416 17325 13444
rect 17276 13404 17282 13416
rect 17313 13413 17325 13416
rect 17359 13413 17371 13447
rect 18506 13444 18512 13456
rect 17313 13407 17371 13413
rect 17512 13416 18512 13444
rect 17512 13317 17540 13416
rect 18506 13404 18512 13416
rect 18564 13404 18570 13456
rect 21818 13444 21824 13456
rect 21731 13416 21824 13444
rect 17678 13376 17684 13388
rect 17639 13348 17684 13376
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 21634 13376 21640 13388
rect 21100 13348 21640 13376
rect 17497 13311 17555 13317
rect 17497 13277 17509 13311
rect 17543 13277 17555 13311
rect 17497 13271 17555 13277
rect 17586 13268 17592 13320
rect 17644 13308 17650 13320
rect 17773 13311 17831 13317
rect 17773 13308 17785 13311
rect 17644 13280 17785 13308
rect 17644 13268 17650 13280
rect 17773 13277 17785 13280
rect 17819 13277 17831 13311
rect 17866 13311 17924 13317
rect 17866 13308 17878 13311
rect 17773 13271 17831 13277
rect 17861 13277 17878 13308
rect 17912 13277 17924 13311
rect 18046 13308 18052 13320
rect 18007 13280 18052 13308
rect 17861 13271 17924 13277
rect 17861 13240 17889 13271
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 21100 13317 21128 13348
rect 21634 13336 21640 13348
rect 21692 13336 21698 13388
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 21505 13311 21563 13317
rect 21505 13277 21517 13311
rect 21551 13308 21563 13311
rect 21744 13308 21772 13416
rect 21818 13404 21824 13416
rect 21876 13444 21882 13456
rect 21876 13416 22232 13444
rect 21876 13404 21882 13416
rect 22204 13320 22232 13416
rect 22738 13404 22744 13456
rect 22796 13444 22802 13456
rect 23952 13444 23980 13484
rect 24121 13481 24133 13484
rect 24167 13512 24179 13515
rect 24486 13512 24492 13524
rect 24167 13484 24492 13512
rect 24167 13481 24179 13484
rect 24121 13475 24179 13481
rect 24486 13472 24492 13484
rect 24544 13472 24550 13524
rect 24949 13515 25007 13521
rect 24949 13481 24961 13515
rect 24995 13512 25007 13515
rect 25038 13512 25044 13524
rect 24995 13484 25044 13512
rect 24995 13481 25007 13484
rect 24949 13475 25007 13481
rect 25038 13472 25044 13484
rect 25096 13472 25102 13524
rect 22796 13416 23980 13444
rect 22796 13404 22802 13416
rect 24026 13404 24032 13456
rect 24084 13444 24090 13456
rect 25317 13447 25375 13453
rect 25317 13444 25329 13447
rect 24084 13416 25329 13444
rect 24084 13404 24090 13416
rect 25317 13413 25329 13416
rect 25363 13413 25375 13447
rect 25317 13407 25375 13413
rect 22370 13336 22376 13388
rect 22428 13376 22434 13388
rect 22557 13379 22615 13385
rect 22557 13376 22569 13379
rect 22428 13348 22569 13376
rect 22428 13336 22434 13348
rect 22557 13345 22569 13348
rect 22603 13345 22615 13379
rect 22557 13339 22615 13345
rect 23308 13348 23980 13376
rect 21551 13280 21772 13308
rect 21551 13277 21563 13280
rect 21505 13271 21563 13277
rect 21818 13268 21824 13320
rect 21876 13308 21882 13320
rect 21876 13280 21921 13308
rect 21876 13268 21882 13280
rect 22002 13268 22008 13320
rect 22060 13308 22066 13320
rect 22060 13280 22105 13308
rect 22060 13268 22066 13280
rect 22186 13268 22192 13320
rect 22244 13317 22250 13320
rect 22244 13308 22252 13317
rect 22244 13280 22337 13308
rect 22244 13271 22252 13280
rect 22244 13268 22250 13271
rect 15120 13212 15516 13240
rect 17144 13212 17889 13240
rect 18325 13243 18383 13249
rect 14660 13184 14688 13212
rect 15488 13184 15516 13212
rect 18325 13209 18337 13243
rect 18371 13240 18383 13243
rect 20254 13240 20260 13252
rect 18371 13212 20260 13240
rect 18371 13209 18383 13212
rect 18325 13203 18383 13209
rect 20254 13200 20260 13212
rect 20312 13240 20318 13252
rect 20809 13243 20867 13249
rect 20809 13240 20821 13243
rect 20312 13212 20821 13240
rect 20312 13200 20318 13212
rect 20809 13209 20821 13212
rect 20855 13209 20867 13243
rect 20809 13203 20867 13209
rect 20990 13200 20996 13252
rect 21048 13240 21054 13252
rect 21269 13243 21327 13249
rect 21269 13240 21281 13243
rect 21048 13212 21281 13240
rect 21048 13200 21054 13212
rect 21269 13209 21281 13212
rect 21315 13209 21327 13243
rect 21269 13203 21327 13209
rect 21361 13243 21419 13249
rect 21361 13209 21373 13243
rect 21407 13209 21419 13243
rect 21361 13203 21419 13209
rect 22097 13243 22155 13249
rect 22097 13209 22109 13243
rect 22143 13240 22155 13243
rect 22388 13240 22416 13336
rect 23308 13317 23336 13348
rect 23952 13320 23980 13348
rect 23293 13311 23351 13317
rect 23293 13277 23305 13311
rect 23339 13277 23351 13311
rect 23569 13311 23627 13317
rect 23569 13308 23581 13311
rect 23293 13271 23351 13277
rect 23400 13280 23581 13308
rect 23400 13240 23428 13280
rect 23569 13277 23581 13280
rect 23615 13277 23627 13311
rect 23569 13271 23627 13277
rect 23713 13311 23771 13317
rect 23713 13277 23725 13311
rect 23759 13308 23771 13311
rect 23759 13280 23888 13308
rect 23759 13277 23771 13280
rect 23713 13271 23771 13277
rect 22143 13212 22416 13240
rect 23308 13212 23428 13240
rect 23477 13243 23535 13249
rect 22143 13209 22155 13212
rect 22097 13203 22155 13209
rect 12989 13175 13047 13181
rect 12989 13141 13001 13175
rect 13035 13172 13047 13175
rect 14550 13172 14556 13184
rect 13035 13144 14556 13172
rect 13035 13141 13047 13144
rect 12989 13135 13047 13141
rect 14550 13132 14556 13144
rect 14608 13132 14614 13184
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 14700 13144 14745 13172
rect 14700 13132 14706 13144
rect 15470 13132 15476 13184
rect 15528 13172 15534 13184
rect 15657 13175 15715 13181
rect 15657 13172 15669 13175
rect 15528 13144 15669 13172
rect 15528 13132 15534 13144
rect 15657 13141 15669 13144
rect 15703 13141 15715 13175
rect 15657 13135 15715 13141
rect 17126 13132 17132 13184
rect 17184 13172 17190 13184
rect 17954 13172 17960 13184
rect 17184 13144 17960 13172
rect 17184 13132 17190 13144
rect 17954 13132 17960 13144
rect 18012 13172 18018 13184
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 18012 13144 18245 13172
rect 18012 13132 18018 13144
rect 18233 13141 18245 13144
rect 18279 13172 18291 13175
rect 19242 13172 19248 13184
rect 18279 13144 19248 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 21376 13172 21404 13203
rect 23308 13184 23336 13212
rect 23477 13209 23489 13243
rect 23523 13209 23535 13243
rect 23860 13240 23888 13280
rect 23934 13268 23940 13320
rect 23992 13308 23998 13320
rect 24397 13311 24455 13317
rect 24397 13308 24409 13311
rect 23992 13280 24409 13308
rect 23992 13268 23998 13280
rect 24397 13277 24409 13280
rect 24443 13277 24455 13311
rect 24397 13271 24455 13277
rect 24486 13268 24492 13320
rect 24544 13308 24550 13320
rect 24770 13311 24828 13317
rect 24770 13308 24782 13311
rect 24544 13280 24782 13308
rect 24544 13268 24550 13280
rect 24770 13277 24782 13280
rect 24816 13277 24828 13311
rect 24770 13271 24828 13277
rect 24578 13240 24584 13252
rect 23860 13212 24164 13240
rect 24539 13212 24584 13240
rect 23477 13203 23535 13209
rect 22738 13172 22744 13184
rect 19392 13144 22744 13172
rect 19392 13132 19398 13144
rect 22738 13132 22744 13144
rect 22796 13132 22802 13184
rect 23201 13175 23259 13181
rect 23201 13141 23213 13175
rect 23247 13172 23259 13175
rect 23290 13172 23296 13184
rect 23247 13144 23296 13172
rect 23247 13141 23259 13144
rect 23201 13135 23259 13141
rect 23290 13132 23296 13144
rect 23348 13132 23354 13184
rect 23492 13172 23520 13203
rect 24026 13172 24032 13184
rect 23492 13144 24032 13172
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 24136 13172 24164 13212
rect 24578 13200 24584 13212
rect 24636 13200 24642 13252
rect 24670 13200 24676 13252
rect 24728 13240 24734 13252
rect 25130 13240 25136 13252
rect 24728 13212 25136 13240
rect 24728 13200 24734 13212
rect 25130 13200 25136 13212
rect 25188 13200 25194 13252
rect 24486 13172 24492 13184
rect 24136 13144 24492 13172
rect 24486 13132 24492 13144
rect 24544 13132 24550 13184
rect 1104 13082 29440 13104
rect 1104 13030 10395 13082
rect 10447 13030 10459 13082
rect 10511 13030 10523 13082
rect 10575 13030 10587 13082
rect 10639 13030 10651 13082
rect 10703 13030 19840 13082
rect 19892 13030 19904 13082
rect 19956 13030 19968 13082
rect 20020 13030 20032 13082
rect 20084 13030 20096 13082
rect 20148 13030 29440 13082
rect 1104 13008 29440 13030
rect 3602 12928 3608 12980
rect 3660 12968 3666 12980
rect 3973 12971 4031 12977
rect 3973 12968 3985 12971
rect 3660 12940 3985 12968
rect 3660 12928 3666 12940
rect 3973 12937 3985 12940
rect 4019 12937 4031 12971
rect 3973 12931 4031 12937
rect 4062 12928 4068 12980
rect 4120 12968 4126 12980
rect 8662 12968 8668 12980
rect 4120 12940 8668 12968
rect 4120 12928 4126 12940
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 8864 12940 10640 12968
rect 8864 12912 8892 12940
rect 2685 12903 2743 12909
rect 2685 12869 2697 12903
rect 2731 12900 2743 12903
rect 3050 12900 3056 12912
rect 2731 12872 3056 12900
rect 2731 12869 2743 12872
rect 2685 12863 2743 12869
rect 3050 12860 3056 12872
rect 3108 12900 3114 12912
rect 3878 12900 3884 12912
rect 3108 12872 3884 12900
rect 3108 12860 3114 12872
rect 3878 12860 3884 12872
rect 3936 12860 3942 12912
rect 5534 12860 5540 12912
rect 5592 12900 5598 12912
rect 6730 12900 6736 12912
rect 5592 12872 6736 12900
rect 5592 12860 5598 12872
rect 6730 12860 6736 12872
rect 6788 12860 6794 12912
rect 6917 12903 6975 12909
rect 6917 12869 6929 12903
rect 6963 12900 6975 12903
rect 8846 12900 8852 12912
rect 6963 12872 8852 12900
rect 6963 12869 6975 12872
rect 6917 12863 6975 12869
rect 8846 12860 8852 12872
rect 8904 12860 8910 12912
rect 9490 12860 9496 12912
rect 9548 12860 9554 12912
rect 10042 12860 10048 12912
rect 10100 12900 10106 12912
rect 10612 12909 10640 12940
rect 12342 12928 12348 12980
rect 12400 12968 12406 12980
rect 12526 12968 12532 12980
rect 12400 12940 12532 12968
rect 12400 12928 12406 12940
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 13262 12928 13268 12980
rect 13320 12928 13326 12980
rect 13538 12928 13544 12980
rect 13596 12968 13602 12980
rect 14369 12971 14427 12977
rect 14369 12968 14381 12971
rect 13596 12940 14381 12968
rect 13596 12928 13602 12940
rect 14369 12937 14381 12940
rect 14415 12937 14427 12971
rect 14369 12931 14427 12937
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 17589 12971 17647 12977
rect 17589 12968 17601 12971
rect 17552 12940 17601 12968
rect 17552 12928 17558 12940
rect 17589 12937 17601 12940
rect 17635 12937 17647 12971
rect 17589 12931 17647 12937
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18322 12968 18328 12980
rect 18095 12940 18328 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18322 12928 18328 12940
rect 18380 12968 18386 12980
rect 18601 12971 18659 12977
rect 18601 12968 18613 12971
rect 18380 12940 18613 12968
rect 18380 12928 18386 12940
rect 18601 12937 18613 12940
rect 18647 12937 18659 12971
rect 18601 12931 18659 12937
rect 19702 12928 19708 12980
rect 19760 12928 19766 12980
rect 20254 12968 20260 12980
rect 20215 12940 20260 12968
rect 20254 12928 20260 12940
rect 20312 12928 20318 12980
rect 20990 12928 20996 12980
rect 21048 12968 21054 12980
rect 22278 12968 22284 12980
rect 21048 12940 22284 12968
rect 21048 12928 21054 12940
rect 22278 12928 22284 12940
rect 22336 12928 22342 12980
rect 22833 12971 22891 12977
rect 22833 12937 22845 12971
rect 22879 12968 22891 12971
rect 23566 12968 23572 12980
rect 22879 12940 23572 12968
rect 22879 12937 22891 12940
rect 22833 12931 22891 12937
rect 23566 12928 23572 12940
rect 23624 12968 23630 12980
rect 23934 12968 23940 12980
rect 23624 12940 23940 12968
rect 23624 12928 23630 12940
rect 23934 12928 23940 12940
rect 23992 12928 23998 12980
rect 10597 12903 10655 12909
rect 10100 12872 10456 12900
rect 10100 12860 10106 12872
rect 4062 12832 4068 12844
rect 4023 12804 4068 12832
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 6638 12832 6644 12844
rect 6599 12804 6644 12832
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 7282 12832 7288 12844
rect 7243 12804 7288 12832
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12801 7619 12835
rect 7561 12795 7619 12801
rect 7687 12835 7745 12841
rect 7687 12801 7699 12835
rect 7733 12832 7745 12835
rect 8754 12832 8760 12844
rect 7733 12804 8760 12832
rect 7733 12801 7745 12804
rect 7687 12795 7745 12801
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 4154 12764 4160 12776
rect 3927 12736 4160 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 4154 12724 4160 12736
rect 4212 12764 4218 12776
rect 4430 12764 4436 12776
rect 4212 12736 4436 12764
rect 4212 12724 4218 12736
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 7576 12764 7604 12795
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 10428 12841 10456 12872
rect 10597 12869 10609 12903
rect 10643 12869 10655 12903
rect 10597 12863 10655 12869
rect 10781 12903 10839 12909
rect 10781 12869 10793 12903
rect 10827 12900 10839 12903
rect 10962 12900 10968 12912
rect 10827 12872 10968 12900
rect 10827 12869 10839 12872
rect 10781 12863 10839 12869
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 10796 12832 10824 12863
rect 10962 12860 10968 12872
rect 11020 12900 11026 12912
rect 12894 12900 12900 12912
rect 11020 12872 12900 12900
rect 11020 12860 11026 12872
rect 11790 12841 11796 12844
rect 11788 12832 11796 12841
rect 10459 12804 10824 12832
rect 11751 12804 11796 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 11788 12795 11796 12804
rect 11790 12792 11796 12795
rect 11848 12792 11854 12844
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12801 11943 12835
rect 11885 12795 11943 12801
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12801 12035 12835
rect 11977 12795 12035 12801
rect 8386 12764 8392 12776
rect 7576 12736 8392 12764
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12764 10195 12767
rect 10183 12736 11652 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12696 2467 12699
rect 2774 12696 2780 12708
rect 2455 12668 2780 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 2774 12656 2780 12668
rect 2832 12656 2838 12708
rect 7926 12696 7932 12708
rect 7887 12668 7932 12696
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 11624 12705 11652 12736
rect 11609 12699 11667 12705
rect 11609 12665 11621 12699
rect 11655 12665 11667 12699
rect 11609 12659 11667 12665
rect 2225 12631 2283 12637
rect 2225 12597 2237 12631
rect 2271 12628 2283 12631
rect 2958 12628 2964 12640
rect 2271 12600 2964 12628
rect 2271 12597 2283 12600
rect 2225 12591 2283 12597
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 4430 12628 4436 12640
rect 4391 12600 4436 12628
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 6420 12600 6561 12628
rect 6420 12588 6426 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 11900 12628 11928 12795
rect 11992 12764 12020 12795
rect 12066 12792 12072 12844
rect 12124 12832 12130 12844
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 12124 12804 12173 12832
rect 12124 12792 12130 12804
rect 12161 12801 12173 12804
rect 12207 12801 12219 12835
rect 12161 12795 12219 12801
rect 12250 12792 12256 12844
rect 12308 12832 12314 12844
rect 12636 12841 12664 12872
rect 12894 12860 12900 12872
rect 12952 12900 12958 12912
rect 13280 12900 13308 12928
rect 12952 12872 13308 12900
rect 12952 12860 12958 12872
rect 14550 12860 14556 12912
rect 14608 12900 14614 12912
rect 19334 12900 19340 12912
rect 14608 12872 19340 12900
rect 14608 12860 14614 12872
rect 19334 12860 19340 12872
rect 19392 12860 19398 12912
rect 19518 12860 19524 12912
rect 19576 12860 19582 12912
rect 19720 12900 19748 12928
rect 20165 12903 20223 12909
rect 20165 12900 20177 12903
rect 19720 12872 20177 12900
rect 20165 12869 20177 12872
rect 20211 12869 20223 12903
rect 22094 12900 22100 12912
rect 22055 12872 22100 12900
rect 20165 12863 20223 12869
rect 22094 12860 22100 12872
rect 22152 12860 22158 12912
rect 23290 12860 23296 12912
rect 23348 12900 23354 12912
rect 23753 12903 23811 12909
rect 23753 12900 23765 12903
rect 23348 12872 23765 12900
rect 23348 12860 23354 12872
rect 23753 12869 23765 12872
rect 23799 12900 23811 12903
rect 24118 12900 24124 12912
rect 23799 12872 24124 12900
rect 23799 12869 23811 12872
rect 23753 12863 23811 12869
rect 24118 12860 24124 12872
rect 24176 12860 24182 12912
rect 24213 12903 24271 12909
rect 24213 12869 24225 12903
rect 24259 12900 24271 12903
rect 24259 12872 24900 12900
rect 24259 12869 24271 12872
rect 24213 12863 24271 12869
rect 12621 12835 12679 12841
rect 12308 12804 12353 12832
rect 12308 12792 12314 12804
rect 12621 12801 12633 12835
rect 12667 12801 12679 12835
rect 12621 12795 12679 12801
rect 13998 12792 14004 12844
rect 14056 12792 14062 12844
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 14737 12835 14795 12841
rect 14737 12832 14749 12835
rect 14332 12804 14749 12832
rect 14332 12792 14338 12804
rect 14737 12801 14749 12804
rect 14783 12801 14795 12835
rect 14737 12795 14795 12801
rect 17034 12792 17040 12844
rect 17092 12832 17098 12844
rect 17957 12835 18015 12841
rect 17957 12832 17969 12835
rect 17092 12804 17969 12832
rect 17092 12792 17098 12804
rect 17957 12801 17969 12804
rect 18003 12801 18015 12835
rect 19536 12832 19564 12860
rect 19714 12835 19772 12841
rect 19714 12832 19726 12835
rect 19536 12804 19726 12832
rect 17957 12795 18015 12801
rect 19714 12801 19726 12804
rect 19760 12801 19772 12835
rect 19714 12795 19772 12801
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 21082 12832 21088 12844
rect 20763 12804 21088 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 22005 12835 22063 12841
rect 22005 12801 22017 12835
rect 22051 12832 22063 12835
rect 22462 12832 22468 12844
rect 22051 12804 22468 12832
rect 22051 12801 22063 12804
rect 22005 12795 22063 12801
rect 22462 12792 22468 12804
rect 22520 12832 22526 12844
rect 22649 12835 22707 12841
rect 22649 12832 22661 12835
rect 22520 12804 22661 12832
rect 22520 12792 22526 12804
rect 22649 12801 22661 12804
rect 22695 12801 22707 12835
rect 23934 12832 23940 12844
rect 23895 12804 23940 12832
rect 22649 12795 22707 12801
rect 23934 12792 23940 12804
rect 23992 12792 23998 12844
rect 24357 12835 24415 12841
rect 24357 12801 24369 12835
rect 24403 12832 24415 12835
rect 24486 12832 24492 12844
rect 24403 12804 24492 12832
rect 24403 12801 24415 12804
rect 24357 12795 24415 12801
rect 24486 12792 24492 12804
rect 24544 12792 24550 12844
rect 24872 12841 24900 12872
rect 24857 12835 24915 12841
rect 24857 12801 24869 12835
rect 24903 12832 24915 12835
rect 25406 12832 25412 12844
rect 24903 12804 25412 12832
rect 24903 12801 24915 12804
rect 24857 12795 24915 12801
rect 25406 12792 25412 12804
rect 25464 12832 25470 12844
rect 25682 12832 25688 12844
rect 25464 12804 25688 12832
rect 25464 12792 25470 12804
rect 25682 12792 25688 12804
rect 25740 12792 25746 12844
rect 12342 12764 12348 12776
rect 11992 12736 12348 12764
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12764 12955 12767
rect 12986 12764 12992 12776
rect 12943 12736 12992 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 18233 12767 18291 12773
rect 18233 12733 18245 12767
rect 18279 12764 18291 12767
rect 18414 12764 18420 12776
rect 18279 12736 18420 12764
rect 18279 12733 18291 12736
rect 18233 12727 18291 12733
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12764 20039 12767
rect 20070 12764 20076 12776
rect 20027 12736 20076 12764
rect 20027 12733 20039 12736
rect 19981 12727 20039 12733
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 23658 12656 23664 12708
rect 23716 12696 23722 12708
rect 24670 12696 24676 12708
rect 23716 12668 24676 12696
rect 23716 12656 23722 12668
rect 24670 12656 24676 12668
rect 24728 12656 24734 12708
rect 14550 12628 14556 12640
rect 8720 12600 11928 12628
rect 14511 12600 14556 12628
rect 8720 12588 8726 12600
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 20438 12588 20444 12640
rect 20496 12628 20502 12640
rect 20533 12631 20591 12637
rect 20533 12628 20545 12631
rect 20496 12600 20545 12628
rect 20496 12588 20502 12600
rect 20533 12597 20545 12600
rect 20579 12597 20591 12631
rect 21818 12628 21824 12640
rect 21779 12600 21824 12628
rect 20533 12591 20591 12597
rect 21818 12588 21824 12600
rect 21876 12588 21882 12640
rect 24486 12628 24492 12640
rect 24447 12600 24492 12628
rect 24486 12588 24492 12600
rect 24544 12588 24550 12640
rect 1104 12538 29440 12560
rect 1104 12486 5672 12538
rect 5724 12486 5736 12538
rect 5788 12486 5800 12538
rect 5852 12486 5864 12538
rect 5916 12486 5928 12538
rect 5980 12486 15118 12538
rect 15170 12486 15182 12538
rect 15234 12486 15246 12538
rect 15298 12486 15310 12538
rect 15362 12486 15374 12538
rect 15426 12486 24563 12538
rect 24615 12486 24627 12538
rect 24679 12486 24691 12538
rect 24743 12486 24755 12538
rect 24807 12486 24819 12538
rect 24871 12486 29440 12538
rect 1104 12464 29440 12486
rect 2590 12384 2596 12436
rect 2648 12424 2654 12436
rect 2777 12427 2835 12433
rect 2777 12424 2789 12427
rect 2648 12396 2789 12424
rect 2648 12384 2654 12396
rect 2777 12393 2789 12396
rect 2823 12393 2835 12427
rect 5258 12424 5264 12436
rect 5219 12396 5264 12424
rect 2777 12387 2835 12393
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 6178 12384 6184 12436
rect 6236 12424 6242 12436
rect 7650 12424 7656 12436
rect 6236 12396 7656 12424
rect 6236 12384 6242 12396
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 8665 12427 8723 12433
rect 8665 12393 8677 12427
rect 8711 12424 8723 12427
rect 8754 12424 8760 12436
rect 8711 12396 8760 12424
rect 8711 12393 8723 12396
rect 8665 12387 8723 12393
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 9490 12424 9496 12436
rect 9451 12396 9496 12424
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 12802 12424 12808 12436
rect 9600 12396 12204 12424
rect 12763 12396 12808 12424
rect 3418 12356 3424 12368
rect 3379 12328 3424 12356
rect 3418 12316 3424 12328
rect 3476 12316 3482 12368
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 3050 12288 3056 12300
rect 3011 12260 3056 12288
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 5534 12288 5540 12300
rect 4908 12260 5540 12288
rect 1412 12220 1440 12248
rect 3881 12223 3939 12229
rect 3881 12220 3893 12223
rect 1412 12192 3893 12220
rect 3881 12189 3893 12192
rect 3927 12220 3939 12223
rect 4908 12220 4936 12260
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 9600 12288 9628 12396
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 10134 12356 10140 12368
rect 9732 12328 10140 12356
rect 9732 12316 9738 12328
rect 10134 12316 10140 12328
rect 10192 12316 10198 12368
rect 11241 12359 11299 12365
rect 11241 12325 11253 12359
rect 11287 12325 11299 12359
rect 11241 12319 11299 12325
rect 11146 12288 11152 12300
rect 8312 12260 9628 12288
rect 11072 12260 11152 12288
rect 3927 12192 4936 12220
rect 3927 12189 3939 12192
rect 3881 12183 3939 12189
rect 5258 12180 5264 12232
rect 5316 12220 5322 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 5316 12192 5457 12220
rect 5316 12180 5322 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 6178 12220 6184 12232
rect 6139 12192 6184 12220
rect 5445 12183 5503 12189
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 6362 12220 6368 12232
rect 6323 12192 6368 12220
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 6730 12180 6736 12232
rect 6788 12220 6794 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 6788 12192 7297 12220
rect 6788 12180 6794 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 7552 12223 7610 12229
rect 7552 12189 7564 12223
rect 7598 12220 7610 12223
rect 7926 12220 7932 12232
rect 7598 12192 7932 12220
rect 7598 12189 7610 12192
rect 7552 12183 7610 12189
rect 7926 12180 7932 12192
rect 7984 12180 7990 12232
rect 1664 12155 1722 12161
rect 1664 12121 1676 12155
rect 1710 12152 1722 12155
rect 1946 12152 1952 12164
rect 1710 12124 1952 12152
rect 1710 12121 1722 12124
rect 1664 12115 1722 12121
rect 1946 12112 1952 12124
rect 2004 12112 2010 12164
rect 4148 12155 4206 12161
rect 4148 12121 4160 12155
rect 4194 12152 4206 12155
rect 4430 12152 4436 12164
rect 4194 12124 4436 12152
rect 4194 12121 4206 12124
rect 4148 12115 4206 12121
rect 4430 12112 4436 12124
rect 4488 12112 4494 12164
rect 8312 12152 8340 12260
rect 11072 12232 11100 12260
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 11256 12288 11284 12319
rect 11330 12288 11336 12300
rect 11243 12260 11336 12288
rect 11330 12248 11336 12260
rect 11388 12288 11394 12300
rect 12066 12288 12072 12300
rect 11388 12260 12072 12288
rect 11388 12248 11394 12260
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12220 9275 12223
rect 9490 12220 9496 12232
rect 9263 12192 9496 12220
rect 9263 12189 9275 12192
rect 9217 12183 9275 12189
rect 9490 12180 9496 12192
rect 9548 12180 9554 12232
rect 9677 12223 9735 12229
rect 9677 12220 9689 12223
rect 9600 12192 9689 12220
rect 4540 12124 8340 12152
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12084 3571 12087
rect 3786 12084 3792 12096
rect 3559 12056 3792 12084
rect 3559 12053 3571 12056
rect 3513 12047 3571 12053
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 3970 12044 3976 12096
rect 4028 12084 4034 12096
rect 4540 12084 4568 12124
rect 4028 12056 4568 12084
rect 4028 12044 4034 12056
rect 4982 12044 4988 12096
rect 5040 12084 5046 12096
rect 5537 12087 5595 12093
rect 5537 12084 5549 12087
rect 5040 12056 5549 12084
rect 5040 12044 5046 12056
rect 5537 12053 5549 12056
rect 5583 12053 5595 12087
rect 5537 12047 5595 12053
rect 5997 12087 6055 12093
rect 5997 12053 6009 12087
rect 6043 12084 6055 12087
rect 6178 12084 6184 12096
rect 6043 12056 6184 12084
rect 6043 12053 6055 12056
rect 5997 12047 6055 12053
rect 6178 12044 6184 12056
rect 6236 12044 6242 12096
rect 6365 12087 6423 12093
rect 6365 12053 6377 12087
rect 6411 12084 6423 12087
rect 6454 12084 6460 12096
rect 6411 12056 6460 12084
rect 6411 12053 6423 12056
rect 6365 12047 6423 12053
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 9600 12084 9628 12192
rect 9677 12189 9689 12192
rect 9723 12189 9735 12223
rect 11054 12220 11060 12232
rect 10967 12192 11060 12220
rect 9677 12183 9735 12189
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11422 12220 11428 12232
rect 11164 12192 11428 12220
rect 9447 12056 9628 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 11164 12084 11192 12192
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 11900 12229 11928 12260
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12176 12288 12204 12396
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 14056 12396 14105 12424
rect 14056 12384 14062 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 14093 12387 14151 12393
rect 17678 12384 17684 12436
rect 17736 12424 17742 12436
rect 18417 12427 18475 12433
rect 17736 12396 18184 12424
rect 17736 12384 17742 12396
rect 12437 12359 12495 12365
rect 12437 12325 12449 12359
rect 12483 12356 12495 12359
rect 15654 12356 15660 12368
rect 12483 12328 15660 12356
rect 12483 12325 12495 12328
rect 12437 12319 12495 12325
rect 15654 12316 15660 12328
rect 15712 12316 15718 12368
rect 17586 12316 17592 12368
rect 17644 12356 17650 12368
rect 18046 12356 18052 12368
rect 17644 12328 18052 12356
rect 17644 12316 17650 12328
rect 18046 12316 18052 12328
rect 18104 12316 18110 12368
rect 14645 12291 14703 12297
rect 14645 12288 14657 12291
rect 12176 12260 14657 12288
rect 14645 12257 14657 12260
rect 14691 12288 14703 12291
rect 15105 12291 15163 12297
rect 14691 12260 14964 12288
rect 14691 12257 14703 12260
rect 14645 12251 14703 12257
rect 11885 12223 11943 12229
rect 11885 12189 11897 12223
rect 11931 12189 11943 12223
rect 12258 12223 12316 12229
rect 12258 12220 12270 12223
rect 11885 12183 11943 12189
rect 11992 12192 12270 12220
rect 11992 12152 12020 12192
rect 12258 12189 12270 12192
rect 12304 12189 12316 12223
rect 12258 12183 12316 12189
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12621 12223 12679 12229
rect 12621 12220 12633 12223
rect 12492 12192 12633 12220
rect 12492 12180 12498 12192
rect 12621 12189 12633 12192
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 14550 12220 14556 12232
rect 14323 12192 14556 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 14826 12220 14832 12232
rect 14787 12192 14832 12220
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 14936 12220 14964 12260
rect 15105 12257 15117 12291
rect 15151 12288 15163 12291
rect 15470 12288 15476 12300
rect 15151 12260 15476 12288
rect 15151 12257 15163 12260
rect 15105 12251 15163 12257
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 18156 12297 18184 12396
rect 18417 12393 18429 12427
rect 18463 12424 18475 12427
rect 19518 12424 19524 12436
rect 18463 12396 19524 12424
rect 18463 12393 18475 12396
rect 18417 12387 18475 12393
rect 19518 12384 19524 12396
rect 19576 12384 19582 12436
rect 21453 12427 21511 12433
rect 21453 12393 21465 12427
rect 21499 12424 21511 12427
rect 21542 12424 21548 12436
rect 21499 12396 21548 12424
rect 21499 12393 21511 12396
rect 21453 12387 21511 12393
rect 21542 12384 21548 12396
rect 21600 12424 21606 12436
rect 22094 12424 22100 12436
rect 21600 12396 22100 12424
rect 21600 12384 21606 12396
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 18322 12316 18328 12368
rect 18380 12356 18386 12368
rect 18380 12328 18460 12356
rect 18380 12316 18386 12328
rect 18141 12291 18199 12297
rect 18141 12257 18153 12291
rect 18187 12257 18199 12291
rect 18141 12251 18199 12257
rect 14994 12223 15052 12229
rect 14994 12220 15006 12223
rect 14936 12192 15006 12220
rect 14994 12189 15006 12192
rect 15040 12189 15052 12223
rect 15194 12220 15200 12232
rect 15155 12192 15200 12220
rect 14994 12183 15052 12189
rect 15194 12180 15200 12192
rect 15252 12180 15258 12232
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12189 15439 12223
rect 15654 12220 15660 12232
rect 15615 12192 15660 12220
rect 15381 12183 15439 12189
rect 11624 12124 12020 12152
rect 12069 12155 12127 12161
rect 11624 12096 11652 12124
rect 12069 12121 12081 12155
rect 12115 12121 12127 12155
rect 12069 12115 12127 12121
rect 12161 12155 12219 12161
rect 12161 12121 12173 12155
rect 12207 12152 12219 12155
rect 12986 12152 12992 12164
rect 12207 12124 12992 12152
rect 12207 12121 12219 12124
rect 12161 12115 12219 12121
rect 11606 12084 11612 12096
rect 9732 12056 11192 12084
rect 11567 12056 11612 12084
rect 9732 12044 9738 12056
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 12084 12084 12112 12115
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 12618 12084 12624 12096
rect 12084 12056 12624 12084
rect 12618 12044 12624 12056
rect 12676 12084 12682 12096
rect 13170 12084 13176 12096
rect 12676 12056 13176 12084
rect 12676 12044 12682 12056
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 15396 12084 15424 12183
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 17770 12220 17776 12232
rect 17731 12192 17776 12220
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 17862 12180 17868 12232
rect 17920 12220 17926 12232
rect 17956 12223 18014 12229
rect 17956 12220 17968 12223
rect 17920 12192 17968 12220
rect 17920 12180 17926 12192
rect 17956 12189 17968 12192
rect 18002 12189 18014 12223
rect 17956 12183 18014 12189
rect 18046 12180 18052 12232
rect 18104 12220 18110 12232
rect 18298 12223 18356 12229
rect 18104 12192 18149 12220
rect 18104 12180 18110 12192
rect 18298 12189 18310 12223
rect 18344 12217 18356 12223
rect 18432 12217 18460 12328
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 19334 12288 19340 12300
rect 19300 12260 19340 12288
rect 19300 12248 19306 12260
rect 19334 12248 19340 12260
rect 19392 12288 19398 12300
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 19392 12260 19441 12288
rect 19392 12248 19398 12260
rect 19429 12257 19441 12260
rect 19475 12288 19487 12291
rect 20070 12288 20076 12300
rect 19475 12260 20076 12288
rect 19475 12257 19487 12260
rect 19429 12251 19487 12257
rect 20070 12248 20076 12260
rect 20128 12248 20134 12300
rect 23382 12288 23388 12300
rect 22848 12260 23388 12288
rect 18344 12189 18460 12217
rect 18298 12183 18356 12189
rect 22738 12180 22744 12232
rect 22796 12220 22802 12232
rect 22848 12229 22876 12260
rect 23382 12248 23388 12260
rect 23440 12288 23446 12300
rect 24581 12291 24639 12297
rect 24581 12288 24593 12291
rect 23440 12260 24593 12288
rect 23440 12248 23446 12260
rect 24581 12257 24593 12260
rect 24627 12257 24639 12291
rect 24581 12251 24639 12257
rect 22833 12223 22891 12229
rect 22833 12220 22845 12223
rect 22796 12192 22845 12220
rect 22796 12180 22802 12192
rect 22833 12189 22845 12192
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 22922 12180 22928 12232
rect 22980 12220 22986 12232
rect 23109 12223 23167 12229
rect 23109 12220 23121 12223
rect 22980 12192 23121 12220
rect 22980 12180 22986 12192
rect 23109 12189 23121 12192
rect 23155 12220 23167 12223
rect 23293 12223 23351 12229
rect 23293 12220 23305 12223
rect 23155 12192 23305 12220
rect 23155 12189 23167 12192
rect 23109 12183 23167 12189
rect 23293 12189 23305 12192
rect 23339 12189 23351 12223
rect 23566 12220 23572 12232
rect 23527 12192 23572 12220
rect 23293 12183 23351 12189
rect 23566 12180 23572 12192
rect 23624 12180 23630 12232
rect 23842 12220 23848 12232
rect 23803 12192 23848 12220
rect 23842 12180 23848 12192
rect 23900 12180 23906 12232
rect 23989 12223 24047 12229
rect 23989 12189 24001 12223
rect 24035 12220 24047 12223
rect 24394 12220 24400 12232
rect 24035 12192 24400 12220
rect 24035 12189 24072 12192
rect 23989 12183 24072 12189
rect 15565 12155 15623 12161
rect 15565 12121 15577 12155
rect 15611 12152 15623 12155
rect 15902 12155 15960 12161
rect 15902 12152 15914 12155
rect 15611 12124 15914 12152
rect 15611 12121 15623 12124
rect 15565 12115 15623 12121
rect 15902 12121 15914 12124
rect 15948 12121 15960 12155
rect 17788 12152 17816 12180
rect 17788 12124 18092 12152
rect 15902 12115 15960 12121
rect 17034 12084 17040 12096
rect 15396 12056 17040 12084
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 17494 12044 17500 12096
rect 17552 12084 17558 12096
rect 17589 12087 17647 12093
rect 17589 12084 17601 12087
rect 17552 12056 17601 12084
rect 17552 12044 17558 12056
rect 17589 12053 17601 12056
rect 17635 12084 17647 12087
rect 17862 12084 17868 12096
rect 17635 12056 17868 12084
rect 17635 12053 17647 12056
rect 17589 12047 17647 12053
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 18064 12084 18092 12124
rect 18598 12112 18604 12164
rect 18656 12152 18662 12164
rect 19705 12155 19763 12161
rect 19705 12152 19717 12155
rect 18656 12124 19717 12152
rect 18656 12112 18662 12124
rect 19705 12121 19717 12124
rect 19751 12121 19763 12155
rect 19705 12115 19763 12121
rect 20438 12112 20444 12164
rect 20496 12112 20502 12164
rect 22370 12112 22376 12164
rect 22428 12152 22434 12164
rect 22566 12155 22624 12161
rect 22566 12152 22578 12155
rect 22428 12124 22578 12152
rect 22428 12112 22434 12124
rect 22566 12121 22578 12124
rect 22612 12121 22624 12155
rect 22566 12115 22624 12121
rect 23658 12112 23664 12164
rect 23716 12152 23722 12164
rect 23753 12155 23811 12161
rect 23753 12152 23765 12155
rect 23716 12124 23765 12152
rect 23716 12112 23722 12124
rect 23753 12121 23765 12124
rect 23799 12121 23811 12155
rect 24044 12152 24072 12183
rect 24394 12180 24400 12192
rect 24452 12180 24458 12232
rect 23753 12115 23811 12121
rect 23952 12124 24072 12152
rect 24138 12155 24196 12161
rect 18138 12084 18144 12096
rect 18064 12056 18144 12084
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 20990 12084 20996 12096
rect 18288 12056 20996 12084
rect 18288 12044 18294 12056
rect 20990 12044 20996 12056
rect 21048 12044 21054 12096
rect 21174 12084 21180 12096
rect 21135 12056 21180 12084
rect 21174 12044 21180 12056
rect 21232 12044 21238 12096
rect 22186 12044 22192 12096
rect 22244 12084 22250 12096
rect 22925 12087 22983 12093
rect 22925 12084 22937 12087
rect 22244 12056 22937 12084
rect 22244 12044 22250 12056
rect 22925 12053 22937 12056
rect 22971 12053 22983 12087
rect 22925 12047 22983 12053
rect 23477 12087 23535 12093
rect 23477 12053 23489 12087
rect 23523 12084 23535 12087
rect 23952 12084 23980 12124
rect 24138 12121 24150 12155
rect 24184 12152 24196 12155
rect 24826 12155 24884 12161
rect 24826 12152 24838 12155
rect 24184 12124 24838 12152
rect 24184 12121 24196 12124
rect 24138 12115 24196 12121
rect 24826 12121 24838 12124
rect 24872 12121 24884 12155
rect 24826 12115 24884 12121
rect 23523 12056 23980 12084
rect 23523 12053 23535 12056
rect 23477 12047 23535 12053
rect 24026 12044 24032 12096
rect 24084 12084 24090 12096
rect 24489 12087 24547 12093
rect 24489 12084 24501 12087
rect 24084 12056 24501 12084
rect 24084 12044 24090 12056
rect 24489 12053 24501 12056
rect 24535 12084 24547 12087
rect 25961 12087 26019 12093
rect 25961 12084 25973 12087
rect 24535 12056 25973 12084
rect 24535 12053 24547 12056
rect 24489 12047 24547 12053
rect 25961 12053 25973 12056
rect 26007 12053 26019 12087
rect 25961 12047 26019 12053
rect 1104 11994 29440 12016
rect 1104 11942 10395 11994
rect 10447 11942 10459 11994
rect 10511 11942 10523 11994
rect 10575 11942 10587 11994
rect 10639 11942 10651 11994
rect 10703 11942 19840 11994
rect 19892 11942 19904 11994
rect 19956 11942 19968 11994
rect 20020 11942 20032 11994
rect 20084 11942 20096 11994
rect 20148 11942 29440 11994
rect 1104 11920 29440 11942
rect 1946 11880 1952 11892
rect 1907 11852 1952 11880
rect 1946 11840 1952 11852
rect 2004 11840 2010 11892
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 2777 11883 2835 11889
rect 2777 11880 2789 11883
rect 2363 11852 2789 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 2777 11849 2789 11852
rect 2823 11849 2835 11883
rect 2777 11843 2835 11849
rect 3973 11883 4031 11889
rect 3973 11849 3985 11883
rect 4019 11880 4031 11883
rect 4062 11880 4068 11892
rect 4019 11852 4068 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 5994 11880 6000 11892
rect 5644 11852 6000 11880
rect 4982 11812 4988 11824
rect 4540 11784 4988 11812
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2774 11744 2780 11756
rect 2455 11716 2780 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 2958 11744 2964 11756
rect 2919 11716 2964 11744
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 3786 11744 3792 11756
rect 3747 11716 3792 11744
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 4540 11753 4568 11784
rect 4982 11772 4988 11784
rect 5040 11772 5046 11824
rect 4505 11747 4568 11753
rect 4505 11713 4517 11747
rect 4551 11716 4568 11747
rect 4551 11713 4563 11716
rect 4505 11707 4563 11713
rect 4614 11704 4620 11756
rect 4672 11744 4678 11756
rect 5644 11753 5672 11852
rect 5994 11840 6000 11852
rect 6052 11880 6058 11892
rect 8754 11880 8760 11892
rect 6052 11852 8760 11880
rect 6052 11840 6058 11852
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 9214 11880 9220 11892
rect 9048 11852 9220 11880
rect 6730 11812 6736 11824
rect 6380 11784 6736 11812
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4672 11716 4905 11744
rect 4672 11704 4678 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 4154 11676 4160 11688
rect 2639 11648 4160 11676
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 6380 11685 6408 11784
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 8846 11812 8852 11824
rect 8807 11784 8852 11812
rect 8846 11772 8852 11784
rect 8904 11772 8910 11824
rect 9048 11821 9076 11852
rect 9214 11840 9220 11852
rect 9272 11880 9278 11892
rect 9309 11883 9367 11889
rect 9309 11880 9321 11883
rect 9272 11852 9321 11880
rect 9272 11840 9278 11852
rect 9309 11849 9321 11852
rect 9355 11880 9367 11883
rect 15010 11880 15016 11892
rect 9355 11852 15016 11880
rect 9355 11849 9367 11852
rect 9309 11843 9367 11849
rect 15010 11840 15016 11852
rect 15068 11840 15074 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15252 11852 15608 11880
rect 15252 11840 15258 11852
rect 9033 11815 9091 11821
rect 9033 11781 9045 11815
rect 9079 11781 9091 11815
rect 11606 11812 11612 11824
rect 9033 11775 9091 11781
rect 9968 11784 10916 11812
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 6621 11747 6679 11753
rect 6621 11744 6633 11747
rect 6512 11716 6633 11744
rect 6512 11704 6518 11716
rect 6621 11713 6633 11716
rect 6667 11713 6679 11747
rect 6621 11707 6679 11713
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 9968 11744 9996 11784
rect 7800 11716 9996 11744
rect 10045 11747 10103 11753
rect 7800 11704 7806 11716
rect 10045 11713 10057 11747
rect 10091 11744 10103 11747
rect 10134 11744 10140 11756
rect 10091 11716 10140 11744
rect 10091 11713 10103 11716
rect 10045 11707 10103 11713
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 10244 11716 10425 11744
rect 6365 11679 6423 11685
rect 6365 11676 6377 11679
rect 5592 11648 6377 11676
rect 5592 11636 5598 11648
rect 6365 11645 6377 11648
rect 6411 11645 6423 11679
rect 6365 11639 6423 11645
rect 3418 11568 3424 11620
rect 3476 11608 3482 11620
rect 10244 11617 10272 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 4341 11611 4399 11617
rect 4341 11608 4353 11611
rect 3476 11580 4353 11608
rect 3476 11568 3482 11580
rect 4341 11577 4353 11580
rect 4387 11577 4399 11611
rect 10229 11611 10287 11617
rect 4341 11571 4399 11577
rect 4448 11580 5672 11608
rect 3878 11500 3884 11552
rect 3936 11540 3942 11552
rect 4448 11540 4476 11580
rect 3936 11512 4476 11540
rect 3936 11500 3942 11512
rect 5166 11500 5172 11552
rect 5224 11540 5230 11552
rect 5537 11543 5595 11549
rect 5537 11540 5549 11543
rect 5224 11512 5549 11540
rect 5224 11500 5230 11512
rect 5537 11509 5549 11512
rect 5583 11509 5595 11543
rect 5644 11540 5672 11580
rect 7300 11580 7880 11608
rect 7300 11540 7328 11580
rect 7742 11540 7748 11552
rect 5644 11512 7328 11540
rect 7703 11512 7748 11540
rect 5537 11503 5595 11509
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 7852 11540 7880 11580
rect 10229 11577 10241 11611
rect 10275 11577 10287 11611
rect 10229 11571 10287 11577
rect 10410 11540 10416 11552
rect 7852 11512 10416 11540
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 10594 11540 10600 11552
rect 10555 11512 10600 11540
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 10778 11540 10784 11552
rect 10739 11512 10784 11540
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 10888 11540 10916 11784
rect 10980 11784 11612 11812
rect 10980 11753 11008 11784
rect 11606 11772 11612 11784
rect 11664 11772 11670 11824
rect 12802 11812 12808 11824
rect 12728 11784 12808 11812
rect 10960 11747 11018 11753
rect 10960 11713 10972 11747
rect 11006 11713 11018 11747
rect 10960 11707 11018 11713
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11713 11115 11747
rect 11057 11707 11115 11713
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11713 11207 11747
rect 11330 11744 11336 11756
rect 11291 11716 11336 11744
rect 11149 11707 11207 11713
rect 11072 11608 11100 11707
rect 11164 11676 11192 11707
rect 11330 11704 11336 11716
rect 11388 11704 11394 11756
rect 11974 11704 11980 11756
rect 12032 11744 12038 11756
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 12032 11716 12173 11744
rect 12032 11704 12038 11716
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12342 11744 12348 11756
rect 12303 11716 12348 11744
rect 12161 11707 12219 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 12581 11747 12639 11753
rect 12581 11713 12593 11747
rect 12627 11744 12639 11747
rect 12728 11744 12756 11784
rect 12802 11772 12808 11784
rect 12860 11772 12866 11824
rect 13906 11772 13912 11824
rect 13964 11772 13970 11824
rect 15470 11812 15476 11824
rect 15396 11784 15476 11812
rect 12894 11744 12900 11756
rect 12627 11716 12756 11744
rect 12855 11716 12900 11744
rect 12627 11713 12639 11716
rect 12581 11707 12639 11713
rect 11609 11679 11667 11685
rect 11609 11676 11621 11679
rect 11164 11648 11621 11676
rect 11609 11645 11621 11648
rect 11655 11676 11667 11679
rect 12360 11676 12388 11704
rect 11655 11648 12388 11676
rect 12452 11676 12480 11707
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 14826 11704 14832 11756
rect 14884 11744 14890 11756
rect 15396 11753 15424 11784
rect 15470 11772 15476 11784
rect 15528 11772 15534 11824
rect 15105 11747 15163 11753
rect 15105 11744 15117 11747
rect 14884 11716 15117 11744
rect 14884 11704 14890 11716
rect 15105 11713 15117 11716
rect 15151 11713 15163 11747
rect 15105 11707 15163 11713
rect 15288 11747 15346 11753
rect 15288 11713 15300 11747
rect 15334 11713 15346 11747
rect 15288 11707 15346 11713
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 13173 11679 13231 11685
rect 13173 11676 13185 11679
rect 12452 11648 12572 11676
rect 11655 11645 11667 11648
rect 11609 11639 11667 11645
rect 11072 11580 11652 11608
rect 11624 11552 11652 11580
rect 11238 11540 11244 11552
rect 10888 11512 11244 11540
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11606 11500 11612 11552
rect 11664 11500 11670 11552
rect 12544 11540 12572 11648
rect 12728 11648 13185 11676
rect 12728 11617 12756 11648
rect 13173 11645 13185 11648
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 13814 11636 13820 11688
rect 13872 11676 13878 11688
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 13872 11648 14933 11676
rect 13872 11636 13878 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 12713 11611 12771 11617
rect 12713 11577 12725 11611
rect 12759 11577 12771 11611
rect 14936 11608 14964 11639
rect 15304 11608 15332 11707
rect 15580 11688 15608 11852
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 17405 11883 17463 11889
rect 17405 11880 17417 11883
rect 17368 11852 17417 11880
rect 17368 11840 17374 11852
rect 17405 11849 17417 11852
rect 17451 11849 17463 11883
rect 17405 11843 17463 11849
rect 17770 11840 17776 11892
rect 17828 11880 17834 11892
rect 18230 11880 18236 11892
rect 17828 11852 18236 11880
rect 17828 11840 17834 11852
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 19426 11880 19432 11892
rect 19387 11852 19432 11880
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 21542 11880 21548 11892
rect 21503 11852 21548 11880
rect 21542 11840 21548 11852
rect 21600 11840 21606 11892
rect 24486 11840 24492 11892
rect 24544 11840 24550 11892
rect 16390 11772 16396 11824
rect 16448 11812 16454 11824
rect 19797 11815 19855 11821
rect 19797 11812 19809 11815
rect 16448 11784 19809 11812
rect 16448 11772 16454 11784
rect 19797 11781 19809 11784
rect 19843 11781 19855 11815
rect 19797 11775 19855 11781
rect 21560 11812 21588 11840
rect 22097 11815 22155 11821
rect 22097 11812 22109 11815
rect 21560 11784 22109 11812
rect 15657 11747 15715 11753
rect 15657 11713 15669 11747
rect 15703 11744 15715 11747
rect 17126 11744 17132 11756
rect 15703 11716 17132 11744
rect 15703 11713 15715 11716
rect 15657 11707 15715 11713
rect 17126 11704 17132 11716
rect 17184 11744 17190 11756
rect 17773 11747 17831 11753
rect 17773 11744 17785 11747
rect 17184 11716 17785 11744
rect 17184 11704 17190 11716
rect 17773 11713 17785 11716
rect 17819 11713 17831 11747
rect 21560 11744 21588 11784
rect 22097 11781 22109 11784
rect 22143 11781 22155 11815
rect 24504 11812 24532 11840
rect 24734 11815 24792 11821
rect 24734 11812 24746 11815
rect 24504 11784 24746 11812
rect 22097 11775 22155 11781
rect 24734 11781 24746 11784
rect 24780 11781 24792 11815
rect 24734 11775 24792 11781
rect 21818 11744 21824 11756
rect 17773 11707 17831 11713
rect 21192 11716 21588 11744
rect 21779 11716 21824 11744
rect 15473 11679 15531 11685
rect 15473 11645 15485 11679
rect 15519 11676 15531 11679
rect 15562 11676 15568 11688
rect 15519 11648 15568 11676
rect 15519 11645 15531 11648
rect 15473 11639 15531 11645
rect 15562 11636 15568 11648
rect 15620 11676 15626 11688
rect 16666 11676 16672 11688
rect 15620 11648 16672 11676
rect 15620 11636 15626 11648
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 17862 11676 17868 11688
rect 17823 11648 17868 11676
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 17957 11679 18015 11685
rect 17957 11645 17969 11679
rect 18003 11676 18015 11679
rect 18414 11676 18420 11688
rect 18003 11648 18420 11676
rect 18003 11645 18015 11648
rect 17957 11639 18015 11645
rect 18414 11636 18420 11648
rect 18472 11676 18478 11688
rect 19886 11676 19892 11688
rect 18472 11648 18828 11676
rect 19847 11648 19892 11676
rect 18472 11636 18478 11648
rect 12713 11571 12771 11577
rect 14200 11580 14780 11608
rect 14936 11580 15332 11608
rect 15396 11580 16068 11608
rect 12986 11540 12992 11552
rect 12544 11512 12992 11540
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 14200 11540 14228 11580
rect 13228 11512 14228 11540
rect 13228 11500 13234 11512
rect 14550 11500 14556 11552
rect 14608 11540 14614 11552
rect 14645 11543 14703 11549
rect 14645 11540 14657 11543
rect 14608 11512 14657 11540
rect 14608 11500 14614 11512
rect 14645 11509 14657 11512
rect 14691 11509 14703 11543
rect 14752 11540 14780 11580
rect 15396 11540 15424 11580
rect 14752 11512 15424 11540
rect 15749 11543 15807 11549
rect 14645 11503 14703 11509
rect 15749 11509 15761 11543
rect 15795 11540 15807 11543
rect 15930 11540 15936 11552
rect 15795 11512 15936 11540
rect 15795 11509 15807 11512
rect 15749 11503 15807 11509
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 16040 11540 16068 11580
rect 16114 11568 16120 11620
rect 16172 11608 16178 11620
rect 17770 11608 17776 11620
rect 16172 11580 17776 11608
rect 16172 11568 16178 11580
rect 17770 11568 17776 11580
rect 17828 11568 17834 11620
rect 18800 11608 18828 11648
rect 19886 11636 19892 11648
rect 19944 11636 19950 11688
rect 19981 11679 20039 11685
rect 19981 11645 19993 11679
rect 20027 11645 20039 11679
rect 19981 11639 20039 11645
rect 19996 11608 20024 11639
rect 17880 11580 18460 11608
rect 18800 11580 20024 11608
rect 17880 11540 17908 11580
rect 18322 11540 18328 11552
rect 16040 11512 17908 11540
rect 18283 11512 18328 11540
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 18432 11540 18460 11580
rect 21192 11540 21220 11716
rect 21818 11704 21824 11716
rect 21876 11704 21882 11756
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 22020 11676 22048 11707
rect 22186 11704 22192 11756
rect 22244 11753 22250 11756
rect 22244 11744 22252 11753
rect 22557 11747 22615 11753
rect 22244 11716 22289 11744
rect 22244 11707 22252 11716
rect 22557 11713 22569 11747
rect 22603 11744 22615 11747
rect 22646 11744 22652 11756
rect 22603 11716 22652 11744
rect 22603 11713 22615 11716
rect 22557 11707 22615 11713
rect 22244 11704 22250 11707
rect 22646 11704 22652 11716
rect 22704 11704 22710 11756
rect 22824 11747 22882 11753
rect 22824 11713 22836 11747
rect 22870 11744 22882 11747
rect 23198 11744 23204 11756
rect 22870 11716 23204 11744
rect 22870 11713 22882 11716
rect 22824 11707 22882 11713
rect 23198 11704 23204 11716
rect 23256 11704 23262 11756
rect 23382 11704 23388 11756
rect 23440 11744 23446 11756
rect 24489 11747 24547 11753
rect 24489 11744 24501 11747
rect 23440 11716 24501 11744
rect 23440 11704 23446 11716
rect 24489 11713 24501 11716
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 21376 11648 22048 11676
rect 21376 11552 21404 11648
rect 22370 11608 22376 11620
rect 22331 11580 22376 11608
rect 22370 11568 22376 11580
rect 22428 11568 22434 11620
rect 21358 11540 21364 11552
rect 18432 11512 21220 11540
rect 21319 11512 21364 11540
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 23934 11540 23940 11552
rect 23895 11512 23940 11540
rect 23934 11500 23940 11512
rect 23992 11500 23998 11552
rect 25406 11500 25412 11552
rect 25464 11540 25470 11552
rect 25866 11540 25872 11552
rect 25464 11512 25872 11540
rect 25464 11500 25470 11512
rect 25866 11500 25872 11512
rect 25924 11500 25930 11552
rect 1104 11450 29440 11472
rect 1104 11398 5672 11450
rect 5724 11398 5736 11450
rect 5788 11398 5800 11450
rect 5852 11398 5864 11450
rect 5916 11398 5928 11450
rect 5980 11398 15118 11450
rect 15170 11398 15182 11450
rect 15234 11398 15246 11450
rect 15298 11398 15310 11450
rect 15362 11398 15374 11450
rect 15426 11398 24563 11450
rect 24615 11398 24627 11450
rect 24679 11398 24691 11450
rect 24743 11398 24755 11450
rect 24807 11398 24819 11450
rect 24871 11398 29440 11450
rect 1104 11376 29440 11398
rect 2593 11339 2651 11345
rect 2593 11305 2605 11339
rect 2639 11336 2651 11339
rect 2682 11336 2688 11348
rect 2639 11308 2688 11336
rect 2639 11305 2651 11308
rect 2593 11299 2651 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 4798 11296 4804 11348
rect 4856 11336 4862 11348
rect 4985 11339 5043 11345
rect 4985 11336 4997 11339
rect 4856 11308 4997 11336
rect 4856 11296 4862 11308
rect 4985 11305 4997 11308
rect 5031 11305 5043 11339
rect 4985 11299 5043 11305
rect 6362 11296 6368 11348
rect 6420 11336 6426 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6420 11308 6745 11336
rect 6420 11296 6426 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 6733 11299 6791 11305
rect 7101 11339 7159 11345
rect 7101 11305 7113 11339
rect 7147 11336 7159 11339
rect 7282 11336 7288 11348
rect 7147 11308 7288 11336
rect 7147 11305 7159 11308
rect 7101 11299 7159 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 10032 11339 10090 11345
rect 10032 11305 10044 11339
rect 10078 11336 10090 11339
rect 10778 11336 10784 11348
rect 10078 11308 10784 11336
rect 10078 11305 10090 11308
rect 10032 11299 10090 11305
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 12161 11339 12219 11345
rect 12161 11336 12173 11339
rect 12032 11308 12173 11336
rect 12032 11296 12038 11308
rect 12161 11305 12173 11308
rect 12207 11305 12219 11339
rect 13906 11336 13912 11348
rect 13867 11308 13912 11336
rect 12161 11299 12219 11305
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 16114 11336 16120 11348
rect 14016 11308 16120 11336
rect 6638 11228 6644 11280
rect 6696 11268 6702 11280
rect 7469 11271 7527 11277
rect 7469 11268 7481 11271
rect 6696 11240 7481 11268
rect 6696 11228 6702 11240
rect 7469 11237 7481 11240
rect 7515 11237 7527 11271
rect 7469 11231 7527 11237
rect 9125 11271 9183 11277
rect 9125 11237 9137 11271
rect 9171 11237 9183 11271
rect 9125 11231 9183 11237
rect 9493 11271 9551 11277
rect 9493 11237 9505 11271
rect 9539 11268 9551 11271
rect 9674 11268 9680 11280
rect 9539 11240 9680 11268
rect 9539 11237 9551 11240
rect 9493 11231 9551 11237
rect 5994 11200 6000 11212
rect 3804 11172 6000 11200
rect 3804 11141 3832 11172
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 2271 11104 3801 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3789 11095 3847 11101
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 5166 11132 5172 11144
rect 5127 11104 5172 11132
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 5552 11141 5580 11172
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 7742 11200 7748 11212
rect 6748 11172 7748 11200
rect 5537 11135 5595 11141
rect 5537 11101 5549 11135
rect 5583 11101 5595 11135
rect 5537 11095 5595 11101
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11132 5779 11135
rect 6362 11132 6368 11144
rect 5767 11104 6368 11132
rect 5767 11101 5779 11104
rect 5721 11095 5779 11101
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 6748 11141 6776 11172
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11132 6883 11135
rect 7285 11135 7343 11141
rect 7285 11132 7297 11135
rect 6871 11104 7297 11132
rect 6871 11101 6883 11104
rect 6825 11095 6883 11101
rect 7285 11101 7297 11104
rect 7331 11101 7343 11135
rect 7285 11095 7343 11101
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11101 8999 11135
rect 9140 11132 9168 11231
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 11238 11228 11244 11280
rect 11296 11268 11302 11280
rect 11296 11240 11744 11268
rect 11296 11228 11302 11240
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11200 9827 11203
rect 10042 11200 10048 11212
rect 9815 11172 10048 11200
rect 9815 11169 9827 11172
rect 9769 11163 9827 11169
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10410 11160 10416 11212
rect 10468 11200 10474 11212
rect 11517 11203 11575 11209
rect 10468 11172 11376 11200
rect 10468 11160 10474 11172
rect 9401 11135 9459 11141
rect 9401 11132 9413 11135
rect 9140 11104 9413 11132
rect 8941 11095 8999 11101
rect 9401 11101 9413 11104
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 1394 11024 1400 11076
rect 1452 11064 1458 11076
rect 2041 11067 2099 11073
rect 2041 11064 2053 11067
rect 1452 11036 2053 11064
rect 1452 11024 1458 11036
rect 2041 11033 2053 11036
rect 2087 11033 2099 11067
rect 2406 11064 2412 11076
rect 2367 11036 2412 11064
rect 2041 11027 2099 11033
rect 2406 11024 2412 11036
rect 2464 11024 2470 11076
rect 5184 11064 5212 11092
rect 6840 11064 6868 11095
rect 5184 11036 6868 11064
rect 8956 11064 8984 11095
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9640 11104 9689 11132
rect 9640 11092 9646 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 10134 11064 10140 11076
rect 8956 11036 10140 11064
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 10594 11024 10600 11076
rect 10652 11024 10658 11076
rect 11348 11064 11376 11172
rect 11517 11169 11529 11203
rect 11563 11200 11575 11203
rect 11606 11200 11612 11212
rect 11563 11172 11612 11200
rect 11563 11169 11575 11172
rect 11517 11163 11575 11169
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 11716 11200 11744 11240
rect 12342 11228 12348 11280
rect 12400 11268 12406 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 12400 11240 13185 11268
rect 12400 11228 12406 11240
rect 13173 11237 13185 11240
rect 13219 11268 13231 11271
rect 14016 11268 14044 11308
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 17126 11336 17132 11348
rect 17087 11308 17132 11336
rect 17126 11296 17132 11308
rect 17184 11296 17190 11348
rect 17236 11308 19288 11336
rect 13219 11240 14044 11268
rect 14093 11271 14151 11277
rect 13219 11237 13231 11240
rect 13173 11231 13231 11237
rect 14093 11237 14105 11271
rect 14139 11237 14151 11271
rect 15470 11268 15476 11280
rect 14093 11231 14151 11237
rect 15212 11240 15476 11268
rect 13906 11200 13912 11212
rect 11716 11172 13912 11200
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 12342 11132 12348 11144
rect 12303 11104 12348 11132
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 14108 11132 14136 11231
rect 15212 11209 15240 11240
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 15197 11203 15255 11209
rect 15197 11169 15209 11203
rect 15243 11169 15255 11203
rect 15197 11163 15255 11169
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15562 11200 15568 11212
rect 15335 11172 15568 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 15654 11160 15660 11212
rect 15712 11200 15718 11212
rect 15749 11203 15807 11209
rect 15749 11200 15761 11203
rect 15712 11172 15761 11200
rect 15712 11160 15718 11172
rect 15749 11169 15761 11172
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 14274 11132 14280 11144
rect 13771 11104 14136 11132
rect 14235 11104 14280 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14826 11092 14832 11144
rect 14884 11132 14890 11144
rect 14921 11135 14979 11141
rect 14921 11132 14933 11135
rect 14884 11104 14933 11132
rect 14884 11092 14890 11104
rect 14921 11101 14933 11104
rect 14967 11101 14979 11135
rect 15086 11135 15144 11141
rect 15086 11132 15098 11135
rect 14921 11095 14979 11101
rect 15028 11104 15098 11132
rect 14737 11067 14795 11073
rect 14737 11064 14749 11067
rect 11348 11036 14749 11064
rect 14737 11033 14749 11036
rect 14783 11064 14795 11067
rect 15028 11064 15056 11104
rect 15086 11101 15098 11104
rect 15132 11101 15144 11135
rect 15086 11095 15144 11101
rect 15473 11135 15531 11141
rect 15473 11101 15485 11135
rect 15519 11132 15531 11135
rect 15764 11132 15792 11163
rect 17236 11132 17264 11308
rect 17678 11228 17684 11280
rect 17736 11268 17742 11280
rect 17736 11240 18552 11268
rect 17736 11228 17742 11240
rect 17586 11200 17592 11212
rect 17547 11172 17592 11200
rect 17586 11160 17592 11172
rect 17644 11200 17650 11212
rect 18524 11209 18552 11240
rect 19260 11212 19288 11308
rect 19886 11296 19892 11348
rect 19944 11336 19950 11348
rect 20625 11339 20683 11345
rect 20625 11336 20637 11339
rect 19944 11308 20637 11336
rect 19944 11296 19950 11308
rect 20625 11305 20637 11308
rect 20671 11305 20683 11339
rect 20625 11299 20683 11305
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 26234 11336 26240 11348
rect 21232 11308 26240 11336
rect 21232 11296 21238 11308
rect 26234 11296 26240 11308
rect 26292 11296 26298 11348
rect 18417 11203 18475 11209
rect 18417 11200 18429 11203
rect 17644 11172 18429 11200
rect 17644 11160 17650 11172
rect 18417 11169 18429 11172
rect 18463 11169 18475 11203
rect 18417 11163 18475 11169
rect 18509 11203 18567 11209
rect 18509 11169 18521 11203
rect 18555 11169 18567 11203
rect 19242 11200 19248 11212
rect 19155 11172 19248 11200
rect 18509 11163 18567 11169
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 15519 11104 15700 11132
rect 15764 11104 17264 11132
rect 17313 11135 17371 11141
rect 15519 11101 15531 11104
rect 15473 11095 15531 11101
rect 14783 11036 15056 11064
rect 14783 11033 14795 11036
rect 14737 11027 14795 11033
rect 4065 10999 4123 11005
rect 4065 10965 4077 10999
rect 4111 10996 4123 10999
rect 4246 10996 4252 11008
rect 4111 10968 4252 10996
rect 4111 10965 4123 10968
rect 4065 10959 4123 10965
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 5718 10996 5724 11008
rect 5679 10968 5724 10996
rect 5718 10956 5724 10968
rect 5776 10956 5782 11008
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9217 10999 9275 11005
rect 9217 10996 9229 10999
rect 9180 10968 9229 10996
rect 9180 10956 9186 10968
rect 9217 10965 9229 10968
rect 9263 10965 9275 10999
rect 12986 10996 12992 11008
rect 12899 10968 12992 10996
rect 9217 10959 9275 10965
rect 12986 10956 12992 10968
rect 13044 10996 13050 11008
rect 14550 10996 14556 11008
rect 13044 10968 14556 10996
rect 13044 10956 13050 10968
rect 14550 10956 14556 10968
rect 14608 10956 14614 11008
rect 15562 10996 15568 11008
rect 15523 10968 15568 10996
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 15672 10996 15700 11104
rect 17313 11101 17325 11135
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 15930 11024 15936 11076
rect 15988 11073 15994 11076
rect 15988 11067 16052 11073
rect 15988 11033 16006 11067
rect 16040 11033 16052 11067
rect 17328 11064 17356 11095
rect 17402 11092 17408 11144
rect 17460 11141 17466 11144
rect 17460 11135 17519 11141
rect 17460 11101 17473 11135
rect 17507 11101 17519 11135
rect 17678 11132 17684 11144
rect 17639 11104 17684 11132
rect 17460 11095 17519 11101
rect 17460 11092 17466 11095
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 17862 11132 17868 11144
rect 17823 11104 17868 11132
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 18138 11132 18144 11144
rect 18064 11106 18144 11132
rect 17972 11104 18144 11106
rect 17972 11078 18092 11104
rect 18138 11092 18144 11104
rect 18196 11092 18202 11144
rect 18322 11092 18328 11144
rect 18380 11132 18386 11144
rect 18693 11135 18751 11141
rect 18380 11104 18424 11132
rect 18380 11092 18386 11104
rect 18693 11101 18705 11135
rect 18739 11132 18751 11135
rect 19886 11132 19892 11144
rect 18739 11104 19892 11132
rect 18739 11101 18751 11104
rect 18693 11095 18751 11101
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 17972 11064 18000 11078
rect 17328 11036 18000 11064
rect 18877 11067 18935 11073
rect 15988 11027 16052 11033
rect 18877 11033 18889 11067
rect 18923 11064 18935 11067
rect 19490 11067 19548 11073
rect 19490 11064 19502 11067
rect 18923 11036 19502 11064
rect 18923 11033 18935 11036
rect 18877 11027 18935 11033
rect 19490 11033 19502 11036
rect 19536 11033 19548 11067
rect 19490 11027 19548 11033
rect 15988 11024 15994 11027
rect 16390 10996 16396 11008
rect 15672 10968 16396 10996
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 17954 10996 17960 11008
rect 17915 10968 17960 10996
rect 17954 10956 17960 10968
rect 18012 10956 18018 11008
rect 1104 10906 29440 10928
rect 1104 10854 10395 10906
rect 10447 10854 10459 10906
rect 10511 10854 10523 10906
rect 10575 10854 10587 10906
rect 10639 10854 10651 10906
rect 10703 10854 19840 10906
rect 19892 10854 19904 10906
rect 19956 10854 19968 10906
rect 20020 10854 20032 10906
rect 20084 10854 20096 10906
rect 20148 10854 29440 10906
rect 1104 10832 29440 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 2133 10795 2191 10801
rect 2133 10792 2145 10795
rect 1627 10764 2145 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 2133 10761 2145 10764
rect 2179 10761 2191 10795
rect 2133 10755 2191 10761
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 2464 10764 2513 10792
rect 2464 10752 2470 10764
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 2501 10755 2559 10761
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 3234 10792 3240 10804
rect 2915 10764 3240 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 3234 10752 3240 10764
rect 3292 10792 3298 10804
rect 3970 10792 3976 10804
rect 3292 10764 3976 10792
rect 3292 10752 3298 10764
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 5537 10795 5595 10801
rect 5537 10761 5549 10795
rect 5583 10792 5595 10795
rect 5718 10792 5724 10804
rect 5583 10764 5724 10792
rect 5583 10761 5595 10764
rect 5537 10755 5595 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12342 10792 12348 10804
rect 12299 10764 12348 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12342 10752 12348 10764
rect 12400 10792 12406 10804
rect 16390 10792 16396 10804
rect 12400 10752 12434 10792
rect 16351 10764 16396 10792
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 17862 10752 17868 10804
rect 17920 10792 17926 10804
rect 18785 10795 18843 10801
rect 18785 10792 18797 10795
rect 17920 10764 18797 10792
rect 17920 10752 17926 10764
rect 18785 10761 18797 10764
rect 18831 10761 18843 10795
rect 18785 10755 18843 10761
rect 22462 10752 22468 10804
rect 22520 10792 22526 10804
rect 22649 10795 22707 10801
rect 22649 10792 22661 10795
rect 22520 10764 22661 10792
rect 22520 10752 22526 10764
rect 22649 10761 22661 10764
rect 22695 10761 22707 10795
rect 22649 10755 22707 10761
rect 2041 10727 2099 10733
rect 2041 10693 2053 10727
rect 2087 10724 2099 10727
rect 2424 10724 2452 10752
rect 5629 10727 5687 10733
rect 5629 10724 5641 10727
rect 2087 10696 2452 10724
rect 4908 10696 5641 10724
rect 2087 10693 2099 10696
rect 2041 10687 2099 10693
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2372 10628 2697 10656
rect 2372 10616 2378 10628
rect 2685 10625 2697 10628
rect 2731 10625 2743 10659
rect 3970 10656 3976 10668
rect 4028 10665 4034 10668
rect 3940 10628 3976 10656
rect 2685 10619 2743 10625
rect 3970 10616 3976 10628
rect 4028 10619 4040 10665
rect 4614 10656 4620 10668
rect 4575 10628 4620 10656
rect 4028 10616 4034 10619
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 4908 10665 4936 10696
rect 5629 10693 5641 10696
rect 5675 10724 5687 10727
rect 6457 10727 6515 10733
rect 6457 10724 6469 10727
rect 5675 10696 6469 10724
rect 5675 10693 5687 10696
rect 5629 10687 5687 10693
rect 6457 10693 6469 10696
rect 6503 10693 6515 10727
rect 9122 10724 9128 10736
rect 9062 10696 9128 10724
rect 6457 10687 6515 10693
rect 9122 10684 9128 10696
rect 9180 10684 9186 10736
rect 9953 10727 10011 10733
rect 9953 10693 9965 10727
rect 9999 10724 10011 10727
rect 12406 10724 12434 10752
rect 17672 10727 17730 10733
rect 9999 10696 10364 10724
rect 12406 10696 12940 10724
rect 9999 10693 10011 10696
rect 9953 10687 10011 10693
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10625 4951 10659
rect 6362 10656 6368 10668
rect 6323 10628 6368 10656
rect 4893 10619 4951 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 7561 10659 7619 10665
rect 7561 10656 7573 10659
rect 6788 10628 7573 10656
rect 6788 10616 6794 10628
rect 7561 10625 7573 10628
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 9674 10616 9680 10668
rect 9732 10665 9738 10668
rect 9732 10659 9775 10665
rect 9763 10625 9775 10659
rect 9732 10619 9775 10625
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10656 10195 10659
rect 10183 10628 10272 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 9732 10616 9738 10619
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2590 10588 2596 10600
rect 2271 10560 2596 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10557 4307 10591
rect 4522 10588 4528 10600
rect 4483 10560 4528 10588
rect 4249 10551 4307 10557
rect 1670 10412 1676 10464
rect 1728 10452 1734 10464
rect 4264 10452 4292 10551
rect 4522 10548 4528 10560
rect 4580 10548 4586 10600
rect 5445 10591 5503 10597
rect 5445 10557 5457 10591
rect 5491 10588 5503 10591
rect 7837 10591 7895 10597
rect 5491 10560 6224 10588
rect 5491 10557 5503 10560
rect 5445 10551 5503 10557
rect 5534 10452 5540 10464
rect 1728 10424 1773 10452
rect 4264 10424 5540 10452
rect 1728 10412 1734 10424
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 5994 10452 6000 10464
rect 5955 10424 6000 10452
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 6196 10461 6224 10560
rect 7837 10557 7849 10591
rect 7883 10588 7895 10591
rect 7883 10560 9628 10588
rect 7883 10557 7895 10560
rect 7837 10551 7895 10557
rect 9600 10529 9628 10560
rect 9585 10523 9643 10529
rect 9585 10489 9597 10523
rect 9631 10489 9643 10523
rect 9585 10483 9643 10489
rect 6181 10455 6239 10461
rect 6181 10421 6193 10455
rect 6227 10452 6239 10455
rect 6914 10452 6920 10464
rect 6227 10424 6920 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 9309 10455 9367 10461
rect 9309 10421 9321 10455
rect 9355 10452 9367 10455
rect 9398 10452 9404 10464
rect 9355 10424 9404 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 9398 10412 9404 10424
rect 9456 10452 9462 10464
rect 9876 10452 9904 10619
rect 10244 10461 10272 10628
rect 10336 10588 10364 10696
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10656 10471 10659
rect 11054 10656 11060 10668
rect 10459 10628 11060 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 12345 10659 12403 10665
rect 12345 10625 12357 10659
rect 12391 10656 12403 10659
rect 12434 10656 12440 10668
rect 12391 10628 12440 10656
rect 12391 10625 12403 10628
rect 12345 10619 12403 10625
rect 12434 10616 12440 10628
rect 12492 10656 12498 10668
rect 12912 10665 12940 10696
rect 15028 10696 17172 10724
rect 12621 10659 12679 10665
rect 12621 10656 12633 10659
rect 12492 10628 12633 10656
rect 12492 10616 12498 10628
rect 12621 10625 12633 10628
rect 12667 10625 12679 10659
rect 12621 10619 12679 10625
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 13633 10659 13691 10665
rect 13633 10625 13645 10659
rect 13679 10656 13691 10659
rect 14274 10656 14280 10668
rect 13679 10628 14280 10656
rect 13679 10625 13691 10628
rect 13633 10619 13691 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 15028 10665 15056 10696
rect 15013 10659 15071 10665
rect 15013 10625 15025 10659
rect 15059 10625 15071 10659
rect 15013 10619 15071 10625
rect 15280 10659 15338 10665
rect 15280 10625 15292 10659
rect 15326 10656 15338 10659
rect 15562 10656 15568 10668
rect 15326 10628 15568 10656
rect 15326 10625 15338 10628
rect 15280 10619 15338 10625
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 17144 10600 17172 10696
rect 17672 10693 17684 10727
rect 17718 10724 17730 10727
rect 17954 10724 17960 10736
rect 17718 10696 17960 10724
rect 17718 10693 17730 10696
rect 17672 10687 17730 10693
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 22480 10724 22508 10752
rect 22388 10696 22508 10724
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 20165 10659 20223 10665
rect 20165 10656 20177 10659
rect 19392 10628 20177 10656
rect 19392 10616 19398 10628
rect 20165 10625 20177 10628
rect 20211 10625 20223 10659
rect 20165 10619 20223 10625
rect 20432 10659 20490 10665
rect 20432 10625 20444 10659
rect 20478 10656 20490 10659
rect 21913 10659 21971 10665
rect 21913 10656 21925 10659
rect 20478 10628 21925 10656
rect 20478 10625 20490 10628
rect 20432 10619 20490 10625
rect 21913 10625 21925 10628
rect 21959 10625 21971 10659
rect 22094 10656 22100 10668
rect 22055 10628 22100 10656
rect 21913 10619 21971 10625
rect 22094 10616 22100 10628
rect 22152 10616 22158 10668
rect 22278 10665 22284 10668
rect 22235 10659 22284 10665
rect 22235 10625 22247 10659
rect 22281 10625 22284 10659
rect 22235 10619 22284 10625
rect 22278 10616 22284 10619
rect 22336 10616 22342 10668
rect 10336 10560 10640 10588
rect 9456 10424 9904 10452
rect 10229 10455 10287 10461
rect 9456 10412 9462 10424
rect 10229 10421 10241 10455
rect 10275 10452 10287 10455
rect 10318 10452 10324 10464
rect 10275 10424 10324 10452
rect 10275 10421 10287 10424
rect 10229 10415 10287 10421
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 10612 10461 10640 10560
rect 17126 10548 17132 10600
rect 17184 10588 17190 10600
rect 22388 10597 22416 10696
rect 22557 10659 22615 10665
rect 22557 10625 22569 10659
rect 22603 10656 22615 10659
rect 22646 10656 22652 10668
rect 22603 10628 22652 10656
rect 22603 10625 22615 10628
rect 22557 10619 22615 10625
rect 22646 10616 22652 10628
rect 22704 10616 22710 10668
rect 22922 10656 22928 10668
rect 22883 10628 22928 10656
rect 22922 10616 22928 10628
rect 22980 10616 22986 10668
rect 23106 10656 23112 10668
rect 23067 10628 23112 10656
rect 23106 10616 23112 10628
rect 23164 10616 23170 10668
rect 23385 10659 23443 10665
rect 23385 10625 23397 10659
rect 23431 10625 23443 10659
rect 23385 10619 23443 10625
rect 23569 10659 23627 10665
rect 23569 10625 23581 10659
rect 23615 10625 23627 10659
rect 23569 10619 23627 10625
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 17184 10560 17417 10588
rect 17184 10548 17190 10560
rect 17405 10557 17417 10560
rect 17451 10557 17463 10591
rect 17405 10551 17463 10557
rect 22373 10591 22431 10597
rect 22373 10557 22385 10591
rect 22419 10557 22431 10591
rect 22373 10551 22431 10557
rect 22462 10548 22468 10600
rect 22520 10588 22526 10600
rect 23198 10588 23204 10600
rect 22520 10560 22565 10588
rect 23159 10560 23204 10588
rect 22520 10548 22526 10560
rect 23198 10548 23204 10560
rect 23256 10548 23262 10600
rect 23400 10588 23428 10619
rect 23474 10588 23480 10600
rect 23400 10560 23480 10588
rect 23474 10548 23480 10560
rect 23532 10548 23538 10600
rect 21545 10523 21603 10529
rect 21545 10489 21557 10523
rect 21591 10520 21603 10523
rect 22480 10520 22508 10548
rect 21591 10492 22508 10520
rect 21591 10489 21603 10492
rect 21545 10483 21603 10489
rect 23014 10480 23020 10532
rect 23072 10520 23078 10532
rect 23584 10520 23612 10619
rect 23934 10616 23940 10668
rect 23992 10656 23998 10668
rect 24946 10656 24952 10668
rect 23992 10628 24037 10656
rect 24907 10628 24952 10656
rect 23992 10616 23998 10628
rect 24946 10616 24952 10628
rect 25004 10616 25010 10668
rect 25041 10659 25099 10665
rect 25041 10625 25053 10659
rect 25087 10656 25099 10659
rect 25498 10656 25504 10668
rect 25087 10628 25504 10656
rect 25087 10625 25099 10628
rect 25041 10619 25099 10625
rect 25498 10616 25504 10628
rect 25556 10616 25562 10668
rect 24486 10548 24492 10600
rect 24544 10588 24550 10600
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 24544 10560 24685 10588
rect 24544 10548 24550 10560
rect 24673 10557 24685 10560
rect 24719 10557 24731 10591
rect 24673 10551 24731 10557
rect 23845 10523 23903 10529
rect 23845 10520 23857 10523
rect 23072 10492 23857 10520
rect 23072 10480 23078 10492
rect 23845 10489 23857 10492
rect 23891 10489 23903 10523
rect 23845 10483 23903 10489
rect 10597 10455 10655 10461
rect 10597 10421 10609 10455
rect 10643 10452 10655 10455
rect 12158 10452 12164 10464
rect 10643 10424 12164 10452
rect 10643 10421 10655 10424
rect 10597 10415 10655 10421
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12710 10452 12716 10464
rect 12492 10424 12537 10452
rect 12671 10424 12716 10452
rect 12492 10412 12498 10424
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 13449 10455 13507 10461
rect 13449 10421 13461 10455
rect 13495 10452 13507 10455
rect 13630 10452 13636 10464
rect 13495 10424 13636 10452
rect 13495 10421 13507 10424
rect 13449 10415 13507 10421
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 17129 10455 17187 10461
rect 17129 10452 17141 10455
rect 16632 10424 17141 10452
rect 16632 10412 16638 10424
rect 17129 10421 17141 10424
rect 17175 10452 17187 10455
rect 17402 10452 17408 10464
rect 17175 10424 17408 10452
rect 17175 10421 17187 10424
rect 17129 10415 17187 10421
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 22186 10412 22192 10464
rect 22244 10452 22250 10464
rect 23290 10452 23296 10464
rect 22244 10424 23296 10452
rect 22244 10412 22250 10424
rect 23290 10412 23296 10424
rect 23348 10412 23354 10464
rect 23750 10412 23756 10464
rect 23808 10452 23814 10464
rect 24765 10455 24823 10461
rect 24765 10452 24777 10455
rect 23808 10424 24777 10452
rect 23808 10412 23814 10424
rect 24765 10421 24777 10424
rect 24811 10421 24823 10455
rect 24765 10415 24823 10421
rect 25038 10412 25044 10464
rect 25096 10452 25102 10464
rect 25225 10455 25283 10461
rect 25225 10452 25237 10455
rect 25096 10424 25237 10452
rect 25096 10412 25102 10424
rect 25225 10421 25237 10424
rect 25271 10421 25283 10455
rect 25225 10415 25283 10421
rect 1104 10362 29440 10384
rect 1104 10310 5672 10362
rect 5724 10310 5736 10362
rect 5788 10310 5800 10362
rect 5852 10310 5864 10362
rect 5916 10310 5928 10362
rect 5980 10310 15118 10362
rect 15170 10310 15182 10362
rect 15234 10310 15246 10362
rect 15298 10310 15310 10362
rect 15362 10310 15374 10362
rect 15426 10310 24563 10362
rect 24615 10310 24627 10362
rect 24679 10310 24691 10362
rect 24743 10310 24755 10362
rect 24807 10310 24819 10362
rect 24871 10310 29440 10362
rect 1104 10288 29440 10310
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 3789 10251 3847 10257
rect 3789 10217 3801 10251
rect 3835 10248 3847 10251
rect 3970 10248 3976 10260
rect 3835 10220 3976 10248
rect 3835 10217 3847 10220
rect 3789 10211 3847 10217
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 13814 10248 13820 10260
rect 4120 10220 13820 10248
rect 4120 10208 4126 10220
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 14185 10251 14243 10257
rect 14185 10248 14197 10251
rect 14148 10220 14197 10248
rect 14148 10208 14154 10220
rect 14185 10217 14197 10220
rect 14231 10217 14243 10251
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 14185 10211 14243 10217
rect 14752 10220 14933 10248
rect 4522 10180 4528 10192
rect 2424 10152 4528 10180
rect 2424 10053 2452 10152
rect 4522 10140 4528 10152
rect 4580 10140 4586 10192
rect 2590 10072 2596 10124
rect 2648 10112 2654 10124
rect 2866 10112 2872 10124
rect 2648 10084 2872 10112
rect 2648 10072 2654 10084
rect 2866 10072 2872 10084
rect 2924 10112 2930 10124
rect 4246 10112 4252 10124
rect 2924 10084 3188 10112
rect 4207 10084 4252 10112
rect 2924 10072 2930 10084
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10013 2467 10047
rect 2409 10007 2467 10013
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 2832 10016 3065 10044
rect 2832 10004 2838 10016
rect 3053 10013 3065 10016
rect 3099 10013 3111 10047
rect 3160 10044 3188 10084
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10112 4491 10115
rect 4479 10084 4752 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 4448 10044 4476 10075
rect 3160 10016 4476 10044
rect 3053 10007 3111 10013
rect 2593 9979 2651 9985
rect 2593 9945 2605 9979
rect 2639 9976 2651 9979
rect 2958 9976 2964 9988
rect 2639 9948 2964 9976
rect 2639 9945 2651 9948
rect 2593 9939 2651 9945
rect 2958 9936 2964 9948
rect 3016 9936 3022 9988
rect 3145 9911 3203 9917
rect 3145 9877 3157 9911
rect 3191 9908 3203 9911
rect 3326 9908 3332 9920
rect 3191 9880 3332 9908
rect 3191 9877 3203 9880
rect 3145 9871 3203 9877
rect 3326 9868 3332 9880
rect 3384 9868 3390 9920
rect 4154 9908 4160 9920
rect 4115 9880 4160 9908
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 4724 9917 4752 10084
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 5813 10115 5871 10121
rect 5813 10112 5825 10115
rect 5592 10084 5825 10112
rect 5592 10072 5598 10084
rect 5813 10081 5825 10084
rect 5859 10081 5871 10115
rect 5813 10075 5871 10081
rect 12250 10072 12256 10124
rect 12308 10112 12314 10124
rect 13909 10115 13967 10121
rect 13909 10112 13921 10115
rect 12308 10084 13921 10112
rect 12308 10072 12314 10084
rect 13909 10081 13921 10084
rect 13955 10081 13967 10115
rect 14458 10112 14464 10124
rect 14419 10084 14464 10112
rect 13909 10075 13967 10081
rect 14458 10072 14464 10084
rect 14516 10072 14522 10124
rect 14642 10112 14648 10124
rect 14603 10084 14648 10112
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 14752 10121 14780 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 14921 10211 14979 10217
rect 15289 10251 15347 10257
rect 15289 10217 15301 10251
rect 15335 10248 15347 10251
rect 16298 10248 16304 10260
rect 15335 10220 16304 10248
rect 15335 10217 15347 10220
rect 15289 10211 15347 10217
rect 16298 10208 16304 10220
rect 16356 10208 16362 10260
rect 19337 10251 19395 10257
rect 19337 10217 19349 10251
rect 19383 10248 19395 10251
rect 19702 10248 19708 10260
rect 19383 10220 19708 10248
rect 19383 10217 19395 10220
rect 19337 10211 19395 10217
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 22094 10208 22100 10260
rect 22152 10248 22158 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 22152 10220 22293 10248
rect 22152 10208 22158 10220
rect 22281 10217 22293 10220
rect 22327 10248 22339 10251
rect 22370 10248 22376 10260
rect 22327 10220 22376 10248
rect 22327 10217 22339 10220
rect 22281 10211 22339 10217
rect 22370 10208 22376 10220
rect 22428 10208 22434 10260
rect 22833 10251 22891 10257
rect 22833 10217 22845 10251
rect 22879 10248 22891 10251
rect 23106 10248 23112 10260
rect 22879 10220 23112 10248
rect 22879 10217 22891 10220
rect 22833 10211 22891 10217
rect 23106 10208 23112 10220
rect 23164 10208 23170 10260
rect 24121 10251 24179 10257
rect 24121 10217 24133 10251
rect 24167 10248 24179 10251
rect 24765 10251 24823 10257
rect 24765 10248 24777 10251
rect 24167 10220 24777 10248
rect 24167 10217 24179 10220
rect 24121 10211 24179 10217
rect 24765 10217 24777 10220
rect 24811 10248 24823 10251
rect 24946 10248 24952 10260
rect 24811 10220 24952 10248
rect 24811 10217 24823 10220
rect 24765 10211 24823 10217
rect 24946 10208 24952 10220
rect 25004 10208 25010 10260
rect 22186 10180 22192 10192
rect 17236 10152 22192 10180
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10112 14795 10115
rect 15470 10112 15476 10124
rect 14783 10084 15476 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 9122 10044 9128 10056
rect 9083 10016 9128 10044
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 14366 10044 14372 10056
rect 14327 10016 14372 10044
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 14918 10044 14924 10056
rect 14879 10016 14924 10044
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 15105 10047 15163 10053
rect 15105 10013 15117 10047
rect 15151 10044 15163 10047
rect 15838 10044 15844 10056
rect 15151 10016 15844 10044
rect 15151 10013 15163 10016
rect 15105 10007 15163 10013
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 5994 9936 6000 9988
rect 6052 9985 6058 9988
rect 6052 9979 6116 9985
rect 6052 9945 6070 9979
rect 6104 9945 6116 9979
rect 6052 9939 6116 9945
rect 6052 9936 6058 9939
rect 11054 9936 11060 9988
rect 11112 9976 11118 9988
rect 11517 9979 11575 9985
rect 11517 9976 11529 9979
rect 11112 9948 11529 9976
rect 11112 9936 11118 9948
rect 11517 9945 11529 9948
rect 11563 9976 11575 9979
rect 11563 9948 12296 9976
rect 11563 9945 11575 9948
rect 11517 9939 11575 9945
rect 4709 9911 4767 9917
rect 4709 9877 4721 9911
rect 4755 9908 4767 9911
rect 4982 9908 4988 9920
rect 4755 9880 4988 9908
rect 4755 9877 4767 9880
rect 4709 9871 4767 9877
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 7190 9908 7196 9920
rect 7151 9880 7196 9908
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 8938 9908 8944 9920
rect 8899 9880 8944 9908
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 12161 9911 12219 9917
rect 12161 9908 12173 9911
rect 12032 9880 12173 9908
rect 12032 9868 12038 9880
rect 12161 9877 12173 9880
rect 12207 9877 12219 9911
rect 12268 9908 12296 9948
rect 13170 9936 13176 9988
rect 13228 9936 13234 9988
rect 13354 9936 13360 9988
rect 13412 9976 13418 9988
rect 13633 9979 13691 9985
rect 13633 9976 13645 9979
rect 13412 9948 13645 9976
rect 13412 9936 13418 9948
rect 13633 9945 13645 9948
rect 13679 9945 13691 9979
rect 13633 9939 13691 9945
rect 14829 9979 14887 9985
rect 14829 9945 14841 9979
rect 14875 9976 14887 9979
rect 15194 9976 15200 9988
rect 14875 9948 15200 9976
rect 14875 9945 14887 9948
rect 14829 9939 14887 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 17236 9908 17264 10152
rect 22186 10140 22192 10152
rect 22244 10140 22250 10192
rect 23198 10140 23204 10192
rect 23256 10180 23262 10192
rect 23256 10152 23704 10180
rect 23256 10140 23262 10152
rect 22646 10112 22652 10124
rect 22112 10084 22652 10112
rect 22112 10056 22140 10084
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10044 21971 10047
rect 22094 10044 22100 10056
rect 21959 10016 22100 10044
rect 21959 10013 21971 10016
rect 21913 10007 21971 10013
rect 22094 10004 22100 10016
rect 22152 10004 22158 10056
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10044 22247 10047
rect 22462 10044 22468 10056
rect 22235 10016 22468 10044
rect 22235 10013 22247 10016
rect 22189 10007 22247 10013
rect 22462 10004 22468 10016
rect 22520 10044 22526 10056
rect 23012 10047 23070 10053
rect 23012 10044 23024 10047
rect 22520 10016 23024 10044
rect 22520 10004 22526 10016
rect 23012 10013 23024 10016
rect 23058 10013 23070 10047
rect 23198 10044 23204 10056
rect 23159 10016 23204 10044
rect 23012 10007 23070 10013
rect 12268 9880 17264 9908
rect 22097 9911 22155 9917
rect 12161 9871 12219 9877
rect 22097 9877 22109 9911
rect 22143 9908 22155 9911
rect 22922 9908 22928 9920
rect 22143 9880 22928 9908
rect 22143 9877 22155 9880
rect 22097 9871 22155 9877
rect 22922 9868 22928 9880
rect 22980 9868 22986 9920
rect 23032 9908 23060 10007
rect 23198 10004 23204 10016
rect 23256 10004 23262 10056
rect 23382 10044 23388 10056
rect 23343 10016 23388 10044
rect 23382 10004 23388 10016
rect 23440 10004 23446 10056
rect 23676 10053 23704 10152
rect 23842 10140 23848 10192
rect 23900 10180 23906 10192
rect 24581 10183 24639 10189
rect 24581 10180 24593 10183
rect 23900 10152 24593 10180
rect 23900 10140 23906 10152
rect 24581 10149 24593 10152
rect 24627 10149 24639 10183
rect 24581 10143 24639 10149
rect 24946 10072 24952 10124
rect 25004 10112 25010 10124
rect 25041 10115 25099 10121
rect 25041 10112 25053 10115
rect 25004 10084 25053 10112
rect 25004 10072 25010 10084
rect 25041 10081 25053 10084
rect 25087 10081 25099 10115
rect 25041 10075 25099 10081
rect 23661 10047 23719 10053
rect 23661 10013 23673 10047
rect 23707 10044 23719 10047
rect 23934 10044 23940 10056
rect 23707 10016 23940 10044
rect 23707 10013 23719 10016
rect 23661 10007 23719 10013
rect 23934 10004 23940 10016
rect 23992 10004 23998 10056
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10013 24087 10047
rect 24029 10007 24087 10013
rect 23106 9936 23112 9988
rect 23164 9976 23170 9988
rect 23477 9979 23535 9985
rect 23164 9948 23209 9976
rect 23164 9936 23170 9948
rect 23477 9945 23489 9979
rect 23523 9945 23535 9979
rect 23477 9939 23535 9945
rect 23492 9908 23520 9939
rect 23750 9936 23756 9988
rect 23808 9976 23814 9988
rect 23845 9979 23903 9985
rect 23845 9976 23857 9979
rect 23808 9948 23857 9976
rect 23808 9936 23814 9948
rect 23845 9945 23857 9948
rect 23891 9976 23903 9979
rect 24044 9976 24072 10007
rect 23891 9948 24072 9976
rect 24949 9979 25007 9985
rect 23891 9945 23903 9948
rect 23845 9939 23903 9945
rect 24949 9945 24961 9979
rect 24995 9945 25007 9979
rect 24949 9939 25007 9945
rect 23032 9880 23520 9908
rect 23566 9868 23572 9920
rect 23624 9908 23630 9920
rect 24762 9908 24768 9920
rect 23624 9880 24768 9908
rect 23624 9868 23630 9880
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 24964 9908 24992 9939
rect 25130 9936 25136 9988
rect 25188 9976 25194 9988
rect 25286 9979 25344 9985
rect 25286 9976 25298 9979
rect 25188 9948 25298 9976
rect 25188 9936 25194 9948
rect 25286 9945 25298 9948
rect 25332 9945 25344 9979
rect 25286 9939 25344 9945
rect 25498 9908 25504 9920
rect 24964 9880 25504 9908
rect 25498 9868 25504 9880
rect 25556 9868 25562 9920
rect 25590 9868 25596 9920
rect 25648 9908 25654 9920
rect 26421 9911 26479 9917
rect 26421 9908 26433 9911
rect 25648 9880 26433 9908
rect 25648 9868 25654 9880
rect 26421 9877 26433 9880
rect 26467 9877 26479 9911
rect 26421 9871 26479 9877
rect 1104 9818 29440 9840
rect 1104 9766 10395 9818
rect 10447 9766 10459 9818
rect 10511 9766 10523 9818
rect 10575 9766 10587 9818
rect 10639 9766 10651 9818
rect 10703 9766 19840 9818
rect 19892 9766 19904 9818
rect 19956 9766 19968 9818
rect 20020 9766 20032 9818
rect 20084 9766 20096 9818
rect 20148 9766 29440 9818
rect 1104 9744 29440 9766
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 4157 9707 4215 9713
rect 2832 9676 2877 9704
rect 2832 9664 2838 9676
rect 4157 9673 4169 9707
rect 4203 9704 4215 9707
rect 4614 9704 4620 9716
rect 4203 9676 4620 9704
rect 4203 9673 4215 9676
rect 4157 9667 4215 9673
rect 4614 9664 4620 9676
rect 4672 9664 4678 9716
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6457 9707 6515 9713
rect 6457 9704 6469 9707
rect 6420 9676 6469 9704
rect 6420 9664 6426 9676
rect 6457 9673 6469 9676
rect 6503 9673 6515 9707
rect 6457 9667 6515 9673
rect 6641 9707 6699 9713
rect 6641 9673 6653 9707
rect 6687 9673 6699 9707
rect 6641 9667 6699 9673
rect 11701 9707 11759 9713
rect 11701 9673 11713 9707
rect 11747 9674 11759 9707
rect 12710 9704 12716 9716
rect 12406 9676 12716 9704
rect 11747 9673 11827 9674
rect 11701 9667 11827 9673
rect 1670 9645 1676 9648
rect 1664 9636 1676 9645
rect 1631 9608 1676 9636
rect 1664 9599 1676 9608
rect 1670 9596 1676 9599
rect 1728 9596 1734 9648
rect 2682 9596 2688 9648
rect 2740 9636 2746 9648
rect 2866 9636 2872 9648
rect 2740 9608 2872 9636
rect 2740 9596 2746 9608
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 3053 9639 3111 9645
rect 3053 9636 3065 9639
rect 3016 9608 3065 9636
rect 3016 9596 3022 9608
rect 3053 9605 3065 9608
rect 3099 9605 3111 9639
rect 6086 9636 6092 9648
rect 3053 9599 3111 9605
rect 3620 9608 4016 9636
rect 3234 9568 3240 9580
rect 3195 9540 3240 9568
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3620 9577 3648 9608
rect 3988 9577 4016 9608
rect 5552 9608 6092 9636
rect 3605 9571 3663 9577
rect 3384 9540 3429 9568
rect 3384 9528 3390 9540
rect 3605 9537 3617 9571
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9568 3755 9571
rect 3973 9571 4031 9577
rect 3743 9540 3924 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 3142 9500 3148 9512
rect 2832 9472 3148 9500
rect 2832 9460 2838 9472
rect 3142 9460 3148 9472
rect 3200 9500 3206 9512
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 3200 9472 3525 9500
rect 3200 9460 3206 9472
rect 3513 9469 3525 9472
rect 3559 9469 3571 9503
rect 3786 9500 3792 9512
rect 3747 9472 3792 9500
rect 3513 9463 3571 9469
rect 3528 9364 3556 9463
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 3896 9500 3924 9540
rect 3973 9537 3985 9571
rect 4019 9568 4031 9571
rect 4154 9568 4160 9580
rect 4019 9540 4160 9568
rect 4019 9537 4031 9540
rect 3973 9531 4031 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4706 9568 4712 9580
rect 4667 9540 4712 9568
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 5552 9577 5580 9608
rect 6086 9596 6092 9608
rect 6144 9596 6150 9648
rect 6656 9636 6684 9667
rect 6564 9608 6684 9636
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 4847 9540 5181 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 5169 9537 5181 9540
rect 5215 9537 5227 9571
rect 5169 9531 5227 9537
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 4614 9500 4620 9512
rect 3896 9472 4620 9500
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 4982 9500 4988 9512
rect 4895 9472 4988 9500
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5276 9500 5304 9531
rect 5132 9472 5304 9500
rect 5132 9460 5138 9472
rect 6086 9460 6092 9512
rect 6144 9500 6150 9512
rect 6564 9500 6592 9608
rect 8938 9596 8944 9648
rect 8996 9596 9002 9648
rect 9674 9596 9680 9648
rect 9732 9596 9738 9648
rect 9766 9596 9772 9648
rect 9824 9636 9830 9648
rect 11716 9646 11827 9667
rect 11900 9648 12112 9674
rect 10137 9639 10195 9645
rect 10137 9636 10149 9639
rect 9824 9608 10149 9636
rect 9824 9596 9830 9608
rect 10137 9605 10149 9608
rect 10183 9605 10195 9639
rect 10137 9599 10195 9605
rect 10704 9608 11468 9636
rect 6639 9571 6697 9577
rect 6639 9537 6651 9571
rect 6685 9568 6697 9571
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6685 9540 7113 9568
rect 6685 9537 6697 9540
rect 6639 9531 6697 9537
rect 7101 9537 7113 9540
rect 7147 9568 7159 9571
rect 7190 9568 7196 9580
rect 7147 9540 7196 9568
rect 7147 9537 7159 9540
rect 7101 9531 7159 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7340 9540 7389 9568
rect 7340 9528 7346 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 9692 9568 9720 9596
rect 9993 9571 10051 9577
rect 9993 9568 10005 9571
rect 9692 9540 10005 9568
rect 7377 9531 7435 9537
rect 9993 9537 10005 9540
rect 10039 9537 10051 9571
rect 9993 9531 10051 9537
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 9401 9503 9459 9509
rect 6144 9472 7052 9500
rect 6144 9460 6150 9472
rect 5000 9432 5028 9460
rect 7024 9441 7052 9472
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9677 9503 9735 9509
rect 9447 9472 9628 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 7009 9435 7067 9441
rect 5000 9404 5764 9432
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3528 9336 3709 9364
rect 3697 9333 3709 9336
rect 3743 9333 3755 9367
rect 4338 9364 4344 9376
rect 4299 9336 4344 9364
rect 3697 9327 3755 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 5736 9373 5764 9404
rect 7009 9401 7021 9435
rect 7055 9401 7067 9435
rect 9600 9432 9628 9472
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 9723 9472 10180 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 9861 9435 9919 9441
rect 9861 9432 9873 9435
rect 9600 9404 9873 9432
rect 7009 9395 7067 9401
rect 9861 9401 9873 9404
rect 9907 9401 9919 9435
rect 9861 9395 9919 9401
rect 5721 9367 5779 9373
rect 5721 9333 5733 9367
rect 5767 9364 5779 9367
rect 6914 9364 6920 9376
rect 5767 9336 6920 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 7156 9336 7205 9364
rect 7156 9324 7162 9336
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 7926 9364 7932 9376
rect 7887 9336 7932 9364
rect 7193 9327 7251 9333
rect 7926 9324 7932 9336
rect 7984 9364 7990 9376
rect 9766 9364 9772 9376
rect 7984 9336 9772 9364
rect 7984 9324 7990 9336
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 10152 9364 10180 9472
rect 10244 9432 10272 9531
rect 10318 9528 10324 9580
rect 10376 9568 10382 9580
rect 10704 9577 10732 9608
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 10376 9540 10425 9568
rect 10376 9528 10382 9540
rect 10413 9537 10425 9540
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9537 10747 9571
rect 10870 9568 10876 9580
rect 10831 9540 10876 9568
rect 10689 9531 10747 9537
rect 10870 9528 10876 9540
rect 10928 9528 10934 9580
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 11109 9571 11167 9577
rect 11109 9537 11121 9571
rect 11155 9537 11167 9571
rect 11109 9531 11167 9537
rect 10980 9444 11008 9531
rect 10597 9435 10655 9441
rect 10597 9432 10609 9435
rect 10244 9404 10609 9432
rect 10597 9401 10609 9404
rect 10643 9432 10655 9435
rect 10870 9432 10876 9444
rect 10643 9404 10876 9432
rect 10643 9401 10655 9404
rect 10597 9395 10655 9401
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 10962 9392 10968 9444
rect 11020 9392 11026 9444
rect 11124 9432 11152 9531
rect 11440 9500 11468 9608
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 11799 9568 11827 9646
rect 11882 9596 11888 9648
rect 11940 9646 12112 9648
rect 11940 9596 11946 9646
rect 12084 9636 12112 9646
rect 12406 9636 12434 9676
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 13170 9664 13176 9716
rect 13228 9704 13234 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 13228 9676 13461 9704
rect 13228 9664 13234 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 13449 9667 13507 9673
rect 13722 9664 13728 9716
rect 13780 9704 13786 9716
rect 14001 9707 14059 9713
rect 14001 9704 14013 9707
rect 13780 9676 14013 9704
rect 13780 9664 13786 9676
rect 14001 9673 14013 9676
rect 14047 9704 14059 9707
rect 14366 9704 14372 9716
rect 14047 9676 14372 9704
rect 14047 9673 14059 9676
rect 14001 9667 14059 9673
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 14918 9664 14924 9716
rect 14976 9704 14982 9716
rect 15013 9707 15071 9713
rect 15013 9704 15025 9707
rect 14976 9676 15025 9704
rect 14976 9664 14982 9676
rect 15013 9673 15025 9676
rect 15059 9673 15071 9707
rect 15013 9667 15071 9673
rect 16117 9707 16175 9713
rect 16117 9673 16129 9707
rect 16163 9673 16175 9707
rect 19150 9704 19156 9716
rect 19063 9676 19156 9704
rect 16117 9667 16175 9673
rect 12084 9608 12434 9636
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11572 9540 11617 9568
rect 11799 9540 11989 9568
rect 11572 9528 11578 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9537 12127 9571
rect 12069 9531 12127 9537
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 11882 9500 11888 9512
rect 11440 9472 11888 9500
rect 11882 9460 11888 9472
rect 11940 9500 11946 9512
rect 12084 9500 12112 9531
rect 11940 9472 12112 9500
rect 12268 9500 12296 9531
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 12526 9577 12532 9580
rect 12483 9571 12532 9577
rect 12400 9540 12445 9568
rect 12400 9528 12406 9540
rect 12483 9537 12495 9571
rect 12529 9537 12532 9571
rect 12483 9531 12532 9537
rect 12526 9528 12532 9531
rect 12584 9528 12590 9580
rect 13630 9568 13636 9580
rect 13591 9540 13636 9568
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9568 14887 9571
rect 14936 9568 14964 9664
rect 15194 9636 15200 9648
rect 15155 9608 15200 9636
rect 15194 9596 15200 9608
rect 15252 9636 15258 9648
rect 15749 9639 15807 9645
rect 15749 9636 15761 9639
rect 15252 9608 15761 9636
rect 15252 9596 15258 9608
rect 15749 9605 15761 9608
rect 15795 9605 15807 9639
rect 16132 9636 16160 9667
rect 19150 9664 19156 9676
rect 19208 9704 19214 9716
rect 19208 9676 19840 9704
rect 19208 9664 19214 9676
rect 18966 9636 18972 9648
rect 16132 9608 18972 9636
rect 15749 9599 15807 9605
rect 18966 9596 18972 9608
rect 19024 9636 19030 9648
rect 19429 9639 19487 9645
rect 19024 9608 19334 9636
rect 19024 9596 19030 9608
rect 15102 9568 15108 9580
rect 14875 9540 14964 9568
rect 15063 9540 15108 9568
rect 14875 9537 14887 9540
rect 14829 9531 14887 9537
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 15381 9571 15439 9577
rect 15381 9537 15393 9571
rect 15427 9537 15439 9571
rect 15838 9568 15844 9580
rect 15799 9540 15844 9568
rect 15381 9531 15439 9537
rect 12894 9500 12900 9512
rect 12268 9472 12900 9500
rect 11940 9460 11946 9472
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 15010 9500 15016 9512
rect 13964 9472 15016 9500
rect 13964 9460 13970 9472
rect 15010 9460 15016 9472
rect 15068 9500 15074 9512
rect 15396 9500 15424 9531
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 15933 9571 15991 9577
rect 15933 9537 15945 9571
rect 15979 9537 15991 9571
rect 15933 9531 15991 9537
rect 17764 9571 17822 9577
rect 17764 9537 17776 9571
rect 17810 9568 17822 9571
rect 18230 9568 18236 9580
rect 17810 9540 18236 9568
rect 17810 9537 17822 9540
rect 17764 9531 17822 9537
rect 15068 9472 15424 9500
rect 15565 9503 15623 9509
rect 15068 9460 15074 9472
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 15948 9500 15976 9531
rect 18230 9528 18236 9540
rect 18288 9528 18294 9580
rect 19306 9568 19334 9608
rect 19429 9605 19441 9639
rect 19475 9636 19487 9639
rect 19702 9636 19708 9648
rect 19475 9608 19708 9636
rect 19475 9605 19487 9608
rect 19429 9599 19487 9605
rect 19702 9596 19708 9608
rect 19760 9596 19766 9648
rect 19812 9636 19840 9676
rect 23474 9664 23480 9716
rect 23532 9704 23538 9716
rect 23569 9707 23627 9713
rect 23569 9704 23581 9707
rect 23532 9676 23581 9704
rect 23532 9664 23538 9676
rect 23569 9673 23581 9676
rect 23615 9673 23627 9707
rect 25498 9704 25504 9716
rect 25459 9676 25504 9704
rect 23569 9667 23627 9673
rect 25498 9664 25504 9676
rect 25556 9664 25562 9716
rect 20165 9639 20223 9645
rect 20165 9636 20177 9639
rect 19812 9608 20177 9636
rect 20165 9605 20177 9608
rect 20211 9636 20223 9639
rect 21174 9636 21180 9648
rect 20211 9608 21180 9636
rect 20211 9605 20223 9608
rect 20165 9599 20223 9605
rect 21174 9596 21180 9608
rect 21232 9636 21238 9648
rect 21821 9639 21879 9645
rect 21821 9636 21833 9639
rect 21232 9608 21833 9636
rect 21232 9596 21238 9608
rect 21821 9605 21833 9608
rect 21867 9605 21879 9639
rect 21821 9599 21879 9605
rect 22278 9596 22284 9648
rect 22336 9636 22342 9648
rect 23290 9636 23296 9648
rect 22336 9608 23296 9636
rect 22336 9596 22342 9608
rect 23290 9596 23296 9608
rect 23348 9636 23354 9648
rect 25516 9636 25544 9664
rect 23348 9608 23520 9636
rect 23348 9596 23354 9608
rect 20073 9571 20131 9577
rect 20073 9568 20085 9571
rect 19306 9540 20085 9568
rect 20073 9537 20085 9540
rect 20119 9568 20131 9571
rect 20622 9568 20628 9580
rect 20119 9540 20628 9568
rect 20119 9537 20131 9540
rect 20073 9531 20131 9537
rect 20622 9528 20628 9540
rect 20680 9568 20686 9580
rect 20901 9571 20959 9577
rect 20901 9568 20913 9571
rect 20680 9540 20913 9568
rect 20680 9528 20686 9540
rect 20901 9537 20913 9540
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 20993 9571 21051 9577
rect 20993 9537 21005 9571
rect 21039 9568 21051 9571
rect 21545 9571 21603 9577
rect 21039 9540 21312 9568
rect 21039 9537 21051 9540
rect 20993 9531 21051 9537
rect 15611 9472 15976 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 17126 9460 17132 9512
rect 17184 9500 17190 9512
rect 17497 9503 17555 9509
rect 17497 9500 17509 9503
rect 17184 9472 17509 9500
rect 17184 9460 17190 9472
rect 17497 9469 17509 9472
rect 17543 9469 17555 9503
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 17497 9463 17555 9469
rect 18524 9472 20269 9500
rect 12526 9432 12532 9444
rect 11124 9404 12532 9432
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 12621 9435 12679 9441
rect 12621 9401 12633 9435
rect 12667 9432 12679 9435
rect 13354 9432 13360 9444
rect 12667 9404 13360 9432
rect 12667 9401 12679 9404
rect 12621 9395 12679 9401
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 11054 9364 11060 9376
rect 10152 9336 11060 9364
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 11238 9364 11244 9376
rect 11199 9336 11244 9364
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 11790 9364 11796 9376
rect 11751 9336 11796 9364
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 14642 9364 14648 9376
rect 14603 9336 14648 9364
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 18524 9364 18552 9472
rect 20257 9469 20269 9472
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 21085 9503 21143 9509
rect 21085 9469 21097 9503
rect 21131 9469 21143 9503
rect 21085 9463 21143 9469
rect 19058 9392 19064 9444
rect 19116 9432 19122 9444
rect 19245 9435 19303 9441
rect 19245 9432 19257 9435
rect 19116 9404 19257 9432
rect 19116 9392 19122 9404
rect 19245 9401 19257 9404
rect 19291 9401 19303 9435
rect 20272 9432 20300 9463
rect 20990 9432 20996 9444
rect 20272 9404 20996 9432
rect 19245 9395 19303 9401
rect 20990 9392 20996 9404
rect 21048 9432 21054 9444
rect 21100 9432 21128 9463
rect 21048 9404 21128 9432
rect 21284 9432 21312 9540
rect 21545 9537 21557 9571
rect 21591 9568 21603 9571
rect 23109 9571 23167 9577
rect 21591 9540 22094 9568
rect 21591 9537 21603 9540
rect 21545 9531 21603 9537
rect 21361 9435 21419 9441
rect 21361 9432 21373 9435
rect 21284 9404 21373 9432
rect 21048 9392 21054 9404
rect 21361 9401 21373 9404
rect 21407 9401 21419 9435
rect 22066 9432 22094 9540
rect 23109 9537 23121 9571
rect 23155 9568 23167 9571
rect 23198 9568 23204 9580
rect 23155 9540 23204 9568
rect 23155 9537 23167 9540
rect 23109 9531 23167 9537
rect 23198 9528 23204 9540
rect 23256 9528 23262 9580
rect 23492 9577 23520 9608
rect 24596 9608 25544 9636
rect 24596 9577 24624 9608
rect 23385 9571 23443 9577
rect 23385 9537 23397 9571
rect 23431 9537 23443 9571
rect 23385 9531 23443 9537
rect 23477 9571 23535 9577
rect 23477 9537 23489 9571
rect 23523 9537 23535 9571
rect 23477 9531 23535 9537
rect 24581 9571 24639 9577
rect 24581 9537 24593 9571
rect 24627 9537 24639 9571
rect 24762 9568 24768 9580
rect 24723 9540 24768 9568
rect 24581 9531 24639 9537
rect 22738 9460 22744 9512
rect 22796 9500 22802 9512
rect 23293 9503 23351 9509
rect 23293 9500 23305 9503
rect 22796 9472 23305 9500
rect 22796 9460 22802 9472
rect 23293 9469 23305 9472
rect 23339 9469 23351 9503
rect 23293 9463 23351 9469
rect 22925 9435 22983 9441
rect 22925 9432 22937 9435
rect 22066 9404 22937 9432
rect 21361 9395 21419 9401
rect 22925 9401 22937 9404
rect 22971 9401 22983 9435
rect 22925 9395 22983 9401
rect 23014 9392 23020 9444
rect 23072 9432 23078 9444
rect 23400 9432 23428 9531
rect 24762 9528 24768 9540
rect 24820 9528 24826 9580
rect 25038 9568 25044 9580
rect 24999 9540 25044 9568
rect 25038 9528 25044 9540
rect 25096 9528 25102 9580
rect 25317 9571 25375 9577
rect 25317 9537 25329 9571
rect 25363 9537 25375 9571
rect 25590 9568 25596 9580
rect 25503 9540 25596 9568
rect 25317 9531 25375 9537
rect 24949 9503 25007 9509
rect 24949 9469 24961 9503
rect 24995 9500 25007 9503
rect 25130 9500 25136 9512
rect 24995 9472 25136 9500
rect 24995 9469 25007 9472
rect 24949 9463 25007 9469
rect 25130 9460 25136 9472
rect 25188 9460 25194 9512
rect 25332 9500 25360 9531
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 25498 9500 25504 9512
rect 25332 9472 25504 9500
rect 25498 9460 25504 9472
rect 25556 9460 25562 9512
rect 24486 9432 24492 9444
rect 23072 9404 24492 9432
rect 23072 9392 23078 9404
rect 24486 9392 24492 9404
rect 24544 9432 24550 9444
rect 25608 9432 25636 9528
rect 24544 9404 25636 9432
rect 24544 9392 24550 9404
rect 17368 9336 18552 9364
rect 17368 9324 17374 9336
rect 18874 9324 18880 9376
rect 18932 9364 18938 9376
rect 19702 9364 19708 9376
rect 18932 9336 18977 9364
rect 19663 9336 19708 9364
rect 18932 9324 18938 9336
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 20346 9324 20352 9376
rect 20404 9364 20410 9376
rect 20533 9367 20591 9373
rect 20533 9364 20545 9367
rect 20404 9336 20545 9364
rect 20404 9324 20410 9336
rect 20533 9333 20545 9336
rect 20579 9333 20591 9367
rect 20533 9327 20591 9333
rect 22370 9324 22376 9376
rect 22428 9364 22434 9376
rect 23109 9367 23167 9373
rect 23109 9364 23121 9367
rect 22428 9336 23121 9364
rect 22428 9324 22434 9336
rect 23109 9333 23121 9336
rect 23155 9364 23167 9367
rect 23382 9364 23388 9376
rect 23155 9336 23388 9364
rect 23155 9333 23167 9336
rect 23109 9327 23167 9333
rect 23382 9324 23388 9336
rect 23440 9324 23446 9376
rect 1104 9274 29440 9296
rect 1104 9222 5672 9274
rect 5724 9222 5736 9274
rect 5788 9222 5800 9274
rect 5852 9222 5864 9274
rect 5916 9222 5928 9274
rect 5980 9222 15118 9274
rect 15170 9222 15182 9274
rect 15234 9222 15246 9274
rect 15298 9222 15310 9274
rect 15362 9222 15374 9274
rect 15426 9222 24563 9274
rect 24615 9222 24627 9274
rect 24679 9222 24691 9274
rect 24743 9222 24755 9274
rect 24807 9222 24819 9274
rect 24871 9222 29440 9274
rect 1104 9200 29440 9222
rect 3881 9163 3939 9169
rect 3881 9129 3893 9163
rect 3927 9160 3939 9163
rect 4154 9160 4160 9172
rect 3927 9132 4160 9160
rect 3927 9129 3939 9132
rect 3881 9123 3939 9129
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 4985 9163 5043 9169
rect 4985 9160 4997 9163
rect 4764 9132 4997 9160
rect 4764 9120 4770 9132
rect 4985 9129 4997 9132
rect 5031 9129 5043 9163
rect 4985 9123 5043 9129
rect 6273 9163 6331 9169
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 7282 9160 7288 9172
rect 6319 9132 7288 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 9122 9160 9128 9172
rect 9083 9132 9128 9160
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 11514 9120 11520 9172
rect 11572 9160 11578 9172
rect 12986 9160 12992 9172
rect 11572 9132 12992 9160
rect 11572 9120 11578 9132
rect 12986 9120 12992 9132
rect 13044 9120 13050 9172
rect 13081 9163 13139 9169
rect 13081 9129 13093 9163
rect 13127 9160 13139 9163
rect 13998 9160 14004 9172
rect 13127 9132 14004 9160
rect 13127 9129 13139 9132
rect 13081 9123 13139 9129
rect 12158 9052 12164 9104
rect 12216 9092 12222 9104
rect 13096 9092 13124 9123
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 15010 9160 15016 9172
rect 14971 9132 15016 9160
rect 15010 9120 15016 9132
rect 15068 9160 15074 9172
rect 15197 9163 15255 9169
rect 15197 9160 15209 9163
rect 15068 9132 15209 9160
rect 15068 9120 15074 9132
rect 15197 9129 15209 9132
rect 15243 9129 15255 9163
rect 18230 9160 18236 9172
rect 18191 9132 18236 9160
rect 15197 9123 15255 9129
rect 12216 9064 13124 9092
rect 15212 9092 15240 9123
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 22278 9160 22284 9172
rect 22239 9132 22284 9160
rect 22278 9120 22284 9132
rect 22336 9120 22342 9172
rect 22922 9120 22928 9172
rect 22980 9160 22986 9172
rect 25498 9160 25504 9172
rect 22980 9132 25504 9160
rect 22980 9120 22986 9132
rect 25498 9120 25504 9132
rect 25556 9120 25562 9172
rect 15378 9092 15384 9104
rect 15212 9064 15384 9092
rect 12216 9052 12222 9064
rect 15378 9052 15384 9064
rect 15436 9052 15442 9104
rect 20441 9095 20499 9101
rect 20441 9092 20453 9095
rect 19904 9064 20453 9092
rect 6638 9024 6644 9036
rect 6599 8996 6644 9024
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 10686 9024 10692 9036
rect 8956 8996 10692 9024
rect 3142 8956 3148 8968
rect 3103 8928 3148 8956
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3329 8959 3387 8965
rect 3329 8956 3341 8959
rect 3292 8928 3341 8956
rect 3292 8916 3298 8928
rect 3329 8925 3341 8928
rect 3375 8956 3387 8959
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3375 8928 3985 8956
rect 3375 8925 3387 8928
rect 3329 8919 3387 8925
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 5074 8956 5080 8968
rect 5035 8928 5080 8956
rect 3973 8919 4031 8925
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 6454 8956 6460 8968
rect 6415 8928 6460 8956
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8294 8956 8300 8968
rect 8251 8928 8300 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 8956 8965 8984 8996
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 11296 8996 11713 9024
rect 11296 8984 11302 8996
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 17770 8984 17776 9036
rect 17828 9024 17834 9036
rect 19904 9033 19932 9064
rect 20441 9061 20453 9064
rect 20487 9061 20499 9095
rect 21542 9092 21548 9104
rect 20441 9055 20499 9061
rect 20916 9064 21548 9092
rect 18049 9027 18107 9033
rect 18049 9024 18061 9027
rect 17828 8996 18061 9024
rect 17828 8984 17834 8996
rect 18049 8993 18061 8996
rect 18095 9024 18107 9027
rect 18785 9027 18843 9033
rect 18785 9024 18797 9027
rect 18095 8996 18797 9024
rect 18095 8993 18107 8996
rect 18049 8987 18107 8993
rect 18785 8993 18797 8996
rect 18831 8993 18843 9027
rect 18785 8987 18843 8993
rect 19889 9027 19947 9033
rect 19889 8993 19901 9027
rect 19935 8993 19947 9027
rect 20916 9024 20944 9064
rect 21542 9052 21548 9064
rect 21600 9052 21606 9104
rect 22738 9092 22744 9104
rect 22651 9064 22744 9092
rect 22738 9052 22744 9064
rect 22796 9092 22802 9104
rect 24213 9095 24271 9101
rect 24213 9092 24225 9095
rect 22796 9064 24225 9092
rect 22796 9052 22802 9064
rect 24213 9061 24225 9064
rect 24259 9061 24271 9095
rect 24213 9055 24271 9061
rect 19889 8987 19947 8993
rect 20088 8996 20944 9024
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8812 8928 8953 8956
rect 8812 8916 8818 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12250 8956 12256 8968
rect 12023 8928 12256 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 13722 8956 13728 8968
rect 13683 8928 13728 8956
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 17126 8916 17132 8968
rect 17184 8956 17190 8968
rect 17221 8959 17279 8965
rect 17221 8956 17233 8959
rect 17184 8928 17233 8956
rect 17184 8916 17190 8928
rect 17221 8925 17233 8928
rect 17267 8925 17279 8959
rect 19334 8956 19340 8968
rect 19295 8928 19340 8956
rect 17221 8919 17279 8925
rect 19334 8916 19340 8928
rect 19392 8916 19398 8968
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8956 19855 8959
rect 20088 8956 20116 8996
rect 20990 8984 20996 9036
rect 21048 9024 21054 9036
rect 21048 8996 21496 9024
rect 21048 8984 21054 8996
rect 19843 8928 20116 8956
rect 20165 8959 20223 8965
rect 19843 8925 19855 8928
rect 19797 8919 19855 8925
rect 20165 8925 20177 8959
rect 20211 8925 20223 8959
rect 20346 8956 20352 8968
rect 20307 8928 20352 8956
rect 20165 8919 20223 8925
rect 3513 8891 3571 8897
rect 3513 8857 3525 8891
rect 3559 8888 3571 8891
rect 3602 8888 3608 8900
rect 3559 8860 3608 8888
rect 3559 8857 3571 8860
rect 3513 8851 3571 8857
rect 3602 8848 3608 8860
rect 3660 8848 3666 8900
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 4120 8860 7512 8888
rect 4120 8848 4126 8860
rect 6822 8820 6828 8832
rect 6783 8792 6828 8820
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 7484 8820 7512 8860
rect 7558 8848 7564 8900
rect 7616 8888 7622 8900
rect 7938 8891 7996 8897
rect 7938 8888 7950 8891
rect 7616 8860 7950 8888
rect 7616 8848 7622 8860
rect 7938 8857 7950 8860
rect 7984 8857 7996 8891
rect 11790 8888 11796 8900
rect 11270 8860 11796 8888
rect 7938 8851 7996 8857
rect 11790 8848 11796 8860
rect 11848 8848 11854 8900
rect 12342 8848 12348 8900
rect 12400 8888 12406 8900
rect 12897 8891 12955 8897
rect 12897 8888 12909 8891
rect 12400 8860 12909 8888
rect 12400 8848 12406 8860
rect 12897 8857 12909 8860
rect 12943 8888 12955 8891
rect 13998 8888 14004 8900
rect 12943 8860 14004 8888
rect 12943 8857 12955 8860
rect 12897 8851 12955 8857
rect 13998 8848 14004 8860
rect 14056 8848 14062 8900
rect 16976 8891 17034 8897
rect 16976 8857 16988 8891
rect 17022 8888 17034 8891
rect 17773 8891 17831 8897
rect 17022 8860 17448 8888
rect 17022 8857 17034 8860
rect 16976 8851 17034 8857
rect 10229 8823 10287 8829
rect 10229 8820 10241 8823
rect 7484 8792 10241 8820
rect 10229 8789 10241 8792
rect 10275 8820 10287 8823
rect 10962 8820 10968 8832
rect 10275 8792 10968 8820
rect 10275 8789 10287 8792
rect 10229 8783 10287 8789
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 13909 8823 13967 8829
rect 13909 8820 13921 8823
rect 13872 8792 13921 8820
rect 13872 8780 13878 8792
rect 13909 8789 13921 8792
rect 13955 8789 13967 8823
rect 13909 8783 13967 8789
rect 15194 8780 15200 8832
rect 15252 8820 15258 8832
rect 15838 8820 15844 8832
rect 15252 8792 15844 8820
rect 15252 8780 15258 8792
rect 15838 8780 15844 8792
rect 15896 8820 15902 8832
rect 16850 8820 16856 8832
rect 15896 8792 16856 8820
rect 15896 8780 15902 8792
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 17420 8829 17448 8860
rect 17773 8857 17785 8891
rect 17819 8888 17831 8891
rect 19429 8891 19487 8897
rect 19429 8888 19441 8891
rect 17819 8860 19441 8888
rect 17819 8857 17831 8860
rect 17773 8851 17831 8857
rect 19429 8857 19441 8860
rect 19475 8857 19487 8891
rect 20180 8888 20208 8919
rect 20346 8916 20352 8928
rect 20404 8916 20410 8968
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 20809 8959 20867 8965
rect 20809 8956 20821 8959
rect 20680 8928 20821 8956
rect 20680 8916 20686 8928
rect 20809 8925 20821 8928
rect 20855 8925 20867 8959
rect 20809 8919 20867 8925
rect 21174 8916 21180 8968
rect 21232 8956 21238 8968
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 21232 8928 21373 8956
rect 21232 8916 21238 8928
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 21266 8888 21272 8900
rect 20180 8860 21272 8888
rect 19429 8851 19487 8857
rect 21266 8848 21272 8860
rect 21324 8848 21330 8900
rect 17405 8823 17463 8829
rect 17405 8789 17417 8823
rect 17451 8789 17463 8823
rect 17405 8783 17463 8789
rect 17865 8823 17923 8829
rect 17865 8789 17877 8823
rect 17911 8820 17923 8823
rect 18046 8820 18052 8832
rect 17911 8792 18052 8820
rect 17911 8789 17923 8792
rect 17865 8783 17923 8789
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 18598 8820 18604 8832
rect 18559 8792 18604 8820
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 18690 8780 18696 8832
rect 18748 8820 18754 8832
rect 18748 8792 18793 8820
rect 18748 8780 18754 8792
rect 18874 8780 18880 8832
rect 18932 8820 18938 8832
rect 20346 8820 20352 8832
rect 18932 8792 20352 8820
rect 18932 8780 18938 8792
rect 20346 8780 20352 8792
rect 20404 8780 20410 8832
rect 20901 8823 20959 8829
rect 20901 8789 20913 8823
rect 20947 8820 20959 8823
rect 21082 8820 21088 8832
rect 20947 8792 21088 8820
rect 20947 8789 20959 8792
rect 20901 8783 20959 8789
rect 21082 8780 21088 8792
rect 21140 8780 21146 8832
rect 21468 8820 21496 8996
rect 21818 8984 21824 9036
rect 21876 9024 21882 9036
rect 23109 9027 23167 9033
rect 21876 8996 22232 9024
rect 21876 8984 21882 8996
rect 21634 8956 21640 8968
rect 21595 8928 21640 8956
rect 21634 8916 21640 8928
rect 21692 8916 21698 8968
rect 22204 8965 22232 8996
rect 23109 8993 23121 9027
rect 23155 9024 23167 9027
rect 23753 9027 23811 9033
rect 23155 8996 23612 9024
rect 23155 8993 23167 8996
rect 23109 8987 23167 8993
rect 21729 8959 21787 8965
rect 21729 8925 21741 8959
rect 21775 8956 21787 8959
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 21775 8928 22017 8956
rect 21775 8925 21787 8928
rect 21729 8919 21787 8925
rect 22005 8925 22017 8928
rect 22051 8925 22063 8959
rect 22005 8919 22063 8925
rect 22189 8959 22247 8965
rect 22189 8925 22201 8959
rect 22235 8956 22247 8959
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 22235 8928 22661 8956
rect 22235 8925 22247 8928
rect 22189 8919 22247 8925
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 22833 8959 22891 8965
rect 22833 8925 22845 8959
rect 22879 8925 22891 8959
rect 22833 8919 22891 8925
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8956 22983 8959
rect 23014 8956 23020 8968
rect 22971 8928 23020 8956
rect 22971 8925 22983 8928
rect 22925 8919 22983 8925
rect 21652 8888 21680 8916
rect 22278 8888 22284 8900
rect 21652 8860 22284 8888
rect 22278 8848 22284 8860
rect 22336 8848 22342 8900
rect 22373 8891 22431 8897
rect 22373 8857 22385 8891
rect 22419 8888 22431 8891
rect 22848 8888 22876 8919
rect 23014 8916 23020 8928
rect 23072 8916 23078 8968
rect 23290 8956 23296 8968
rect 23251 8928 23296 8956
rect 23290 8916 23296 8928
rect 23348 8916 23354 8968
rect 23584 8965 23612 8996
rect 23753 8993 23765 9027
rect 23799 9024 23811 9027
rect 23799 8996 24624 9024
rect 23799 8993 23811 8996
rect 23753 8987 23811 8993
rect 23569 8959 23627 8965
rect 23569 8925 23581 8959
rect 23615 8925 23627 8959
rect 23842 8956 23848 8968
rect 23803 8928 23848 8956
rect 23569 8919 23627 8925
rect 23842 8916 23848 8928
rect 23900 8916 23906 8968
rect 24026 8956 24032 8968
rect 23987 8928 24032 8956
rect 24026 8916 24032 8928
rect 24084 8916 24090 8968
rect 23750 8888 23756 8900
rect 22419 8860 22453 8888
rect 22848 8860 23756 8888
rect 22419 8857 22431 8860
rect 22373 8851 22431 8857
rect 22388 8820 22416 8851
rect 23750 8848 23756 8860
rect 23808 8848 23814 8900
rect 23106 8820 23112 8832
rect 21468 8792 23112 8820
rect 23106 8780 23112 8792
rect 23164 8780 23170 8832
rect 24118 8780 24124 8832
rect 24176 8820 24182 8832
rect 24213 8823 24271 8829
rect 24213 8820 24225 8823
rect 24176 8792 24225 8820
rect 24176 8780 24182 8792
rect 24213 8789 24225 8792
rect 24259 8820 24271 8823
rect 24489 8823 24547 8829
rect 24489 8820 24501 8823
rect 24259 8792 24501 8820
rect 24259 8789 24271 8792
rect 24213 8783 24271 8789
rect 24489 8789 24501 8792
rect 24535 8789 24547 8823
rect 24596 8820 24624 8996
rect 25869 8959 25927 8965
rect 25869 8956 25881 8959
rect 24964 8928 25881 8956
rect 24964 8900 24992 8928
rect 25869 8925 25881 8928
rect 25915 8925 25927 8959
rect 25869 8919 25927 8925
rect 24946 8848 24952 8900
rect 25004 8848 25010 8900
rect 25602 8891 25660 8897
rect 25602 8888 25614 8891
rect 25056 8860 25614 8888
rect 25056 8820 25084 8860
rect 25602 8857 25614 8860
rect 25648 8857 25660 8891
rect 25602 8851 25660 8857
rect 24596 8792 25084 8820
rect 24489 8783 24547 8789
rect 1104 8730 29440 8752
rect 1104 8678 10395 8730
rect 10447 8678 10459 8730
rect 10511 8678 10523 8730
rect 10575 8678 10587 8730
rect 10639 8678 10651 8730
rect 10703 8678 19840 8730
rect 19892 8678 19904 8730
rect 19956 8678 19968 8730
rect 20020 8678 20032 8730
rect 20084 8678 20096 8730
rect 20148 8678 29440 8730
rect 1104 8656 29440 8678
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 5132 8588 5273 8616
rect 5132 8576 5138 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 6086 8616 6092 8628
rect 6047 8588 6092 8616
rect 5261 8579 5319 8585
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 7098 8616 7104 8628
rect 7059 8588 7104 8616
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7558 8616 7564 8628
rect 7519 8588 7564 8616
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 9876 8588 11529 8616
rect 5276 8520 5856 8548
rect 5276 8492 5304 8520
rect 2222 8440 2228 8492
rect 2280 8480 2286 8492
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 2280 8452 2329 8480
rect 2280 8440 2286 8452
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 5258 8480 5264 8492
rect 5219 8452 5264 8480
rect 2317 8443 2375 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5828 8489 5856 8520
rect 6454 8508 6460 8560
rect 6512 8548 6518 8560
rect 7193 8551 7251 8557
rect 7193 8548 7205 8551
rect 6512 8520 7205 8548
rect 6512 8508 6518 8520
rect 7193 8517 7205 8520
rect 7239 8517 7251 8551
rect 9214 8548 9220 8560
rect 9175 8520 9220 8548
rect 7193 8511 7251 8517
rect 9214 8508 9220 8520
rect 9272 8508 9278 8560
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5460 8452 5733 8480
rect 5460 8424 5488 8452
rect 5721 8449 5733 8452
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6822 8480 6828 8492
rect 6595 8452 6828 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 5442 8412 5448 8424
rect 5123 8384 5448 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 5534 8372 5540 8424
rect 5592 8412 5598 8424
rect 5629 8415 5687 8421
rect 5629 8412 5641 8415
rect 5592 8384 5641 8412
rect 5592 8372 5598 8384
rect 5629 8381 5641 8384
rect 5675 8381 5687 8415
rect 6564 8412 6592 8443
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 8754 8480 8760 8492
rect 8715 8452 8760 8480
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 9674 8489 9680 8492
rect 9672 8480 9680 8489
rect 9635 8452 9680 8480
rect 9672 8443 9680 8452
rect 9674 8440 9680 8443
rect 9732 8440 9738 8492
rect 9876 8489 9904 8588
rect 11517 8585 11529 8588
rect 11563 8616 11575 8619
rect 11563 8588 11831 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 9950 8508 9956 8560
rect 10008 8548 10014 8560
rect 11803 8548 11831 8588
rect 12250 8576 12256 8628
rect 12308 8616 12314 8628
rect 12308 8588 12848 8616
rect 12308 8576 12314 8588
rect 12158 8548 12164 8560
rect 10008 8520 10180 8548
rect 11803 8520 12164 8548
rect 10008 8508 10014 8520
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 10045 8483 10103 8489
rect 10045 8449 10057 8483
rect 10091 8449 10103 8483
rect 10152 8480 10180 8520
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 12342 8548 12348 8560
rect 12303 8520 12348 8548
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 10361 8483 10419 8489
rect 10361 8480 10373 8483
rect 10152 8452 10373 8480
rect 10045 8443 10103 8449
rect 10361 8449 10373 8452
rect 10407 8449 10419 8483
rect 10361 8443 10419 8449
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 5629 8375 5687 8381
rect 5736 8384 6592 8412
rect 6733 8415 6791 8421
rect 2130 8276 2136 8288
rect 2091 8248 2136 8276
rect 2130 8236 2136 8248
rect 2188 8236 2194 8288
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 5736 8285 5764 8384
rect 6733 8381 6745 8415
rect 6779 8412 6791 8415
rect 6914 8412 6920 8424
rect 6779 8384 6920 8412
rect 6779 8381 6791 8384
rect 6733 8375 6791 8381
rect 6914 8372 6920 8384
rect 6972 8412 6978 8424
rect 7009 8415 7067 8421
rect 7009 8412 7021 8415
rect 6972 8384 7021 8412
rect 6972 8372 6978 8384
rect 7009 8381 7021 8384
rect 7055 8412 7067 8415
rect 7098 8412 7104 8424
rect 7055 8384 7104 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 8110 8372 8116 8424
rect 8168 8412 8174 8424
rect 9784 8412 9812 8443
rect 8168 8384 9812 8412
rect 8168 8372 8174 8384
rect 9033 8347 9091 8353
rect 9033 8313 9045 8347
rect 9079 8344 9091 8347
rect 9306 8344 9312 8356
rect 9079 8316 9312 8344
rect 9079 8313 9091 8316
rect 9033 8307 9091 8313
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 10060 8344 10088 8443
rect 10226 8372 10232 8424
rect 10284 8412 10290 8424
rect 10520 8412 10548 8443
rect 10284 8384 10548 8412
rect 10284 8372 10290 8384
rect 10502 8344 10508 8356
rect 10060 8316 10508 8344
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 5721 8279 5779 8285
rect 5721 8276 5733 8279
rect 4212 8248 5733 8276
rect 4212 8236 4218 8248
rect 5721 8245 5733 8248
rect 5767 8245 5779 8279
rect 5721 8239 5779 8245
rect 6270 8236 6276 8288
rect 6328 8276 6334 8288
rect 6457 8279 6515 8285
rect 6457 8276 6469 8279
rect 6328 8248 6469 8276
rect 6328 8236 6334 8248
rect 6457 8245 6469 8248
rect 6503 8245 6515 8279
rect 6457 8239 6515 8245
rect 8941 8279 8999 8285
rect 8941 8245 8953 8279
rect 8987 8276 8999 8279
rect 9122 8276 9128 8288
rect 8987 8248 9128 8276
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 9493 8279 9551 8285
rect 9493 8245 9505 8279
rect 9539 8276 9551 8279
rect 9582 8276 9588 8288
rect 9539 8248 9588 8276
rect 9539 8245 9551 8248
rect 9493 8239 9551 8245
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 10229 8279 10287 8285
rect 10229 8245 10241 8279
rect 10275 8276 10287 8279
rect 10318 8276 10324 8288
rect 10275 8248 10324 8276
rect 10275 8245 10287 8248
rect 10229 8239 10287 8245
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 10612 8276 10640 8443
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 10744 8452 10793 8480
rect 10744 8440 10750 8452
rect 10781 8449 10793 8452
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 10928 8452 10973 8480
rect 11072 8452 11161 8480
rect 10928 8440 10934 8452
rect 11072 8353 11100 8452
rect 11149 8449 11161 8452
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12176 8480 12204 8508
rect 12526 8489 12532 8492
rect 12253 8483 12311 8489
rect 12253 8480 12265 8483
rect 12176 8452 12265 8480
rect 12069 8443 12127 8449
rect 12253 8449 12265 8452
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12489 8483 12532 8489
rect 12489 8449 12501 8483
rect 12489 8443 12532 8449
rect 12084 8412 12112 8443
rect 12526 8440 12532 8443
rect 12584 8440 12590 8492
rect 12820 8489 12848 8588
rect 14918 8576 14924 8628
rect 14976 8616 14982 8628
rect 15013 8619 15071 8625
rect 15013 8616 15025 8619
rect 14976 8588 15025 8616
rect 14976 8576 14982 8588
rect 15013 8585 15025 8588
rect 15059 8616 15071 8619
rect 16206 8616 16212 8628
rect 15059 8588 16212 8616
rect 15059 8585 15071 8588
rect 15013 8579 15071 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16669 8619 16727 8625
rect 16669 8585 16681 8619
rect 16715 8585 16727 8619
rect 19150 8616 19156 8628
rect 16669 8579 16727 8585
rect 16776 8588 19012 8616
rect 19111 8588 19156 8616
rect 13814 8508 13820 8560
rect 13872 8508 13878 8560
rect 15194 8548 15200 8560
rect 15155 8520 15200 8548
rect 15194 8508 15200 8520
rect 15252 8508 15258 8560
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 15289 8483 15347 8489
rect 15289 8480 15301 8483
rect 14700 8452 15301 8480
rect 14700 8440 14706 8452
rect 15289 8449 15301 8452
rect 15335 8449 15347 8483
rect 15289 8443 15347 8449
rect 12342 8412 12348 8424
rect 12084 8384 12348 8412
rect 12342 8372 12348 8384
rect 12400 8412 12406 8424
rect 12710 8412 12716 8424
rect 12400 8384 12716 8412
rect 12400 8372 12406 8384
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 13078 8412 13084 8424
rect 13039 8384 13084 8412
rect 13078 8372 13084 8384
rect 13136 8372 13142 8424
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 14826 8412 14832 8424
rect 14599 8384 14832 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 15304 8412 15332 8443
rect 15378 8440 15384 8492
rect 15436 8480 15442 8492
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 15436 8452 15485 8480
rect 15436 8440 15442 8452
rect 15473 8449 15485 8452
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 15654 8440 15660 8492
rect 15712 8480 15718 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15712 8452 15945 8480
rect 15712 8440 15718 8452
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 16209 8483 16267 8489
rect 16209 8449 16221 8483
rect 16255 8480 16267 8483
rect 16684 8480 16712 8579
rect 16255 8452 16712 8480
rect 16255 8449 16267 8452
rect 16209 8443 16267 8449
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 15304 8384 16037 8412
rect 16025 8381 16037 8384
rect 16071 8412 16083 8415
rect 16776 8412 16804 8588
rect 17126 8508 17132 8560
rect 17184 8548 17190 8560
rect 17589 8551 17647 8557
rect 17589 8548 17601 8551
rect 17184 8520 17601 8548
rect 17184 8508 17190 8520
rect 17589 8517 17601 8520
rect 17635 8517 17647 8551
rect 17589 8511 17647 8517
rect 17773 8551 17831 8557
rect 17773 8517 17785 8551
rect 17819 8548 17831 8551
rect 18230 8548 18236 8560
rect 17819 8520 18236 8548
rect 17819 8517 17831 8520
rect 17773 8511 17831 8517
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 17034 8480 17040 8492
rect 16995 8452 17040 8480
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17954 8480 17960 8492
rect 17915 8452 17960 8480
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8449 18475 8483
rect 18417 8443 18475 8449
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8449 18843 8483
rect 18984 8480 19012 8588
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 19334 8616 19340 8628
rect 19295 8588 19340 8616
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 23014 8616 23020 8628
rect 19444 8588 23020 8616
rect 19444 8548 19472 8588
rect 23014 8576 23020 8588
rect 23072 8576 23078 8628
rect 24026 8616 24032 8628
rect 23987 8588 24032 8616
rect 24026 8576 24032 8588
rect 24084 8576 24090 8628
rect 20346 8548 20352 8560
rect 19352 8520 19472 8548
rect 19628 8520 20352 8548
rect 19352 8480 19380 8520
rect 18984 8452 19380 8480
rect 18785 8443 18843 8449
rect 16071 8384 16804 8412
rect 16071 8381 16083 8384
rect 16025 8375 16083 8381
rect 16942 8372 16948 8424
rect 17000 8412 17006 8424
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 17000 8384 17141 8412
rect 17000 8372 17006 8384
rect 17129 8381 17141 8384
rect 17175 8381 17187 8415
rect 17310 8412 17316 8424
rect 17271 8384 17316 8412
rect 17129 8375 17187 8381
rect 17310 8372 17316 8384
rect 17368 8372 17374 8424
rect 11057 8347 11115 8353
rect 11057 8313 11069 8347
rect 11103 8313 11115 8347
rect 11330 8344 11336 8356
rect 11291 8316 11336 8344
rect 11057 8307 11115 8313
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 15657 8347 15715 8353
rect 15657 8313 15669 8347
rect 15703 8344 15715 8347
rect 15930 8344 15936 8356
rect 15703 8316 15936 8344
rect 15703 8313 15715 8316
rect 15657 8307 15715 8313
rect 15930 8304 15936 8316
rect 15988 8304 15994 8356
rect 16206 8304 16212 8356
rect 16264 8344 16270 8356
rect 16393 8347 16451 8353
rect 16264 8316 16344 8344
rect 16264 8304 16270 8316
rect 11793 8279 11851 8285
rect 11793 8276 11805 8279
rect 10612 8248 11805 8276
rect 11793 8245 11805 8248
rect 11839 8276 11851 8279
rect 11882 8276 11888 8288
rect 11839 8248 11888 8276
rect 11839 8245 11851 8248
rect 11793 8239 11851 8245
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 12618 8276 12624 8288
rect 12579 8248 12624 8276
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 14829 8279 14887 8285
rect 14829 8245 14841 8279
rect 14875 8276 14887 8279
rect 14918 8276 14924 8288
rect 14875 8248 14924 8276
rect 14875 8245 14887 8248
rect 14829 8239 14887 8245
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 15013 8279 15071 8285
rect 15013 8245 15025 8279
rect 15059 8276 15071 8279
rect 15470 8276 15476 8288
rect 15059 8248 15476 8276
rect 15059 8245 15071 8248
rect 15013 8239 15071 8245
rect 15470 8236 15476 8248
rect 15528 8276 15534 8288
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 15528 8248 15853 8276
rect 15528 8236 15534 8248
rect 15841 8245 15853 8248
rect 15887 8245 15899 8279
rect 16316 8276 16344 8316
rect 16393 8313 16405 8347
rect 16439 8344 16451 8347
rect 18432 8344 18460 8443
rect 18506 8372 18512 8424
rect 18564 8412 18570 8424
rect 18693 8415 18751 8421
rect 18564 8384 18609 8412
rect 18564 8372 18570 8384
rect 18693 8381 18705 8415
rect 18739 8381 18751 8415
rect 18800 8412 18828 8443
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19628 8489 19656 8520
rect 20346 8508 20352 8520
rect 20404 8508 20410 8560
rect 21358 8508 21364 8560
rect 21416 8548 21422 8560
rect 21416 8520 21864 8548
rect 21416 8508 21422 8520
rect 19521 8483 19579 8489
rect 19521 8480 19533 8483
rect 19484 8452 19533 8480
rect 19484 8440 19490 8452
rect 19521 8449 19533 8452
rect 19567 8449 19579 8483
rect 19521 8443 19579 8449
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 19702 8440 19708 8492
rect 19760 8480 19766 8492
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 19760 8452 19901 8480
rect 19760 8440 19766 8452
rect 19889 8449 19901 8452
rect 19935 8449 19947 8483
rect 19889 8443 19947 8449
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8478 21235 8483
rect 21269 8483 21327 8489
rect 21269 8478 21281 8483
rect 21223 8450 21281 8478
rect 21223 8449 21235 8450
rect 21177 8443 21235 8449
rect 21269 8449 21281 8450
rect 21315 8449 21327 8483
rect 21450 8480 21456 8492
rect 21411 8452 21456 8480
rect 21269 8443 21327 8449
rect 21450 8440 21456 8452
rect 21508 8440 21514 8492
rect 21836 8489 21864 8520
rect 21821 8483 21879 8489
rect 21821 8449 21833 8483
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 21910 8440 21916 8492
rect 21968 8480 21974 8492
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21968 8452 22017 8480
rect 21968 8440 21974 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22094 8440 22100 8492
rect 22152 8480 22158 8492
rect 22189 8483 22247 8489
rect 22189 8480 22201 8483
rect 22152 8452 22201 8480
rect 22152 8440 22158 8452
rect 22189 8449 22201 8452
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 22278 8440 22284 8492
rect 22336 8480 22342 8492
rect 24118 8480 24124 8492
rect 22336 8452 22381 8480
rect 24079 8452 24124 8480
rect 22336 8440 22342 8452
rect 24118 8440 24124 8452
rect 24176 8440 24182 8492
rect 24486 8440 24492 8492
rect 24544 8480 24550 8492
rect 25317 8483 25375 8489
rect 25317 8480 25329 8483
rect 24544 8452 25329 8480
rect 24544 8440 24550 8452
rect 25317 8449 25329 8452
rect 25363 8449 25375 8483
rect 25317 8443 25375 8449
rect 19797 8415 19855 8421
rect 19797 8412 19809 8415
rect 18800 8384 19809 8412
rect 18693 8375 18751 8381
rect 18598 8344 18604 8356
rect 16439 8316 18460 8344
rect 18559 8316 18604 8344
rect 16439 8313 16451 8316
rect 16393 8307 16451 8313
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 18708 8344 18736 8375
rect 19720 8356 19748 8384
rect 19797 8381 19809 8384
rect 19843 8381 19855 8415
rect 21634 8412 21640 8424
rect 21595 8384 21640 8412
rect 19797 8375 19855 8381
rect 21634 8372 21640 8384
rect 21692 8372 21698 8424
rect 19334 8344 19340 8356
rect 18708 8316 19340 8344
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 19702 8304 19708 8356
rect 19760 8304 19766 8356
rect 21542 8304 21548 8356
rect 21600 8344 21606 8356
rect 22002 8344 22008 8356
rect 21600 8316 22008 8344
rect 21600 8304 21606 8316
rect 22002 8304 22008 8316
rect 22060 8344 22066 8356
rect 22465 8347 22523 8353
rect 22465 8344 22477 8347
rect 22060 8316 22477 8344
rect 22060 8304 22066 8316
rect 22465 8313 22477 8316
rect 22511 8313 22523 8347
rect 22465 8307 22523 8313
rect 23106 8304 23112 8356
rect 23164 8344 23170 8356
rect 25409 8347 25467 8353
rect 25409 8344 25421 8347
rect 23164 8316 25421 8344
rect 23164 8304 23170 8316
rect 25409 8313 25421 8316
rect 25455 8313 25467 8347
rect 25409 8307 25467 8313
rect 17678 8276 17684 8288
rect 16316 8248 17684 8276
rect 15841 8239 15899 8245
rect 17678 8236 17684 8248
rect 17736 8276 17742 8288
rect 18874 8276 18880 8288
rect 17736 8248 18880 8276
rect 17736 8236 17742 8248
rect 18874 8236 18880 8248
rect 18932 8236 18938 8288
rect 20990 8236 20996 8288
rect 21048 8276 21054 8288
rect 21177 8279 21235 8285
rect 21177 8276 21189 8279
rect 21048 8248 21189 8276
rect 21048 8236 21054 8248
rect 21177 8245 21189 8248
rect 21223 8276 21235 8279
rect 23198 8276 23204 8288
rect 21223 8248 23204 8276
rect 21223 8245 21235 8248
rect 21177 8239 21235 8245
rect 23198 8236 23204 8248
rect 23256 8236 23262 8288
rect 1104 8186 29440 8208
rect 1104 8134 5672 8186
rect 5724 8134 5736 8186
rect 5788 8134 5800 8186
rect 5852 8134 5864 8186
rect 5916 8134 5928 8186
rect 5980 8134 15118 8186
rect 15170 8134 15182 8186
rect 15234 8134 15246 8186
rect 15298 8134 15310 8186
rect 15362 8134 15374 8186
rect 15426 8134 24563 8186
rect 24615 8134 24627 8186
rect 24679 8134 24691 8186
rect 24743 8134 24755 8186
rect 24807 8134 24819 8186
rect 24871 8134 29440 8186
rect 1104 8112 29440 8134
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6454 8072 6460 8084
rect 6411 8044 6460 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 9214 8032 9220 8084
rect 9272 8072 9278 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 9272 8044 9413 8072
rect 9272 8032 9278 8044
rect 9401 8041 9413 8044
rect 9447 8041 9459 8075
rect 9401 8035 9459 8041
rect 12805 8075 12863 8081
rect 12805 8041 12817 8075
rect 12851 8072 12863 8075
rect 13078 8072 13084 8084
rect 12851 8044 13084 8072
rect 12851 8041 12863 8044
rect 12805 8035 12863 8041
rect 13078 8032 13084 8044
rect 13136 8032 13142 8084
rect 13722 8072 13728 8084
rect 13683 8044 13728 8072
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 15010 8072 15016 8084
rect 14971 8044 15016 8072
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 16669 8075 16727 8081
rect 16669 8072 16681 8075
rect 15712 8044 16681 8072
rect 15712 8032 15718 8044
rect 16669 8041 16681 8044
rect 16715 8041 16727 8075
rect 16669 8035 16727 8041
rect 17129 8075 17187 8081
rect 17129 8041 17141 8075
rect 17175 8072 17187 8075
rect 17954 8072 17960 8084
rect 17175 8044 17960 8072
rect 17175 8041 17187 8044
rect 17129 8035 17187 8041
rect 17954 8032 17960 8044
rect 18012 8032 18018 8084
rect 20530 8032 20536 8084
rect 20588 8072 20594 8084
rect 21174 8072 21180 8084
rect 20588 8044 21180 8072
rect 20588 8032 20594 8044
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 21266 8032 21272 8084
rect 21324 8072 21330 8084
rect 21361 8075 21419 8081
rect 21361 8072 21373 8075
rect 21324 8044 21373 8072
rect 21324 8032 21330 8044
rect 21361 8041 21373 8044
rect 21407 8041 21419 8075
rect 21361 8035 21419 8041
rect 21729 8075 21787 8081
rect 21729 8041 21741 8075
rect 21775 8072 21787 8075
rect 21818 8072 21824 8084
rect 21775 8044 21824 8072
rect 21775 8041 21787 8044
rect 21729 8035 21787 8041
rect 5534 7964 5540 8016
rect 5592 8004 5598 8016
rect 5721 8007 5779 8013
rect 5721 8004 5733 8007
rect 5592 7976 5733 8004
rect 5592 7964 5598 7976
rect 5721 7973 5733 7976
rect 5767 8004 5779 8007
rect 6086 8004 6092 8016
rect 5767 7976 6092 8004
rect 5767 7973 5779 7976
rect 5721 7967 5779 7973
rect 6086 7964 6092 7976
rect 6144 7964 6150 8016
rect 12526 7964 12532 8016
rect 12584 7964 12590 8016
rect 13170 8004 13176 8016
rect 13131 7976 13176 8004
rect 13170 7964 13176 7976
rect 13228 7964 13234 8016
rect 13909 8007 13967 8013
rect 13909 8004 13921 8007
rect 13280 7976 13921 8004
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 5368 7908 7389 7936
rect 1394 7828 1400 7880
rect 1452 7868 1458 7880
rect 1489 7871 1547 7877
rect 1489 7868 1501 7871
rect 1452 7840 1501 7868
rect 1452 7828 1458 7840
rect 1489 7837 1501 7840
rect 1535 7868 1547 7871
rect 3881 7871 3939 7877
rect 3881 7868 3893 7871
rect 1535 7840 3893 7868
rect 1535 7837 1547 7840
rect 1489 7831 1547 7837
rect 3881 7837 3893 7840
rect 3927 7868 3939 7871
rect 5368 7868 5396 7908
rect 7377 7905 7389 7908
rect 7423 7936 7435 7939
rect 8294 7936 8300 7948
rect 7423 7908 8300 7936
rect 7423 7905 7435 7908
rect 7377 7899 7435 7905
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 10045 7939 10103 7945
rect 10045 7905 10057 7939
rect 10091 7936 10103 7939
rect 11054 7936 11060 7948
rect 10091 7908 11060 7936
rect 10091 7905 10103 7908
rect 10045 7899 10103 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 12544 7936 12572 7964
rect 13280 7936 13308 7976
rect 13909 7973 13921 7976
rect 13955 8004 13967 8007
rect 14826 8004 14832 8016
rect 13955 7976 14832 8004
rect 13955 7973 13967 7976
rect 13909 7967 13967 7973
rect 14826 7964 14832 7976
rect 14884 7964 14890 8016
rect 15028 8004 15056 8032
rect 15378 8004 15384 8016
rect 15028 7976 15384 8004
rect 15378 7964 15384 7976
rect 15436 7964 15442 8016
rect 16117 8007 16175 8013
rect 16117 7973 16129 8007
rect 16163 8004 16175 8007
rect 17034 8004 17040 8016
rect 16163 7976 17040 8004
rect 16163 7973 16175 7976
rect 16117 7967 16175 7973
rect 12544 7908 12669 7936
rect 3927 7840 5396 7868
rect 5445 7871 5503 7877
rect 3927 7837 3939 7840
rect 3881 7831 3939 7837
rect 5445 7837 5457 7871
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 1762 7809 1768 7812
rect 1756 7763 1768 7809
rect 1820 7800 1826 7812
rect 4148 7803 4206 7809
rect 1820 7772 1856 7800
rect 1762 7760 1768 7763
rect 1820 7760 1826 7772
rect 4148 7769 4160 7803
rect 4194 7800 4206 7803
rect 4338 7800 4344 7812
rect 4194 7772 4344 7800
rect 4194 7769 4206 7772
rect 4148 7763 4206 7769
rect 4338 7760 4344 7772
rect 4396 7760 4402 7812
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 3510 7732 3516 7744
rect 2915 7704 3516 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 5258 7732 5264 7744
rect 4028 7704 5264 7732
rect 4028 7692 4034 7704
rect 5258 7692 5264 7704
rect 5316 7732 5322 7744
rect 5460 7732 5488 7831
rect 5534 7828 5540 7880
rect 5592 7868 5598 7880
rect 5629 7871 5687 7877
rect 5629 7868 5641 7871
rect 5592 7840 5641 7868
rect 5592 7828 5598 7840
rect 5629 7837 5641 7840
rect 5675 7837 5687 7871
rect 6086 7868 6092 7880
rect 6047 7840 6092 7868
rect 5629 7831 5687 7837
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6270 7868 6276 7880
rect 6231 7840 6276 7868
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 6880 7840 7941 7868
rect 6880 7828 6886 7840
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 9122 7868 9128 7880
rect 9083 7840 9128 7868
rect 7929 7831 7987 7837
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7868 12311 7871
rect 12342 7868 12348 7880
rect 12299 7840 12348 7868
rect 12299 7837 12311 7840
rect 12253 7831 12311 7837
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 12641 7877 12669 7908
rect 12820 7908 13308 7936
rect 12529 7871 12587 7877
rect 12529 7837 12541 7871
rect 12575 7837 12587 7871
rect 12529 7831 12587 7837
rect 12626 7871 12684 7877
rect 12626 7837 12638 7871
rect 12672 7837 12684 7871
rect 12626 7831 12684 7837
rect 6178 7760 6184 7812
rect 6236 7800 6242 7812
rect 6457 7803 6515 7809
rect 6457 7800 6469 7803
rect 6236 7772 6469 7800
rect 6236 7760 6242 7772
rect 6457 7769 6469 7772
rect 6503 7769 6515 7803
rect 6457 7763 6515 7769
rect 7561 7803 7619 7809
rect 7561 7769 7573 7803
rect 7607 7800 7619 7803
rect 9306 7800 9312 7812
rect 7607 7772 9312 7800
rect 7607 7769 7619 7772
rect 7561 7763 7619 7769
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 10318 7800 10324 7812
rect 10279 7772 10324 7800
rect 10318 7760 10324 7772
rect 10376 7760 10382 7812
rect 11330 7760 11336 7812
rect 11388 7760 11394 7812
rect 11882 7760 11888 7812
rect 11940 7800 11946 7812
rect 12437 7803 12495 7809
rect 12437 7800 12449 7803
rect 11940 7772 12449 7800
rect 11940 7760 11946 7772
rect 12437 7769 12449 7772
rect 12483 7769 12495 7803
rect 12544 7800 12572 7831
rect 12820 7800 12848 7908
rect 13354 7896 13360 7948
rect 13412 7936 13418 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 13412 7908 14197 7936
rect 13412 7896 13418 7908
rect 14185 7905 14197 7908
rect 14231 7936 14243 7939
rect 14274 7936 14280 7948
rect 14231 7908 14280 7936
rect 14231 7905 14243 7908
rect 14185 7899 14243 7905
rect 14274 7896 14280 7908
rect 14332 7896 14338 7948
rect 16776 7945 16804 7976
rect 17034 7964 17040 7976
rect 17092 7964 17098 8016
rect 17770 8004 17776 8016
rect 17731 7976 17776 8004
rect 17770 7964 17776 7976
rect 17828 7964 17834 8016
rect 21376 8004 21404 8035
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 25866 8072 25872 8084
rect 22066 8044 25872 8072
rect 21910 8004 21916 8016
rect 21376 7976 21916 8004
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7936 15623 7939
rect 16761 7939 16819 7945
rect 15611 7908 16252 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 12986 7868 12992 7880
rect 12947 7840 12992 7868
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 13170 7828 13176 7880
rect 13228 7868 13234 7880
rect 13265 7871 13323 7877
rect 13265 7868 13277 7871
rect 13228 7840 13277 7868
rect 13228 7828 13234 7840
rect 13265 7837 13277 7840
rect 13311 7837 13323 7871
rect 13265 7831 13323 7837
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7837 13599 7871
rect 14918 7868 14924 7880
rect 14879 7840 14924 7868
rect 13541 7831 13599 7837
rect 12544 7772 12848 7800
rect 13004 7800 13032 7828
rect 13556 7800 13584 7831
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 15197 7871 15255 7877
rect 15197 7837 15209 7871
rect 15243 7868 15255 7871
rect 15470 7868 15476 7880
rect 15243 7840 15476 7868
rect 15243 7837 15255 7840
rect 15197 7831 15255 7837
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 15930 7868 15936 7880
rect 15891 7840 15936 7868
rect 15930 7828 15936 7840
rect 15988 7828 15994 7880
rect 16224 7877 16252 7908
rect 16761 7905 16773 7939
rect 16807 7905 16819 7939
rect 16761 7899 16819 7905
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7837 16267 7871
rect 16209 7831 16267 7837
rect 16850 7828 16856 7880
rect 16908 7868 16914 7880
rect 16945 7871 17003 7877
rect 16945 7868 16957 7871
rect 16908 7840 16957 7868
rect 16908 7828 16914 7840
rect 16945 7837 16957 7840
rect 16991 7837 17003 7871
rect 17052 7868 17080 7964
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 22066 7936 22094 8044
rect 25866 8032 25872 8044
rect 25924 8032 25930 8084
rect 24397 8007 24455 8013
rect 24397 7973 24409 8007
rect 24443 7973 24455 8007
rect 24397 7967 24455 7973
rect 23014 7936 23020 7948
rect 17276 7908 22094 7936
rect 22975 7908 23020 7936
rect 17276 7896 17282 7908
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 17497 7871 17555 7877
rect 17497 7868 17509 7871
rect 17052 7840 17509 7868
rect 16945 7831 17003 7837
rect 17497 7837 17509 7840
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17920 7840 17969 7868
rect 17920 7828 17926 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 18230 7828 18236 7880
rect 18288 7868 18294 7880
rect 19058 7868 19064 7880
rect 18288 7840 19064 7868
rect 18288 7828 18294 7840
rect 19058 7828 19064 7840
rect 19116 7868 19122 7880
rect 20625 7871 20683 7877
rect 20625 7868 20637 7871
rect 19116 7840 20637 7868
rect 19116 7828 19122 7840
rect 20625 7837 20637 7840
rect 20671 7837 20683 7871
rect 21174 7868 21180 7880
rect 21135 7840 21180 7868
rect 20625 7831 20683 7837
rect 21174 7828 21180 7840
rect 21232 7868 21238 7880
rect 21637 7871 21695 7877
rect 21637 7868 21649 7871
rect 21232 7840 21649 7868
rect 21232 7828 21238 7840
rect 21637 7837 21649 7840
rect 21683 7837 21695 7871
rect 21637 7831 21695 7837
rect 23201 7871 23259 7877
rect 23201 7837 23213 7871
rect 23247 7868 23259 7871
rect 24412 7868 24440 7967
rect 24486 7896 24492 7948
rect 24544 7936 24550 7948
rect 24949 7939 25007 7945
rect 24949 7936 24961 7939
rect 24544 7908 24961 7936
rect 24544 7896 24550 7908
rect 24949 7905 24961 7908
rect 24995 7905 25007 7939
rect 24949 7899 25007 7905
rect 23247 7840 24440 7868
rect 23247 7837 23259 7840
rect 23201 7831 23259 7837
rect 24670 7828 24676 7880
rect 24728 7868 24734 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 24728 7840 24869 7868
rect 24728 7828 24734 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 15378 7800 15384 7812
rect 13004 7772 13584 7800
rect 15339 7772 15384 7800
rect 12437 7763 12495 7769
rect 5316 7704 5488 7732
rect 5316 7692 5322 7704
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 7745 7735 7803 7741
rect 7745 7732 7757 7735
rect 7340 7704 7757 7732
rect 7340 7692 7346 7704
rect 7745 7701 7757 7704
rect 7791 7701 7803 7735
rect 8938 7732 8944 7744
rect 8899 7704 8944 7732
rect 7745 7695 7803 7701
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 10226 7692 10232 7744
rect 10284 7732 10290 7744
rect 11793 7735 11851 7741
rect 11793 7732 11805 7735
rect 10284 7704 11805 7732
rect 10284 7692 10290 7704
rect 11793 7701 11805 7704
rect 11839 7701 11851 7735
rect 12452 7732 12480 7763
rect 15378 7760 15384 7772
rect 15436 7760 15442 7812
rect 16669 7803 16727 7809
rect 16669 7769 16681 7803
rect 16715 7800 16727 7803
rect 16715 7772 16835 7800
rect 16715 7769 16727 7772
rect 16669 7763 16727 7769
rect 13354 7732 13360 7744
rect 12452 7704 13360 7732
rect 11793 7695 11851 7701
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 13449 7735 13507 7741
rect 13449 7701 13461 7735
rect 13495 7732 13507 7735
rect 13538 7732 13544 7744
rect 13495 7704 13544 7732
rect 13495 7701 13507 7704
rect 13449 7695 13507 7701
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 14734 7732 14740 7744
rect 14695 7704 14740 7732
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 16390 7732 16396 7744
rect 16351 7704 16396 7732
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 16807 7732 16835 7772
rect 18506 7760 18512 7812
rect 18564 7800 18570 7812
rect 20809 7803 20867 7809
rect 18564 7772 18828 7800
rect 18564 7760 18570 7772
rect 17310 7732 17316 7744
rect 16807 7704 17316 7732
rect 17310 7692 17316 7704
rect 17368 7692 17374 7744
rect 17589 7735 17647 7741
rect 17589 7701 17601 7735
rect 17635 7732 17647 7735
rect 18690 7732 18696 7744
rect 17635 7704 18696 7732
rect 17635 7701 17647 7704
rect 17589 7695 17647 7701
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 18800 7732 18828 7772
rect 20809 7769 20821 7803
rect 20855 7800 20867 7803
rect 24946 7800 24952 7812
rect 20855 7772 24952 7800
rect 20855 7769 20867 7772
rect 20809 7763 20867 7769
rect 24946 7760 24952 7772
rect 25004 7760 25010 7812
rect 20990 7732 20996 7744
rect 18800 7704 20996 7732
rect 20990 7692 20996 7704
rect 21048 7692 21054 7744
rect 23382 7732 23388 7744
rect 23343 7704 23388 7732
rect 23382 7692 23388 7704
rect 23440 7692 23446 7744
rect 24762 7732 24768 7744
rect 24723 7704 24768 7732
rect 24762 7692 24768 7704
rect 24820 7692 24826 7744
rect 1104 7642 29440 7664
rect 1104 7590 10395 7642
rect 10447 7590 10459 7642
rect 10511 7590 10523 7642
rect 10575 7590 10587 7642
rect 10639 7590 10651 7642
rect 10703 7590 19840 7642
rect 19892 7590 19904 7642
rect 19956 7590 19968 7642
rect 20020 7590 20032 7642
rect 20084 7590 20096 7642
rect 20148 7590 29440 7642
rect 1104 7568 29440 7590
rect 1762 7528 1768 7540
rect 1723 7500 1768 7528
rect 1762 7488 1768 7500
rect 1820 7488 1826 7540
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 2225 7531 2283 7537
rect 2225 7528 2237 7531
rect 2188 7500 2237 7528
rect 2188 7488 2194 7500
rect 2225 7497 2237 7500
rect 2271 7497 2283 7531
rect 3786 7528 3792 7540
rect 3747 7500 3792 7528
rect 2225 7491 2283 7497
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 4163 7500 4476 7528
rect 3602 7420 3608 7472
rect 3660 7460 3666 7472
rect 4163 7460 4191 7500
rect 3660 7432 4191 7460
rect 3660 7420 3666 7432
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 4448 7460 4476 7500
rect 6638 7488 6644 7540
rect 6696 7488 6702 7540
rect 6822 7528 6828 7540
rect 6783 7500 6828 7528
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7282 7528 7288 7540
rect 7243 7500 7288 7528
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 11146 7488 11152 7540
rect 11204 7528 11210 7540
rect 11422 7528 11428 7540
rect 11204 7500 11428 7528
rect 11204 7488 11210 7500
rect 11422 7488 11428 7500
rect 11480 7528 11486 7540
rect 14734 7528 14740 7540
rect 11480 7500 14740 7528
rect 11480 7488 11486 7500
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 17236 7500 17908 7528
rect 4893 7463 4951 7469
rect 4893 7460 4905 7463
rect 4304 7432 4349 7460
rect 4448 7432 4905 7460
rect 4304 7420 4310 7432
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2823 7364 2973 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 3203 7395 3261 7401
rect 3203 7361 3215 7395
rect 3249 7361 3261 7395
rect 3510 7392 3516 7404
rect 3471 7364 3516 7392
rect 3203 7355 3261 7361
rect 2148 7256 2176 7355
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7324 2375 7327
rect 2682 7324 2688 7336
rect 2363 7296 2688 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 2406 7256 2412 7268
rect 2148 7228 2412 7256
rect 2406 7216 2412 7228
rect 2464 7256 2470 7268
rect 2593 7259 2651 7265
rect 2593 7256 2605 7259
rect 2464 7228 2605 7256
rect 2464 7216 2470 7228
rect 2593 7225 2605 7228
rect 2639 7225 2651 7259
rect 3218 7256 3246 7355
rect 3510 7352 3516 7364
rect 3568 7392 3574 7404
rect 3568 7364 3924 7392
rect 3568 7352 3574 7364
rect 3602 7324 3608 7336
rect 3563 7296 3608 7324
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 3896 7324 3924 7364
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4341 7395 4399 7401
rect 4028 7364 4073 7392
rect 4028 7352 4034 7364
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4448 7392 4476 7432
rect 4893 7429 4905 7432
rect 4939 7429 4951 7463
rect 6656 7460 6684 7488
rect 4893 7423 4951 7429
rect 6564 7432 6684 7460
rect 4387 7364 4476 7392
rect 5077 7395 5135 7401
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5994 7392 6000 7404
rect 5955 7364 6000 7392
rect 5077 7355 5135 7361
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 3896 7296 4077 7324
rect 4065 7293 4077 7296
rect 4111 7324 4123 7327
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 4111 7296 4445 7324
rect 4111 7293 4123 7296
rect 4065 7287 4123 7293
rect 4433 7293 4445 7296
rect 4479 7324 4491 7327
rect 5092 7324 5120 7355
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 6564 7401 6592 7432
rect 8938 7420 8944 7472
rect 8996 7420 9002 7472
rect 9306 7420 9312 7472
rect 9364 7460 9370 7472
rect 10965 7463 11023 7469
rect 10965 7460 10977 7463
rect 9364 7432 10977 7460
rect 9364 7420 9370 7432
rect 10965 7429 10977 7432
rect 11011 7429 11023 7463
rect 10965 7423 11023 7429
rect 12529 7463 12587 7469
rect 12529 7429 12541 7463
rect 12575 7460 12587 7463
rect 12618 7460 12624 7472
rect 12575 7432 12624 7460
rect 12575 7429 12587 7432
rect 12529 7423 12587 7429
rect 12618 7420 12624 7432
rect 12676 7420 12682 7472
rect 13538 7420 13544 7472
rect 13596 7420 13602 7472
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 6687 7364 7389 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 4479 7296 5120 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 4522 7256 4528 7268
rect 3218 7228 4528 7256
rect 2593 7219 2651 7225
rect 4522 7216 4528 7228
rect 4580 7256 4586 7268
rect 6181 7259 6239 7265
rect 4580 7228 5212 7256
rect 4580 7216 4586 7228
rect 4062 7148 4068 7200
rect 4120 7188 4126 7200
rect 4157 7191 4215 7197
rect 4157 7188 4169 7191
rect 4120 7160 4169 7188
rect 4120 7148 4126 7160
rect 4157 7157 4169 7160
rect 4203 7157 4215 7191
rect 4338 7188 4344 7200
rect 4299 7160 4344 7188
rect 4157 7151 4215 7157
rect 4338 7148 4344 7160
rect 4396 7148 4402 7200
rect 4709 7191 4767 7197
rect 4709 7157 4721 7191
rect 4755 7188 4767 7191
rect 4890 7188 4896 7200
rect 4755 7160 4896 7188
rect 4755 7157 4767 7160
rect 4709 7151 4767 7157
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 5184 7197 5212 7228
rect 6181 7225 6193 7259
rect 6227 7256 6239 7259
rect 6656 7256 6684 7355
rect 16390 7352 16396 7404
rect 16448 7392 16454 7404
rect 17236 7401 17264 7500
rect 17497 7463 17555 7469
rect 17497 7429 17509 7463
rect 17543 7429 17555 7463
rect 17678 7460 17684 7472
rect 17639 7432 17684 7460
rect 17497 7423 17555 7429
rect 17221 7395 17279 7401
rect 17221 7392 17233 7395
rect 16448 7364 17233 7392
rect 16448 7352 16454 7364
rect 17221 7361 17233 7364
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 17313 7395 17371 7401
rect 17313 7361 17325 7395
rect 17359 7392 17371 7395
rect 17512 7392 17540 7423
rect 17678 7420 17684 7432
rect 17736 7420 17742 7472
rect 17880 7460 17908 7500
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 19061 7531 19119 7537
rect 18012 7500 19012 7528
rect 18012 7488 18018 7500
rect 18984 7472 19012 7500
rect 19061 7497 19073 7531
rect 19107 7528 19119 7531
rect 21174 7528 21180 7540
rect 19107 7500 21180 7528
rect 19107 7497 19119 7500
rect 19061 7491 19119 7497
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 24762 7528 24768 7540
rect 24723 7500 24768 7528
rect 24762 7488 24768 7500
rect 24820 7488 24826 7540
rect 17880 7432 18736 7460
rect 17359 7364 17816 7392
rect 17359 7361 17371 7364
rect 17313 7355 17371 7361
rect 7098 7324 7104 7336
rect 7059 7296 7104 7324
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 9582 7324 9588 7336
rect 9543 7296 9588 7324
rect 9582 7284 9588 7296
rect 9640 7284 9646 7336
rect 9861 7327 9919 7333
rect 9861 7293 9873 7327
rect 9907 7324 9919 7327
rect 12250 7324 12256 7336
rect 9907 7296 12256 7324
rect 9907 7293 9919 7296
rect 9861 7287 9919 7293
rect 6227 7228 6684 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 11072 7200 11100 7296
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 17788 7324 17816 7364
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18049 7395 18107 7401
rect 18049 7392 18061 7395
rect 18012 7364 18061 7392
rect 18012 7352 18018 7364
rect 18049 7361 18061 7364
rect 18095 7361 18107 7395
rect 18230 7392 18236 7404
rect 18191 7364 18236 7392
rect 18049 7355 18107 7361
rect 18230 7352 18236 7364
rect 18288 7352 18294 7404
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7392 18475 7395
rect 18506 7392 18512 7404
rect 18463 7364 18512 7392
rect 18463 7361 18475 7364
rect 18417 7355 18475 7361
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 18708 7401 18736 7432
rect 18966 7420 18972 7472
rect 19024 7460 19030 7472
rect 21358 7460 21364 7472
rect 19024 7432 19472 7460
rect 19024 7420 19030 7432
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7361 18751 7395
rect 18693 7355 18751 7361
rect 18248 7324 18276 7352
rect 17788 7296 18276 7324
rect 18708 7324 18736 7355
rect 18782 7352 18788 7404
rect 18840 7392 18846 7404
rect 19444 7401 19472 7432
rect 19536 7432 21364 7460
rect 19536 7401 19564 7432
rect 21358 7420 21364 7432
rect 21416 7420 21422 7472
rect 21818 7420 21824 7472
rect 21876 7460 21882 7472
rect 21913 7463 21971 7469
rect 21913 7460 21925 7463
rect 21876 7432 21925 7460
rect 21876 7420 21882 7432
rect 21913 7429 21925 7432
rect 21959 7429 21971 7463
rect 24670 7460 24676 7472
rect 21913 7423 21971 7429
rect 24136 7432 24676 7460
rect 18877 7395 18935 7401
rect 18877 7392 18889 7395
rect 18840 7364 18889 7392
rect 18840 7352 18846 7364
rect 18877 7361 18889 7364
rect 18923 7392 18935 7395
rect 19337 7395 19395 7401
rect 19337 7392 19349 7395
rect 18923 7364 19349 7392
rect 18923 7361 18935 7364
rect 18877 7355 18935 7361
rect 19337 7361 19349 7364
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 19521 7395 19579 7401
rect 19521 7361 19533 7395
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 19702 7352 19708 7404
rect 19760 7392 19766 7404
rect 19981 7395 20039 7401
rect 19981 7392 19993 7395
rect 19760 7364 19993 7392
rect 19760 7352 19766 7364
rect 19981 7361 19993 7364
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 19794 7324 19800 7336
rect 18708 7296 19800 7324
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 20073 7327 20131 7333
rect 20073 7293 20085 7327
rect 20119 7293 20131 7327
rect 20254 7324 20260 7336
rect 20215 7296 20260 7324
rect 20073 7287 20131 7293
rect 17862 7256 17868 7268
rect 17823 7228 17868 7256
rect 17862 7216 17868 7228
rect 17920 7216 17926 7268
rect 17954 7216 17960 7268
rect 18012 7256 18018 7268
rect 19613 7259 19671 7265
rect 19613 7256 19625 7259
rect 18012 7228 19625 7256
rect 18012 7216 18018 7228
rect 19613 7225 19625 7228
rect 19659 7225 19671 7259
rect 20088 7256 20116 7287
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 20364 7324 20392 7355
rect 20438 7352 20444 7404
rect 20496 7392 20502 7404
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20496 7364 21005 7392
rect 20496 7352 20502 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 21082 7352 21088 7404
rect 21140 7392 21146 7404
rect 22281 7395 22339 7401
rect 22281 7392 22293 7395
rect 21140 7364 21185 7392
rect 21284 7364 22293 7392
rect 21140 7352 21146 7364
rect 21284 7336 21312 7364
rect 22281 7361 22293 7364
rect 22327 7392 22339 7395
rect 23014 7392 23020 7404
rect 22327 7364 23020 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 23198 7392 23204 7404
rect 23159 7364 23204 7392
rect 23198 7352 23204 7364
rect 23256 7352 23262 7404
rect 23382 7392 23388 7404
rect 23343 7364 23388 7392
rect 23382 7352 23388 7364
rect 23440 7352 23446 7404
rect 23661 7395 23719 7401
rect 23661 7392 23673 7395
rect 23584 7364 23673 7392
rect 20364 7296 21036 7324
rect 20625 7259 20683 7265
rect 20625 7256 20637 7259
rect 20088 7228 20637 7256
rect 19613 7219 19671 7225
rect 20625 7225 20637 7228
rect 20671 7225 20683 7259
rect 21008 7256 21036 7296
rect 21266 7284 21272 7336
rect 21324 7324 21330 7336
rect 22465 7327 22523 7333
rect 21324 7296 21417 7324
rect 21324 7284 21330 7296
rect 22465 7293 22477 7327
rect 22511 7324 22523 7327
rect 22646 7324 22652 7336
rect 22511 7296 22652 7324
rect 22511 7293 22523 7296
rect 22465 7287 22523 7293
rect 22646 7284 22652 7296
rect 22704 7284 22710 7336
rect 23474 7324 23480 7336
rect 23435 7296 23480 7324
rect 23474 7284 23480 7296
rect 23532 7284 23538 7336
rect 21634 7256 21640 7268
rect 21008 7228 21640 7256
rect 20625 7219 20683 7225
rect 21634 7216 21640 7228
rect 21692 7216 21698 7268
rect 22186 7256 22192 7268
rect 22147 7228 22192 7256
rect 22186 7216 22192 7228
rect 22244 7216 22250 7268
rect 22278 7216 22284 7268
rect 22336 7256 22342 7268
rect 23382 7256 23388 7268
rect 22336 7228 23388 7256
rect 22336 7216 22342 7228
rect 23382 7216 23388 7228
rect 23440 7256 23446 7268
rect 23584 7256 23612 7364
rect 23661 7361 23673 7364
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 23845 7395 23903 7401
rect 23845 7361 23857 7395
rect 23891 7392 23903 7395
rect 23934 7392 23940 7404
rect 23891 7364 23940 7392
rect 23891 7361 23903 7364
rect 23845 7355 23903 7361
rect 23934 7352 23940 7364
rect 23992 7392 23998 7404
rect 24136 7401 24164 7432
rect 24670 7420 24676 7432
rect 24728 7420 24734 7472
rect 24121 7395 24179 7401
rect 24121 7392 24133 7395
rect 23992 7364 24133 7392
rect 23992 7352 23998 7364
rect 24121 7361 24133 7364
rect 24167 7361 24179 7395
rect 24302 7392 24308 7404
rect 24263 7364 24308 7392
rect 24121 7355 24179 7361
rect 24302 7352 24308 7364
rect 24360 7352 24366 7404
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 24581 7395 24639 7401
rect 24581 7392 24593 7395
rect 24535 7364 24593 7392
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 24581 7361 24593 7364
rect 24627 7361 24639 7395
rect 25774 7392 25780 7404
rect 25735 7364 25780 7392
rect 24581 7355 24639 7361
rect 25774 7352 25780 7364
rect 25832 7352 25838 7404
rect 23440 7228 23612 7256
rect 23440 7216 23446 7228
rect 5169 7191 5227 7197
rect 5169 7157 5181 7191
rect 5215 7157 5227 7191
rect 7742 7188 7748 7200
rect 7703 7160 7748 7188
rect 5169 7151 5227 7157
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 8110 7188 8116 7200
rect 8071 7160 8116 7188
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 11054 7188 11060 7200
rect 11015 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 13998 7188 14004 7200
rect 13911 7160 14004 7188
rect 13998 7148 14004 7160
rect 14056 7188 14062 7200
rect 14734 7188 14740 7200
rect 14056 7160 14740 7188
rect 14056 7148 14062 7160
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 17681 7191 17739 7197
rect 17681 7157 17693 7191
rect 17727 7188 17739 7191
rect 18046 7188 18052 7200
rect 17727 7160 18052 7188
rect 17727 7157 17739 7160
rect 17681 7151 17739 7157
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18690 7188 18696 7200
rect 18651 7160 18696 7188
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 25958 7188 25964 7200
rect 25919 7160 25964 7188
rect 25958 7148 25964 7160
rect 26016 7148 26022 7200
rect 1104 7098 29440 7120
rect 1104 7046 5672 7098
rect 5724 7046 5736 7098
rect 5788 7046 5800 7098
rect 5852 7046 5864 7098
rect 5916 7046 5928 7098
rect 5980 7046 15118 7098
rect 15170 7046 15182 7098
rect 15234 7046 15246 7098
rect 15298 7046 15310 7098
rect 15362 7046 15374 7098
rect 15426 7046 24563 7098
rect 24615 7046 24627 7098
rect 24679 7046 24691 7098
rect 24743 7046 24755 7098
rect 24807 7046 24819 7098
rect 24871 7046 29440 7098
rect 1104 7024 29440 7046
rect 2682 6984 2688 6996
rect 2643 6956 2688 6984
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 5629 6987 5687 6993
rect 5629 6953 5641 6987
rect 5675 6984 5687 6987
rect 5994 6984 6000 6996
rect 5675 6956 6000 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 11974 6984 11980 6996
rect 10376 6956 11980 6984
rect 10376 6944 10382 6956
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 15654 6984 15660 6996
rect 15615 6956 15660 6984
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 18046 6944 18052 6996
rect 18104 6984 18110 6996
rect 18598 6984 18604 6996
rect 18104 6956 18604 6984
rect 18104 6944 18110 6956
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 18966 6944 18972 6996
rect 19024 6984 19030 6996
rect 19521 6987 19579 6993
rect 19521 6984 19533 6987
rect 19024 6956 19533 6984
rect 19024 6944 19030 6956
rect 19521 6953 19533 6956
rect 19567 6953 19579 6987
rect 20254 6984 20260 6996
rect 20215 6956 20260 6984
rect 19521 6947 19579 6953
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 22094 6944 22100 6996
rect 22152 6984 22158 6996
rect 25774 6984 25780 6996
rect 22152 6956 22324 6984
rect 25735 6956 25780 6984
rect 22152 6944 22158 6956
rect 4522 6916 4528 6928
rect 4448 6888 4528 6916
rect 2133 6851 2191 6857
rect 2133 6817 2145 6851
rect 2179 6848 2191 6851
rect 2222 6848 2228 6860
rect 2179 6820 2228 6848
rect 2179 6817 2191 6820
rect 2133 6811 2191 6817
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 4448 6857 4476 6888
rect 4522 6876 4528 6888
rect 4580 6876 4586 6928
rect 19337 6919 19395 6925
rect 19337 6885 19349 6919
rect 19383 6916 19395 6919
rect 19702 6916 19708 6928
rect 19383 6888 19708 6916
rect 19383 6885 19395 6888
rect 19337 6879 19395 6885
rect 19702 6876 19708 6888
rect 19760 6876 19766 6928
rect 20070 6876 20076 6928
rect 20128 6916 20134 6928
rect 21082 6916 21088 6928
rect 20128 6888 21088 6916
rect 20128 6876 20134 6888
rect 21082 6876 21088 6888
rect 21140 6876 21146 6928
rect 21928 6888 22232 6916
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12124 6820 12541 6848
rect 12124 6808 12130 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 12713 6851 12771 6857
rect 12713 6817 12725 6851
rect 12759 6848 12771 6851
rect 13906 6848 13912 6860
rect 12759 6820 13912 6848
rect 12759 6817 12771 6820
rect 12713 6811 12771 6817
rect 13906 6808 13912 6820
rect 13964 6848 13970 6860
rect 15013 6851 15071 6857
rect 15013 6848 15025 6851
rect 13964 6820 15025 6848
rect 13964 6808 13970 6820
rect 15013 6817 15025 6820
rect 15059 6817 15071 6851
rect 17770 6848 17776 6860
rect 15013 6811 15071 6817
rect 16960 6820 17448 6848
rect 17731 6820 17776 6848
rect 16960 6792 16988 6820
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 2406 6780 2412 6792
rect 2363 6752 2412 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 4031 6783 4089 6789
rect 4031 6749 4043 6783
rect 4077 6780 4089 6783
rect 4077 6752 4292 6780
rect 4077 6749 4089 6752
rect 4031 6743 4089 6749
rect 2516 6712 2544 6743
rect 4264 6724 4292 6752
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4396 6752 4441 6780
rect 4396 6740 4402 6752
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 4709 6783 4767 6789
rect 4709 6780 4721 6783
rect 4672 6752 4721 6780
rect 4672 6740 4678 6752
rect 4709 6749 4721 6752
rect 4755 6749 4767 6783
rect 4890 6780 4896 6792
rect 4851 6752 4896 6780
rect 4709 6743 4767 6749
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5534 6780 5540 6792
rect 5123 6752 5540 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 5534 6740 5540 6752
rect 5592 6780 5598 6792
rect 5722 6783 5780 6789
rect 5722 6780 5734 6783
rect 5592 6752 5734 6780
rect 5592 6740 5598 6752
rect 5722 6749 5734 6752
rect 5768 6749 5780 6783
rect 5722 6743 5780 6749
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 4154 6712 4160 6724
rect 2516 6684 4160 6712
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 4246 6672 4252 6724
rect 4304 6712 4310 6724
rect 4908 6712 4936 6740
rect 4304 6684 4936 6712
rect 4304 6672 4310 6684
rect 5994 6672 6000 6724
rect 6052 6712 6058 6724
rect 6104 6712 6132 6743
rect 6178 6740 6184 6792
rect 6236 6780 6242 6792
rect 6917 6783 6975 6789
rect 6236 6752 6281 6780
rect 6236 6740 6242 6752
rect 6917 6749 6929 6783
rect 6963 6780 6975 6783
rect 7098 6780 7104 6792
rect 6963 6752 7104 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 8214 6783 8272 6789
rect 8214 6780 8226 6783
rect 7800 6752 8226 6780
rect 7800 6740 7806 6752
rect 8214 6749 8226 6752
rect 8260 6749 8272 6783
rect 8214 6743 8272 6749
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 8444 6752 8493 6780
rect 8444 6740 8450 6752
rect 8481 6749 8493 6752
rect 8527 6749 8539 6783
rect 9490 6780 9496 6792
rect 9451 6752 9496 6780
rect 8481 6743 8539 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 9585 6783 9643 6789
rect 9585 6749 9597 6783
rect 9631 6749 9643 6783
rect 9585 6743 9643 6749
rect 6052 6684 7144 6712
rect 6052 6672 6058 6684
rect 3234 6604 3240 6656
rect 3292 6644 3298 6656
rect 7116 6653 7144 6684
rect 8846 6672 8852 6724
rect 8904 6712 8910 6724
rect 9309 6715 9367 6721
rect 9309 6712 9321 6715
rect 8904 6684 9321 6712
rect 8904 6672 8910 6684
rect 9309 6681 9321 6684
rect 9355 6681 9367 6715
rect 9309 6675 9367 6681
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3292 6616 3893 6644
rect 3292 6604 3298 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 3881 6607 3939 6613
rect 7101 6647 7159 6653
rect 7101 6613 7113 6647
rect 7147 6613 7159 6647
rect 7101 6607 7159 6613
rect 9125 6647 9183 6653
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 9214 6644 9220 6656
rect 9171 6616 9220 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 9214 6604 9220 6616
rect 9272 6644 9278 6656
rect 9600 6644 9628 6743
rect 11882 6740 11888 6792
rect 11940 6780 11946 6792
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11940 6752 11989 6780
rect 11940 6740 11946 6752
rect 11977 6749 11989 6752
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 16942 6740 16948 6792
rect 17000 6740 17006 6792
rect 17037 6783 17095 6789
rect 17037 6749 17049 6783
rect 17083 6780 17095 6783
rect 17126 6780 17132 6792
rect 17083 6752 17132 6780
rect 17083 6749 17095 6752
rect 17037 6743 17095 6749
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 11732 6715 11790 6721
rect 11732 6681 11744 6715
rect 11778 6712 11790 6715
rect 16792 6715 16850 6721
rect 11778 6684 12112 6712
rect 11778 6681 11790 6684
rect 11732 6675 11790 6681
rect 9272 6616 9628 6644
rect 10597 6647 10655 6653
rect 9272 6604 9278 6616
rect 10597 6613 10609 6647
rect 10643 6644 10655 6647
rect 11238 6644 11244 6656
rect 10643 6616 11244 6644
rect 10643 6613 10655 6616
rect 10597 6607 10655 6613
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 12084 6653 12112 6684
rect 16792 6681 16804 6715
rect 16838 6712 16850 6715
rect 17420 6712 17448 6820
rect 17770 6808 17776 6820
rect 17828 6808 17834 6860
rect 19613 6851 19671 6857
rect 19613 6817 19625 6851
rect 19659 6848 19671 6851
rect 19794 6848 19800 6860
rect 19659 6820 19800 6848
rect 19659 6817 19671 6820
rect 19613 6811 19671 6817
rect 19794 6808 19800 6820
rect 19852 6848 19858 6860
rect 20438 6848 20444 6860
rect 19852 6820 20444 6848
rect 19852 6808 19858 6820
rect 20438 6808 20444 6820
rect 20496 6808 20502 6860
rect 20530 6808 20536 6860
rect 20588 6848 20594 6860
rect 20717 6851 20775 6857
rect 20717 6848 20729 6851
rect 20588 6820 20729 6848
rect 20588 6808 20594 6820
rect 20717 6817 20729 6820
rect 20763 6817 20775 6851
rect 20717 6811 20775 6817
rect 20901 6851 20959 6857
rect 20901 6817 20913 6851
rect 20947 6848 20959 6851
rect 21266 6848 21272 6860
rect 20947 6820 21272 6848
rect 20947 6817 20959 6820
rect 20901 6811 20959 6817
rect 21266 6808 21272 6820
rect 21324 6808 21330 6860
rect 21358 6808 21364 6860
rect 21416 6848 21422 6860
rect 21729 6851 21787 6857
rect 21416 6820 21461 6848
rect 21416 6808 21422 6820
rect 21729 6817 21741 6851
rect 21775 6848 21787 6851
rect 21928 6848 21956 6888
rect 22094 6848 22100 6860
rect 21775 6820 21956 6848
rect 21775 6817 21787 6820
rect 21729 6811 21787 6817
rect 22066 6808 22100 6848
rect 22152 6808 22158 6860
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6780 17555 6783
rect 17954 6780 17960 6792
rect 17543 6752 17960 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 18782 6780 18788 6792
rect 18743 6752 18788 6780
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 18874 6740 18880 6792
rect 18932 6780 18938 6792
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 18932 6752 19717 6780
rect 18932 6740 18938 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 20456 6780 20484 6808
rect 21542 6780 21548 6792
rect 20456 6774 20576 6780
rect 20456 6752 20668 6774
rect 21503 6752 21548 6780
rect 19705 6743 19763 6749
rect 20548 6746 20668 6752
rect 20070 6712 20076 6724
rect 16838 6684 17172 6712
rect 17420 6684 20076 6712
rect 16838 6681 16850 6684
rect 16792 6675 16850 6681
rect 12069 6647 12127 6653
rect 12069 6613 12081 6647
rect 12115 6613 12127 6647
rect 12069 6607 12127 6613
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 12308 6616 12449 6644
rect 12308 6604 12314 6616
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 14458 6644 14464 6656
rect 14419 6616 14464 6644
rect 12437 6607 12495 6613
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 14826 6644 14832 6656
rect 14787 6616 14832 6644
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 14918 6604 14924 6656
rect 14976 6644 14982 6656
rect 17144 6653 17172 6684
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 17129 6647 17187 6653
rect 14976 6616 15021 6644
rect 14976 6604 14982 6616
rect 17129 6613 17141 6647
rect 17175 6613 17187 6647
rect 17129 6607 17187 6613
rect 17589 6647 17647 6653
rect 17589 6613 17601 6647
rect 17635 6644 17647 6647
rect 17954 6644 17960 6656
rect 17635 6616 17960 6644
rect 17635 6613 17647 6616
rect 17589 6607 17647 6613
rect 17954 6604 17960 6616
rect 18012 6644 18018 6656
rect 18230 6644 18236 6656
rect 18012 6616 18236 6644
rect 18012 6604 18018 6616
rect 18230 6604 18236 6616
rect 18288 6604 18294 6656
rect 20165 6647 20223 6653
rect 20165 6613 20177 6647
rect 20211 6644 20223 6647
rect 20254 6644 20260 6656
rect 20211 6616 20260 6644
rect 20211 6613 20223 6616
rect 20165 6607 20223 6613
rect 20254 6604 20260 6616
rect 20312 6644 20318 6656
rect 20530 6644 20536 6656
rect 20312 6616 20536 6644
rect 20312 6604 20318 6616
rect 20530 6604 20536 6616
rect 20588 6604 20594 6656
rect 20640 6653 20668 6746
rect 21542 6740 21548 6752
rect 21600 6740 21606 6792
rect 21913 6783 21971 6789
rect 21913 6749 21925 6783
rect 21959 6780 21971 6783
rect 22066 6780 22094 6808
rect 21959 6752 22094 6780
rect 22204 6780 22232 6888
rect 22296 6848 22324 6956
rect 25774 6944 25780 6956
rect 25832 6944 25838 6996
rect 22646 6876 22652 6928
rect 22704 6916 22710 6928
rect 23201 6919 23259 6925
rect 23201 6916 23213 6919
rect 22704 6888 23213 6916
rect 22704 6876 22710 6888
rect 23201 6885 23213 6888
rect 23247 6885 23259 6919
rect 23201 6879 23259 6885
rect 23382 6876 23388 6928
rect 23440 6916 23446 6928
rect 23440 6888 24808 6916
rect 23440 6876 23446 6888
rect 22465 6851 22523 6857
rect 22296 6820 22416 6848
rect 22278 6780 22284 6792
rect 22204 6752 22284 6780
rect 21959 6749 21971 6752
rect 21913 6743 21971 6749
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 22388 6789 22416 6820
rect 22465 6817 22477 6851
rect 22511 6848 22523 6851
rect 22922 6848 22928 6860
rect 22511 6820 22928 6848
rect 22511 6817 22523 6820
rect 22465 6811 22523 6817
rect 22922 6808 22928 6820
rect 22980 6808 22986 6860
rect 22373 6783 22431 6789
rect 22373 6749 22385 6783
rect 22419 6749 22431 6783
rect 22373 6743 22431 6749
rect 22741 6783 22799 6789
rect 22741 6749 22753 6783
rect 22787 6749 22799 6783
rect 22741 6743 22799 6749
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6780 22891 6783
rect 23198 6780 23204 6792
rect 22879 6752 23204 6780
rect 22879 6749 22891 6752
rect 22833 6743 22891 6749
rect 22005 6715 22063 6721
rect 22005 6681 22017 6715
rect 22051 6712 22063 6715
rect 22462 6712 22468 6724
rect 22051 6684 22468 6712
rect 22051 6681 22063 6684
rect 22005 6675 22063 6681
rect 22462 6672 22468 6684
rect 22520 6672 22526 6724
rect 20625 6647 20683 6653
rect 20625 6613 20637 6647
rect 20671 6613 20683 6647
rect 20625 6607 20683 6613
rect 21542 6604 21548 6656
rect 21600 6644 21606 6656
rect 22756 6644 22784 6743
rect 23198 6740 23204 6752
rect 23256 6740 23262 6792
rect 24673 6783 24731 6789
rect 24673 6749 24685 6783
rect 24719 6749 24731 6783
rect 24780 6780 24808 6888
rect 24854 6876 24860 6928
rect 24912 6876 24918 6928
rect 24872 6848 24900 6876
rect 24949 6851 25007 6857
rect 24949 6848 24961 6851
rect 24872 6820 24961 6848
rect 24949 6817 24961 6820
rect 24995 6817 25007 6851
rect 24949 6811 25007 6817
rect 24857 6783 24915 6789
rect 24857 6780 24869 6783
rect 24780 6752 24869 6780
rect 24673 6743 24731 6749
rect 24857 6749 24869 6752
rect 24903 6749 24915 6783
rect 24857 6743 24915 6749
rect 24688 6712 24716 6743
rect 25038 6740 25044 6792
rect 25096 6780 25102 6792
rect 25133 6783 25191 6789
rect 25133 6780 25145 6783
rect 25096 6752 25145 6780
rect 25096 6740 25102 6752
rect 25133 6749 25145 6752
rect 25179 6749 25191 6783
rect 25314 6780 25320 6792
rect 25275 6752 25320 6780
rect 25133 6743 25191 6749
rect 25314 6740 25320 6752
rect 25372 6740 25378 6792
rect 25961 6783 26019 6789
rect 25961 6780 25973 6783
rect 25424 6752 25973 6780
rect 24688 6684 24900 6712
rect 24872 6656 24900 6684
rect 24946 6672 24952 6724
rect 25004 6712 25010 6724
rect 25424 6712 25452 6752
rect 25961 6749 25973 6752
rect 26007 6749 26019 6783
rect 25961 6743 26019 6749
rect 25004 6684 25452 6712
rect 25004 6672 25010 6684
rect 25498 6672 25504 6724
rect 25556 6712 25562 6724
rect 25556 6684 25601 6712
rect 25556 6672 25562 6684
rect 25682 6672 25688 6724
rect 25740 6712 25746 6724
rect 26206 6715 26264 6721
rect 26206 6712 26218 6715
rect 25740 6684 25785 6712
rect 25884 6684 26218 6712
rect 25740 6672 25746 6684
rect 21600 6616 22784 6644
rect 21600 6604 21606 6616
rect 24854 6604 24860 6656
rect 24912 6604 24918 6656
rect 25130 6604 25136 6656
rect 25188 6644 25194 6656
rect 25884 6644 25912 6684
rect 26206 6681 26218 6684
rect 26252 6681 26264 6715
rect 26206 6675 26264 6681
rect 25188 6616 25912 6644
rect 27341 6647 27399 6653
rect 25188 6604 25194 6616
rect 27341 6613 27353 6647
rect 27387 6644 27399 6647
rect 27706 6644 27712 6656
rect 27387 6616 27712 6644
rect 27387 6613 27399 6616
rect 27341 6607 27399 6613
rect 27706 6604 27712 6616
rect 27764 6604 27770 6656
rect 1104 6554 29440 6576
rect 1104 6502 10395 6554
rect 10447 6502 10459 6554
rect 10511 6502 10523 6554
rect 10575 6502 10587 6554
rect 10639 6502 10651 6554
rect 10703 6502 19840 6554
rect 19892 6502 19904 6554
rect 19956 6502 19968 6554
rect 20020 6502 20032 6554
rect 20084 6502 20096 6554
rect 20148 6502 29440 6554
rect 1104 6480 29440 6502
rect 2869 6443 2927 6449
rect 2869 6409 2881 6443
rect 2915 6440 2927 6443
rect 4338 6440 4344 6452
rect 2915 6412 4344 6440
rect 2915 6409 2927 6412
rect 2869 6403 2927 6409
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 5537 6443 5595 6449
rect 5537 6440 5549 6443
rect 4672 6412 5549 6440
rect 4672 6400 4678 6412
rect 5537 6409 5549 6412
rect 5583 6409 5595 6443
rect 10226 6440 10232 6452
rect 5537 6403 5595 6409
rect 5828 6412 10232 6440
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 5828 6372 5856 6412
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6440 12035 6443
rect 12066 6440 12072 6452
rect 12023 6412 12072 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 12250 6440 12256 6452
rect 12211 6412 12256 6440
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 14918 6400 14924 6452
rect 14976 6440 14982 6452
rect 15841 6443 15899 6449
rect 15841 6440 15853 6443
rect 14976 6412 15853 6440
rect 14976 6400 14982 6412
rect 15841 6409 15853 6412
rect 15887 6409 15899 6443
rect 15841 6403 15899 6409
rect 18877 6443 18935 6449
rect 18877 6409 18889 6443
rect 18923 6440 18935 6443
rect 20346 6440 20352 6452
rect 18923 6412 20352 6440
rect 18923 6409 18935 6412
rect 18877 6403 18935 6409
rect 20088 6384 20116 6412
rect 20346 6400 20352 6412
rect 20404 6440 20410 6452
rect 22462 6440 22468 6452
rect 20404 6412 20668 6440
rect 22423 6412 22468 6440
rect 20404 6400 20410 6412
rect 5994 6372 6000 6384
rect 4120 6344 5856 6372
rect 5955 6344 6000 6372
rect 4120 6332 4126 6344
rect 5994 6332 6000 6344
rect 6052 6332 6058 6384
rect 11054 6372 11060 6384
rect 9140 6344 11060 6372
rect 1756 6307 1814 6313
rect 1756 6273 1768 6307
rect 1802 6304 1814 6307
rect 2222 6304 2228 6316
rect 1802 6276 2228 6304
rect 1802 6273 1814 6276
rect 1756 6267 1814 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 3234 6304 3240 6316
rect 3195 6276 3240 6304
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 4304 6276 4353 6304
rect 4304 6264 4310 6276
rect 4341 6273 4353 6276
rect 4387 6304 4399 6307
rect 4614 6304 4620 6316
rect 4387 6276 4620 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 4800 6307 4858 6313
rect 4800 6273 4812 6307
rect 4846 6304 4858 6307
rect 4890 6304 4896 6316
rect 4846 6276 4896 6304
rect 4846 6273 4858 6276
rect 4800 6267 4858 6273
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 6178 6304 6184 6316
rect 5767 6276 6184 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 6178 6264 6184 6276
rect 6236 6304 6242 6316
rect 6236 6276 6316 6304
rect 6236 6264 6242 6276
rect 1486 6236 1492 6248
rect 1447 6208 1492 6236
rect 1486 6196 1492 6208
rect 1544 6196 1550 6248
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 5813 6239 5871 6245
rect 5813 6236 5825 6239
rect 4479 6208 5825 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4816 6180 4844 6208
rect 5813 6205 5825 6208
rect 5859 6205 5871 6239
rect 6288 6236 6316 6276
rect 6362 6264 6368 6316
rect 6420 6304 6426 6316
rect 8846 6304 8852 6316
rect 6420 6276 6465 6304
rect 8807 6276 8852 6304
rect 6420 6264 6426 6276
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 9140 6313 9168 6344
rect 11054 6332 11060 6344
rect 11112 6372 11118 6384
rect 11882 6372 11888 6384
rect 11112 6344 11888 6372
rect 11112 6332 11118 6344
rect 11882 6332 11888 6344
rect 11940 6372 11946 6384
rect 14458 6381 14464 6384
rect 14452 6372 14464 6381
rect 11940 6344 14228 6372
rect 14419 6344 14464 6372
rect 11940 6332 11946 6344
rect 9398 6313 9404 6316
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9392 6267 9404 6313
rect 9456 6304 9462 6316
rect 9456 6276 9492 6304
rect 9398 6264 9404 6267
rect 9456 6264 9462 6276
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 11793 6307 11851 6313
rect 11793 6304 11805 6307
rect 11756 6276 11805 6304
rect 11756 6264 11762 6276
rect 11793 6273 11805 6276
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 6288 6208 6469 6236
rect 5813 6199 5871 6205
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 4798 6128 4804 6180
rect 4856 6128 4862 6180
rect 5442 6128 5448 6180
rect 5500 6168 5506 6180
rect 5500 6140 5764 6168
rect 5500 6128 5506 6140
rect 3053 6103 3111 6109
rect 3053 6069 3065 6103
rect 3099 6100 3111 6103
rect 3326 6100 3332 6112
rect 3099 6072 3332 6100
rect 3099 6069 3111 6072
rect 3053 6063 3111 6069
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 4893 6103 4951 6109
rect 4893 6069 4905 6103
rect 4939 6100 4951 6103
rect 5258 6100 5264 6112
rect 4939 6072 5264 6100
rect 4939 6069 4951 6072
rect 4893 6063 4951 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5736 6109 5764 6140
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 6733 6171 6791 6177
rect 6733 6168 6745 6171
rect 6052 6140 6745 6168
rect 6052 6128 6058 6140
rect 6733 6137 6745 6140
rect 6779 6137 6791 6171
rect 11992 6168 12020 6267
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12216 6276 12261 6304
rect 12216 6264 12222 6276
rect 12406 6248 12434 6344
rect 12894 6313 12900 6316
rect 12888 6267 12900 6313
rect 12952 6304 12958 6316
rect 14200 6313 14228 6344
rect 14452 6335 14464 6344
rect 14458 6332 14464 6335
rect 14516 6332 14522 6384
rect 18049 6375 18107 6381
rect 15396 6344 16068 6372
rect 14185 6307 14243 6313
rect 12952 6276 12988 6304
rect 12894 6264 12900 6267
rect 12952 6264 12958 6276
rect 14185 6273 14197 6307
rect 14231 6273 14243 6307
rect 15396 6304 15424 6344
rect 14185 6267 14243 6273
rect 14292 6276 15424 6304
rect 12342 6196 12348 6248
rect 12400 6236 12434 6248
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12400 6208 12633 6236
rect 12400 6196 12406 6208
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 14292 6236 14320 6276
rect 15470 6264 15476 6316
rect 15528 6304 15534 6316
rect 16040 6313 16068 6344
rect 18049 6341 18061 6375
rect 18095 6372 18107 6375
rect 18690 6372 18696 6384
rect 18095 6344 18696 6372
rect 18095 6341 18107 6344
rect 18049 6335 18107 6341
rect 18690 6332 18696 6344
rect 18748 6332 18754 6384
rect 20070 6332 20076 6384
rect 20128 6332 20134 6384
rect 20640 6381 20668 6412
rect 22462 6400 22468 6412
rect 22520 6400 22526 6452
rect 22557 6443 22615 6449
rect 22557 6409 22569 6443
rect 22603 6440 22615 6443
rect 22646 6440 22652 6452
rect 22603 6412 22652 6440
rect 22603 6409 22615 6412
rect 22557 6403 22615 6409
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 22922 6440 22928 6452
rect 22883 6412 22928 6440
rect 22922 6400 22928 6412
rect 22980 6400 22986 6452
rect 24762 6440 24768 6452
rect 24723 6412 24768 6440
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 25130 6440 25136 6452
rect 25091 6412 25136 6440
rect 25130 6400 25136 6412
rect 25188 6400 25194 6452
rect 25314 6400 25320 6452
rect 25372 6440 25378 6452
rect 25501 6443 25559 6449
rect 25501 6440 25513 6443
rect 25372 6412 25513 6440
rect 25372 6400 25378 6412
rect 25501 6409 25513 6412
rect 25547 6409 25559 6443
rect 25501 6403 25559 6409
rect 25869 6443 25927 6449
rect 25869 6409 25881 6443
rect 25915 6440 25927 6443
rect 25958 6440 25964 6452
rect 25915 6412 25964 6440
rect 25915 6409 25927 6412
rect 25869 6403 25927 6409
rect 25958 6400 25964 6412
rect 26016 6400 26022 6452
rect 20625 6375 20683 6381
rect 20625 6341 20637 6375
rect 20671 6341 20683 6375
rect 20625 6335 20683 6341
rect 20993 6375 21051 6381
rect 20993 6341 21005 6375
rect 21039 6372 21051 6375
rect 21542 6372 21548 6384
rect 21039 6344 21548 6372
rect 21039 6341 21051 6344
rect 20993 6335 21051 6341
rect 21542 6332 21548 6344
rect 21600 6332 21606 6384
rect 26234 6372 26240 6384
rect 22066 6344 26240 6372
rect 15841 6307 15899 6313
rect 15841 6304 15853 6307
rect 15528 6276 15853 6304
rect 15528 6264 15534 6276
rect 15841 6273 15853 6276
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6304 16083 6307
rect 16942 6304 16948 6316
rect 16071 6276 16948 6304
rect 16071 6273 16083 6276
rect 16025 6267 16083 6273
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 17954 6304 17960 6316
rect 17867 6276 17960 6304
rect 17954 6264 17960 6276
rect 18012 6304 18018 6316
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 18012 6276 18521 6304
rect 18012 6264 18018 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 18598 6264 18604 6316
rect 18656 6304 18662 6316
rect 19886 6304 19892 6316
rect 18656 6276 18701 6304
rect 19847 6276 19892 6304
rect 18656 6264 18662 6276
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 20806 6304 20812 6316
rect 20767 6276 20812 6304
rect 20806 6264 20812 6276
rect 20864 6264 20870 6316
rect 22066 6304 22094 6344
rect 26234 6332 26240 6344
rect 26292 6332 26298 6384
rect 20916 6276 22094 6304
rect 12621 6199 12679 6205
rect 13924 6208 14320 6236
rect 17865 6239 17923 6245
rect 11992 6140 12434 6168
rect 6733 6131 6791 6137
rect 5721 6103 5779 6109
rect 5721 6069 5733 6103
rect 5767 6100 5779 6103
rect 6365 6103 6423 6109
rect 6365 6100 6377 6103
rect 5767 6072 6377 6100
rect 5767 6069 5779 6072
rect 5721 6063 5779 6069
rect 6365 6069 6377 6072
rect 6411 6069 6423 6103
rect 6365 6063 6423 6069
rect 9033 6103 9091 6109
rect 9033 6069 9045 6103
rect 9079 6100 9091 6103
rect 9766 6100 9772 6112
rect 9079 6072 9772 6100
rect 9079 6069 9091 6072
rect 9033 6063 9091 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10505 6103 10563 6109
rect 10505 6069 10517 6103
rect 10551 6100 10563 6103
rect 11146 6100 11152 6112
rect 10551 6072 11152 6100
rect 10551 6069 10563 6072
rect 10505 6063 10563 6069
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11698 6060 11704 6112
rect 11756 6100 11762 6112
rect 12158 6100 12164 6112
rect 11756 6072 12164 6100
rect 11756 6060 11762 6072
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12406 6100 12434 6140
rect 13924 6100 13952 6208
rect 17865 6205 17877 6239
rect 17911 6236 17923 6239
rect 18046 6236 18052 6248
rect 17911 6208 18052 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 20916 6236 20944 6276
rect 23198 6264 23204 6316
rect 23256 6304 23262 6316
rect 23293 6307 23351 6313
rect 23293 6304 23305 6307
rect 23256 6276 23305 6304
rect 23256 6264 23262 6276
rect 23293 6273 23305 6276
rect 23339 6273 23351 6307
rect 23293 6267 23351 6273
rect 24854 6264 24860 6316
rect 24912 6304 24918 6316
rect 25409 6307 25467 6313
rect 25409 6304 25421 6307
rect 24912 6276 25421 6304
rect 24912 6264 24918 6276
rect 25409 6273 25421 6276
rect 25455 6304 25467 6307
rect 25498 6304 25504 6316
rect 25455 6276 25504 6304
rect 25455 6273 25467 6276
rect 25409 6267 25467 6273
rect 25498 6264 25504 6276
rect 25556 6304 25562 6316
rect 25556 6276 26004 6304
rect 25556 6264 25562 6276
rect 25976 6248 26004 6276
rect 22649 6239 22707 6245
rect 22649 6236 22661 6239
rect 18156 6208 20944 6236
rect 22066 6208 22661 6236
rect 18156 6168 18184 6208
rect 15120 6140 18184 6168
rect 18417 6171 18475 6177
rect 12406 6072 13952 6100
rect 14001 6103 14059 6109
rect 14001 6069 14013 6103
rect 14047 6100 14059 6103
rect 14366 6100 14372 6112
rect 14047 6072 14372 6100
rect 14047 6069 14059 6072
rect 14001 6063 14059 6069
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 14550 6060 14556 6112
rect 14608 6100 14614 6112
rect 15120 6100 15148 6140
rect 18417 6137 18429 6171
rect 18463 6168 18475 6171
rect 19334 6168 19340 6180
rect 18463 6140 19340 6168
rect 18463 6137 18475 6140
rect 18417 6131 18475 6137
rect 19334 6128 19340 6140
rect 19392 6168 19398 6180
rect 22066 6168 22094 6208
rect 22649 6205 22661 6208
rect 22695 6205 22707 6239
rect 23382 6236 23388 6248
rect 23343 6208 23388 6236
rect 22649 6199 22707 6205
rect 23382 6196 23388 6208
rect 23440 6196 23446 6248
rect 23477 6239 23535 6245
rect 23477 6205 23489 6239
rect 23523 6205 23535 6239
rect 24486 6236 24492 6248
rect 24447 6208 24492 6236
rect 23477 6199 23535 6205
rect 19392 6140 22094 6168
rect 19392 6128 19398 6140
rect 23014 6128 23020 6180
rect 23072 6168 23078 6180
rect 23492 6168 23520 6199
rect 24486 6196 24492 6208
rect 24544 6196 24550 6248
rect 24673 6239 24731 6245
rect 24673 6205 24685 6239
rect 24719 6236 24731 6239
rect 25317 6239 25375 6245
rect 25317 6236 25329 6239
rect 24719 6208 25329 6236
rect 24719 6205 24731 6208
rect 24673 6199 24731 6205
rect 25317 6205 25329 6208
rect 25363 6205 25375 6239
rect 25958 6236 25964 6248
rect 25919 6208 25964 6236
rect 25317 6199 25375 6205
rect 23072 6140 23520 6168
rect 23072 6128 23078 6140
rect 24118 6128 24124 6180
rect 24176 6168 24182 6180
rect 24688 6168 24716 6199
rect 25958 6196 25964 6208
rect 26016 6196 26022 6248
rect 26053 6239 26111 6245
rect 26053 6205 26065 6239
rect 26099 6205 26111 6239
rect 26053 6199 26111 6205
rect 26068 6168 26096 6199
rect 24176 6140 24716 6168
rect 25976 6140 26096 6168
rect 24176 6128 24182 6140
rect 15562 6100 15568 6112
rect 14608 6072 15148 6100
rect 15523 6072 15568 6100
rect 14608 6060 14614 6072
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 18782 6100 18788 6112
rect 18739 6072 18788 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 18782 6060 18788 6072
rect 18840 6060 18846 6112
rect 19702 6100 19708 6112
rect 19663 6072 19708 6100
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 22097 6103 22155 6109
rect 22097 6069 22109 6103
rect 22143 6100 22155 6103
rect 22186 6100 22192 6112
rect 22143 6072 22192 6100
rect 22143 6069 22155 6072
rect 22097 6063 22155 6069
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 24394 6060 24400 6112
rect 24452 6100 24458 6112
rect 25976 6100 26004 6140
rect 24452 6072 26004 6100
rect 24452 6060 24458 6072
rect 1104 6010 29440 6032
rect 1104 5958 5672 6010
rect 5724 5958 5736 6010
rect 5788 5958 5800 6010
rect 5852 5958 5864 6010
rect 5916 5958 5928 6010
rect 5980 5958 15118 6010
rect 15170 5958 15182 6010
rect 15234 5958 15246 6010
rect 15298 5958 15310 6010
rect 15362 5958 15374 6010
rect 15426 5958 24563 6010
rect 24615 5958 24627 6010
rect 24679 5958 24691 6010
rect 24743 5958 24755 6010
rect 24807 5958 24819 6010
rect 24871 5958 29440 6010
rect 1104 5936 29440 5958
rect 2222 5896 2228 5908
rect 2183 5868 2228 5896
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 4890 5896 4896 5908
rect 4851 5868 4896 5896
rect 4890 5856 4896 5868
rect 4948 5896 4954 5908
rect 6086 5896 6092 5908
rect 4948 5868 6092 5896
rect 4948 5856 4954 5868
rect 5828 5840 5856 5868
rect 6086 5856 6092 5868
rect 6144 5896 6150 5908
rect 6362 5896 6368 5908
rect 6144 5868 6368 5896
rect 6144 5856 6150 5868
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 9309 5899 9367 5905
rect 9309 5865 9321 5899
rect 9355 5896 9367 5899
rect 9398 5896 9404 5908
rect 9355 5868 9404 5896
rect 9355 5865 9367 5868
rect 9309 5859 9367 5865
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 14826 5856 14832 5908
rect 14884 5896 14890 5908
rect 15381 5899 15439 5905
rect 15381 5896 15393 5899
rect 14884 5868 15393 5896
rect 14884 5856 14890 5868
rect 15381 5865 15393 5868
rect 15427 5865 15439 5899
rect 18690 5896 18696 5908
rect 18651 5868 18696 5896
rect 15381 5859 15439 5865
rect 18690 5856 18696 5868
rect 18748 5856 18754 5908
rect 18800 5868 19748 5896
rect 2590 5788 2596 5840
rect 2648 5828 2654 5840
rect 3605 5831 3663 5837
rect 2648 5800 2774 5828
rect 2648 5788 2654 5800
rect 2746 5760 2774 5800
rect 3605 5797 3617 5831
rect 3651 5828 3663 5831
rect 4154 5828 4160 5840
rect 3651 5800 4160 5828
rect 3651 5797 3663 5800
rect 3605 5791 3663 5797
rect 3988 5769 4016 5800
rect 4154 5788 4160 5800
rect 4212 5788 4218 5840
rect 5810 5788 5816 5840
rect 5868 5788 5874 5840
rect 6178 5788 6184 5840
rect 6236 5828 6242 5840
rect 7193 5831 7251 5837
rect 7193 5828 7205 5831
rect 6236 5800 7205 5828
rect 6236 5788 6242 5800
rect 7193 5797 7205 5800
rect 7239 5797 7251 5831
rect 15286 5828 15292 5840
rect 7193 5791 7251 5797
rect 14844 5800 15292 5828
rect 2869 5763 2927 5769
rect 2869 5760 2881 5763
rect 2746 5732 2881 5760
rect 2869 5729 2881 5732
rect 2915 5760 2927 5763
rect 3973 5763 4031 5769
rect 2915 5732 3924 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 3326 5692 3332 5704
rect 2639 5664 3332 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5692 3571 5695
rect 3605 5695 3663 5701
rect 3605 5692 3617 5695
rect 3559 5664 3617 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 3605 5661 3617 5664
rect 3651 5661 3663 5695
rect 3605 5655 3663 5661
rect 2682 5516 2688 5568
rect 2740 5556 2746 5568
rect 3142 5556 3148 5568
rect 2740 5528 2785 5556
rect 3103 5528 3148 5556
rect 2740 5516 2746 5528
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 3896 5565 3924 5732
rect 3973 5729 3985 5763
rect 4019 5760 4031 5763
rect 4706 5760 4712 5772
rect 4019 5732 4712 5760
rect 4019 5729 4031 5732
rect 3973 5723 4031 5729
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5760 5411 5763
rect 6270 5760 6276 5772
rect 5399 5732 6276 5760
rect 5399 5729 5411 5732
rect 5353 5723 5411 5729
rect 6270 5720 6276 5732
rect 6328 5760 6334 5772
rect 9766 5760 9772 5772
rect 6328 5732 6408 5760
rect 9727 5732 9772 5760
rect 6328 5720 6334 5732
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5692 4215 5695
rect 4246 5692 4252 5704
rect 4203 5664 4252 5692
rect 4203 5661 4215 5664
rect 4157 5655 4215 5661
rect 4246 5652 4252 5664
rect 4304 5692 4310 5704
rect 5258 5692 5264 5704
rect 4304 5664 5120 5692
rect 5219 5664 5264 5692
rect 4304 5652 4310 5664
rect 4614 5624 4620 5636
rect 4575 5596 4620 5624
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 4798 5624 4804 5636
rect 4759 5596 4804 5624
rect 4798 5584 4804 5596
rect 4856 5584 4862 5636
rect 3881 5559 3939 5565
rect 3881 5525 3893 5559
rect 3927 5556 3939 5559
rect 4062 5556 4068 5568
rect 3927 5528 4068 5556
rect 3927 5525 3939 5528
rect 3881 5519 3939 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4341 5559 4399 5565
rect 4341 5525 4353 5559
rect 4387 5556 4399 5559
rect 4890 5556 4896 5568
rect 4387 5528 4896 5556
rect 4387 5525 4399 5528
rect 4341 5519 4399 5525
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 5092 5565 5120 5664
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5442 5692 5448 5704
rect 5403 5664 5448 5692
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5812 5695 5870 5701
rect 5812 5661 5824 5695
rect 5858 5692 5870 5695
rect 5902 5692 5908 5704
rect 5858 5664 5908 5692
rect 5858 5661 5870 5664
rect 5812 5655 5870 5661
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6086 5692 6092 5704
rect 6047 5664 6092 5692
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6178 5652 6184 5704
rect 6236 5692 6242 5704
rect 6380 5692 6408 5732
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 9858 5720 9864 5772
rect 9916 5760 9922 5772
rect 9916 5732 9961 5760
rect 9916 5720 9922 5732
rect 6491 5695 6549 5701
rect 6491 5692 6503 5695
rect 6236 5664 6281 5692
rect 6380 5664 6503 5692
rect 6236 5652 6242 5664
rect 6491 5661 6503 5664
rect 6537 5661 6549 5695
rect 6491 5655 6549 5661
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5692 6791 5695
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 6779 5664 6837 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 6825 5661 6837 5664
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 8478 5652 8484 5704
rect 8536 5692 8542 5704
rect 8573 5695 8631 5701
rect 8573 5692 8585 5695
rect 8536 5664 8585 5692
rect 8536 5652 8542 5664
rect 8573 5661 8585 5664
rect 8619 5661 8631 5695
rect 11238 5692 11244 5704
rect 11199 5664 11244 5692
rect 8573 5655 8631 5661
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 11514 5692 11520 5704
rect 11475 5664 11520 5692
rect 11514 5652 11520 5664
rect 11572 5652 11578 5704
rect 12986 5692 12992 5704
rect 12947 5664 12992 5692
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 13814 5692 13820 5704
rect 13587 5664 13820 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 14550 5652 14556 5704
rect 14608 5692 14614 5704
rect 14844 5701 14872 5800
rect 15286 5788 15292 5800
rect 15344 5828 15350 5840
rect 15562 5828 15568 5840
rect 15344 5800 15568 5828
rect 15344 5788 15350 5800
rect 15562 5788 15568 5800
rect 15620 5788 15626 5840
rect 18800 5828 18828 5868
rect 19610 5828 19616 5840
rect 18524 5800 18828 5828
rect 19571 5800 19616 5828
rect 15105 5763 15163 5769
rect 15105 5729 15117 5763
rect 15151 5760 15163 5763
rect 15151 5732 15516 5760
rect 15151 5729 15163 5732
rect 15105 5723 15163 5729
rect 15488 5704 15516 5732
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 14608 5664 14657 5692
rect 14608 5652 14614 5664
rect 14645 5661 14657 5664
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5661 14887 5695
rect 15194 5692 15200 5704
rect 15155 5664 15200 5692
rect 14829 5655 14887 5661
rect 15194 5652 15200 5664
rect 15252 5652 15258 5704
rect 15470 5692 15476 5704
rect 15431 5664 15476 5692
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 17586 5692 17592 5704
rect 17547 5664 17592 5692
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5692 17831 5695
rect 18414 5692 18420 5704
rect 17819 5664 18420 5692
rect 17819 5661 17831 5664
rect 17773 5655 17831 5661
rect 18414 5652 18420 5664
rect 18472 5652 18478 5704
rect 18524 5701 18552 5800
rect 19610 5788 19616 5800
rect 19668 5788 19674 5840
rect 19720 5828 19748 5868
rect 19886 5856 19892 5908
rect 19944 5896 19950 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 19944 5868 20637 5896
rect 19944 5856 19950 5868
rect 20625 5865 20637 5868
rect 20671 5865 20683 5899
rect 20625 5859 20683 5865
rect 20806 5856 20812 5908
rect 20864 5896 20870 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20864 5868 20913 5896
rect 20864 5856 20870 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 21082 5896 21088 5908
rect 21043 5868 21088 5896
rect 20901 5859 20959 5865
rect 20070 5828 20076 5840
rect 19720 5800 20076 5828
rect 20070 5788 20076 5800
rect 20128 5788 20134 5840
rect 19426 5760 19432 5772
rect 18616 5732 19432 5760
rect 18616 5701 18644 5732
rect 19426 5720 19432 5732
rect 19484 5760 19490 5772
rect 19484 5732 20392 5760
rect 19484 5720 19490 5732
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5661 18567 5695
rect 18509 5655 18567 5661
rect 18601 5695 18659 5701
rect 18601 5661 18613 5695
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 18690 5652 18696 5704
rect 18748 5692 18754 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 18748 5664 18793 5692
rect 18984 5664 19257 5692
rect 18748 5652 18754 5664
rect 5994 5624 6000 5636
rect 5955 5596 6000 5624
rect 5994 5584 6000 5596
rect 6052 5584 6058 5636
rect 8294 5624 8300 5636
rect 8352 5633 8358 5636
rect 8264 5596 8300 5624
rect 8294 5584 8300 5596
rect 8352 5587 8364 5633
rect 11609 5627 11667 5633
rect 11609 5593 11621 5627
rect 11655 5624 11667 5627
rect 12066 5624 12072 5636
rect 11655 5596 12072 5624
rect 11655 5593 11667 5596
rect 11609 5587 11667 5593
rect 8352 5584 8358 5587
rect 12066 5584 12072 5596
rect 12124 5584 12130 5636
rect 5077 5559 5135 5565
rect 5077 5525 5089 5559
rect 5123 5525 5135 5559
rect 7006 5556 7012 5568
rect 6967 5528 7012 5556
rect 5077 5519 5135 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 9677 5559 9735 5565
rect 9677 5556 9689 5559
rect 9548 5528 9689 5556
rect 9548 5516 9554 5528
rect 9677 5525 9689 5528
rect 9723 5556 9735 5559
rect 12618 5556 12624 5568
rect 9723 5528 12624 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 13170 5556 13176 5568
rect 13131 5528 13176 5556
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 13262 5516 13268 5568
rect 13320 5556 13326 5568
rect 13357 5559 13415 5565
rect 13357 5556 13369 5559
rect 13320 5528 13369 5556
rect 13320 5516 13326 5528
rect 13357 5525 13369 5528
rect 13403 5525 13415 5559
rect 17678 5556 17684 5568
rect 17639 5528 17684 5556
rect 13357 5519 13415 5525
rect 17678 5516 17684 5528
rect 17736 5516 17742 5568
rect 18046 5516 18052 5568
rect 18104 5556 18110 5568
rect 18984 5565 19012 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19518 5692 19524 5704
rect 19479 5664 19524 5692
rect 19245 5655 19303 5661
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 19705 5695 19763 5701
rect 19705 5661 19717 5695
rect 19751 5661 19763 5695
rect 20070 5692 20076 5704
rect 20031 5664 20076 5692
rect 19705 5655 19763 5661
rect 18417 5559 18475 5565
rect 18417 5556 18429 5559
rect 18104 5528 18429 5556
rect 18104 5516 18110 5528
rect 18417 5525 18429 5528
rect 18463 5525 18475 5559
rect 18417 5519 18475 5525
rect 18969 5559 19027 5565
rect 18969 5525 18981 5559
rect 19015 5525 19027 5559
rect 19720 5556 19748 5655
rect 20070 5652 20076 5664
rect 20128 5652 20134 5704
rect 20254 5692 20260 5704
rect 20215 5664 20260 5692
rect 20254 5652 20260 5664
rect 20312 5652 20318 5704
rect 20364 5701 20392 5732
rect 20349 5695 20407 5701
rect 20349 5661 20361 5695
rect 20395 5661 20407 5695
rect 20809 5695 20867 5701
rect 20809 5692 20821 5695
rect 20349 5655 20407 5661
rect 20456 5664 20821 5692
rect 20272 5624 20300 5652
rect 20456 5624 20484 5664
rect 20809 5661 20821 5664
rect 20855 5661 20867 5695
rect 20916 5692 20944 5859
rect 21082 5856 21088 5868
rect 21140 5856 21146 5908
rect 21634 5896 21640 5908
rect 21595 5868 21640 5896
rect 21634 5856 21640 5868
rect 21692 5896 21698 5908
rect 22370 5896 22376 5908
rect 21692 5868 22376 5896
rect 21692 5856 21698 5868
rect 22370 5856 22376 5868
rect 22428 5856 22434 5908
rect 23290 5856 23296 5908
rect 23348 5896 23354 5908
rect 24118 5896 24124 5908
rect 23348 5868 23980 5896
rect 24079 5868 24124 5896
rect 23348 5856 23354 5868
rect 20990 5788 20996 5840
rect 21048 5828 21054 5840
rect 22002 5828 22008 5840
rect 21048 5800 22008 5828
rect 21048 5788 21054 5800
rect 22002 5788 22008 5800
rect 22060 5788 22066 5840
rect 22649 5831 22707 5837
rect 22649 5797 22661 5831
rect 22695 5828 22707 5831
rect 23382 5828 23388 5840
rect 22695 5800 23388 5828
rect 22695 5797 22707 5800
rect 22649 5791 22707 5797
rect 23382 5788 23388 5800
rect 23440 5788 23446 5840
rect 23952 5828 23980 5868
rect 24118 5856 24124 5868
rect 24176 5856 24182 5908
rect 24394 5856 24400 5908
rect 24452 5896 24458 5908
rect 24581 5899 24639 5905
rect 24581 5896 24593 5899
rect 24452 5868 24593 5896
rect 24452 5856 24458 5868
rect 24581 5865 24593 5868
rect 24627 5865 24639 5899
rect 24581 5859 24639 5865
rect 24762 5828 24768 5840
rect 23952 5800 24768 5828
rect 24762 5788 24768 5800
rect 24820 5788 24826 5840
rect 24302 5760 24308 5772
rect 21468 5732 24308 5760
rect 21269 5695 21327 5701
rect 21269 5692 21281 5695
rect 20916 5664 21281 5692
rect 20809 5655 20867 5661
rect 21269 5661 21281 5664
rect 21315 5692 21327 5695
rect 21361 5695 21419 5701
rect 21361 5692 21373 5695
rect 21315 5664 21373 5692
rect 21315 5661 21327 5664
rect 21269 5655 21327 5661
rect 21361 5661 21373 5664
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 20272 5596 20484 5624
rect 20533 5627 20591 5633
rect 20533 5593 20545 5627
rect 20579 5624 20591 5627
rect 20622 5624 20628 5636
rect 20579 5596 20628 5624
rect 20579 5593 20591 5596
rect 20533 5587 20591 5593
rect 20622 5584 20628 5596
rect 20680 5624 20686 5636
rect 21468 5624 21496 5732
rect 24302 5720 24308 5732
rect 24360 5760 24366 5772
rect 25682 5760 25688 5772
rect 24360 5732 24532 5760
rect 24360 5720 24366 5732
rect 21821 5695 21879 5701
rect 21821 5661 21833 5695
rect 21867 5692 21879 5695
rect 22002 5692 22008 5704
rect 21867 5664 22008 5692
rect 21867 5661 21879 5664
rect 21821 5655 21879 5661
rect 22002 5652 22008 5664
rect 22060 5652 22066 5704
rect 22373 5695 22431 5701
rect 22373 5661 22385 5695
rect 22419 5661 22431 5695
rect 22646 5692 22652 5704
rect 22607 5664 22652 5692
rect 22373 5655 22431 5661
rect 20680 5596 21496 5624
rect 20680 5584 20686 5596
rect 20990 5556 20996 5568
rect 19720 5528 20996 5556
rect 18969 5519 19027 5525
rect 20990 5516 20996 5528
rect 21048 5516 21054 5568
rect 21450 5516 21456 5568
rect 21508 5556 21514 5568
rect 21545 5559 21603 5565
rect 21545 5556 21557 5559
rect 21508 5528 21557 5556
rect 21508 5516 21514 5528
rect 21545 5525 21557 5528
rect 21591 5556 21603 5559
rect 22002 5556 22008 5568
rect 21591 5528 22008 5556
rect 21591 5525 21603 5528
rect 21545 5519 21603 5525
rect 22002 5516 22008 5528
rect 22060 5556 22066 5568
rect 22388 5556 22416 5655
rect 22646 5652 22652 5664
rect 22704 5692 22710 5704
rect 23937 5695 23995 5701
rect 23937 5692 23949 5695
rect 22704 5664 23949 5692
rect 22704 5652 22710 5664
rect 23937 5661 23949 5664
rect 23983 5661 23995 5695
rect 23937 5655 23995 5661
rect 24118 5652 24124 5704
rect 24176 5692 24182 5704
rect 24394 5692 24400 5704
rect 24176 5664 24221 5692
rect 24355 5664 24400 5692
rect 24176 5652 24182 5664
rect 24394 5652 24400 5664
rect 24452 5652 24458 5704
rect 24504 5624 24532 5732
rect 25240 5732 25688 5760
rect 25240 5624 25268 5732
rect 25682 5720 25688 5732
rect 25740 5720 25746 5772
rect 25317 5695 25375 5701
rect 25317 5661 25329 5695
rect 25363 5692 25375 5695
rect 25590 5692 25596 5704
rect 25363 5664 25596 5692
rect 25363 5661 25375 5664
rect 25317 5655 25375 5661
rect 25590 5652 25596 5664
rect 25648 5652 25654 5704
rect 25501 5627 25559 5633
rect 25501 5624 25513 5627
rect 24504 5596 25513 5624
rect 25501 5593 25513 5596
rect 25547 5593 25559 5627
rect 25501 5587 25559 5593
rect 25685 5627 25743 5633
rect 25685 5593 25697 5627
rect 25731 5624 25743 5627
rect 26418 5624 26424 5636
rect 25731 5596 26424 5624
rect 25731 5593 25743 5596
rect 25685 5587 25743 5593
rect 26418 5584 26424 5596
rect 26476 5584 26482 5636
rect 23750 5556 23756 5568
rect 22060 5528 22416 5556
rect 23711 5528 23756 5556
rect 22060 5516 22066 5528
rect 23750 5516 23756 5528
rect 23808 5516 23814 5568
rect 1104 5466 29440 5488
rect 1104 5414 10395 5466
rect 10447 5414 10459 5466
rect 10511 5414 10523 5466
rect 10575 5414 10587 5466
rect 10639 5414 10651 5466
rect 10703 5414 19840 5466
rect 19892 5414 19904 5466
rect 19956 5414 19968 5466
rect 20020 5414 20032 5466
rect 20084 5414 20096 5466
rect 20148 5414 29440 5466
rect 1104 5392 29440 5414
rect 2593 5355 2651 5361
rect 2593 5321 2605 5355
rect 2639 5352 2651 5355
rect 2682 5352 2688 5364
rect 2639 5324 2688 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 4246 5352 4252 5364
rect 4207 5324 4252 5352
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 4709 5355 4767 5361
rect 4709 5352 4721 5355
rect 4387 5324 4721 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 4709 5321 4721 5324
rect 4755 5321 4767 5355
rect 4709 5315 4767 5321
rect 7469 5355 7527 5361
rect 7469 5321 7481 5355
rect 7515 5352 7527 5355
rect 8021 5355 8079 5361
rect 8021 5352 8033 5355
rect 7515 5324 8033 5352
rect 7515 5321 7527 5324
rect 7469 5315 7527 5321
rect 8021 5321 8033 5324
rect 8067 5321 8079 5355
rect 11422 5352 11428 5364
rect 8021 5315 8079 5321
rect 11164 5324 11428 5352
rect 5810 5284 5816 5296
rect 5771 5256 5816 5284
rect 5810 5244 5816 5256
rect 5868 5244 5874 5296
rect 5997 5287 6055 5293
rect 5997 5253 6009 5287
rect 6043 5284 6055 5287
rect 6086 5284 6092 5296
rect 6043 5256 6092 5284
rect 6043 5253 6055 5256
rect 5997 5247 6055 5253
rect 6086 5244 6092 5256
rect 6144 5244 6150 5296
rect 6181 5287 6239 5293
rect 6181 5253 6193 5287
rect 6227 5284 6239 5287
rect 6270 5284 6276 5296
rect 6227 5256 6276 5284
rect 6227 5253 6239 5256
rect 6181 5247 6239 5253
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 11164 5284 11192 5324
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 11698 5352 11704 5364
rect 11659 5324 11704 5352
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 12805 5355 12863 5361
rect 12805 5321 12817 5355
rect 12851 5352 12863 5355
rect 12894 5352 12900 5364
rect 12851 5324 12900 5352
rect 12851 5321 12863 5324
rect 12805 5315 12863 5321
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 13265 5355 13323 5361
rect 13265 5352 13277 5355
rect 13228 5324 13277 5352
rect 13228 5312 13234 5324
rect 13265 5321 13277 5324
rect 13311 5321 13323 5355
rect 13265 5315 13323 5321
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 15252 5324 15301 5352
rect 15252 5312 15258 5324
rect 15289 5321 15301 5324
rect 15335 5352 15347 5355
rect 17313 5355 17371 5361
rect 15335 5324 16804 5352
rect 15335 5321 15347 5324
rect 15289 5315 15347 5321
rect 6748 5256 11192 5284
rect 11241 5287 11299 5293
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5216 2835 5219
rect 3142 5216 3148 5228
rect 2823 5188 3148 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 4890 5216 4896 5228
rect 4851 5188 4896 5216
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 6638 5216 6644 5228
rect 6599 5188 6644 5216
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4525 5151 4583 5157
rect 4525 5148 4537 5151
rect 4120 5120 4537 5148
rect 4120 5108 4126 5120
rect 4525 5117 4537 5120
rect 4571 5148 4583 5151
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 4571 5120 4997 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 4985 5117 4997 5120
rect 5031 5117 5043 5151
rect 4985 5111 5043 5117
rect 3970 5040 3976 5092
rect 4028 5080 4034 5092
rect 6748 5080 6776 5256
rect 11241 5253 11253 5287
rect 11287 5284 11299 5287
rect 12618 5284 12624 5296
rect 11287 5256 12204 5284
rect 12579 5256 12624 5284
rect 11287 5253 11299 5256
rect 11241 5247 11299 5253
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 7006 5216 7012 5228
rect 6871 5188 7012 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 7006 5176 7012 5188
rect 7064 5216 7070 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 7064 5188 7573 5216
rect 7064 5176 7070 5188
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 8205 5219 8263 5225
rect 8205 5216 8217 5219
rect 7561 5179 7619 5185
rect 7668 5188 8217 5216
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 7285 5151 7343 5157
rect 7285 5148 7297 5151
rect 7156 5120 7297 5148
rect 7156 5108 7162 5120
rect 7285 5117 7297 5120
rect 7331 5117 7343 5151
rect 7285 5111 7343 5117
rect 4028 5052 6776 5080
rect 7009 5083 7067 5089
rect 4028 5040 4034 5052
rect 7009 5049 7021 5083
rect 7055 5080 7067 5083
rect 7668 5080 7696 5188
rect 8205 5185 8217 5188
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5216 9183 5219
rect 9677 5219 9735 5225
rect 9171 5188 9536 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 8757 5151 8815 5157
rect 8757 5117 8769 5151
rect 8803 5148 8815 5151
rect 9214 5148 9220 5160
rect 8803 5120 9220 5148
rect 8803 5117 8815 5120
rect 8757 5111 8815 5117
rect 9214 5108 9220 5120
rect 9272 5148 9278 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 9272 5120 9321 5148
rect 9272 5108 9278 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 9508 5092 9536 5188
rect 9677 5185 9689 5219
rect 9723 5216 9735 5219
rect 10594 5216 10600 5228
rect 9723 5188 10600 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 10594 5176 10600 5188
rect 10652 5176 10658 5228
rect 10870 5216 10876 5228
rect 10831 5188 10876 5216
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11054 5216 11060 5228
rect 11015 5188 11060 5216
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 11204 5188 11249 5216
rect 11204 5176 11210 5188
rect 11422 5176 11428 5228
rect 11480 5216 11486 5228
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11480 5188 11713 5216
rect 11480 5176 11486 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 12066 5216 12072 5228
rect 12027 5188 12072 5216
rect 11701 5179 11759 5185
rect 12066 5176 12072 5188
rect 12124 5176 12130 5228
rect 12176 5225 12204 5256
rect 12618 5244 12624 5256
rect 12676 5244 12682 5296
rect 13814 5284 13820 5296
rect 13775 5256 13820 5284
rect 13814 5244 13820 5256
rect 13872 5244 13878 5296
rect 14366 5244 14372 5296
rect 14424 5284 14430 5296
rect 16776 5293 16804 5324
rect 17313 5321 17325 5355
rect 17359 5321 17371 5355
rect 17313 5315 17371 5321
rect 16761 5287 16819 5293
rect 14424 5256 15516 5284
rect 14424 5244 14430 5256
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5185 12219 5219
rect 12161 5179 12219 5185
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5185 12403 5219
rect 12710 5216 12716 5228
rect 12671 5188 12716 5216
rect 12345 5179 12403 5185
rect 10686 5148 10692 5160
rect 10599 5120 10692 5148
rect 10686 5108 10692 5120
rect 10744 5148 10750 5160
rect 11514 5148 11520 5160
rect 10744 5120 11520 5148
rect 10744 5108 10750 5120
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 12084 5148 12112 5176
rect 12360 5148 12388 5179
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5216 13231 5219
rect 13262 5216 13268 5228
rect 13219 5188 13268 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 14059 5219 14117 5225
rect 14059 5185 14071 5219
rect 14105 5216 14117 5219
rect 14550 5216 14556 5228
rect 14105 5188 14556 5216
rect 14105 5185 14117 5188
rect 14059 5179 14117 5185
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5185 14887 5219
rect 15010 5216 15016 5228
rect 14971 5188 15016 5216
rect 14829 5179 14887 5185
rect 12084 5120 12388 5148
rect 13449 5151 13507 5157
rect 13449 5117 13461 5151
rect 13495 5148 13507 5151
rect 13814 5148 13820 5160
rect 13495 5120 13820 5148
rect 13495 5117 13507 5120
rect 13449 5111 13507 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14366 5148 14372 5160
rect 14327 5120 14372 5148
rect 14366 5108 14372 5120
rect 14424 5108 14430 5160
rect 14458 5108 14464 5160
rect 14516 5148 14522 5160
rect 14516 5120 14561 5148
rect 14516 5108 14522 5120
rect 7055 5052 7696 5080
rect 7929 5083 7987 5089
rect 7055 5049 7067 5052
rect 7009 5043 7067 5049
rect 7929 5049 7941 5083
rect 7975 5080 7987 5083
rect 8294 5080 8300 5092
rect 7975 5052 8300 5080
rect 7975 5049 7987 5052
rect 7929 5043 7987 5049
rect 8294 5040 8300 5052
rect 8352 5040 8358 5092
rect 9490 5080 9496 5092
rect 9403 5052 9496 5080
rect 9490 5040 9496 5052
rect 9548 5040 9554 5092
rect 13538 5040 13544 5092
rect 13596 5080 13602 5092
rect 14844 5080 14872 5179
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 15286 5216 15292 5228
rect 15247 5188 15292 5216
rect 15286 5176 15292 5188
rect 15344 5176 15350 5228
rect 15488 5225 15516 5256
rect 16761 5253 16773 5287
rect 16807 5284 16819 5287
rect 17328 5284 17356 5315
rect 17678 5312 17684 5364
rect 17736 5352 17742 5364
rect 17957 5355 18015 5361
rect 17957 5352 17969 5355
rect 17736 5324 17969 5352
rect 17736 5312 17742 5324
rect 17957 5321 17969 5324
rect 18003 5321 18015 5355
rect 17957 5315 18015 5321
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 19702 5352 19708 5364
rect 19659 5324 19708 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 19981 5355 20039 5361
rect 19981 5321 19993 5355
rect 20027 5321 20039 5355
rect 20622 5352 20628 5364
rect 20583 5324 20628 5352
rect 19981 5315 20039 5321
rect 17586 5284 17592 5296
rect 16807 5256 17080 5284
rect 17328 5256 17592 5284
rect 16807 5253 16819 5256
rect 16761 5247 16819 5253
rect 17052 5225 17080 5256
rect 17586 5244 17592 5256
rect 17644 5284 17650 5296
rect 17644 5256 17724 5284
rect 17644 5244 17650 5256
rect 15473 5219 15531 5225
rect 15473 5185 15485 5219
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5185 17095 5219
rect 17696 5216 17724 5256
rect 17770 5244 17776 5296
rect 17828 5284 17834 5296
rect 17865 5287 17923 5293
rect 17865 5284 17877 5287
rect 17828 5256 17877 5284
rect 17828 5244 17834 5256
rect 17865 5253 17877 5256
rect 17911 5284 17923 5287
rect 18417 5287 18475 5293
rect 18417 5284 18429 5287
rect 17911 5256 18429 5284
rect 17911 5253 17923 5256
rect 17865 5247 17923 5253
rect 18417 5253 18429 5256
rect 18463 5253 18475 5287
rect 18417 5247 18475 5253
rect 19518 5244 19524 5296
rect 19576 5284 19582 5296
rect 19996 5284 20024 5315
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 24029 5355 24087 5361
rect 22066 5324 23888 5352
rect 22066 5284 22094 5324
rect 19576 5256 20024 5284
rect 20088 5256 22094 5284
rect 19576 5244 19582 5256
rect 18325 5219 18383 5225
rect 18325 5216 18337 5219
rect 17696 5188 18337 5216
rect 17037 5179 17095 5185
rect 18325 5185 18337 5188
rect 18371 5185 18383 5219
rect 18325 5179 18383 5185
rect 19702 5176 19708 5228
rect 19760 5216 19766 5228
rect 20088 5225 20116 5256
rect 22278 5244 22284 5296
rect 22336 5284 22342 5296
rect 23109 5287 23167 5293
rect 23109 5284 23121 5287
rect 22336 5256 23121 5284
rect 22336 5244 22342 5256
rect 23109 5253 23121 5256
rect 23155 5253 23167 5287
rect 23109 5247 23167 5253
rect 20073 5219 20131 5225
rect 20073 5216 20085 5219
rect 19760 5188 20085 5216
rect 19760 5176 19766 5188
rect 20073 5185 20085 5188
rect 20119 5185 20131 5219
rect 20806 5216 20812 5228
rect 20767 5188 20812 5216
rect 20073 5179 20131 5185
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 21910 5216 21916 5228
rect 21871 5188 21916 5216
rect 21910 5176 21916 5188
rect 21968 5176 21974 5228
rect 22094 5176 22100 5228
rect 22152 5216 22158 5228
rect 22370 5216 22376 5228
rect 22152 5188 22197 5216
rect 22283 5188 22376 5216
rect 22152 5176 22158 5188
rect 22370 5176 22376 5188
rect 22428 5176 22434 5228
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5216 22615 5219
rect 22603 5188 22784 5216
rect 22603 5185 22615 5188
rect 22557 5179 22615 5185
rect 15838 5108 15844 5160
rect 15896 5148 15902 5160
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 15896 5120 16681 5148
rect 15896 5108 15902 5120
rect 16669 5117 16681 5120
rect 16715 5117 16727 5151
rect 17149 5151 17207 5157
rect 17149 5148 17161 5151
rect 16669 5111 16727 5117
rect 16868 5120 17161 5148
rect 13596 5052 14872 5080
rect 16684 5080 16712 5111
rect 16868 5080 16896 5120
rect 17149 5117 17161 5120
rect 17195 5117 17207 5151
rect 18046 5148 18052 5160
rect 18007 5120 18052 5148
rect 17149 5111 17207 5117
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 18969 5151 19027 5157
rect 18969 5148 18981 5151
rect 18340 5120 18981 5148
rect 18340 5080 18368 5120
rect 18969 5117 18981 5120
rect 19015 5148 19027 5151
rect 19061 5151 19119 5157
rect 19061 5148 19073 5151
rect 19015 5120 19073 5148
rect 19015 5117 19027 5120
rect 18969 5111 19027 5117
rect 19061 5117 19073 5120
rect 19107 5117 19119 5151
rect 19061 5111 19119 5117
rect 19242 5108 19248 5160
rect 19300 5148 19306 5160
rect 19337 5151 19395 5157
rect 19337 5148 19349 5151
rect 19300 5120 19349 5148
rect 19300 5108 19306 5120
rect 19337 5117 19349 5120
rect 19383 5117 19395 5151
rect 19337 5111 19395 5117
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 19521 5151 19579 5157
rect 19521 5148 19533 5151
rect 19484 5120 19533 5148
rect 19484 5108 19490 5120
rect 19521 5117 19533 5120
rect 19567 5148 19579 5151
rect 20165 5151 20223 5157
rect 20165 5148 20177 5151
rect 19567 5120 20177 5148
rect 19567 5117 19579 5120
rect 19521 5111 19579 5117
rect 20165 5117 20177 5120
rect 20211 5117 20223 5151
rect 20165 5111 20223 5117
rect 21358 5108 21364 5160
rect 21416 5148 21422 5160
rect 22189 5151 22247 5157
rect 22189 5148 22201 5151
rect 21416 5120 22201 5148
rect 21416 5108 21422 5120
rect 22189 5117 22201 5120
rect 22235 5117 22247 5151
rect 22189 5111 22247 5117
rect 16684 5052 16896 5080
rect 17328 5052 18368 5080
rect 13596 5040 13602 5052
rect 3878 5012 3884 5024
rect 3839 4984 3884 5012
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 8754 4972 8760 5024
rect 8812 5012 8818 5024
rect 8941 5015 8999 5021
rect 8941 5012 8953 5015
rect 8812 4984 8953 5012
rect 8812 4972 8818 4984
rect 8941 4981 8953 4984
rect 8987 4981 8999 5015
rect 8941 4975 8999 4981
rect 13354 4972 13360 5024
rect 13412 5012 13418 5024
rect 17328 5012 17356 5052
rect 18414 5040 18420 5092
rect 18472 5080 18478 5092
rect 21450 5080 21456 5092
rect 18472 5052 21456 5080
rect 18472 5040 18478 5052
rect 21450 5040 21456 5052
rect 21508 5040 21514 5092
rect 13412 4984 17356 5012
rect 13412 4972 13418 4984
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 17460 4984 17509 5012
rect 17460 4972 17466 4984
rect 17497 4981 17509 4984
rect 17543 4981 17555 5015
rect 17497 4975 17555 4981
rect 18969 5015 19027 5021
rect 18969 4981 18981 5015
rect 19015 5012 19027 5015
rect 20254 5012 20260 5024
rect 19015 4984 20260 5012
rect 19015 4981 19027 4984
rect 18969 4975 19027 4981
rect 20254 4972 20260 4984
rect 20312 5012 20318 5024
rect 20901 5015 20959 5021
rect 20901 5012 20913 5015
rect 20312 4984 20913 5012
rect 20312 4972 20318 4984
rect 20901 4981 20913 4984
rect 20947 4981 20959 5015
rect 22388 5012 22416 5176
rect 22756 5089 22784 5188
rect 23382 5176 23388 5228
rect 23440 5216 23446 5228
rect 23569 5219 23627 5225
rect 23569 5216 23581 5219
rect 23440 5188 23581 5216
rect 23440 5176 23446 5188
rect 23569 5185 23581 5188
rect 23615 5185 23627 5219
rect 23750 5216 23756 5228
rect 23711 5188 23756 5216
rect 23569 5179 23627 5185
rect 23750 5176 23756 5188
rect 23808 5176 23814 5228
rect 23860 5225 23888 5324
rect 24029 5321 24041 5355
rect 24075 5352 24087 5355
rect 24394 5352 24400 5364
rect 24075 5324 24400 5352
rect 24075 5321 24087 5324
rect 24029 5315 24087 5321
rect 24394 5312 24400 5324
rect 24452 5312 24458 5364
rect 25409 5355 25467 5361
rect 25409 5321 25421 5355
rect 25455 5321 25467 5355
rect 25409 5315 25467 5321
rect 25869 5355 25927 5361
rect 25869 5321 25881 5355
rect 25915 5352 25927 5355
rect 26237 5355 26295 5361
rect 26237 5352 26249 5355
rect 25915 5324 26249 5352
rect 25915 5321 25927 5324
rect 25869 5315 25927 5321
rect 26237 5321 26249 5324
rect 26283 5321 26295 5355
rect 26237 5315 26295 5321
rect 24118 5244 24124 5296
rect 24176 5284 24182 5296
rect 24305 5287 24363 5293
rect 24305 5284 24317 5287
rect 24176 5256 24317 5284
rect 24176 5244 24182 5256
rect 24305 5253 24317 5256
rect 24351 5253 24363 5287
rect 24305 5247 24363 5253
rect 24596 5256 24992 5284
rect 24596 5225 24624 5256
rect 23845 5219 23903 5225
rect 23845 5185 23857 5219
rect 23891 5185 23903 5219
rect 23845 5179 23903 5185
rect 24397 5219 24455 5225
rect 24397 5185 24409 5219
rect 24443 5216 24455 5219
rect 24581 5219 24639 5225
rect 24581 5216 24593 5219
rect 24443 5188 24593 5216
rect 24443 5185 24455 5188
rect 24397 5179 24455 5185
rect 24581 5185 24593 5188
rect 24627 5185 24639 5219
rect 24762 5216 24768 5228
rect 24723 5188 24768 5216
rect 24581 5179 24639 5185
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 22830 5108 22836 5160
rect 22888 5148 22894 5160
rect 23201 5151 23259 5157
rect 23201 5148 23213 5151
rect 22888 5120 23213 5148
rect 22888 5108 22894 5120
rect 23201 5117 23213 5120
rect 23247 5117 23259 5151
rect 23201 5111 23259 5117
rect 23293 5151 23351 5157
rect 23293 5117 23305 5151
rect 23339 5148 23351 5151
rect 24857 5151 24915 5157
rect 24857 5148 24869 5151
rect 23339 5120 23704 5148
rect 23339 5117 23351 5120
rect 23293 5111 23351 5117
rect 22741 5083 22799 5089
rect 22741 5049 22753 5083
rect 22787 5049 22799 5083
rect 22741 5043 22799 5049
rect 23014 5040 23020 5092
rect 23072 5080 23078 5092
rect 23308 5080 23336 5111
rect 23072 5052 23336 5080
rect 23072 5040 23078 5052
rect 22922 5012 22928 5024
rect 22388 4984 22928 5012
rect 20901 4975 20959 4981
rect 22922 4972 22928 4984
rect 22980 4972 22986 5024
rect 23566 5012 23572 5024
rect 23527 4984 23572 5012
rect 23566 4972 23572 4984
rect 23624 4972 23630 5024
rect 23676 5012 23704 5120
rect 24504 5120 24869 5148
rect 24504 5092 24532 5120
rect 24857 5117 24869 5120
rect 24903 5117 24915 5151
rect 24964 5148 24992 5256
rect 25038 5176 25044 5228
rect 25096 5216 25102 5228
rect 25225 5219 25283 5225
rect 25096 5188 25141 5216
rect 25096 5176 25102 5188
rect 25225 5185 25237 5219
rect 25271 5216 25283 5219
rect 25424 5216 25452 5315
rect 27246 5312 27252 5364
rect 27304 5352 27310 5364
rect 27525 5355 27583 5361
rect 27525 5352 27537 5355
rect 27304 5324 27537 5352
rect 27304 5312 27310 5324
rect 27525 5321 27537 5324
rect 27571 5321 27583 5355
rect 27525 5315 27583 5321
rect 27893 5287 27951 5293
rect 27893 5284 27905 5287
rect 27448 5256 27905 5284
rect 27448 5228 27476 5256
rect 27893 5253 27905 5256
rect 27939 5253 27951 5287
rect 27893 5247 27951 5253
rect 25271 5188 25452 5216
rect 25271 5185 25283 5188
rect 25225 5179 25283 5185
rect 25590 5176 25596 5228
rect 25648 5216 25654 5228
rect 25777 5219 25835 5225
rect 25777 5216 25789 5219
rect 25648 5188 25789 5216
rect 25648 5176 25654 5188
rect 25777 5185 25789 5188
rect 25823 5185 25835 5219
rect 26418 5216 26424 5228
rect 26379 5188 26424 5216
rect 25777 5179 25835 5185
rect 26418 5176 26424 5188
rect 26476 5176 26482 5228
rect 27430 5225 27436 5228
rect 27157 5219 27215 5225
rect 27157 5185 27169 5219
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27413 5219 27436 5225
rect 27413 5185 27425 5219
rect 27413 5179 27436 5185
rect 25608 5148 25636 5176
rect 24964 5120 25636 5148
rect 25961 5151 26019 5157
rect 24857 5111 24915 5117
rect 25961 5117 25973 5151
rect 26007 5117 26019 5151
rect 27172 5148 27200 5179
rect 27430 5176 27436 5179
rect 27488 5176 27494 5228
rect 27706 5216 27712 5228
rect 27667 5188 27712 5216
rect 27706 5176 27712 5188
rect 27764 5216 27770 5228
rect 27801 5219 27859 5225
rect 27801 5216 27813 5219
rect 27764 5188 27813 5216
rect 27764 5176 27770 5188
rect 27801 5185 27813 5188
rect 27847 5185 27859 5219
rect 27801 5179 27859 5185
rect 27522 5148 27528 5160
rect 27172 5120 27528 5148
rect 25961 5111 26019 5117
rect 24486 5040 24492 5092
rect 24544 5040 24550 5092
rect 25976 5012 26004 5111
rect 27522 5108 27528 5120
rect 27580 5108 27586 5160
rect 27617 5151 27675 5157
rect 27617 5117 27629 5151
rect 27663 5117 27675 5151
rect 27617 5111 27675 5117
rect 27338 5040 27344 5092
rect 27396 5080 27402 5092
rect 27632 5080 27660 5111
rect 27396 5052 27660 5080
rect 27396 5040 27402 5052
rect 23676 4984 26004 5012
rect 26878 4972 26884 5024
rect 26936 5012 26942 5024
rect 26973 5015 27031 5021
rect 26973 5012 26985 5015
rect 26936 4984 26985 5012
rect 26936 4972 26942 4984
rect 26973 4981 26985 4984
rect 27019 4981 27031 5015
rect 26973 4975 27031 4981
rect 1104 4922 29440 4944
rect 1104 4870 5672 4922
rect 5724 4870 5736 4922
rect 5788 4870 5800 4922
rect 5852 4870 5864 4922
rect 5916 4870 5928 4922
rect 5980 4870 15118 4922
rect 15170 4870 15182 4922
rect 15234 4870 15246 4922
rect 15298 4870 15310 4922
rect 15362 4870 15374 4922
rect 15426 4870 24563 4922
rect 24615 4870 24627 4922
rect 24679 4870 24691 4922
rect 24743 4870 24755 4922
rect 24807 4870 24819 4922
rect 24871 4870 29440 4922
rect 1104 4848 29440 4870
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 4856 4780 5181 4808
rect 4856 4768 4862 4780
rect 5169 4777 5181 4780
rect 5215 4777 5227 4811
rect 10594 4808 10600 4820
rect 10555 4780 10600 4808
rect 5169 4771 5227 4777
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 11241 4811 11299 4817
rect 11241 4777 11253 4811
rect 11287 4777 11299 4811
rect 11241 4771 11299 4777
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 12986 4808 12992 4820
rect 12943 4780 12992 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 10321 4743 10379 4749
rect 10321 4709 10333 4743
rect 10367 4740 10379 4743
rect 10870 4740 10876 4752
rect 10367 4712 10876 4740
rect 10367 4709 10379 4712
rect 10321 4703 10379 4709
rect 10870 4700 10876 4712
rect 10928 4740 10934 4752
rect 11256 4740 11284 4771
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 15381 4811 15439 4817
rect 15381 4777 15393 4811
rect 15427 4808 15439 4811
rect 15470 4808 15476 4820
rect 15427 4780 15476 4808
rect 15427 4777 15439 4780
rect 15381 4771 15439 4777
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 15838 4808 15844 4820
rect 15799 4780 15844 4808
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 21821 4811 21879 4817
rect 15948 4780 21496 4808
rect 14550 4740 14556 4752
rect 10928 4712 11284 4740
rect 12268 4712 14320 4740
rect 14511 4712 14556 4740
rect 10928 4700 10934 4712
rect 1486 4632 1492 4684
rect 1544 4672 1550 4684
rect 1544 4644 2774 4672
rect 1544 4632 1550 4644
rect 1578 4604 1584 4616
rect 1412 4576 1584 4604
rect 1412 4480 1440 4576
rect 1578 4564 1584 4576
rect 1636 4604 1642 4616
rect 1857 4607 1915 4613
rect 1857 4604 1869 4607
rect 1636 4576 1869 4604
rect 1636 4564 1642 4576
rect 1857 4573 1869 4576
rect 1903 4573 1915 4607
rect 2746 4604 2774 4644
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 11072 4681 11100 4712
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 8536 4644 8953 4672
rect 8536 4632 8542 4644
rect 8941 4641 8953 4644
rect 8987 4641 8999 4675
rect 8941 4635 8999 4641
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4641 11115 4675
rect 11330 4672 11336 4684
rect 11291 4644 11336 4672
rect 11057 4635 11115 4641
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 3786 4604 3792 4616
rect 2746 4576 3792 4604
rect 1857 4567 1915 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 4045 4607 4103 4613
rect 4045 4604 4057 4607
rect 3936 4576 4057 4604
rect 3936 4564 3942 4576
rect 4045 4573 4057 4576
rect 4091 4573 4103 4607
rect 5994 4604 6000 4616
rect 5955 4576 6000 4604
rect 4045 4567 4103 4573
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 8754 4604 8760 4616
rect 8619 4576 8760 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 11149 4607 11207 4613
rect 11149 4604 11161 4607
rect 10744 4576 10789 4604
rect 11072 4576 11161 4604
rect 10744 4564 10750 4576
rect 11072 4548 11100 4576
rect 11149 4573 11161 4576
rect 11195 4573 11207 4607
rect 11149 4567 11207 4573
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 11517 4607 11575 4613
rect 11296 4576 11341 4604
rect 11296 4564 11302 4576
rect 11517 4573 11529 4607
rect 11563 4573 11575 4607
rect 11517 4567 11575 4573
rect 8938 4496 8944 4548
rect 8996 4536 9002 4548
rect 9186 4539 9244 4545
rect 9186 4536 9198 4539
rect 8996 4508 9198 4536
rect 8996 4496 9002 4508
rect 9186 4505 9198 4508
rect 9232 4505 9244 4539
rect 9186 4499 9244 4505
rect 11054 4496 11060 4548
rect 11112 4496 11118 4548
rect 11532 4536 11560 4567
rect 12268 4545 12296 4712
rect 12621 4675 12679 4681
rect 12621 4641 12633 4675
rect 12667 4672 12679 4675
rect 12710 4672 12716 4684
rect 12667 4644 12716 4672
rect 12667 4641 12679 4644
rect 12621 4635 12679 4641
rect 12710 4632 12716 4644
rect 12768 4672 12774 4684
rect 14292 4672 14320 4712
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 14734 4700 14740 4752
rect 14792 4740 14798 4752
rect 15948 4740 15976 4780
rect 14792 4712 15976 4740
rect 14792 4700 14798 4712
rect 19334 4700 19340 4752
rect 19392 4740 19398 4752
rect 21468 4740 21496 4780
rect 21821 4777 21833 4811
rect 21867 4808 21879 4811
rect 22462 4808 22468 4820
rect 21867 4780 22468 4808
rect 21867 4777 21879 4780
rect 21821 4771 21879 4777
rect 22462 4768 22468 4780
rect 22520 4768 22526 4820
rect 22830 4808 22836 4820
rect 22791 4780 22836 4808
rect 22830 4768 22836 4780
rect 22888 4768 22894 4820
rect 22922 4768 22928 4820
rect 22980 4808 22986 4820
rect 25038 4808 25044 4820
rect 22980 4780 25044 4808
rect 22980 4768 22986 4780
rect 25038 4768 25044 4780
rect 25096 4768 25102 4820
rect 25590 4808 25596 4820
rect 25551 4780 25596 4808
rect 25590 4768 25596 4780
rect 25648 4768 25654 4820
rect 25958 4768 25964 4820
rect 26016 4808 26022 4820
rect 26421 4811 26479 4817
rect 26421 4808 26433 4811
rect 26016 4780 26433 4808
rect 26016 4768 26022 4780
rect 26421 4777 26433 4780
rect 26467 4777 26479 4811
rect 26421 4771 26479 4777
rect 26234 4740 26240 4752
rect 19392 4712 19840 4740
rect 21468 4712 26240 4740
rect 19392 4700 19398 4712
rect 15010 4672 15016 4684
rect 12768 4644 14228 4672
rect 14292 4644 15016 4672
rect 12768 4632 12774 4644
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4604 13139 4607
rect 13170 4604 13176 4616
rect 13127 4576 13176 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 13265 4607 13323 4613
rect 13265 4573 13277 4607
rect 13311 4604 13323 4607
rect 13354 4604 13360 4616
rect 13311 4576 13360 4604
rect 13311 4573 13323 4576
rect 13265 4567 13323 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 14200 4613 14228 4644
rect 15010 4632 15016 4644
rect 15068 4672 15074 4684
rect 15197 4675 15255 4681
rect 15197 4672 15209 4675
rect 15068 4644 15209 4672
rect 15068 4632 15074 4644
rect 15197 4641 15209 4644
rect 15243 4641 15255 4675
rect 19702 4672 19708 4684
rect 19663 4644 19708 4672
rect 15197 4635 15255 4641
rect 19702 4632 19708 4644
rect 19760 4632 19766 4684
rect 19812 4681 19840 4712
rect 26234 4700 26240 4712
rect 26292 4700 26298 4752
rect 27338 4740 27344 4752
rect 26712 4712 27016 4740
rect 27299 4712 27344 4740
rect 19797 4675 19855 4681
rect 19797 4641 19809 4675
rect 19843 4672 19855 4675
rect 21545 4675 21603 4681
rect 21545 4672 21557 4675
rect 19843 4644 21557 4672
rect 19843 4641 19855 4644
rect 19797 4635 19855 4641
rect 21545 4641 21557 4644
rect 21591 4672 21603 4675
rect 22281 4675 22339 4681
rect 21591 4644 22232 4672
rect 21591 4641 21603 4644
rect 21545 4635 21603 4641
rect 14185 4607 14243 4613
rect 14185 4573 14197 4607
rect 14231 4604 14243 4607
rect 14458 4604 14464 4616
rect 14231 4576 14464 4604
rect 14231 4573 14243 4576
rect 14185 4567 14243 4573
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 14752 4576 15393 4604
rect 11164 4508 11560 4536
rect 12253 4539 12311 4545
rect 11164 4480 11192 4508
rect 12253 4505 12265 4539
rect 12299 4505 12311 4539
rect 12253 4499 12311 4505
rect 1394 4468 1400 4480
rect 1355 4440 1400 4468
rect 1394 4428 1400 4440
rect 1452 4428 1458 4480
rect 6181 4471 6239 4477
rect 6181 4437 6193 4471
rect 6227 4468 6239 4471
rect 6914 4468 6920 4480
rect 6227 4440 6920 4468
rect 6227 4437 6239 4440
rect 6181 4431 6239 4437
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 8757 4471 8815 4477
rect 7064 4440 7109 4468
rect 7064 4428 7070 4440
rect 8757 4437 8769 4471
rect 8803 4468 8815 4471
rect 9398 4468 9404 4480
rect 8803 4440 9404 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 11146 4428 11152 4480
rect 11204 4428 11210 4480
rect 11701 4471 11759 4477
rect 11701 4437 11713 4471
rect 11747 4468 11759 4471
rect 12268 4468 12296 4499
rect 12434 4496 12440 4548
rect 12492 4536 12498 4548
rect 14366 4536 14372 4548
rect 12492 4508 12585 4536
rect 14327 4508 14372 4536
rect 12492 4496 12498 4508
rect 14366 4496 14372 4508
rect 14424 4536 14430 4548
rect 14752 4536 14780 4576
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 15381 4567 15439 4573
rect 16666 4564 16672 4616
rect 16724 4604 16730 4616
rect 17126 4604 17132 4616
rect 16724 4576 17132 4604
rect 16724 4564 16730 4576
rect 17126 4564 17132 4576
rect 17184 4604 17190 4616
rect 17221 4607 17279 4613
rect 17221 4604 17233 4607
rect 17184 4576 17233 4604
rect 17184 4564 17190 4576
rect 17221 4573 17233 4576
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 17313 4607 17371 4613
rect 17313 4573 17325 4607
rect 17359 4604 17371 4607
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 17359 4576 17509 4604
rect 17359 4573 17371 4576
rect 17313 4567 17371 4573
rect 17497 4573 17509 4576
rect 17543 4573 17555 4607
rect 17770 4604 17776 4616
rect 17731 4576 17776 4604
rect 17497 4567 17555 4573
rect 17770 4564 17776 4576
rect 17828 4564 17834 4616
rect 19610 4604 19616 4616
rect 19571 4576 19616 4604
rect 19610 4564 19616 4576
rect 19668 4564 19674 4616
rect 21358 4604 21364 4616
rect 21319 4576 21364 4604
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 22002 4564 22008 4616
rect 22060 4604 22066 4616
rect 22097 4607 22155 4613
rect 22097 4604 22109 4607
rect 22060 4576 22109 4604
rect 22060 4564 22066 4576
rect 22097 4573 22109 4576
rect 22143 4573 22155 4607
rect 22204 4604 22232 4644
rect 22281 4641 22293 4675
rect 22327 4672 22339 4675
rect 23385 4675 23443 4681
rect 22327 4644 22692 4672
rect 22327 4641 22339 4644
rect 22281 4635 22339 4641
rect 22370 4604 22376 4616
rect 22204 4576 22376 4604
rect 22097 4567 22155 4573
rect 22370 4564 22376 4576
rect 22428 4564 22434 4616
rect 22664 4613 22692 4644
rect 23385 4641 23397 4675
rect 23431 4641 23443 4675
rect 23566 4672 23572 4684
rect 23527 4644 23572 4672
rect 23385 4635 23443 4641
rect 22557 4607 22615 4613
rect 22557 4604 22569 4607
rect 22480 4576 22569 4604
rect 14424 4508 14780 4536
rect 15105 4539 15163 4545
rect 14424 4496 14430 4508
rect 15105 4505 15117 4539
rect 15151 4536 15163 4539
rect 15470 4536 15476 4548
rect 15151 4508 15476 4536
rect 15151 4505 15163 4508
rect 15105 4499 15163 4505
rect 15470 4496 15476 4508
rect 15528 4496 15534 4548
rect 16976 4539 17034 4545
rect 16976 4505 16988 4539
rect 17022 4536 17034 4539
rect 17402 4536 17408 4548
rect 17022 4508 17408 4536
rect 17022 4505 17034 4508
rect 16976 4499 17034 4505
rect 17402 4496 17408 4508
rect 17460 4496 17466 4548
rect 21910 4536 21916 4548
rect 21823 4508 21916 4536
rect 21910 4496 21916 4508
rect 21968 4536 21974 4548
rect 22278 4536 22284 4548
rect 21968 4508 22284 4536
rect 21968 4496 21974 4508
rect 22278 4496 22284 4508
rect 22336 4536 22342 4548
rect 22480 4536 22508 4576
rect 22557 4573 22569 4576
rect 22603 4573 22615 4607
rect 22557 4567 22615 4573
rect 22649 4607 22707 4613
rect 22649 4573 22661 4607
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 22336 4508 22508 4536
rect 23400 4536 23428 4635
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 24394 4672 24400 4684
rect 23768 4644 24400 4672
rect 23474 4564 23480 4616
rect 23532 4604 23538 4616
rect 23661 4607 23719 4613
rect 23661 4604 23673 4607
rect 23532 4576 23673 4604
rect 23532 4564 23538 4576
rect 23661 4573 23673 4576
rect 23707 4573 23719 4607
rect 23661 4567 23719 4573
rect 23768 4536 23796 4644
rect 24394 4632 24400 4644
rect 24452 4672 24458 4684
rect 24489 4675 24547 4681
rect 24489 4672 24501 4675
rect 24452 4644 24501 4672
rect 24452 4632 24458 4644
rect 24489 4641 24501 4644
rect 24535 4641 24547 4675
rect 24489 4635 24547 4641
rect 25866 4632 25872 4684
rect 25924 4672 25930 4684
rect 26145 4675 26203 4681
rect 26145 4672 26157 4675
rect 25924 4644 26157 4672
rect 25924 4632 25930 4644
rect 26145 4641 26157 4644
rect 26191 4672 26203 4675
rect 26712 4672 26740 4712
rect 26878 4672 26884 4684
rect 26191 4644 26740 4672
rect 26839 4644 26884 4672
rect 26191 4641 26203 4644
rect 26145 4635 26203 4641
rect 26878 4632 26884 4644
rect 26936 4632 26942 4684
rect 26988 4681 27016 4712
rect 27338 4700 27344 4712
rect 27396 4700 27402 4752
rect 26973 4675 27031 4681
rect 26973 4641 26985 4675
rect 27019 4641 27031 4675
rect 27430 4672 27436 4684
rect 26973 4635 27031 4641
rect 27172 4644 27436 4672
rect 24118 4564 24124 4616
rect 24176 4604 24182 4616
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 24176 4576 24685 4604
rect 24176 4564 24182 4576
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 26789 4607 26847 4613
rect 26789 4573 26801 4607
rect 26835 4604 26847 4607
rect 27172 4604 27200 4644
rect 27430 4632 27436 4644
rect 27488 4632 27494 4684
rect 26835 4576 27200 4604
rect 26835 4573 26847 4576
rect 26789 4567 26847 4573
rect 27246 4564 27252 4616
rect 27304 4604 27310 4616
rect 27522 4604 27528 4616
rect 27304 4576 27349 4604
rect 27483 4576 27528 4604
rect 27304 4564 27310 4576
rect 27522 4564 27528 4576
rect 27580 4564 27586 4616
rect 23400 4508 23796 4536
rect 22336 4496 22342 4508
rect 11747 4440 12296 4468
rect 12457 4468 12485 4496
rect 23492 4480 23520 4508
rect 24486 4496 24492 4548
rect 24544 4536 24550 4548
rect 24765 4539 24823 4545
rect 24765 4536 24777 4539
rect 24544 4508 24777 4536
rect 24544 4496 24550 4508
rect 24765 4505 24777 4508
rect 24811 4505 24823 4539
rect 24765 4499 24823 4505
rect 26053 4539 26111 4545
rect 26053 4505 26065 4539
rect 26099 4536 26111 4539
rect 27709 4539 27767 4545
rect 27709 4536 27721 4539
rect 26099 4508 27721 4536
rect 26099 4505 26111 4508
rect 26053 4499 26111 4505
rect 27709 4505 27721 4508
rect 27755 4505 27767 4539
rect 27709 4499 27767 4505
rect 13262 4468 13268 4480
rect 12457 4440 13268 4468
rect 11747 4437 11759 4440
rect 11701 4431 11759 4437
rect 13262 4428 13268 4440
rect 13320 4468 13326 4480
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 13320 4440 13369 4468
rect 13320 4428 13326 4440
rect 13357 4437 13369 4440
rect 13403 4437 13415 4471
rect 13357 4431 13415 4437
rect 15565 4471 15623 4477
rect 15565 4437 15577 4471
rect 15611 4468 15623 4471
rect 17313 4471 17371 4477
rect 17313 4468 17325 4471
rect 15611 4440 17325 4468
rect 15611 4437 15623 4440
rect 15565 4431 15623 4437
rect 17313 4437 17325 4440
rect 17359 4437 17371 4471
rect 17313 4431 17371 4437
rect 17681 4471 17739 4477
rect 17681 4437 17693 4471
rect 17727 4468 17739 4471
rect 17954 4468 17960 4480
rect 17727 4440 17960 4468
rect 17727 4437 17739 4440
rect 17681 4431 17739 4437
rect 17954 4428 17960 4440
rect 18012 4468 18018 4480
rect 19058 4468 19064 4480
rect 18012 4440 19064 4468
rect 18012 4428 18018 4440
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 19245 4471 19303 4477
rect 19245 4437 19257 4471
rect 19291 4468 19303 4471
rect 19518 4468 19524 4480
rect 19291 4440 19524 4468
rect 19291 4437 19303 4440
rect 19245 4431 19303 4437
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 20990 4468 20996 4480
rect 20951 4440 20996 4468
rect 20990 4428 20996 4440
rect 21048 4428 21054 4480
rect 21453 4471 21511 4477
rect 21453 4437 21465 4471
rect 21499 4468 21511 4471
rect 21821 4471 21879 4477
rect 21821 4468 21833 4471
rect 21499 4440 21833 4468
rect 21499 4437 21511 4440
rect 21453 4431 21511 4437
rect 21821 4437 21833 4440
rect 21867 4437 21879 4471
rect 22462 4468 22468 4480
rect 22375 4440 22468 4468
rect 21821 4431 21879 4437
rect 22462 4428 22468 4440
rect 22520 4468 22526 4480
rect 23382 4468 23388 4480
rect 22520 4440 23388 4468
rect 22520 4428 22526 4440
rect 23382 4428 23388 4440
rect 23440 4428 23446 4480
rect 23474 4428 23480 4480
rect 23532 4428 23538 4480
rect 24029 4471 24087 4477
rect 24029 4437 24041 4471
rect 24075 4468 24087 4471
rect 24118 4468 24124 4480
rect 24075 4440 24124 4468
rect 24075 4437 24087 4440
rect 24029 4431 24087 4437
rect 24118 4428 24124 4440
rect 24176 4428 24182 4480
rect 25130 4468 25136 4480
rect 25091 4440 25136 4468
rect 25130 4428 25136 4440
rect 25188 4428 25194 4480
rect 25961 4471 26019 4477
rect 25961 4437 25973 4471
rect 26007 4468 26019 4471
rect 26234 4468 26240 4480
rect 26007 4440 26240 4468
rect 26007 4437 26019 4440
rect 25961 4431 26019 4437
rect 26234 4428 26240 4440
rect 26292 4428 26298 4480
rect 1104 4378 29440 4400
rect 1104 4326 10395 4378
rect 10447 4326 10459 4378
rect 10511 4326 10523 4378
rect 10575 4326 10587 4378
rect 10639 4326 10651 4378
rect 10703 4326 19840 4378
rect 19892 4326 19904 4378
rect 19956 4326 19968 4378
rect 20020 4326 20032 4378
rect 20084 4326 20096 4378
rect 20148 4326 29440 4378
rect 1104 4304 29440 4326
rect 6733 4267 6791 4273
rect 6733 4233 6745 4267
rect 6779 4264 6791 4267
rect 6914 4264 6920 4276
rect 6779 4236 6920 4264
rect 6779 4233 6791 4236
rect 6733 4227 6791 4233
rect 6914 4224 6920 4236
rect 6972 4224 6978 4276
rect 8938 4264 8944 4276
rect 8899 4236 8944 4264
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 9398 4264 9404 4276
rect 9359 4236 9404 4264
rect 9398 4224 9404 4236
rect 9456 4224 9462 4276
rect 13538 4224 13544 4276
rect 13596 4224 13602 4276
rect 18693 4267 18751 4273
rect 18693 4264 18705 4267
rect 18616 4236 18705 4264
rect 3786 4156 3792 4208
rect 3844 4196 3850 4208
rect 3844 4168 6040 4196
rect 3844 4156 3850 4168
rect 5902 4128 5908 4140
rect 5960 4137 5966 4140
rect 5872 4100 5908 4128
rect 5902 4088 5908 4100
rect 5960 4091 5972 4137
rect 6012 4128 6040 4168
rect 6181 4131 6239 4137
rect 6181 4128 6193 4131
rect 6012 4100 6193 4128
rect 6181 4097 6193 4100
rect 6227 4097 6239 4131
rect 6932 4128 6960 4224
rect 9309 4199 9367 4205
rect 9309 4165 9321 4199
rect 9355 4196 9367 4199
rect 9490 4196 9496 4208
rect 9355 4168 9496 4196
rect 9355 4165 9367 4168
rect 9309 4159 9367 4165
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 11238 4196 11244 4208
rect 11151 4168 11244 4196
rect 11238 4156 11244 4168
rect 11296 4196 11302 4208
rect 12434 4196 12440 4208
rect 11296 4168 12440 4196
rect 11296 4156 11302 4168
rect 12434 4156 12440 4168
rect 12492 4156 12498 4208
rect 13357 4199 13415 4205
rect 13357 4165 13369 4199
rect 13403 4196 13415 4199
rect 13556 4196 13584 4224
rect 13403 4168 13584 4196
rect 15289 4199 15347 4205
rect 13403 4165 13415 4168
rect 13357 4159 13415 4165
rect 15289 4165 15301 4199
rect 15335 4196 15347 4199
rect 15654 4196 15660 4208
rect 15335 4168 15660 4196
rect 15335 4165 15347 4168
rect 15289 4159 15347 4165
rect 15654 4156 15660 4168
rect 15712 4156 15718 4208
rect 17773 4199 17831 4205
rect 17773 4165 17785 4199
rect 17819 4196 17831 4199
rect 17954 4196 17960 4208
rect 17819 4168 17960 4196
rect 17819 4165 17831 4168
rect 17773 4159 17831 4165
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 18414 4196 18420 4208
rect 18375 4168 18420 4196
rect 18414 4156 18420 4168
rect 18472 4156 18478 4208
rect 18506 4156 18512 4208
rect 18564 4196 18570 4208
rect 18616 4205 18644 4236
rect 18693 4233 18705 4236
rect 18739 4233 18751 4267
rect 18693 4227 18751 4233
rect 19702 4224 19708 4276
rect 19760 4264 19766 4276
rect 20349 4267 20407 4273
rect 20349 4264 20361 4267
rect 19760 4236 20361 4264
rect 19760 4224 19766 4236
rect 20349 4233 20361 4236
rect 20395 4233 20407 4267
rect 20349 4227 20407 4233
rect 21545 4267 21603 4273
rect 21545 4233 21557 4267
rect 21591 4264 21603 4267
rect 21910 4264 21916 4276
rect 21591 4236 21916 4264
rect 21591 4233 21603 4236
rect 21545 4227 21603 4233
rect 21910 4224 21916 4236
rect 21968 4224 21974 4276
rect 22370 4224 22376 4276
rect 22428 4264 22434 4276
rect 23474 4264 23480 4276
rect 22428 4236 23480 4264
rect 22428 4224 22434 4236
rect 23474 4224 23480 4236
rect 23532 4224 23538 4276
rect 23566 4224 23572 4276
rect 23624 4264 23630 4276
rect 23753 4267 23811 4273
rect 23753 4264 23765 4267
rect 23624 4236 23765 4264
rect 23624 4224 23630 4236
rect 23753 4233 23765 4236
rect 23799 4233 23811 4267
rect 23753 4227 23811 4233
rect 26234 4224 26240 4276
rect 26292 4264 26298 4276
rect 27246 4264 27252 4276
rect 26292 4236 27252 4264
rect 26292 4224 26298 4236
rect 27246 4224 27252 4236
rect 27304 4224 27310 4276
rect 18601 4199 18659 4205
rect 18601 4196 18613 4199
rect 18564 4168 18613 4196
rect 18564 4156 18570 4168
rect 18601 4165 18613 4168
rect 18647 4165 18659 4199
rect 18601 4159 18659 4165
rect 19058 4156 19064 4208
rect 19116 4196 19122 4208
rect 24848 4199 24906 4205
rect 19116 4168 19288 4196
rect 19116 4156 19122 4168
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 6932 4100 7481 4128
rect 6181 4091 6239 4097
rect 7469 4097 7481 4100
rect 7515 4097 7527 4131
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 7469 4091 7527 4097
rect 7576 4100 7757 4128
rect 5960 4088 5966 4091
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6696 4032 6837 4060
rect 6696 4020 6702 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 7006 4020 7012 4072
rect 7064 4060 7070 4072
rect 7576 4060 7604 4100
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 9858 4128 9864 4140
rect 7745 4091 7803 4097
rect 9508 4100 9864 4128
rect 9508 4069 9536 4100
rect 9858 4088 9864 4100
rect 9916 4128 9922 4140
rect 10134 4128 10140 4140
rect 9916 4100 10140 4128
rect 9916 4088 9922 4100
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4128 11115 4131
rect 11146 4128 11152 4140
rect 11103 4100 11152 4128
rect 11103 4097 11115 4100
rect 11057 4091 11115 4097
rect 11146 4088 11152 4100
rect 11204 4088 11210 4140
rect 12345 4131 12403 4137
rect 12345 4097 12357 4131
rect 12391 4128 12403 4131
rect 13170 4128 13176 4140
rect 12391 4100 13176 4128
rect 12391 4097 12403 4100
rect 12345 4091 12403 4097
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 13538 4128 13544 4140
rect 13499 4100 13544 4128
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 13722 4128 13728 4140
rect 13683 4100 13728 4128
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 15473 4131 15531 4137
rect 15473 4097 15485 4131
rect 15519 4128 15531 4131
rect 15562 4128 15568 4140
rect 15519 4100 15568 4128
rect 15519 4097 15531 4100
rect 15473 4091 15531 4097
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 15746 4088 15752 4140
rect 15804 4128 15810 4140
rect 16761 4131 16819 4137
rect 16761 4128 16773 4131
rect 15804 4100 16773 4128
rect 15804 4088 15810 4100
rect 16761 4097 16773 4100
rect 16807 4097 16819 4131
rect 16942 4128 16948 4140
rect 16903 4100 16948 4128
rect 16761 4091 16819 4097
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17586 4128 17592 4140
rect 17547 4100 17592 4128
rect 17586 4088 17592 4100
rect 17644 4088 17650 4140
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4097 18935 4131
rect 19153 4131 19211 4137
rect 19153 4128 19165 4131
rect 18877 4091 18935 4097
rect 18984 4100 19165 4128
rect 7064 4032 7604 4060
rect 7653 4063 7711 4069
rect 7064 4020 7070 4032
rect 7653 4029 7665 4063
rect 7699 4029 7711 4063
rect 7653 4023 7711 4029
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4029 9551 4063
rect 9493 4023 9551 4029
rect 6730 3952 6736 4004
rect 6788 3992 6794 4004
rect 7668 3992 7696 4023
rect 9582 4020 9588 4072
rect 9640 4060 9646 4072
rect 14642 4060 14648 4072
rect 9640 4032 14648 4060
rect 9640 4020 9646 4032
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 16632 4032 16681 4060
rect 16632 4020 16638 4032
rect 16669 4029 16681 4032
rect 16715 4029 16727 4063
rect 16669 4023 16727 4029
rect 17957 4063 18015 4069
rect 17957 4029 17969 4063
rect 18003 4060 18015 4063
rect 18892 4060 18920 4091
rect 18003 4032 18920 4060
rect 18003 4029 18015 4032
rect 17957 4023 18015 4029
rect 6788 3964 7696 3992
rect 6788 3952 6794 3964
rect 12802 3952 12808 4004
rect 12860 3992 12866 4004
rect 18138 3992 18144 4004
rect 12860 3964 18144 3992
rect 12860 3952 12866 3964
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18233 3995 18291 4001
rect 18233 3961 18245 3995
rect 18279 3992 18291 3995
rect 18984 3992 19012 4100
rect 19153 4097 19165 4100
rect 19199 4097 19211 4131
rect 19260 4128 19288 4168
rect 20548 4168 20852 4196
rect 20548 4128 20576 4168
rect 20714 4128 20720 4140
rect 19260 4100 20576 4128
rect 20675 4100 20720 4128
rect 19153 4091 19211 4097
rect 20714 4088 20720 4100
rect 20772 4088 20778 4140
rect 20824 4128 20852 4168
rect 24848 4165 24860 4199
rect 24894 4196 24906 4199
rect 25130 4196 25136 4208
rect 24894 4168 25136 4196
rect 24894 4165 24906 4168
rect 24848 4159 24906 4165
rect 25130 4156 25136 4168
rect 25188 4156 25194 4208
rect 26789 4199 26847 4205
rect 26789 4165 26801 4199
rect 26835 4196 26847 4199
rect 27522 4196 27528 4208
rect 26835 4168 27528 4196
rect 26835 4165 26847 4168
rect 26789 4159 26847 4165
rect 27522 4156 27528 4168
rect 27580 4156 27586 4208
rect 20824 4100 20944 4128
rect 20916 4069 20944 4100
rect 21266 4088 21272 4140
rect 21324 4128 21330 4140
rect 21361 4131 21419 4137
rect 21361 4128 21373 4131
rect 21324 4100 21373 4128
rect 21324 4088 21330 4100
rect 21361 4097 21373 4100
rect 21407 4097 21419 4131
rect 21361 4091 21419 4097
rect 23845 4131 23903 4137
rect 23845 4097 23857 4131
rect 23891 4128 23903 4131
rect 23934 4128 23940 4140
rect 23891 4100 23940 4128
rect 23891 4097 23903 4100
rect 23845 4091 23903 4097
rect 23934 4088 23940 4100
rect 23992 4088 23998 4140
rect 26421 4131 26479 4137
rect 26421 4097 26433 4131
rect 26467 4128 26479 4131
rect 26510 4128 26516 4140
rect 26467 4100 26516 4128
rect 26467 4097 26479 4100
rect 26421 4091 26479 4097
rect 26510 4088 26516 4100
rect 26568 4088 26574 4140
rect 26605 4131 26663 4137
rect 26605 4097 26617 4131
rect 26651 4128 26663 4131
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 26651 4100 26985 4128
rect 26651 4097 26663 4100
rect 26605 4091 26663 4097
rect 26973 4097 26985 4100
rect 27019 4097 27031 4131
rect 26973 4091 27031 4097
rect 29549 4131 29607 4137
rect 29549 4097 29561 4131
rect 29595 4128 29607 4131
rect 29822 4128 29828 4140
rect 29595 4100 29828 4128
rect 29595 4097 29607 4100
rect 29549 4091 29607 4097
rect 20809 4063 20867 4069
rect 20809 4029 20821 4063
rect 20855 4029 20867 4063
rect 20809 4023 20867 4029
rect 20901 4063 20959 4069
rect 20901 4029 20913 4063
rect 20947 4060 20959 4063
rect 21542 4060 21548 4072
rect 20947 4032 21548 4060
rect 20947 4029 20959 4032
rect 20901 4023 20959 4029
rect 18279 3964 19012 3992
rect 20824 3992 20852 4023
rect 21542 4020 21548 4032
rect 21600 4020 21606 4072
rect 24581 4063 24639 4069
rect 24581 4029 24593 4063
rect 24627 4029 24639 4063
rect 24581 4023 24639 4029
rect 22462 3992 22468 4004
rect 20824 3964 22468 3992
rect 18279 3961 18291 3964
rect 18233 3955 18291 3961
rect 22462 3952 22468 3964
rect 22520 3952 22526 4004
rect 4801 3927 4859 3933
rect 4801 3893 4813 3927
rect 4847 3924 4859 3927
rect 5442 3924 5448 3936
rect 4847 3896 5448 3924
rect 4847 3893 4859 3896
rect 4801 3887 4859 3893
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 5994 3884 6000 3936
rect 6052 3924 6058 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6052 3896 6377 3924
rect 6052 3884 6058 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 7285 3927 7343 3933
rect 7285 3924 7297 3927
rect 6512 3896 7297 3924
rect 6512 3884 6518 3896
rect 7285 3893 7297 3896
rect 7331 3893 7343 3927
rect 7285 3887 7343 3893
rect 10965 3927 11023 3933
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 11054 3924 11060 3936
rect 11011 3896 11060 3924
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 12158 3924 12164 3936
rect 12119 3896 12164 3924
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 12710 3924 12716 3936
rect 12671 3896 12716 3924
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 15197 3927 15255 3933
rect 15197 3924 15209 3927
rect 15068 3896 15209 3924
rect 15068 3884 15074 3896
rect 15197 3893 15209 3896
rect 15243 3893 15255 3927
rect 15197 3887 15255 3893
rect 18414 3884 18420 3936
rect 18472 3924 18478 3936
rect 18969 3927 19027 3933
rect 18969 3924 18981 3927
rect 18472 3896 18981 3924
rect 18472 3884 18478 3896
rect 18969 3893 18981 3896
rect 19015 3893 19027 3927
rect 18969 3887 19027 3893
rect 19058 3884 19064 3936
rect 19116 3924 19122 3936
rect 22738 3924 22744 3936
rect 19116 3896 22744 3924
rect 19116 3884 19122 3896
rect 22738 3884 22744 3896
rect 22796 3884 22802 3936
rect 24596 3924 24624 4023
rect 25961 3995 26019 4001
rect 25961 3961 25973 3995
rect 26007 3992 26019 3995
rect 26620 3992 26648 4091
rect 29822 4088 29828 4100
rect 29880 4088 29886 4140
rect 26007 3964 26648 3992
rect 26007 3961 26019 3964
rect 25961 3955 26019 3961
rect 24946 3924 24952 3936
rect 24596 3896 24952 3924
rect 24946 3884 24952 3896
rect 25004 3884 25010 3936
rect 1104 3834 29440 3856
rect 1104 3782 5672 3834
rect 5724 3782 5736 3834
rect 5788 3782 5800 3834
rect 5852 3782 5864 3834
rect 5916 3782 5928 3834
rect 5980 3782 15118 3834
rect 15170 3782 15182 3834
rect 15234 3782 15246 3834
rect 15298 3782 15310 3834
rect 15362 3782 15374 3834
rect 15426 3782 24563 3834
rect 24615 3782 24627 3834
rect 24679 3782 24691 3834
rect 24743 3782 24755 3834
rect 24807 3782 24819 3834
rect 24871 3782 29440 3834
rect 1104 3760 29440 3782
rect 6638 3720 6644 3732
rect 6599 3692 6644 3720
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 9214 3680 9220 3732
rect 9272 3720 9278 3732
rect 9398 3720 9404 3732
rect 9272 3692 9404 3720
rect 9272 3680 9278 3692
rect 9398 3680 9404 3692
rect 9456 3720 9462 3732
rect 9493 3723 9551 3729
rect 9493 3720 9505 3723
rect 9456 3692 9505 3720
rect 9456 3680 9462 3692
rect 9493 3689 9505 3692
rect 9539 3720 9551 3723
rect 12710 3720 12716 3732
rect 9539 3692 12716 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 9582 3652 9588 3664
rect 4212 3624 9588 3652
rect 4212 3612 4218 3624
rect 9582 3612 9588 3624
rect 9640 3612 9646 3664
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 6362 3584 6368 3596
rect 1820 3556 6368 3584
rect 1820 3544 1826 3556
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 6638 3544 6644 3596
rect 6696 3584 6702 3596
rect 8110 3584 8116 3596
rect 6696 3556 8116 3584
rect 6696 3544 6702 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 10060 3593 10088 3692
rect 12710 3680 12716 3692
rect 12768 3720 12774 3732
rect 13170 3720 13176 3732
rect 12768 3692 12848 3720
rect 13131 3692 13176 3720
rect 12768 3680 12774 3692
rect 11054 3652 11060 3664
rect 10980 3624 11060 3652
rect 10045 3587 10103 3593
rect 10045 3553 10057 3587
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 6454 3516 6460 3528
rect 6415 3488 6460 3516
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 9861 3519 9919 3525
rect 9861 3485 9873 3519
rect 9907 3516 9919 3519
rect 10321 3519 10379 3525
rect 9907 3488 9996 3516
rect 9907 3485 9919 3488
rect 9861 3479 9919 3485
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 7926 3448 7932 3460
rect 5500 3420 7932 3448
rect 5500 3408 5506 3420
rect 7926 3408 7932 3420
rect 7984 3408 7990 3460
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 9677 3451 9735 3457
rect 9677 3448 9689 3451
rect 9088 3420 9689 3448
rect 9088 3408 9094 3420
rect 9677 3417 9689 3420
rect 9723 3417 9735 3451
rect 9677 3411 9735 3417
rect 9968 3392 9996 3488
rect 10321 3485 10333 3519
rect 10367 3516 10379 3519
rect 10505 3519 10563 3525
rect 10505 3516 10517 3519
rect 10367 3488 10517 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 10505 3485 10517 3488
rect 10551 3485 10563 3519
rect 10505 3479 10563 3485
rect 10747 3519 10805 3525
rect 10747 3485 10759 3519
rect 10793 3516 10805 3519
rect 10980 3516 11008 3624
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11238 3584 11244 3596
rect 11195 3556 11244 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 12820 3584 12848 3692
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 15470 3680 15476 3732
rect 15528 3720 15534 3732
rect 15565 3723 15623 3729
rect 15565 3720 15577 3723
rect 15528 3692 15577 3720
rect 15528 3680 15534 3692
rect 15565 3689 15577 3692
rect 15611 3689 15623 3723
rect 15565 3683 15623 3689
rect 15749 3723 15807 3729
rect 15749 3689 15761 3723
rect 15795 3689 15807 3723
rect 15749 3683 15807 3689
rect 16117 3723 16175 3729
rect 16117 3689 16129 3723
rect 16163 3720 16175 3723
rect 17586 3720 17592 3732
rect 16163 3692 17448 3720
rect 17547 3692 17592 3720
rect 16163 3689 16175 3692
rect 16117 3683 16175 3689
rect 12897 3655 12955 3661
rect 12897 3621 12909 3655
rect 12943 3652 12955 3655
rect 13538 3652 13544 3664
rect 12943 3624 13544 3652
rect 12943 3621 12955 3624
rect 12897 3615 12955 3621
rect 13538 3612 13544 3624
rect 13596 3652 13602 3664
rect 15764 3652 15792 3683
rect 13596 3624 15792 3652
rect 13596 3612 13602 3624
rect 15838 3612 15844 3664
rect 15896 3652 15902 3664
rect 17420 3652 17448 3692
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 21266 3720 21272 3732
rect 21227 3692 21272 3720
rect 21266 3680 21272 3692
rect 21324 3680 21330 3732
rect 21542 3680 21548 3732
rect 21600 3720 21606 3732
rect 22462 3720 22468 3732
rect 21600 3692 22094 3720
rect 22423 3692 22468 3720
rect 21600 3680 21606 3692
rect 18046 3652 18052 3664
rect 15896 3624 17356 3652
rect 17420 3624 18052 3652
rect 15896 3612 15902 3624
rect 13354 3584 13360 3596
rect 12820 3556 13360 3584
rect 13354 3544 13360 3556
rect 13412 3544 13418 3596
rect 10793 3488 11008 3516
rect 10793 3485 10805 3488
rect 10747 3479 10805 3485
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11514 3516 11520 3528
rect 11112 3488 11157 3516
rect 11475 3488 11520 3516
rect 11112 3476 11118 3488
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 13556 3516 13584 3612
rect 13722 3584 13728 3596
rect 13635 3556 13728 3584
rect 13722 3544 13728 3556
rect 13780 3584 13786 3596
rect 15654 3584 15660 3596
rect 13780 3556 14412 3584
rect 13780 3544 13786 3556
rect 13633 3519 13691 3525
rect 13633 3516 13645 3519
rect 13320 3488 13365 3516
rect 13556 3488 13645 3516
rect 13320 3476 13326 3488
rect 13633 3485 13645 3488
rect 13679 3485 13691 3519
rect 14274 3516 14280 3528
rect 14235 3488 14280 3516
rect 13633 3479 13691 3485
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 14384 3516 14412 3556
rect 15304 3556 15660 3584
rect 15304 3528 15332 3556
rect 15654 3544 15660 3556
rect 15712 3584 15718 3596
rect 16117 3587 16175 3593
rect 15712 3556 15792 3584
rect 15712 3544 15718 3556
rect 15010 3525 15016 3528
rect 14979 3519 15016 3525
rect 14979 3516 14991 3519
rect 14384 3488 14991 3516
rect 14979 3485 14991 3488
rect 14979 3479 15016 3485
rect 15010 3476 15016 3479
rect 15068 3476 15074 3528
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3516 15439 3519
rect 15562 3516 15568 3528
rect 15427 3488 15568 3516
rect 15427 3485 15439 3488
rect 15381 3479 15439 3485
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 15764 3525 15792 3556
rect 16117 3553 16129 3587
rect 16163 3584 16175 3587
rect 16301 3587 16359 3593
rect 16301 3584 16313 3587
rect 16163 3556 16313 3584
rect 16163 3553 16175 3556
rect 16117 3547 16175 3553
rect 16301 3553 16313 3556
rect 16347 3553 16359 3587
rect 16301 3547 16359 3553
rect 16485 3587 16543 3593
rect 16485 3553 16497 3587
rect 16531 3584 16543 3587
rect 16574 3584 16580 3596
rect 16531 3556 16580 3584
rect 16531 3553 16543 3556
rect 16485 3547 16543 3553
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 17126 3584 17132 3596
rect 17087 3556 17132 3584
rect 17126 3544 17132 3556
rect 17184 3544 17190 3596
rect 17328 3584 17356 3624
rect 18046 3612 18052 3624
rect 18104 3652 18110 3664
rect 20625 3655 20683 3661
rect 18104 3624 18276 3652
rect 18104 3612 18110 3624
rect 18248 3593 18276 3624
rect 20625 3621 20637 3655
rect 20671 3652 20683 3655
rect 20714 3652 20720 3664
rect 20671 3624 20720 3652
rect 20671 3621 20683 3624
rect 20625 3615 20683 3621
rect 20714 3612 20720 3624
rect 20772 3652 20778 3664
rect 21818 3652 21824 3664
rect 20772 3624 21824 3652
rect 20772 3612 20778 3624
rect 21818 3612 21824 3624
rect 21876 3612 21882 3664
rect 18233 3587 18291 3593
rect 17328 3556 17448 3584
rect 15749 3519 15807 3525
rect 15749 3485 15761 3519
rect 15795 3485 15807 3519
rect 15749 3479 15807 3485
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3516 15899 3519
rect 17037 3519 17095 3525
rect 15887 3488 16620 3516
rect 15887 3485 15899 3488
rect 15841 3479 15899 3485
rect 11790 3457 11796 3460
rect 11784 3411 11796 3457
rect 11848 3448 11854 3460
rect 11848 3420 11884 3448
rect 11790 3408 11796 3411
rect 11848 3408 11854 3420
rect 13814 3408 13820 3460
rect 13872 3448 13878 3460
rect 13872 3420 14412 3448
rect 13872 3408 13878 3420
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 10137 3383 10195 3389
rect 10137 3380 10149 3383
rect 10008 3352 10149 3380
rect 10008 3340 10014 3352
rect 10137 3349 10149 3352
rect 10183 3349 10195 3383
rect 10137 3343 10195 3349
rect 11514 3340 11520 3392
rect 11572 3380 11578 3392
rect 12342 3380 12348 3392
rect 11572 3352 12348 3380
rect 11572 3340 11578 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 13262 3340 13268 3392
rect 13320 3380 13326 3392
rect 14093 3383 14151 3389
rect 14093 3380 14105 3383
rect 13320 3352 14105 3380
rect 13320 3340 13326 3352
rect 14093 3349 14105 3352
rect 14139 3349 14151 3383
rect 14384 3380 14412 3420
rect 14458 3408 14464 3460
rect 14516 3448 14522 3460
rect 14737 3451 14795 3457
rect 14737 3448 14749 3451
rect 14516 3420 14749 3448
rect 14516 3408 14522 3420
rect 14737 3417 14749 3420
rect 14783 3417 14795 3451
rect 16022 3448 16028 3460
rect 15983 3420 16028 3448
rect 14737 3411 14795 3417
rect 16022 3408 16028 3420
rect 16080 3408 16086 3460
rect 16592 3457 16620 3488
rect 17037 3485 17049 3519
rect 17083 3485 17095 3519
rect 17310 3516 17316 3528
rect 17271 3488 17316 3516
rect 17037 3479 17095 3485
rect 16577 3451 16635 3457
rect 16577 3417 16589 3451
rect 16623 3448 16635 3451
rect 17052 3448 17080 3479
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17420 3525 17448 3556
rect 18233 3553 18245 3587
rect 18279 3553 18291 3587
rect 18414 3584 18420 3596
rect 18375 3556 18420 3584
rect 18233 3547 18291 3553
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 21433 3587 21491 3593
rect 21433 3584 21445 3587
rect 21376 3556 21445 3584
rect 17405 3519 17463 3525
rect 17405 3485 17417 3519
rect 17451 3516 17463 3519
rect 17957 3519 18015 3525
rect 17957 3516 17969 3519
rect 17451 3488 17969 3516
rect 17451 3485 17463 3488
rect 17405 3479 17463 3485
rect 17957 3485 17969 3488
rect 18003 3516 18015 3519
rect 18046 3516 18052 3528
rect 18003 3488 18052 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 18506 3516 18512 3528
rect 18467 3488 18512 3516
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3516 19303 3519
rect 19291 3488 19748 3516
rect 19291 3485 19303 3488
rect 19245 3479 19303 3485
rect 19720 3460 19748 3488
rect 19518 3457 19524 3460
rect 17865 3451 17923 3457
rect 17865 3448 17877 3451
rect 16623 3420 17877 3448
rect 16623 3417 16635 3420
rect 16577 3411 16635 3417
rect 17865 3417 17877 3420
rect 17911 3417 17923 3451
rect 19512 3448 19524 3457
rect 19479 3420 19524 3448
rect 17865 3411 17923 3417
rect 19512 3411 19524 3420
rect 19518 3408 19524 3411
rect 19576 3408 19582 3460
rect 19702 3408 19708 3460
rect 19760 3408 19766 3460
rect 21266 3408 21272 3460
rect 21324 3448 21330 3460
rect 21376 3448 21404 3556
rect 21433 3553 21445 3556
rect 21479 3553 21491 3587
rect 22066 3584 22094 3692
rect 22462 3680 22468 3692
rect 22520 3680 22526 3732
rect 23198 3720 23204 3732
rect 23159 3692 23204 3720
rect 23198 3680 23204 3692
rect 23256 3680 23262 3732
rect 26605 3723 26663 3729
rect 26605 3689 26617 3723
rect 26651 3720 26663 3723
rect 26786 3720 26792 3732
rect 26651 3692 26792 3720
rect 26651 3689 26663 3692
rect 26605 3683 26663 3689
rect 26786 3680 26792 3692
rect 26844 3720 26850 3732
rect 27338 3720 27344 3732
rect 26844 3692 27344 3720
rect 26844 3680 26850 3692
rect 27338 3680 27344 3692
rect 27396 3680 27402 3732
rect 23753 3587 23811 3593
rect 23753 3584 23765 3587
rect 22066 3556 23765 3584
rect 21433 3547 21491 3553
rect 23753 3553 23765 3556
rect 23799 3584 23811 3587
rect 25866 3584 25872 3596
rect 23799 3556 25872 3584
rect 23799 3553 23811 3556
rect 23753 3547 23811 3553
rect 25866 3544 25872 3556
rect 25924 3544 25930 3596
rect 21542 3516 21548 3528
rect 21503 3488 21548 3516
rect 21542 3476 21548 3488
rect 21600 3516 21606 3528
rect 21821 3519 21879 3525
rect 21821 3516 21833 3519
rect 21600 3488 21833 3516
rect 21600 3476 21606 3488
rect 21821 3485 21833 3488
rect 21867 3485 21879 3519
rect 22002 3516 22008 3528
rect 21963 3488 22008 3516
rect 21821 3479 21879 3485
rect 22002 3476 22008 3488
rect 22060 3476 22066 3528
rect 22281 3519 22339 3525
rect 22281 3485 22293 3519
rect 22327 3516 22339 3519
rect 23566 3516 23572 3528
rect 22327 3488 23572 3516
rect 22327 3485 22339 3488
rect 22281 3479 22339 3485
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 23842 3476 23848 3528
rect 23900 3516 23906 3528
rect 24029 3519 24087 3525
rect 24029 3516 24041 3519
rect 23900 3488 24041 3516
rect 23900 3476 23906 3488
rect 24029 3485 24041 3488
rect 24075 3485 24087 3519
rect 26510 3516 26516 3528
rect 26471 3488 26516 3516
rect 24029 3479 24087 3485
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 21913 3451 21971 3457
rect 21913 3448 21925 3451
rect 21324 3420 21925 3448
rect 21324 3408 21330 3420
rect 21913 3417 21925 3420
rect 21959 3417 21971 3451
rect 23750 3448 23756 3460
rect 21913 3411 21971 3417
rect 23584 3420 23756 3448
rect 16117 3383 16175 3389
rect 16117 3380 16129 3383
rect 14384 3352 16129 3380
rect 14093 3343 14151 3349
rect 16117 3349 16129 3352
rect 16163 3349 16175 3383
rect 16942 3380 16948 3392
rect 16903 3352 16948 3380
rect 16117 3343 16175 3349
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 18874 3380 18880 3392
rect 18835 3352 18880 3380
rect 18874 3340 18880 3352
rect 18932 3340 18938 3392
rect 21928 3380 21956 3411
rect 22002 3380 22008 3392
rect 21928 3352 22008 3380
rect 22002 3340 22008 3352
rect 22060 3380 22066 3392
rect 23584 3389 23612 3420
rect 23750 3408 23756 3420
rect 23808 3448 23814 3460
rect 24121 3451 24179 3457
rect 24121 3448 24133 3451
rect 23808 3420 24133 3448
rect 23808 3408 23814 3420
rect 24121 3417 24133 3420
rect 24167 3417 24179 3451
rect 24121 3411 24179 3417
rect 22097 3383 22155 3389
rect 22097 3380 22109 3383
rect 22060 3352 22109 3380
rect 22060 3340 22066 3352
rect 22097 3349 22109 3352
rect 22143 3349 22155 3383
rect 22097 3343 22155 3349
rect 23569 3383 23627 3389
rect 23569 3349 23581 3383
rect 23615 3349 23627 3383
rect 23569 3343 23627 3349
rect 23658 3340 23664 3392
rect 23716 3380 23722 3392
rect 23716 3352 23761 3380
rect 23716 3340 23722 3352
rect 1104 3290 29440 3312
rect 1104 3238 10395 3290
rect 10447 3238 10459 3290
rect 10511 3238 10523 3290
rect 10575 3238 10587 3290
rect 10639 3238 10651 3290
rect 10703 3238 19840 3290
rect 19892 3238 19904 3290
rect 19956 3238 19968 3290
rect 20020 3238 20032 3290
rect 20084 3238 20096 3290
rect 20148 3238 29440 3290
rect 1104 3216 29440 3238
rect 10689 3179 10747 3185
rect 10689 3145 10701 3179
rect 10735 3176 10747 3179
rect 11054 3176 11060 3188
rect 10735 3148 11060 3176
rect 10735 3145 10747 3148
rect 10689 3139 10747 3145
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 11701 3179 11759 3185
rect 11701 3145 11713 3179
rect 11747 3176 11759 3179
rect 11790 3176 11796 3188
rect 11747 3148 11796 3176
rect 11747 3145 11759 3148
rect 11701 3139 11759 3145
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 12069 3179 12127 3185
rect 12069 3145 12081 3179
rect 12115 3176 12127 3179
rect 12158 3176 12164 3188
rect 12115 3148 12164 3176
rect 12115 3145 12127 3148
rect 12069 3139 12127 3145
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 12529 3179 12587 3185
rect 12529 3176 12541 3179
rect 12268 3148 12541 3176
rect 11514 3108 11520 3120
rect 9324 3080 11520 3108
rect 9030 3040 9036 3052
rect 8991 3012 9036 3040
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9324 3049 9352 3080
rect 11514 3068 11520 3080
rect 11572 3068 11578 3120
rect 9582 3049 9588 3052
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 9576 3003 9588 3049
rect 9640 3040 9646 3052
rect 9640 3012 9676 3040
rect 9582 3000 9588 3003
rect 9640 3000 9646 3012
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 12161 3043 12219 3049
rect 10192 3012 11560 3040
rect 10192 3000 10198 3012
rect 2958 2972 2964 2984
rect 2919 2944 2964 2972
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 7834 2972 7840 2984
rect 7795 2944 7840 2972
rect 7834 2932 7840 2944
rect 7892 2932 7898 2984
rect 11532 2972 11560 3012
rect 12161 3009 12173 3043
rect 12207 3040 12219 3043
rect 12268 3040 12296 3148
rect 12529 3145 12541 3148
rect 12575 3145 12587 3179
rect 12529 3139 12587 3145
rect 13173 3179 13231 3185
rect 13173 3145 13185 3179
rect 13219 3176 13231 3179
rect 13262 3176 13268 3188
rect 13219 3148 13268 3176
rect 13219 3145 13231 3148
rect 13173 3139 13231 3145
rect 13262 3136 13268 3148
rect 13320 3136 13326 3188
rect 13633 3179 13691 3185
rect 13633 3145 13645 3179
rect 13679 3176 13691 3179
rect 15105 3179 15163 3185
rect 13679 3148 13860 3176
rect 13679 3145 13691 3148
rect 13633 3139 13691 3145
rect 13832 3108 13860 3148
rect 15105 3145 15117 3179
rect 15151 3176 15163 3179
rect 15286 3176 15292 3188
rect 15151 3148 15292 3176
rect 15151 3145 15163 3148
rect 15105 3139 15163 3145
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 16022 3176 16028 3188
rect 15935 3148 16028 3176
rect 13970 3111 14028 3117
rect 13970 3108 13982 3111
rect 12406 3080 13768 3108
rect 13832 3080 13982 3108
rect 12406 3052 12434 3080
rect 12207 3012 12296 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12342 3000 12348 3052
rect 12400 3012 12434 3052
rect 12710 3040 12716 3052
rect 12671 3012 12716 3040
rect 12400 3000 12406 3012
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3040 13323 3043
rect 13630 3040 13636 3052
rect 13311 3012 13636 3040
rect 13311 3009 13323 3012
rect 13265 3003 13323 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 13740 3049 13768 3080
rect 13970 3077 13982 3080
rect 14016 3077 14028 3111
rect 15562 3108 15568 3120
rect 15523 3080 15568 3108
rect 13970 3071 14028 3077
rect 15562 3068 15568 3080
rect 15620 3068 15626 3120
rect 15746 3108 15752 3120
rect 15707 3080 15752 3108
rect 15746 3068 15752 3080
rect 15804 3068 15810 3120
rect 15948 3117 15976 3148
rect 16022 3136 16028 3148
rect 16080 3176 16086 3188
rect 17126 3176 17132 3188
rect 16080 3148 17132 3176
rect 16080 3136 16086 3148
rect 17126 3136 17132 3148
rect 17184 3176 17190 3188
rect 17402 3176 17408 3188
rect 17184 3148 17408 3176
rect 17184 3136 17190 3148
rect 17402 3136 17408 3148
rect 17460 3176 17466 3188
rect 18325 3179 18383 3185
rect 18325 3176 18337 3179
rect 17460 3148 18337 3176
rect 17460 3136 17466 3148
rect 18325 3145 18337 3148
rect 18371 3145 18383 3179
rect 21266 3176 21272 3188
rect 21227 3148 21272 3176
rect 18325 3139 18383 3145
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 23566 3176 23572 3188
rect 23527 3148 23572 3176
rect 23566 3136 23572 3148
rect 23624 3136 23630 3188
rect 23934 3136 23940 3188
rect 23992 3176 23998 3188
rect 25409 3179 25467 3185
rect 25409 3176 25421 3179
rect 23992 3148 25421 3176
rect 23992 3136 23998 3148
rect 25409 3145 25421 3148
rect 25455 3145 25467 3179
rect 25409 3139 25467 3145
rect 25869 3179 25927 3185
rect 25869 3145 25881 3179
rect 25915 3176 25927 3179
rect 26421 3179 26479 3185
rect 26421 3176 26433 3179
rect 25915 3148 26433 3176
rect 25915 3145 25927 3148
rect 25869 3139 25927 3145
rect 26421 3145 26433 3148
rect 26467 3145 26479 3179
rect 26421 3139 26479 3145
rect 16942 3117 16948 3120
rect 15933 3111 15991 3117
rect 15933 3077 15945 3111
rect 15979 3077 15991 3111
rect 16936 3108 16948 3117
rect 16903 3080 16948 3108
rect 15933 3071 15991 3077
rect 16936 3071 16948 3080
rect 16942 3068 16948 3071
rect 17000 3068 17006 3120
rect 18874 3068 18880 3120
rect 18932 3108 18938 3120
rect 19438 3111 19496 3117
rect 19438 3108 19450 3111
rect 18932 3080 19450 3108
rect 18932 3068 18938 3080
rect 19438 3077 19450 3080
rect 19484 3077 19496 3111
rect 24946 3108 24952 3120
rect 19438 3071 19496 3077
rect 19904 3080 24952 3108
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 13814 3000 13820 3052
rect 13872 3000 13878 3052
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 19702 3040 19708 3052
rect 16776 3012 18460 3040
rect 19663 3012 19708 3040
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 11532 2944 12265 2972
rect 12253 2941 12265 2944
rect 12299 2972 12311 2975
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12299 2944 13001 2972
rect 12299 2941 12311 2944
rect 12253 2935 12311 2941
rect 12989 2941 13001 2944
rect 13035 2972 13047 2975
rect 13832 2972 13860 3000
rect 13035 2944 13860 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 14918 2932 14924 2984
rect 14976 2972 14982 2984
rect 16776 2972 16804 3012
rect 14976 2944 16804 2972
rect 14976 2932 14982 2944
rect 18046 2904 18052 2916
rect 18007 2876 18052 2904
rect 18046 2864 18052 2876
rect 18104 2864 18110 2916
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2836 9275 2839
rect 10042 2836 10048 2848
rect 9263 2808 10048 2836
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 15470 2796 15476 2848
rect 15528 2836 15534 2848
rect 18322 2836 18328 2848
rect 15528 2808 18328 2836
rect 15528 2796 15534 2808
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 18432 2836 18460 3012
rect 19702 3000 19708 3012
rect 19760 3040 19766 3052
rect 19904 3049 19932 3080
rect 19889 3043 19947 3049
rect 19889 3040 19901 3043
rect 19760 3012 19901 3040
rect 19760 3000 19766 3012
rect 19889 3009 19901 3012
rect 19935 3009 19947 3043
rect 19889 3003 19947 3009
rect 20156 3043 20214 3049
rect 20156 3009 20168 3043
rect 20202 3040 20214 3043
rect 20990 3040 20996 3052
rect 20202 3012 20996 3040
rect 20202 3009 20214 3012
rect 20156 3003 20214 3009
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 21928 3049 21956 3080
rect 22186 3049 22192 3052
rect 21913 3043 21971 3049
rect 21913 3009 21925 3043
rect 21959 3009 21971 3043
rect 22180 3040 22192 3049
rect 22147 3012 22192 3040
rect 21913 3003 21971 3009
rect 22180 3003 22192 3012
rect 22186 3000 22192 3003
rect 22244 3000 22250 3052
rect 23566 3000 23572 3052
rect 23624 3040 23630 3052
rect 23860 3049 23888 3080
rect 24946 3068 24952 3080
rect 25004 3068 25010 3120
rect 24118 3049 24124 3052
rect 23661 3043 23719 3049
rect 23661 3040 23673 3043
rect 23624 3012 23673 3040
rect 23624 3000 23630 3012
rect 23661 3009 23673 3012
rect 23707 3009 23719 3043
rect 23661 3003 23719 3009
rect 23845 3043 23903 3049
rect 23845 3009 23857 3043
rect 23891 3009 23903 3043
rect 24112 3040 24124 3049
rect 24079 3012 24124 3040
rect 23845 3003 23903 3009
rect 24112 3003 24124 3012
rect 24118 3000 24124 3003
rect 24176 3000 24182 3052
rect 25774 3040 25780 3052
rect 25735 3012 25780 3040
rect 25774 3000 25780 3012
rect 25832 3000 25838 3052
rect 26050 3000 26056 3052
rect 26108 3040 26114 3052
rect 26421 3043 26479 3049
rect 26421 3040 26433 3043
rect 26108 3012 26433 3040
rect 26108 3000 26114 3012
rect 26421 3009 26433 3012
rect 26467 3009 26479 3043
rect 26786 3040 26792 3052
rect 26747 3012 26792 3040
rect 26421 3003 26479 3009
rect 26786 3000 26792 3012
rect 26844 3000 26850 3052
rect 25866 2932 25872 2984
rect 25924 2972 25930 2984
rect 25961 2975 26019 2981
rect 25961 2972 25973 2975
rect 25924 2944 25973 2972
rect 25924 2932 25930 2944
rect 25961 2941 25973 2944
rect 26007 2941 26019 2975
rect 25961 2935 26019 2941
rect 26142 2932 26148 2984
rect 26200 2972 26206 2984
rect 26237 2975 26295 2981
rect 26237 2972 26249 2975
rect 26200 2944 26249 2972
rect 26200 2932 26206 2944
rect 26237 2941 26249 2944
rect 26283 2941 26295 2975
rect 26237 2935 26295 2941
rect 23293 2907 23351 2913
rect 23293 2873 23305 2907
rect 23339 2904 23351 2907
rect 23842 2904 23848 2916
rect 23339 2876 23848 2904
rect 23339 2873 23351 2876
rect 23293 2867 23351 2873
rect 23842 2864 23848 2876
rect 23900 2864 23906 2916
rect 26326 2904 26332 2916
rect 25056 2876 26332 2904
rect 25056 2836 25084 2876
rect 26326 2864 26332 2876
rect 26384 2864 26390 2916
rect 25222 2836 25228 2848
rect 18432 2808 25084 2836
rect 25183 2808 25228 2836
rect 25222 2796 25228 2808
rect 25280 2796 25286 2848
rect 1104 2746 29440 2768
rect 1104 2694 5672 2746
rect 5724 2694 5736 2746
rect 5788 2694 5800 2746
rect 5852 2694 5864 2746
rect 5916 2694 5928 2746
rect 5980 2694 15118 2746
rect 15170 2694 15182 2746
rect 15234 2694 15246 2746
rect 15298 2694 15310 2746
rect 15362 2694 15374 2746
rect 15426 2694 24563 2746
rect 24615 2694 24627 2746
rect 24679 2694 24691 2746
rect 24743 2694 24755 2746
rect 24807 2694 24819 2746
rect 24871 2694 29440 2746
rect 1104 2672 29440 2694
rect 3050 2592 3056 2644
rect 3108 2632 3114 2644
rect 9398 2632 9404 2644
rect 3108 2604 9404 2632
rect 3108 2592 3114 2604
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 12069 2635 12127 2641
rect 12069 2601 12081 2635
rect 12115 2632 12127 2635
rect 12710 2632 12716 2644
rect 12115 2604 12716 2632
rect 12115 2601 12127 2604
rect 12069 2595 12127 2601
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 13354 2632 13360 2644
rect 13315 2604 13360 2632
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 13817 2635 13875 2641
rect 13817 2601 13829 2635
rect 13863 2632 13875 2635
rect 14274 2632 14280 2644
rect 13863 2604 14280 2632
rect 13863 2601 13875 2604
rect 13817 2595 13875 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 17310 2592 17316 2644
rect 17368 2632 17374 2644
rect 17497 2635 17555 2641
rect 17497 2632 17509 2635
rect 17368 2604 17509 2632
rect 17368 2592 17374 2604
rect 17497 2601 17509 2604
rect 17543 2601 17555 2635
rect 17497 2595 17555 2601
rect 25685 2635 25743 2641
rect 25685 2601 25697 2635
rect 25731 2632 25743 2635
rect 25774 2632 25780 2644
rect 25731 2604 25780 2632
rect 25731 2601 25743 2604
rect 25685 2595 25743 2601
rect 25774 2592 25780 2604
rect 25832 2592 25838 2644
rect 26145 2635 26203 2641
rect 26145 2601 26157 2635
rect 26191 2632 26203 2635
rect 26510 2632 26516 2644
rect 26191 2604 26516 2632
rect 26191 2601 26203 2604
rect 26145 2595 26203 2601
rect 26510 2592 26516 2604
rect 26568 2592 26574 2644
rect 10042 2496 10048 2508
rect 10003 2468 10048 2496
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 10134 2456 10140 2508
rect 10192 2496 10198 2508
rect 11609 2499 11667 2505
rect 10192 2468 10237 2496
rect 10192 2456 10198 2468
rect 11609 2465 11621 2499
rect 11655 2496 11667 2499
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11655 2468 11713 2496
rect 11655 2465 11667 2468
rect 11609 2459 11667 2465
rect 11701 2465 11713 2468
rect 11747 2496 11759 2499
rect 13372 2496 13400 2592
rect 23474 2524 23480 2576
rect 23532 2564 23538 2576
rect 23661 2567 23719 2573
rect 23661 2564 23673 2567
rect 23532 2536 23673 2564
rect 23532 2524 23538 2536
rect 23661 2533 23673 2536
rect 23707 2533 23719 2567
rect 23661 2527 23719 2533
rect 23768 2536 24256 2564
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 11747 2468 13461 2496
rect 11747 2465 11759 2468
rect 11701 2459 11759 2465
rect 13449 2465 13461 2468
rect 13495 2465 13507 2499
rect 23768 2496 23796 2536
rect 13449 2459 13507 2465
rect 23492 2468 23796 2496
rect 9950 2428 9956 2440
rect 9911 2400 9956 2428
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 12066 2428 12072 2440
rect 11931 2400 12072 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 13630 2428 13636 2440
rect 13591 2400 13636 2428
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 14458 2428 14464 2440
rect 14419 2400 14464 2428
rect 14458 2388 14464 2400
rect 14516 2388 14522 2440
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17460 2400 17601 2428
rect 17460 2388 17466 2400
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 21818 2428 21824 2440
rect 21779 2400 21824 2428
rect 17589 2391 17647 2397
rect 21818 2388 21824 2400
rect 21876 2388 21882 2440
rect 22002 2428 22008 2440
rect 21963 2400 22008 2428
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 23492 2437 23520 2468
rect 23842 2456 23848 2508
rect 23900 2496 23906 2508
rect 23900 2468 24072 2496
rect 23900 2456 23906 2468
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 23750 2388 23756 2440
rect 23808 2428 23814 2440
rect 24044 2437 24072 2468
rect 24029 2431 24087 2437
rect 23808 2400 23853 2428
rect 23808 2388 23814 2400
rect 24029 2397 24041 2431
rect 24075 2397 24087 2431
rect 24029 2391 24087 2397
rect 13648 2292 13676 2388
rect 22189 2363 22247 2369
rect 22189 2329 22201 2363
rect 22235 2360 22247 2363
rect 23566 2360 23572 2372
rect 22235 2332 23572 2360
rect 22235 2329 22247 2332
rect 22189 2323 22247 2329
rect 23566 2320 23572 2332
rect 23624 2360 23630 2372
rect 24228 2369 24256 2536
rect 25222 2524 25228 2576
rect 25280 2564 25286 2576
rect 26050 2564 26056 2576
rect 25280 2536 26056 2564
rect 25280 2524 25286 2536
rect 25608 2437 25636 2536
rect 26050 2524 26056 2536
rect 26108 2524 26114 2576
rect 26068 2437 26096 2524
rect 25593 2431 25651 2437
rect 25593 2397 25605 2431
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 26053 2431 26111 2437
rect 26053 2397 26065 2431
rect 26099 2397 26111 2431
rect 26053 2391 26111 2397
rect 23845 2363 23903 2369
rect 23845 2360 23857 2363
rect 23624 2332 23857 2360
rect 23624 2320 23630 2332
rect 23845 2329 23857 2332
rect 23891 2329 23903 2363
rect 23845 2323 23903 2329
rect 24213 2363 24271 2369
rect 24213 2329 24225 2363
rect 24259 2360 24271 2363
rect 25869 2363 25927 2369
rect 25869 2360 25881 2363
rect 24259 2332 25881 2360
rect 24259 2329 24271 2332
rect 24213 2323 24271 2329
rect 25869 2329 25881 2332
rect 25915 2360 25927 2363
rect 26142 2360 26148 2372
rect 25915 2332 26148 2360
rect 25915 2329 25927 2332
rect 25869 2323 25927 2329
rect 26142 2320 26148 2332
rect 26200 2320 26206 2372
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13648 2264 14289 2292
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 23293 2295 23351 2301
rect 23293 2261 23305 2295
rect 23339 2292 23351 2295
rect 23658 2292 23664 2304
rect 23339 2264 23664 2292
rect 23339 2261 23351 2264
rect 23293 2255 23351 2261
rect 23658 2252 23664 2264
rect 23716 2252 23722 2304
rect 1104 2202 29440 2224
rect 1104 2150 10395 2202
rect 10447 2150 10459 2202
rect 10511 2150 10523 2202
rect 10575 2150 10587 2202
rect 10639 2150 10651 2202
rect 10703 2150 19840 2202
rect 19892 2150 19904 2202
rect 19956 2150 19968 2202
rect 20020 2150 20032 2202
rect 20084 2150 20096 2202
rect 20148 2150 29440 2202
rect 1104 2128 29440 2150
rect 3326 1300 3332 1352
rect 3384 1340 3390 1352
rect 6546 1340 6552 1352
rect 3384 1312 6552 1340
rect 3384 1300 3390 1312
rect 6546 1300 6552 1312
rect 6604 1300 6610 1352
rect 8570 1300 8576 1352
rect 8628 1340 8634 1352
rect 26234 1340 26240 1352
rect 8628 1312 26240 1340
rect 8628 1300 8634 1312
rect 26234 1300 26240 1312
rect 26292 1300 26298 1352
<< via1 >>
rect 4068 30540 4120 30592
rect 19616 30540 19668 30592
rect 10395 30438 10447 30490
rect 10459 30438 10511 30490
rect 10523 30438 10575 30490
rect 10587 30438 10639 30490
rect 10651 30438 10703 30490
rect 19840 30438 19892 30490
rect 19904 30438 19956 30490
rect 19968 30438 20020 30490
rect 20032 30438 20084 30490
rect 20096 30438 20148 30490
rect 3976 30336 4028 30388
rect 22192 30336 22244 30388
rect 11152 30200 11204 30252
rect 14924 30243 14976 30252
rect 14924 30209 14933 30243
rect 14933 30209 14967 30243
rect 14967 30209 14976 30243
rect 14924 30200 14976 30209
rect 18604 30200 18656 30252
rect 26240 30268 26292 30320
rect 20352 30200 20404 30252
rect 20720 30243 20772 30252
rect 20720 30209 20729 30243
rect 20729 30209 20763 30243
rect 20763 30209 20772 30243
rect 20720 30200 20772 30209
rect 22008 30243 22060 30252
rect 22008 30209 22057 30243
rect 22057 30209 22060 30243
rect 22008 30200 22060 30209
rect 22468 30243 22520 30252
rect 18696 30132 18748 30184
rect 19064 30064 19116 30116
rect 12256 29996 12308 30048
rect 14648 29996 14700 30048
rect 19340 30039 19392 30048
rect 19340 30005 19349 30039
rect 19349 30005 19383 30039
rect 19383 30005 19392 30039
rect 19340 29996 19392 30005
rect 19616 29996 19668 30048
rect 21732 30132 21784 30184
rect 21088 30064 21140 30116
rect 20536 30039 20588 30048
rect 20536 30005 20545 30039
rect 20545 30005 20579 30039
rect 20579 30005 20588 30039
rect 20536 29996 20588 30005
rect 21732 29996 21784 30048
rect 22468 30209 22477 30243
rect 22477 30209 22511 30243
rect 22511 30209 22520 30243
rect 22468 30200 22520 30209
rect 22836 30243 22888 30252
rect 22836 30209 22845 30243
rect 22845 30209 22879 30243
rect 22879 30209 22888 30243
rect 22836 30200 22888 30209
rect 22652 30039 22704 30048
rect 22652 30005 22661 30039
rect 22661 30005 22695 30039
rect 22695 30005 22704 30039
rect 22652 29996 22704 30005
rect 23112 29996 23164 30048
rect 5672 29894 5724 29946
rect 5736 29894 5788 29946
rect 5800 29894 5852 29946
rect 5864 29894 5916 29946
rect 5928 29894 5980 29946
rect 15118 29894 15170 29946
rect 15182 29894 15234 29946
rect 15246 29894 15298 29946
rect 15310 29894 15362 29946
rect 15374 29894 15426 29946
rect 24563 29894 24615 29946
rect 24627 29894 24679 29946
rect 24691 29894 24743 29946
rect 24755 29894 24807 29946
rect 24819 29894 24871 29946
rect 4068 29792 4120 29844
rect 17040 29792 17092 29844
rect 3240 29656 3292 29708
rect 4620 29699 4672 29708
rect 4620 29665 4629 29699
rect 4629 29665 4663 29699
rect 4663 29665 4672 29699
rect 4620 29656 4672 29665
rect 7104 29656 7156 29708
rect 12532 29656 12584 29708
rect 15660 29656 15712 29708
rect 17960 29656 18012 29708
rect 18696 29724 18748 29776
rect 5172 29588 5224 29640
rect 11152 29631 11204 29640
rect 11152 29597 11161 29631
rect 11161 29597 11195 29631
rect 11195 29597 11204 29631
rect 11152 29588 11204 29597
rect 13636 29588 13688 29640
rect 26148 29792 26200 29844
rect 19616 29767 19668 29776
rect 19616 29733 19625 29767
rect 19625 29733 19659 29767
rect 19659 29733 19668 29767
rect 19616 29724 19668 29733
rect 5632 29520 5684 29572
rect 9312 29563 9364 29572
rect 9312 29529 9321 29563
rect 9321 29529 9355 29563
rect 9355 29529 9364 29563
rect 9312 29520 9364 29529
rect 10324 29520 10376 29572
rect 6920 29495 6972 29504
rect 6920 29461 6929 29495
rect 6929 29461 6963 29495
rect 6963 29461 6972 29495
rect 6920 29452 6972 29461
rect 7380 29452 7432 29504
rect 10784 29495 10836 29504
rect 10784 29461 10793 29495
rect 10793 29461 10827 29495
rect 10827 29461 10836 29495
rect 10784 29452 10836 29461
rect 10968 29495 11020 29504
rect 10968 29461 10977 29495
rect 10977 29461 11011 29495
rect 11011 29461 11020 29495
rect 10968 29452 11020 29461
rect 12256 29520 12308 29572
rect 12992 29563 13044 29572
rect 12992 29529 13001 29563
rect 13001 29529 13035 29563
rect 13035 29529 13044 29563
rect 12992 29520 13044 29529
rect 14648 29520 14700 29572
rect 15384 29520 15436 29572
rect 11612 29452 11664 29504
rect 14372 29452 14424 29504
rect 15844 29452 15896 29504
rect 18144 29452 18196 29504
rect 18972 29631 19024 29640
rect 18972 29597 18981 29631
rect 18981 29597 19015 29631
rect 19015 29597 19024 29631
rect 20352 29656 20404 29708
rect 21088 29699 21140 29708
rect 21088 29665 21097 29699
rect 21097 29665 21131 29699
rect 21131 29665 21140 29699
rect 21088 29656 21140 29665
rect 18972 29588 19024 29597
rect 21732 29588 21784 29640
rect 19064 29520 19116 29572
rect 20536 29520 20588 29572
rect 22100 29563 22152 29572
rect 22100 29529 22109 29563
rect 22109 29529 22143 29563
rect 22143 29529 22152 29563
rect 22100 29520 22152 29529
rect 23112 29520 23164 29572
rect 22928 29452 22980 29504
rect 10395 29350 10447 29402
rect 10459 29350 10511 29402
rect 10523 29350 10575 29402
rect 10587 29350 10639 29402
rect 10651 29350 10703 29402
rect 19840 29350 19892 29402
rect 19904 29350 19956 29402
rect 19968 29350 20020 29402
rect 20032 29350 20084 29402
rect 20096 29350 20148 29402
rect 5632 29291 5684 29300
rect 5632 29257 5641 29291
rect 5641 29257 5675 29291
rect 5675 29257 5684 29291
rect 5632 29248 5684 29257
rect 9312 29291 9364 29300
rect 9312 29257 9321 29291
rect 9321 29257 9355 29291
rect 9355 29257 9364 29291
rect 9312 29248 9364 29257
rect 10324 29248 10376 29300
rect 12532 29248 12584 29300
rect 5172 29180 5224 29232
rect 3976 29112 4028 29164
rect 6920 29180 6972 29232
rect 10784 29180 10836 29232
rect 12992 29180 13044 29232
rect 15384 29248 15436 29300
rect 18604 29291 18656 29300
rect 5908 29155 5960 29164
rect 5908 29121 5917 29155
rect 5917 29121 5951 29155
rect 5951 29121 5960 29155
rect 5908 29112 5960 29121
rect 4160 28908 4212 28960
rect 6092 29019 6144 29028
rect 6092 28985 6101 29019
rect 6101 28985 6135 29019
rect 6135 28985 6144 29019
rect 7104 29044 7156 29096
rect 10968 29112 11020 29164
rect 11612 29155 11664 29164
rect 10140 29087 10192 29096
rect 10140 29053 10149 29087
rect 10149 29053 10183 29087
rect 10183 29053 10192 29087
rect 10140 29044 10192 29053
rect 10876 29044 10928 29096
rect 11612 29121 11621 29155
rect 11621 29121 11655 29155
rect 11655 29121 11664 29155
rect 11612 29112 11664 29121
rect 6092 28976 6144 28985
rect 12532 29112 12584 29164
rect 12900 29155 12952 29164
rect 12900 29121 12909 29155
rect 12909 29121 12943 29155
rect 12943 29121 12952 29155
rect 12900 29112 12952 29121
rect 12164 29044 12216 29096
rect 13268 29155 13320 29164
rect 13268 29121 13282 29155
rect 13282 29121 13316 29155
rect 13316 29121 13320 29155
rect 14372 29180 14424 29232
rect 18604 29257 18613 29291
rect 18613 29257 18647 29291
rect 18647 29257 18656 29291
rect 18604 29248 18656 29257
rect 20720 29248 20772 29300
rect 22836 29291 22888 29300
rect 22836 29257 22845 29291
rect 22845 29257 22879 29291
rect 22879 29257 22888 29291
rect 22836 29248 22888 29257
rect 22192 29223 22244 29232
rect 15936 29155 15988 29164
rect 13268 29112 13320 29121
rect 15936 29121 15945 29155
rect 15945 29121 15979 29155
rect 15979 29121 15988 29155
rect 15936 29112 15988 29121
rect 13636 29044 13688 29096
rect 14096 29044 14148 29096
rect 15660 29044 15712 29096
rect 17408 29112 17460 29164
rect 19340 29112 19392 29164
rect 22192 29189 22201 29223
rect 22201 29189 22235 29223
rect 22235 29189 22244 29223
rect 22928 29223 22980 29232
rect 22192 29180 22244 29189
rect 22928 29189 22937 29223
rect 22937 29189 22971 29223
rect 22971 29189 22980 29223
rect 22928 29180 22980 29189
rect 20260 29112 20312 29164
rect 20352 29112 20404 29164
rect 20536 29112 20588 29164
rect 20720 29155 20772 29164
rect 20720 29121 20729 29155
rect 20729 29121 20763 29155
rect 20763 29121 20772 29155
rect 20720 29112 20772 29121
rect 22008 29155 22060 29164
rect 22008 29121 22057 29155
rect 22057 29121 22060 29155
rect 22008 29112 22060 29121
rect 22192 29044 22244 29096
rect 18236 28976 18288 29028
rect 22100 28976 22152 29028
rect 22560 29112 22612 29164
rect 22744 29112 22796 29164
rect 24400 29112 24452 29164
rect 23848 28976 23900 29028
rect 13728 28908 13780 28960
rect 19248 28908 19300 28960
rect 20812 28908 20864 28960
rect 23940 28908 23992 28960
rect 25872 28908 25924 28960
rect 5672 28806 5724 28858
rect 5736 28806 5788 28858
rect 5800 28806 5852 28858
rect 5864 28806 5916 28858
rect 5928 28806 5980 28858
rect 15118 28806 15170 28858
rect 15182 28806 15234 28858
rect 15246 28806 15298 28858
rect 15310 28806 15362 28858
rect 15374 28806 15426 28858
rect 24563 28806 24615 28858
rect 24627 28806 24679 28858
rect 24691 28806 24743 28858
rect 24755 28806 24807 28858
rect 24819 28806 24871 28858
rect 3976 28747 4028 28756
rect 3976 28713 3985 28747
rect 3985 28713 4019 28747
rect 4019 28713 4028 28747
rect 3976 28704 4028 28713
rect 4344 28704 4396 28756
rect 6092 28704 6144 28756
rect 13728 28747 13780 28756
rect 13728 28713 13737 28747
rect 13737 28713 13771 28747
rect 13771 28713 13780 28747
rect 13728 28704 13780 28713
rect 14924 28704 14976 28756
rect 15936 28704 15988 28756
rect 17040 28704 17092 28756
rect 18052 28704 18104 28756
rect 25228 28704 25280 28756
rect 5172 28611 5224 28620
rect 5172 28577 5181 28611
rect 5181 28577 5215 28611
rect 5215 28577 5224 28611
rect 5172 28568 5224 28577
rect 4160 28543 4212 28552
rect 4160 28509 4169 28543
rect 4169 28509 4203 28543
rect 4203 28509 4212 28543
rect 4160 28500 4212 28509
rect 4252 28543 4304 28552
rect 4252 28509 4261 28543
rect 4261 28509 4295 28543
rect 4295 28509 4304 28543
rect 4528 28543 4580 28552
rect 4252 28500 4304 28509
rect 4528 28509 4537 28543
rect 4537 28509 4571 28543
rect 4571 28509 4580 28543
rect 4528 28500 4580 28509
rect 15476 28636 15528 28688
rect 16212 28636 16264 28688
rect 17408 28679 17460 28688
rect 17408 28645 17417 28679
rect 17417 28645 17451 28679
rect 17451 28645 17460 28679
rect 17408 28636 17460 28645
rect 7380 28611 7432 28620
rect 7380 28577 7389 28611
rect 7389 28577 7423 28611
rect 7423 28577 7432 28611
rect 7380 28568 7432 28577
rect 7012 28543 7064 28552
rect 7012 28509 7021 28543
rect 7021 28509 7055 28543
rect 7055 28509 7064 28543
rect 7012 28500 7064 28509
rect 8576 28543 8628 28552
rect 6000 28364 6052 28416
rect 8576 28509 8585 28543
rect 8585 28509 8619 28543
rect 8619 28509 8628 28543
rect 8576 28500 8628 28509
rect 10232 28543 10284 28552
rect 10232 28509 10241 28543
rect 10241 28509 10275 28543
rect 10275 28509 10284 28543
rect 10232 28500 10284 28509
rect 11152 28568 11204 28620
rect 11244 28568 11296 28620
rect 11980 28568 12032 28620
rect 18696 28568 18748 28620
rect 29828 28636 29880 28688
rect 8392 28407 8444 28416
rect 8392 28373 8401 28407
rect 8401 28373 8435 28407
rect 8435 28373 8444 28407
rect 8392 28364 8444 28373
rect 9772 28364 9824 28416
rect 12900 28500 12952 28552
rect 13268 28500 13320 28552
rect 15476 28500 15528 28552
rect 17868 28543 17920 28552
rect 11152 28407 11204 28416
rect 11152 28373 11161 28407
rect 11161 28373 11195 28407
rect 11195 28373 11204 28407
rect 13912 28432 13964 28484
rect 17868 28509 17877 28543
rect 17877 28509 17911 28543
rect 17911 28509 17920 28543
rect 17868 28500 17920 28509
rect 18052 28500 18104 28552
rect 18972 28500 19024 28552
rect 18236 28432 18288 28484
rect 20720 28432 20772 28484
rect 21732 28432 21784 28484
rect 22468 28568 22520 28620
rect 22284 28543 22336 28552
rect 22284 28509 22333 28543
rect 22333 28509 22336 28543
rect 22284 28500 22336 28509
rect 23204 28543 23256 28552
rect 23204 28509 23218 28543
rect 23218 28509 23252 28543
rect 23252 28509 23256 28543
rect 23204 28500 23256 28509
rect 23388 28500 23440 28552
rect 24400 28543 24452 28552
rect 24400 28509 24409 28543
rect 24409 28509 24443 28543
rect 24443 28509 24452 28543
rect 24400 28500 24452 28509
rect 11152 28364 11204 28373
rect 14004 28364 14056 28416
rect 15936 28407 15988 28416
rect 15936 28373 15945 28407
rect 15945 28373 15979 28407
rect 15979 28373 15988 28407
rect 15936 28364 15988 28373
rect 22560 28475 22612 28484
rect 22560 28441 22569 28475
rect 22569 28441 22603 28475
rect 22603 28441 22612 28475
rect 22560 28432 22612 28441
rect 22928 28432 22980 28484
rect 23664 28432 23716 28484
rect 22284 28364 22336 28416
rect 23204 28364 23256 28416
rect 23572 28364 23624 28416
rect 24032 28364 24084 28416
rect 24676 28407 24728 28416
rect 24676 28373 24685 28407
rect 24685 28373 24719 28407
rect 24719 28373 24728 28407
rect 24676 28364 24728 28373
rect 10395 28262 10447 28314
rect 10459 28262 10511 28314
rect 10523 28262 10575 28314
rect 10587 28262 10639 28314
rect 10651 28262 10703 28314
rect 19840 28262 19892 28314
rect 19904 28262 19956 28314
rect 19968 28262 20020 28314
rect 20032 28262 20084 28314
rect 20096 28262 20148 28314
rect 4528 28160 4580 28212
rect 7012 28203 7064 28212
rect 7012 28169 7021 28203
rect 7021 28169 7055 28203
rect 7055 28169 7064 28203
rect 7012 28160 7064 28169
rect 10048 28160 10100 28212
rect 19248 28160 19300 28212
rect 20720 28160 20772 28212
rect 22468 28203 22520 28212
rect 22468 28169 22477 28203
rect 22477 28169 22511 28203
rect 22511 28169 22520 28203
rect 22468 28160 22520 28169
rect 8392 28092 8444 28144
rect 9772 28135 9824 28144
rect 9772 28101 9781 28135
rect 9781 28101 9815 28135
rect 9815 28101 9824 28135
rect 9772 28092 9824 28101
rect 11152 28092 11204 28144
rect 13820 28092 13872 28144
rect 4252 27956 4304 28008
rect 7104 27999 7156 28008
rect 7104 27965 7113 27999
rect 7113 27965 7147 27999
rect 7147 27965 7156 27999
rect 7104 27956 7156 27965
rect 6552 27863 6604 27872
rect 6552 27829 6561 27863
rect 6561 27829 6595 27863
rect 6595 27829 6604 27863
rect 6552 27820 6604 27829
rect 12440 28067 12492 28076
rect 12440 28033 12449 28067
rect 12449 28033 12483 28067
rect 12483 28033 12492 28067
rect 12440 28024 12492 28033
rect 14096 28024 14148 28076
rect 9036 27999 9088 28008
rect 9036 27965 9045 27999
rect 9045 27965 9079 27999
rect 9079 27965 9088 27999
rect 9036 27956 9088 27965
rect 9312 27999 9364 28008
rect 9312 27965 9321 27999
rect 9321 27965 9355 27999
rect 9355 27965 9364 27999
rect 9312 27956 9364 27965
rect 14556 27888 14608 27940
rect 15936 28092 15988 28144
rect 23388 28160 23440 28212
rect 23664 28160 23716 28212
rect 28540 28160 28592 28212
rect 23572 28135 23624 28144
rect 16396 28024 16448 28076
rect 17960 28067 18012 28076
rect 17960 28033 17969 28067
rect 17969 28033 18003 28067
rect 18003 28033 18012 28067
rect 17960 28024 18012 28033
rect 19432 28024 19484 28076
rect 20260 28067 20312 28076
rect 20260 28033 20269 28067
rect 20269 28033 20303 28067
rect 20303 28033 20312 28067
rect 20260 28024 20312 28033
rect 16580 27956 16632 28008
rect 17592 27956 17644 28008
rect 18328 27956 18380 28008
rect 8944 27820 8996 27872
rect 12624 27863 12676 27872
rect 12624 27829 12633 27863
rect 12633 27829 12667 27863
rect 12667 27829 12676 27863
rect 12624 27820 12676 27829
rect 14464 27863 14516 27872
rect 14464 27829 14473 27863
rect 14473 27829 14507 27863
rect 14507 27829 14516 27863
rect 14464 27820 14516 27829
rect 15752 27820 15804 27872
rect 22192 28024 22244 28076
rect 23572 28101 23581 28135
rect 23581 28101 23615 28135
rect 23615 28101 23624 28135
rect 23572 28092 23624 28101
rect 26792 28092 26844 28144
rect 24676 28024 24728 28076
rect 25228 28067 25280 28076
rect 25228 28033 25237 28067
rect 25237 28033 25271 28067
rect 25271 28033 25280 28067
rect 25228 28024 25280 28033
rect 25412 28067 25464 28076
rect 25412 28033 25421 28067
rect 25421 28033 25455 28067
rect 25455 28033 25464 28067
rect 25412 28024 25464 28033
rect 21272 27956 21324 28008
rect 21732 27956 21784 28008
rect 23664 27956 23716 28008
rect 21824 27888 21876 27940
rect 22468 27888 22520 27940
rect 25412 27888 25464 27940
rect 22008 27863 22060 27872
rect 22008 27829 22017 27863
rect 22017 27829 22051 27863
rect 22051 27829 22060 27863
rect 22008 27820 22060 27829
rect 22284 27820 22336 27872
rect 23388 27820 23440 27872
rect 25780 27863 25832 27872
rect 25780 27829 25789 27863
rect 25789 27829 25823 27863
rect 25823 27829 25832 27863
rect 25780 27820 25832 27829
rect 5672 27718 5724 27770
rect 5736 27718 5788 27770
rect 5800 27718 5852 27770
rect 5864 27718 5916 27770
rect 5928 27718 5980 27770
rect 15118 27718 15170 27770
rect 15182 27718 15234 27770
rect 15246 27718 15298 27770
rect 15310 27718 15362 27770
rect 15374 27718 15426 27770
rect 24563 27718 24615 27770
rect 24627 27718 24679 27770
rect 24691 27718 24743 27770
rect 24755 27718 24807 27770
rect 24819 27718 24871 27770
rect 4068 27616 4120 27668
rect 10232 27659 10284 27668
rect 4344 27591 4396 27600
rect 4344 27557 4353 27591
rect 4353 27557 4387 27591
rect 4387 27557 4396 27591
rect 4344 27548 4396 27557
rect 8576 27548 8628 27600
rect 9036 27548 9088 27600
rect 10232 27625 10241 27659
rect 10241 27625 10275 27659
rect 10275 27625 10284 27659
rect 10232 27616 10284 27625
rect 16304 27616 16356 27668
rect 17224 27616 17276 27668
rect 17776 27616 17828 27668
rect 4252 27480 4304 27532
rect 8944 27523 8996 27532
rect 8944 27489 8953 27523
rect 8953 27489 8987 27523
rect 8987 27489 8996 27523
rect 8944 27480 8996 27489
rect 9312 27480 9364 27532
rect 11336 27548 11388 27600
rect 12348 27548 12400 27600
rect 4160 27455 4212 27464
rect 4160 27421 4169 27455
rect 4169 27421 4203 27455
rect 4203 27421 4212 27455
rect 4436 27455 4488 27464
rect 4160 27412 4212 27421
rect 4436 27421 4445 27455
rect 4445 27421 4479 27455
rect 4479 27421 4488 27455
rect 4436 27412 4488 27421
rect 7840 27412 7892 27464
rect 8300 27412 8352 27464
rect 9404 27412 9456 27464
rect 10784 27480 10836 27532
rect 11244 27480 11296 27532
rect 12716 27480 12768 27532
rect 10876 27344 10928 27396
rect 13636 27455 13688 27464
rect 13636 27421 13645 27455
rect 13645 27421 13679 27455
rect 13679 27421 13688 27455
rect 14096 27455 14148 27464
rect 13636 27412 13688 27421
rect 14096 27421 14105 27455
rect 14105 27421 14139 27455
rect 14139 27421 14148 27455
rect 14096 27412 14148 27421
rect 14556 27455 14608 27464
rect 3884 27319 3936 27328
rect 3884 27285 3893 27319
rect 3893 27285 3927 27319
rect 3927 27285 3936 27319
rect 3884 27276 3936 27285
rect 8208 27319 8260 27328
rect 8208 27285 8217 27319
rect 8217 27285 8251 27319
rect 8251 27285 8260 27319
rect 8208 27276 8260 27285
rect 10048 27276 10100 27328
rect 11612 27276 11664 27328
rect 12624 27344 12676 27396
rect 13360 27387 13412 27396
rect 13360 27353 13369 27387
rect 13369 27353 13403 27387
rect 13403 27353 13412 27387
rect 13360 27344 13412 27353
rect 12992 27276 13044 27328
rect 13084 27276 13136 27328
rect 13728 27344 13780 27396
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 15660 27455 15712 27464
rect 15660 27421 15669 27455
rect 15669 27421 15703 27455
rect 15703 27421 15712 27455
rect 15660 27412 15712 27421
rect 18696 27548 18748 27600
rect 19432 27616 19484 27668
rect 21548 27616 21600 27668
rect 23664 27659 23716 27668
rect 23664 27625 23673 27659
rect 23673 27625 23707 27659
rect 23707 27625 23716 27659
rect 23664 27616 23716 27625
rect 25780 27616 25832 27668
rect 19708 27548 19760 27600
rect 22008 27548 22060 27600
rect 22560 27548 22612 27600
rect 22928 27548 22980 27600
rect 23296 27591 23348 27600
rect 23296 27557 23305 27591
rect 23305 27557 23339 27591
rect 23339 27557 23348 27591
rect 23296 27548 23348 27557
rect 26792 27591 26844 27600
rect 26792 27557 26801 27591
rect 26801 27557 26835 27591
rect 26835 27557 26844 27591
rect 26792 27548 26844 27557
rect 18052 27412 18104 27464
rect 16672 27344 16724 27396
rect 17868 27344 17920 27396
rect 18328 27480 18380 27532
rect 18420 27412 18472 27464
rect 18696 27412 18748 27464
rect 18972 27412 19024 27464
rect 19248 27412 19300 27464
rect 16856 27276 16908 27328
rect 18144 27276 18196 27328
rect 19064 27276 19116 27328
rect 19340 27276 19392 27328
rect 22744 27455 22796 27464
rect 22744 27421 22753 27455
rect 22753 27421 22787 27455
rect 22787 27421 22796 27455
rect 22744 27412 22796 27421
rect 23020 27455 23072 27464
rect 23020 27421 23029 27455
rect 23029 27421 23063 27455
rect 23063 27421 23072 27455
rect 23020 27412 23072 27421
rect 23664 27480 23716 27532
rect 24032 27480 24084 27532
rect 23480 27455 23532 27464
rect 23480 27421 23489 27455
rect 23489 27421 23523 27455
rect 23523 27421 23532 27455
rect 23480 27412 23532 27421
rect 23572 27412 23624 27464
rect 21456 27344 21508 27396
rect 22560 27344 22612 27396
rect 22836 27344 22888 27396
rect 20168 27319 20220 27328
rect 20168 27285 20177 27319
rect 20177 27285 20211 27319
rect 20211 27285 20220 27319
rect 20168 27276 20220 27285
rect 20352 27319 20404 27328
rect 20352 27285 20361 27319
rect 20361 27285 20395 27319
rect 20395 27285 20404 27319
rect 20352 27276 20404 27285
rect 24400 27344 24452 27396
rect 24952 27412 25004 27464
rect 25872 27344 25924 27396
rect 24032 27319 24084 27328
rect 24032 27285 24041 27319
rect 24041 27285 24075 27319
rect 24075 27285 24084 27319
rect 24032 27276 24084 27285
rect 25688 27276 25740 27328
rect 10395 27174 10447 27226
rect 10459 27174 10511 27226
rect 10523 27174 10575 27226
rect 10587 27174 10639 27226
rect 10651 27174 10703 27226
rect 19840 27174 19892 27226
rect 19904 27174 19956 27226
rect 19968 27174 20020 27226
rect 20032 27174 20084 27226
rect 20096 27174 20148 27226
rect 4252 27072 4304 27124
rect 4436 27115 4488 27124
rect 4436 27081 4445 27115
rect 4445 27081 4479 27115
rect 4479 27081 4488 27115
rect 4436 27072 4488 27081
rect 3884 27004 3936 27056
rect 3332 26936 3384 26988
rect 8208 27004 8260 27056
rect 4988 26936 5040 26988
rect 2688 26868 2740 26920
rect 6000 26936 6052 26988
rect 6552 26936 6604 26988
rect 6644 26868 6696 26920
rect 7104 26911 7156 26920
rect 7104 26877 7113 26911
rect 7113 26877 7147 26911
rect 7147 26877 7156 26911
rect 9312 26936 9364 26988
rect 9404 26979 9456 26988
rect 9404 26945 9413 26979
rect 9413 26945 9447 26979
rect 9447 26945 9456 26979
rect 9404 26936 9456 26945
rect 10968 27004 11020 27056
rect 11244 27072 11296 27124
rect 12624 27072 12676 27124
rect 11612 27004 11664 27056
rect 12992 27072 13044 27124
rect 14464 27072 14516 27124
rect 14556 27072 14608 27124
rect 13360 27004 13412 27056
rect 10324 26936 10376 26988
rect 10876 26936 10928 26988
rect 11060 26936 11112 26988
rect 12164 26936 12216 26988
rect 7104 26868 7156 26877
rect 12716 26936 12768 26988
rect 13544 26979 13596 26988
rect 13544 26945 13553 26979
rect 13553 26945 13587 26979
rect 13587 26945 13596 26979
rect 13544 26936 13596 26945
rect 14096 26936 14148 26988
rect 14464 26979 14516 26988
rect 14464 26945 14473 26979
rect 14473 26945 14507 26979
rect 14507 26945 14516 26979
rect 14924 27072 14976 27124
rect 15752 27004 15804 27056
rect 16304 27072 16356 27124
rect 21456 27072 21508 27124
rect 18512 27047 18564 27056
rect 18512 27013 18521 27047
rect 18521 27013 18555 27047
rect 18555 27013 18564 27047
rect 18512 27004 18564 27013
rect 18788 27004 18840 27056
rect 19340 27004 19392 27056
rect 23020 27072 23072 27124
rect 23480 27072 23532 27124
rect 24492 27072 24544 27124
rect 25872 27115 25924 27124
rect 25872 27081 25881 27115
rect 25881 27081 25915 27115
rect 25915 27081 25924 27115
rect 25872 27072 25924 27081
rect 23296 27004 23348 27056
rect 24032 27004 24084 27056
rect 14464 26936 14516 26945
rect 4068 26800 4120 26852
rect 4344 26732 4396 26784
rect 5540 26732 5592 26784
rect 6092 26775 6144 26784
rect 6092 26741 6101 26775
rect 6101 26741 6135 26775
rect 6135 26741 6144 26775
rect 6092 26732 6144 26741
rect 6460 26775 6512 26784
rect 6460 26741 6469 26775
rect 6469 26741 6503 26775
rect 6503 26741 6512 26775
rect 6460 26732 6512 26741
rect 7564 26800 7616 26852
rect 14096 26800 14148 26852
rect 15200 26936 15252 26988
rect 16028 26936 16080 26988
rect 16672 26979 16724 26988
rect 16672 26945 16681 26979
rect 16681 26945 16715 26979
rect 16715 26945 16724 26979
rect 16672 26936 16724 26945
rect 16764 26936 16816 26988
rect 17224 26979 17276 26988
rect 17224 26945 17234 26979
rect 17234 26945 17268 26979
rect 17268 26945 17276 26979
rect 17224 26936 17276 26945
rect 17408 26979 17460 26988
rect 17408 26945 17417 26979
rect 17417 26945 17451 26979
rect 17451 26945 17460 26979
rect 17408 26936 17460 26945
rect 19156 26979 19208 26988
rect 17040 26911 17092 26920
rect 17040 26877 17049 26911
rect 17049 26877 17083 26911
rect 17083 26877 17092 26911
rect 17040 26868 17092 26877
rect 17132 26911 17184 26920
rect 17132 26877 17141 26911
rect 17141 26877 17175 26911
rect 17175 26877 17184 26911
rect 17132 26868 17184 26877
rect 18604 26911 18656 26920
rect 18604 26877 18613 26911
rect 18613 26877 18647 26911
rect 18647 26877 18656 26911
rect 18604 26868 18656 26877
rect 19156 26945 19164 26979
rect 19164 26945 19198 26979
rect 19198 26945 19208 26979
rect 19156 26936 19208 26945
rect 19524 26979 19576 26988
rect 19524 26945 19533 26979
rect 19533 26945 19567 26979
rect 19567 26945 19576 26979
rect 19524 26936 19576 26945
rect 21640 26936 21692 26988
rect 25688 26979 25740 26988
rect 25688 26945 25697 26979
rect 25697 26945 25731 26979
rect 25731 26945 25740 26979
rect 25688 26936 25740 26945
rect 14924 26800 14976 26852
rect 15752 26800 15804 26852
rect 10048 26732 10100 26784
rect 12532 26732 12584 26784
rect 14464 26732 14516 26784
rect 14832 26732 14884 26784
rect 15476 26775 15528 26784
rect 15476 26741 15485 26775
rect 15485 26741 15519 26775
rect 15519 26741 15528 26775
rect 15476 26732 15528 26741
rect 16488 26732 16540 26784
rect 18696 26800 18748 26852
rect 19064 26868 19116 26920
rect 19248 26911 19300 26920
rect 19248 26877 19257 26911
rect 19257 26877 19291 26911
rect 19291 26877 19300 26911
rect 19248 26868 19300 26877
rect 21272 26911 21324 26920
rect 18880 26800 18932 26852
rect 21272 26877 21281 26911
rect 21281 26877 21315 26911
rect 21315 26877 21324 26911
rect 21272 26868 21324 26877
rect 24952 26868 25004 26920
rect 25320 26911 25372 26920
rect 25320 26877 25329 26911
rect 25329 26877 25363 26911
rect 25363 26877 25372 26911
rect 25320 26868 25372 26877
rect 19524 26732 19576 26784
rect 22652 26732 22704 26784
rect 23020 26732 23072 26784
rect 24952 26732 25004 26784
rect 5672 26630 5724 26682
rect 5736 26630 5788 26682
rect 5800 26630 5852 26682
rect 5864 26630 5916 26682
rect 5928 26630 5980 26682
rect 15118 26630 15170 26682
rect 15182 26630 15234 26682
rect 15246 26630 15298 26682
rect 15310 26630 15362 26682
rect 15374 26630 15426 26682
rect 24563 26630 24615 26682
rect 24627 26630 24679 26682
rect 24691 26630 24743 26682
rect 24755 26630 24807 26682
rect 24819 26630 24871 26682
rect 4160 26528 4212 26580
rect 6644 26571 6696 26580
rect 6644 26537 6653 26571
rect 6653 26537 6687 26571
rect 6687 26537 6696 26571
rect 6644 26528 6696 26537
rect 8300 26571 8352 26580
rect 8300 26537 8309 26571
rect 8309 26537 8343 26571
rect 8343 26537 8352 26571
rect 8300 26528 8352 26537
rect 10324 26571 10376 26580
rect 10324 26537 10333 26571
rect 10333 26537 10367 26571
rect 10367 26537 10376 26571
rect 10324 26528 10376 26537
rect 10784 26571 10836 26580
rect 10784 26537 10793 26571
rect 10793 26537 10827 26571
rect 10827 26537 10836 26571
rect 10784 26528 10836 26537
rect 10968 26528 11020 26580
rect 13176 26528 13228 26580
rect 14556 26528 14608 26580
rect 15752 26528 15804 26580
rect 16396 26571 16448 26580
rect 16396 26537 16405 26571
rect 16405 26537 16439 26571
rect 16439 26537 16448 26571
rect 16396 26528 16448 26537
rect 21640 26571 21692 26580
rect 21640 26537 21649 26571
rect 21649 26537 21683 26571
rect 21683 26537 21692 26571
rect 21640 26528 21692 26537
rect 23572 26528 23624 26580
rect 25320 26528 25372 26580
rect 5172 26392 5224 26444
rect 11060 26392 11112 26444
rect 2780 26324 2832 26376
rect 3332 26324 3384 26376
rect 4896 26324 4948 26376
rect 5540 26367 5592 26376
rect 5540 26333 5574 26367
rect 5574 26333 5592 26367
rect 5540 26324 5592 26333
rect 8024 26367 8076 26376
rect 8024 26333 8033 26367
rect 8033 26333 8067 26367
rect 8067 26333 8076 26367
rect 8024 26324 8076 26333
rect 9588 26324 9640 26376
rect 10968 26256 11020 26308
rect 13544 26392 13596 26444
rect 13176 26367 13228 26376
rect 13176 26333 13185 26367
rect 13185 26333 13219 26367
rect 13219 26333 13228 26367
rect 13176 26324 13228 26333
rect 14924 26460 14976 26512
rect 15016 26460 15068 26512
rect 16488 26392 16540 26444
rect 16856 26435 16908 26444
rect 16856 26401 16865 26435
rect 16865 26401 16899 26435
rect 16899 26401 16908 26435
rect 16856 26392 16908 26401
rect 17224 26392 17276 26444
rect 18696 26460 18748 26512
rect 18788 26460 18840 26512
rect 19248 26503 19300 26512
rect 19248 26469 19257 26503
rect 19257 26469 19291 26503
rect 19291 26469 19300 26503
rect 19248 26460 19300 26469
rect 20168 26460 20220 26512
rect 18604 26392 18656 26444
rect 18972 26392 19024 26444
rect 19156 26392 19208 26444
rect 23940 26392 23992 26444
rect 14832 26367 14884 26376
rect 14832 26333 14841 26367
rect 14841 26333 14875 26367
rect 14875 26333 14884 26367
rect 14832 26324 14884 26333
rect 15476 26324 15528 26376
rect 17316 26324 17368 26376
rect 18144 26324 18196 26376
rect 18420 26324 18472 26376
rect 3056 26231 3108 26240
rect 3056 26197 3065 26231
rect 3065 26197 3099 26231
rect 3099 26197 3108 26231
rect 3056 26188 3108 26197
rect 7840 26231 7892 26240
rect 7840 26197 7849 26231
rect 7849 26197 7883 26231
rect 7883 26197 7892 26231
rect 7840 26188 7892 26197
rect 11428 26188 11480 26240
rect 12164 26231 12216 26240
rect 12164 26197 12173 26231
rect 12173 26197 12207 26231
rect 12207 26197 12216 26231
rect 14556 26299 14608 26308
rect 14556 26265 14565 26299
rect 14565 26265 14599 26299
rect 14599 26265 14608 26299
rect 14556 26256 14608 26265
rect 12164 26188 12216 26197
rect 14004 26188 14056 26240
rect 14464 26188 14516 26240
rect 15660 26256 15712 26308
rect 18696 26299 18748 26308
rect 18696 26265 18705 26299
rect 18705 26265 18739 26299
rect 18739 26265 18748 26299
rect 18696 26256 18748 26265
rect 19616 26299 19668 26308
rect 19616 26265 19625 26299
rect 19625 26265 19659 26299
rect 19659 26265 19668 26299
rect 19616 26256 19668 26265
rect 21732 26256 21784 26308
rect 22744 26324 22796 26376
rect 23204 26367 23256 26376
rect 23204 26333 23213 26367
rect 23213 26333 23247 26367
rect 23247 26333 23256 26367
rect 23204 26324 23256 26333
rect 23480 26367 23532 26376
rect 23480 26333 23489 26367
rect 23489 26333 23523 26367
rect 23523 26333 23532 26367
rect 23480 26324 23532 26333
rect 23664 26367 23716 26376
rect 23664 26333 23667 26367
rect 23667 26333 23716 26367
rect 23664 26324 23716 26333
rect 23112 26299 23164 26308
rect 23112 26265 23121 26299
rect 23121 26265 23155 26299
rect 23155 26265 23164 26299
rect 23112 26256 23164 26265
rect 14740 26188 14792 26240
rect 17868 26231 17920 26240
rect 17868 26197 17877 26231
rect 17877 26197 17911 26231
rect 17911 26197 17920 26231
rect 17868 26188 17920 26197
rect 18144 26188 18196 26240
rect 18880 26188 18932 26240
rect 10395 26086 10447 26138
rect 10459 26086 10511 26138
rect 10523 26086 10575 26138
rect 10587 26086 10639 26138
rect 10651 26086 10703 26138
rect 19840 26086 19892 26138
rect 19904 26086 19956 26138
rect 19968 26086 20020 26138
rect 20032 26086 20084 26138
rect 20096 26086 20148 26138
rect 5172 25984 5224 26036
rect 6000 25984 6052 26036
rect 1400 25848 1452 25900
rect 2688 25916 2740 25968
rect 2596 25848 2648 25900
rect 3884 25891 3936 25900
rect 3884 25857 3918 25891
rect 3918 25857 3936 25891
rect 3884 25848 3936 25857
rect 4896 25848 4948 25900
rect 6460 25848 6512 25900
rect 10140 25984 10192 26036
rect 15568 26027 15620 26036
rect 15568 25993 15577 26027
rect 15577 25993 15611 26027
rect 15611 25993 15620 26027
rect 15568 25984 15620 25993
rect 9220 25916 9272 25968
rect 12164 25916 12216 25968
rect 6736 25891 6788 25900
rect 6736 25857 6745 25891
rect 6745 25857 6779 25891
rect 6779 25857 6788 25891
rect 6736 25848 6788 25857
rect 6092 25712 6144 25764
rect 10876 25848 10928 25900
rect 11796 25891 11848 25900
rect 11796 25857 11805 25891
rect 11805 25857 11839 25891
rect 11839 25857 11848 25891
rect 15476 25916 15528 25968
rect 11796 25848 11848 25857
rect 12532 25848 12584 25900
rect 14464 25848 14516 25900
rect 14740 25848 14792 25900
rect 15016 25891 15068 25900
rect 15016 25857 15020 25891
rect 15020 25857 15054 25891
rect 15054 25857 15068 25891
rect 15016 25848 15068 25857
rect 15108 25891 15160 25900
rect 15108 25857 15117 25891
rect 15117 25857 15151 25891
rect 15151 25857 15160 25891
rect 15108 25848 15160 25857
rect 15752 25891 15804 25900
rect 9404 25823 9456 25832
rect 9404 25789 9413 25823
rect 9413 25789 9447 25823
rect 9447 25789 9456 25823
rect 9404 25780 9456 25789
rect 9588 25780 9640 25832
rect 10140 25780 10192 25832
rect 10968 25780 11020 25832
rect 11704 25823 11756 25832
rect 11704 25789 11713 25823
rect 11713 25789 11747 25823
rect 11747 25789 11756 25823
rect 11704 25780 11756 25789
rect 11336 25755 11388 25764
rect 11336 25721 11345 25755
rect 11345 25721 11379 25755
rect 11379 25721 11388 25755
rect 11336 25712 11388 25721
rect 14096 25780 14148 25832
rect 14832 25780 14884 25832
rect 15752 25857 15761 25891
rect 15761 25857 15795 25891
rect 15795 25857 15804 25891
rect 15752 25848 15804 25857
rect 17132 25984 17184 26036
rect 18788 25984 18840 26036
rect 19616 25984 19668 26036
rect 26240 25984 26292 26036
rect 17040 25916 17092 25968
rect 18144 25823 18196 25832
rect 13176 25755 13228 25764
rect 2780 25644 2832 25696
rect 3976 25644 4028 25696
rect 6920 25687 6972 25696
rect 6920 25653 6929 25687
rect 6929 25653 6963 25687
rect 6963 25653 6972 25687
rect 6920 25644 6972 25653
rect 7748 25644 7800 25696
rect 13176 25721 13185 25755
rect 13185 25721 13219 25755
rect 13219 25721 13228 25755
rect 13176 25712 13228 25721
rect 13820 25712 13872 25764
rect 14556 25712 14608 25764
rect 15016 25712 15068 25764
rect 18144 25789 18153 25823
rect 18153 25789 18187 25823
rect 18187 25789 18196 25823
rect 18144 25780 18196 25789
rect 12072 25644 12124 25696
rect 12256 25687 12308 25696
rect 12256 25653 12265 25687
rect 12265 25653 12299 25687
rect 12299 25653 12308 25687
rect 12256 25644 12308 25653
rect 12532 25687 12584 25696
rect 12532 25653 12541 25687
rect 12541 25653 12575 25687
rect 12575 25653 12584 25687
rect 12532 25644 12584 25653
rect 12992 25644 13044 25696
rect 13636 25644 13688 25696
rect 14372 25687 14424 25696
rect 14372 25653 14381 25687
rect 14381 25653 14415 25687
rect 14415 25653 14424 25687
rect 14372 25644 14424 25653
rect 16764 25687 16816 25696
rect 16764 25653 16773 25687
rect 16773 25653 16807 25687
rect 16807 25653 16816 25687
rect 16764 25644 16816 25653
rect 20260 25916 20312 25968
rect 22008 25891 22060 25900
rect 18788 25823 18840 25832
rect 18788 25789 18797 25823
rect 18797 25789 18831 25823
rect 18831 25789 18840 25823
rect 18788 25780 18840 25789
rect 18880 25823 18932 25832
rect 18880 25789 18889 25823
rect 18889 25789 18923 25823
rect 18923 25789 18932 25823
rect 22008 25857 22017 25891
rect 22017 25857 22051 25891
rect 22051 25857 22060 25891
rect 22008 25848 22060 25857
rect 23296 25891 23348 25900
rect 23296 25857 23305 25891
rect 23305 25857 23339 25891
rect 23339 25857 23348 25891
rect 23296 25848 23348 25857
rect 27160 25891 27212 25900
rect 27160 25857 27169 25891
rect 27169 25857 27203 25891
rect 27203 25857 27212 25891
rect 27160 25848 27212 25857
rect 24952 25823 25004 25832
rect 18880 25780 18932 25789
rect 19340 25712 19392 25764
rect 24952 25789 24961 25823
rect 24961 25789 24995 25823
rect 24995 25789 25004 25823
rect 24952 25780 25004 25789
rect 25228 25823 25280 25832
rect 25228 25789 25237 25823
rect 25237 25789 25271 25823
rect 25271 25789 25280 25823
rect 25228 25780 25280 25789
rect 27068 25780 27120 25832
rect 19432 25687 19484 25696
rect 19432 25653 19441 25687
rect 19441 25653 19475 25687
rect 19475 25653 19484 25687
rect 19432 25644 19484 25653
rect 21824 25687 21876 25696
rect 21824 25653 21833 25687
rect 21833 25653 21867 25687
rect 21867 25653 21876 25687
rect 21824 25644 21876 25653
rect 22192 25644 22244 25696
rect 22652 25644 22704 25696
rect 25412 25644 25464 25696
rect 5672 25542 5724 25594
rect 5736 25542 5788 25594
rect 5800 25542 5852 25594
rect 5864 25542 5916 25594
rect 5928 25542 5980 25594
rect 15118 25542 15170 25594
rect 15182 25542 15234 25594
rect 15246 25542 15298 25594
rect 15310 25542 15362 25594
rect 15374 25542 15426 25594
rect 24563 25542 24615 25594
rect 24627 25542 24679 25594
rect 24691 25542 24743 25594
rect 24755 25542 24807 25594
rect 24819 25542 24871 25594
rect 2596 25440 2648 25492
rect 3056 25440 3108 25492
rect 3884 25483 3936 25492
rect 3884 25449 3893 25483
rect 3893 25449 3927 25483
rect 3927 25449 3936 25483
rect 3884 25440 3936 25449
rect 6736 25440 6788 25492
rect 2780 25236 2832 25288
rect 4988 25372 5040 25424
rect 4160 25304 4212 25356
rect 4068 25279 4120 25288
rect 4068 25245 4072 25279
rect 4072 25245 4106 25279
rect 4106 25245 4120 25279
rect 4068 25236 4120 25245
rect 5172 25304 5224 25356
rect 9404 25440 9456 25492
rect 7564 25304 7616 25356
rect 4436 25279 4488 25288
rect 4436 25245 4445 25279
rect 4445 25245 4479 25279
rect 4479 25245 4488 25279
rect 4436 25236 4488 25245
rect 6920 25236 6972 25288
rect 7840 25236 7892 25288
rect 10968 25304 11020 25356
rect 11796 25440 11848 25492
rect 12256 25483 12308 25492
rect 12256 25449 12265 25483
rect 12265 25449 12299 25483
rect 12299 25449 12308 25483
rect 12256 25440 12308 25449
rect 14740 25440 14792 25492
rect 14924 25440 14976 25492
rect 17868 25440 17920 25492
rect 19064 25440 19116 25492
rect 22468 25440 22520 25492
rect 23020 25440 23072 25492
rect 12992 25372 13044 25424
rect 13452 25415 13504 25424
rect 13452 25381 13461 25415
rect 13461 25381 13495 25415
rect 13495 25381 13504 25415
rect 13452 25372 13504 25381
rect 7380 25168 7432 25220
rect 7472 25168 7524 25220
rect 10876 25168 10928 25220
rect 12072 25236 12124 25288
rect 12716 25236 12768 25288
rect 13268 25279 13320 25288
rect 13268 25245 13282 25279
rect 13282 25245 13316 25279
rect 13316 25245 13320 25279
rect 13268 25236 13320 25245
rect 13636 25236 13688 25288
rect 14280 25236 14332 25288
rect 15568 25279 15620 25288
rect 15568 25245 15577 25279
rect 15577 25245 15611 25279
rect 15611 25245 15620 25279
rect 15568 25236 15620 25245
rect 15108 25211 15160 25220
rect 3976 25100 4028 25152
rect 6828 25143 6880 25152
rect 6828 25109 6837 25143
rect 6837 25109 6871 25143
rect 6871 25109 6880 25143
rect 6828 25100 6880 25109
rect 8392 25100 8444 25152
rect 8760 25100 8812 25152
rect 10324 25100 10376 25152
rect 11796 25143 11848 25152
rect 11796 25109 11805 25143
rect 11805 25109 11839 25143
rect 11839 25109 11848 25143
rect 11796 25100 11848 25109
rect 12624 25143 12676 25152
rect 12624 25109 12633 25143
rect 12633 25109 12667 25143
rect 12667 25109 12676 25143
rect 12624 25100 12676 25109
rect 12808 25100 12860 25152
rect 15108 25177 15117 25211
rect 15117 25177 15151 25211
rect 15151 25177 15160 25211
rect 15108 25168 15160 25177
rect 14648 25100 14700 25152
rect 14832 25100 14884 25152
rect 16764 25304 16816 25356
rect 17132 25347 17184 25356
rect 17132 25313 17141 25347
rect 17141 25313 17175 25347
rect 17175 25313 17184 25347
rect 17132 25304 17184 25313
rect 19432 25304 19484 25356
rect 20260 25304 20312 25356
rect 16304 25236 16356 25288
rect 19524 25236 19576 25288
rect 15752 25168 15804 25220
rect 19340 25168 19392 25220
rect 16948 25143 17000 25152
rect 16948 25109 16957 25143
rect 16957 25109 16991 25143
rect 16991 25109 17000 25143
rect 16948 25100 17000 25109
rect 17040 25100 17092 25152
rect 18236 25143 18288 25152
rect 18236 25109 18245 25143
rect 18245 25109 18279 25143
rect 18279 25109 18288 25143
rect 18236 25100 18288 25109
rect 19524 25100 19576 25152
rect 19708 25100 19760 25152
rect 20352 25236 20404 25288
rect 20628 25143 20680 25152
rect 20628 25109 20637 25143
rect 20637 25109 20671 25143
rect 20671 25109 20680 25143
rect 20628 25100 20680 25109
rect 21824 25168 21876 25220
rect 22744 25279 22796 25288
rect 22744 25245 22753 25279
rect 22753 25245 22787 25279
rect 22787 25245 22796 25279
rect 22744 25236 22796 25245
rect 22836 25236 22888 25288
rect 25044 25440 25096 25492
rect 25228 25483 25280 25492
rect 25228 25449 25237 25483
rect 25237 25449 25271 25483
rect 25271 25449 25280 25483
rect 25228 25440 25280 25449
rect 27160 25440 27212 25492
rect 24032 25415 24084 25424
rect 24032 25381 24041 25415
rect 24041 25381 24075 25415
rect 24075 25381 24084 25415
rect 24032 25372 24084 25381
rect 23756 25304 23808 25356
rect 24400 25279 24452 25288
rect 24400 25245 24409 25279
rect 24409 25245 24443 25279
rect 24443 25245 24452 25279
rect 24400 25236 24452 25245
rect 24676 25415 24728 25424
rect 24676 25381 24685 25415
rect 24685 25381 24719 25415
rect 24719 25381 24728 25415
rect 24676 25372 24728 25381
rect 25780 25372 25832 25424
rect 27068 25304 27120 25356
rect 25780 25279 25832 25288
rect 22652 25168 22704 25220
rect 23020 25211 23072 25220
rect 23020 25177 23029 25211
rect 23029 25177 23063 25211
rect 23063 25177 23072 25211
rect 23020 25168 23072 25177
rect 23388 25168 23440 25220
rect 23756 25211 23808 25220
rect 23756 25177 23765 25211
rect 23765 25177 23799 25211
rect 23799 25177 23808 25211
rect 23756 25168 23808 25177
rect 25780 25245 25789 25279
rect 25789 25245 25823 25279
rect 25823 25245 25832 25279
rect 25780 25236 25832 25245
rect 25872 25279 25924 25288
rect 25872 25245 25881 25279
rect 25881 25245 25915 25279
rect 25915 25245 25924 25279
rect 25872 25236 25924 25245
rect 25596 25211 25648 25220
rect 25596 25177 25605 25211
rect 25605 25177 25639 25211
rect 25639 25177 25648 25211
rect 25596 25168 25648 25177
rect 25688 25100 25740 25152
rect 10395 24998 10447 25050
rect 10459 24998 10511 25050
rect 10523 24998 10575 25050
rect 10587 24998 10639 25050
rect 10651 24998 10703 25050
rect 19840 24998 19892 25050
rect 19904 24998 19956 25050
rect 19968 24998 20020 25050
rect 20032 24998 20084 25050
rect 20096 24998 20148 25050
rect 2780 24828 2832 24880
rect 2872 24803 2924 24812
rect 2872 24769 2881 24803
rect 2881 24769 2915 24803
rect 2915 24769 2924 24803
rect 2872 24760 2924 24769
rect 4712 24760 4764 24812
rect 4896 24760 4948 24812
rect 8392 24896 8444 24948
rect 9220 24939 9272 24948
rect 9220 24905 9229 24939
rect 9229 24905 9263 24939
rect 9263 24905 9272 24939
rect 9220 24896 9272 24905
rect 7748 24871 7800 24880
rect 7748 24837 7757 24871
rect 7757 24837 7791 24871
rect 7791 24837 7800 24871
rect 7748 24828 7800 24837
rect 8760 24828 8812 24880
rect 10416 24828 10468 24880
rect 7380 24803 7432 24812
rect 7380 24769 7389 24803
rect 7389 24769 7423 24803
rect 7423 24769 7432 24803
rect 7380 24760 7432 24769
rect 9772 24803 9824 24812
rect 3240 24692 3292 24744
rect 5172 24692 5224 24744
rect 7472 24735 7524 24744
rect 7472 24701 7481 24735
rect 7481 24701 7515 24735
rect 7515 24701 7524 24735
rect 7472 24692 7524 24701
rect 9772 24769 9781 24803
rect 9781 24769 9815 24803
rect 9815 24769 9824 24803
rect 10600 24828 10652 24880
rect 18972 24896 19024 24948
rect 22008 24939 22060 24948
rect 22008 24905 22017 24939
rect 22017 24905 22051 24939
rect 22051 24905 22060 24939
rect 22008 24896 22060 24905
rect 23296 24939 23348 24948
rect 23296 24905 23305 24939
rect 23305 24905 23339 24939
rect 23339 24905 23348 24939
rect 23296 24896 23348 24905
rect 12532 24828 12584 24880
rect 13268 24828 13320 24880
rect 13452 24828 13504 24880
rect 14372 24828 14424 24880
rect 14648 24828 14700 24880
rect 9772 24760 9824 24769
rect 10784 24760 10836 24812
rect 12164 24803 12216 24812
rect 10140 24692 10192 24744
rect 10968 24692 11020 24744
rect 11520 24692 11572 24744
rect 12164 24769 12173 24803
rect 12173 24769 12207 24803
rect 12207 24769 12216 24803
rect 12164 24760 12216 24769
rect 12716 24803 12768 24812
rect 12716 24769 12725 24803
rect 12725 24769 12759 24803
rect 12759 24769 12768 24803
rect 12716 24760 12768 24769
rect 14832 24760 14884 24812
rect 15292 24871 15344 24880
rect 15292 24837 15301 24871
rect 15301 24837 15335 24871
rect 15335 24837 15344 24871
rect 15292 24828 15344 24837
rect 16120 24828 16172 24880
rect 18880 24828 18932 24880
rect 20260 24828 20312 24880
rect 12808 24692 12860 24744
rect 13084 24735 13136 24744
rect 13084 24701 13093 24735
rect 13093 24701 13127 24735
rect 13127 24701 13136 24735
rect 13084 24692 13136 24701
rect 17040 24760 17092 24812
rect 20628 24828 20680 24880
rect 24400 24896 24452 24948
rect 25872 24896 25924 24948
rect 24676 24828 24728 24880
rect 26700 24828 26752 24880
rect 4068 24624 4120 24676
rect 6092 24624 6144 24676
rect 6920 24624 6972 24676
rect 2596 24556 2648 24608
rect 4344 24556 4396 24608
rect 7288 24556 7340 24608
rect 9496 24556 9548 24608
rect 10416 24556 10468 24608
rect 12624 24624 12676 24676
rect 12900 24667 12952 24676
rect 12900 24633 12909 24667
rect 12909 24633 12943 24667
rect 12943 24633 12952 24667
rect 12900 24624 12952 24633
rect 11520 24599 11572 24608
rect 11520 24565 11529 24599
rect 11529 24565 11563 24599
rect 11563 24565 11572 24599
rect 11520 24556 11572 24565
rect 12440 24556 12492 24608
rect 12992 24556 13044 24608
rect 14372 24556 14424 24608
rect 15844 24599 15896 24608
rect 15844 24565 15853 24599
rect 15853 24565 15887 24599
rect 15887 24565 15896 24599
rect 15844 24556 15896 24565
rect 16304 24556 16356 24608
rect 18052 24692 18104 24744
rect 18328 24692 18380 24744
rect 18788 24735 18840 24744
rect 18788 24701 18797 24735
rect 18797 24701 18831 24735
rect 18831 24701 18840 24735
rect 18788 24692 18840 24701
rect 19708 24692 19760 24744
rect 19156 24624 19208 24676
rect 19248 24624 19300 24676
rect 21732 24760 21784 24812
rect 25136 24760 25188 24812
rect 24032 24692 24084 24744
rect 25044 24735 25096 24744
rect 25044 24701 25053 24735
rect 25053 24701 25087 24735
rect 25087 24701 25096 24735
rect 25044 24692 25096 24701
rect 25688 24803 25740 24812
rect 25688 24769 25691 24803
rect 25691 24769 25740 24803
rect 25688 24760 25740 24769
rect 25872 24760 25924 24812
rect 19064 24556 19116 24608
rect 20904 24556 20956 24608
rect 20996 24556 21048 24608
rect 21272 24556 21324 24608
rect 24124 24556 24176 24608
rect 25780 24599 25832 24608
rect 25780 24565 25789 24599
rect 25789 24565 25823 24599
rect 25823 24565 25832 24599
rect 25780 24556 25832 24565
rect 26516 24599 26568 24608
rect 26516 24565 26525 24599
rect 26525 24565 26559 24599
rect 26559 24565 26568 24599
rect 26516 24556 26568 24565
rect 26700 24599 26752 24608
rect 26700 24565 26709 24599
rect 26709 24565 26743 24599
rect 26743 24565 26752 24599
rect 26700 24556 26752 24565
rect 5672 24454 5724 24506
rect 5736 24454 5788 24506
rect 5800 24454 5852 24506
rect 5864 24454 5916 24506
rect 5928 24454 5980 24506
rect 15118 24454 15170 24506
rect 15182 24454 15234 24506
rect 15246 24454 15298 24506
rect 15310 24454 15362 24506
rect 15374 24454 15426 24506
rect 24563 24454 24615 24506
rect 24627 24454 24679 24506
rect 24691 24454 24743 24506
rect 24755 24454 24807 24506
rect 24819 24454 24871 24506
rect 2872 24352 2924 24404
rect 4712 24395 4764 24404
rect 4712 24361 4721 24395
rect 4721 24361 4755 24395
rect 4755 24361 4764 24395
rect 4712 24352 4764 24361
rect 10784 24395 10836 24404
rect 10784 24361 10793 24395
rect 10793 24361 10827 24395
rect 10827 24361 10836 24395
rect 10784 24352 10836 24361
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 3056 24259 3108 24268
rect 3056 24225 3065 24259
rect 3065 24225 3099 24259
rect 3099 24225 3108 24259
rect 3056 24216 3108 24225
rect 4252 24259 4304 24268
rect 4252 24225 4261 24259
rect 4261 24225 4295 24259
rect 4295 24225 4304 24259
rect 11520 24352 11572 24404
rect 15568 24352 15620 24404
rect 15844 24352 15896 24404
rect 17868 24352 17920 24404
rect 18328 24352 18380 24404
rect 19708 24395 19760 24404
rect 19708 24361 19717 24395
rect 19717 24361 19751 24395
rect 19751 24361 19760 24395
rect 19708 24352 19760 24361
rect 22652 24352 22704 24404
rect 23388 24352 23440 24404
rect 6920 24259 6972 24268
rect 4252 24216 4304 24225
rect 6920 24225 6929 24259
rect 6929 24225 6963 24259
rect 6963 24225 6972 24259
rect 6920 24216 6972 24225
rect 9496 24259 9548 24268
rect 9496 24225 9505 24259
rect 9505 24225 9539 24259
rect 9539 24225 9548 24259
rect 9496 24216 9548 24225
rect 10416 24259 10468 24268
rect 10416 24225 10425 24259
rect 10425 24225 10459 24259
rect 10459 24225 10468 24259
rect 10416 24216 10468 24225
rect 11336 24216 11388 24268
rect 13084 24216 13136 24268
rect 3240 24191 3292 24200
rect 1952 24080 2004 24132
rect 3240 24157 3249 24191
rect 3249 24157 3283 24191
rect 3283 24157 3292 24191
rect 3240 24148 3292 24157
rect 3148 24080 3200 24132
rect 3424 24148 3476 24200
rect 4344 24191 4396 24200
rect 4344 24157 4353 24191
rect 4353 24157 4387 24191
rect 4387 24157 4396 24191
rect 4344 24148 4396 24157
rect 3608 24080 3660 24132
rect 4896 24148 4948 24200
rect 5172 24148 5224 24200
rect 9588 24191 9640 24200
rect 9588 24157 9597 24191
rect 9597 24157 9631 24191
rect 9631 24157 9640 24191
rect 9588 24148 9640 24157
rect 11152 24148 11204 24200
rect 14372 24191 14424 24200
rect 14372 24157 14381 24191
rect 14381 24157 14415 24191
rect 14415 24157 14424 24191
rect 14372 24148 14424 24157
rect 16856 24191 16908 24200
rect 16856 24157 16865 24191
rect 16865 24157 16899 24191
rect 16899 24157 16908 24191
rect 16856 24148 16908 24157
rect 18144 24148 18196 24200
rect 18696 24284 18748 24336
rect 19248 24327 19300 24336
rect 19248 24293 19257 24327
rect 19257 24293 19291 24327
rect 19291 24293 19300 24327
rect 19248 24284 19300 24293
rect 22468 24327 22520 24336
rect 22468 24293 22477 24327
rect 22477 24293 22511 24327
rect 22511 24293 22520 24327
rect 22468 24284 22520 24293
rect 20352 24148 20404 24200
rect 20996 24148 21048 24200
rect 22744 24216 22796 24268
rect 22928 24216 22980 24268
rect 22192 24191 22244 24200
rect 22192 24157 22201 24191
rect 22201 24157 22235 24191
rect 22235 24157 22244 24191
rect 22192 24148 22244 24157
rect 22836 24148 22888 24200
rect 23204 24148 23256 24200
rect 26240 24352 26292 24404
rect 25780 24259 25832 24268
rect 25780 24225 25789 24259
rect 25789 24225 25823 24259
rect 25823 24225 25832 24259
rect 25780 24216 25832 24225
rect 23664 24191 23716 24200
rect 23664 24157 23678 24191
rect 23678 24157 23712 24191
rect 23712 24157 23716 24191
rect 24400 24191 24452 24200
rect 23664 24148 23716 24157
rect 24400 24157 24409 24191
rect 24409 24157 24443 24191
rect 24443 24157 24452 24191
rect 24400 24148 24452 24157
rect 5540 24080 5592 24132
rect 7196 24123 7248 24132
rect 7196 24089 7205 24123
rect 7205 24089 7239 24123
rect 7239 24089 7248 24123
rect 7196 24080 7248 24089
rect 7288 24080 7340 24132
rect 3332 24012 3384 24064
rect 6460 24055 6512 24064
rect 6460 24021 6469 24055
rect 6469 24021 6503 24055
rect 6503 24021 6512 24055
rect 6460 24012 6512 24021
rect 6736 24012 6788 24064
rect 11060 24080 11112 24132
rect 12716 24080 12768 24132
rect 17776 24080 17828 24132
rect 8760 24012 8812 24064
rect 9864 24012 9916 24064
rect 12624 24012 12676 24064
rect 14556 24055 14608 24064
rect 14556 24021 14565 24055
rect 14565 24021 14599 24055
rect 14599 24021 14608 24055
rect 14556 24012 14608 24021
rect 20168 24080 20220 24132
rect 22652 24080 22704 24132
rect 19340 24012 19392 24064
rect 23020 24012 23072 24064
rect 25044 24080 25096 24132
rect 26516 24080 26568 24132
rect 23388 24012 23440 24064
rect 23572 24012 23624 24064
rect 23756 24012 23808 24064
rect 24032 24012 24084 24064
rect 24584 24055 24636 24064
rect 24584 24021 24593 24055
rect 24593 24021 24627 24055
rect 24627 24021 24636 24055
rect 24584 24012 24636 24021
rect 26700 24012 26752 24064
rect 27620 24012 27672 24064
rect 10395 23910 10447 23962
rect 10459 23910 10511 23962
rect 10523 23910 10575 23962
rect 10587 23910 10639 23962
rect 10651 23910 10703 23962
rect 19840 23910 19892 23962
rect 19904 23910 19956 23962
rect 19968 23910 20020 23962
rect 20032 23910 20084 23962
rect 20096 23910 20148 23962
rect 1952 23783 2004 23792
rect 1952 23749 1961 23783
rect 1961 23749 1995 23783
rect 1995 23749 2004 23783
rect 1952 23740 2004 23749
rect 2596 23851 2648 23860
rect 2596 23817 2605 23851
rect 2605 23817 2639 23851
rect 2639 23817 2648 23851
rect 2596 23808 2648 23817
rect 3240 23808 3292 23860
rect 3608 23851 3660 23860
rect 3608 23817 3617 23851
rect 3617 23817 3651 23851
rect 3651 23817 3660 23851
rect 3608 23808 3660 23817
rect 4344 23808 4396 23860
rect 5540 23851 5592 23860
rect 2872 23740 2924 23792
rect 3148 23740 3200 23792
rect 2780 23715 2832 23724
rect 2780 23681 2789 23715
rect 2789 23681 2823 23715
rect 2823 23681 2832 23715
rect 2780 23672 2832 23681
rect 2780 23536 2832 23588
rect 3056 23604 3108 23656
rect 3792 23672 3844 23724
rect 4252 23672 4304 23724
rect 5540 23817 5549 23851
rect 5549 23817 5583 23851
rect 5583 23817 5592 23851
rect 5540 23808 5592 23817
rect 6736 23851 6788 23860
rect 6736 23817 6745 23851
rect 6745 23817 6779 23851
rect 6779 23817 6788 23851
rect 6736 23808 6788 23817
rect 7196 23808 7248 23860
rect 10876 23808 10928 23860
rect 12164 23808 12216 23860
rect 12716 23851 12768 23860
rect 12716 23817 12725 23851
rect 12725 23817 12759 23851
rect 12759 23817 12768 23851
rect 12716 23808 12768 23817
rect 4804 23715 4856 23724
rect 3884 23604 3936 23656
rect 4804 23681 4813 23715
rect 4813 23681 4847 23715
rect 4847 23681 4856 23715
rect 4804 23672 4856 23681
rect 4988 23715 5040 23724
rect 4988 23681 4991 23715
rect 4991 23681 5040 23715
rect 4988 23672 5040 23681
rect 6460 23740 6512 23792
rect 6552 23672 6604 23724
rect 6828 23604 6880 23656
rect 7472 23672 7524 23724
rect 8760 23672 8812 23724
rect 9772 23672 9824 23724
rect 10784 23672 10836 23724
rect 12624 23672 12676 23724
rect 11704 23647 11756 23656
rect 11704 23613 11713 23647
rect 11713 23613 11747 23647
rect 11747 23613 11756 23647
rect 11704 23604 11756 23613
rect 4068 23536 4120 23588
rect 17776 23851 17828 23860
rect 14556 23740 14608 23792
rect 13176 23715 13228 23724
rect 13176 23681 13185 23715
rect 13185 23681 13219 23715
rect 13219 23681 13228 23715
rect 13176 23672 13228 23681
rect 15568 23672 15620 23724
rect 15844 23715 15896 23724
rect 15844 23681 15853 23715
rect 15853 23681 15887 23715
rect 15887 23681 15896 23715
rect 15844 23672 15896 23681
rect 13084 23604 13136 23656
rect 13728 23647 13780 23656
rect 13728 23613 13737 23647
rect 13737 23613 13771 23647
rect 13771 23613 13780 23647
rect 13728 23604 13780 23613
rect 15752 23604 15804 23656
rect 16304 23672 16356 23724
rect 17776 23817 17785 23851
rect 17785 23817 17819 23851
rect 17819 23817 17828 23851
rect 17776 23808 17828 23817
rect 19156 23808 19208 23860
rect 17868 23715 17920 23724
rect 17868 23681 17877 23715
rect 17877 23681 17911 23715
rect 17911 23681 17920 23715
rect 17868 23672 17920 23681
rect 18052 23672 18104 23724
rect 18328 23672 18380 23724
rect 18972 23740 19024 23792
rect 20168 23808 20220 23860
rect 20352 23808 20404 23860
rect 22376 23808 22428 23860
rect 22560 23808 22612 23860
rect 23388 23808 23440 23860
rect 24400 23808 24452 23860
rect 26240 23808 26292 23860
rect 24032 23783 24084 23792
rect 18604 23672 18656 23724
rect 19156 23672 19208 23724
rect 18328 23536 18380 23588
rect 4988 23468 5040 23520
rect 5540 23468 5592 23520
rect 6092 23468 6144 23520
rect 10232 23511 10284 23520
rect 10232 23477 10241 23511
rect 10241 23477 10275 23511
rect 10275 23477 10284 23511
rect 10232 23468 10284 23477
rect 11428 23468 11480 23520
rect 11796 23468 11848 23520
rect 15476 23511 15528 23520
rect 15476 23477 15485 23511
rect 15485 23477 15519 23511
rect 15519 23477 15528 23511
rect 15476 23468 15528 23477
rect 16672 23511 16724 23520
rect 16672 23477 16681 23511
rect 16681 23477 16715 23511
rect 16715 23477 16724 23511
rect 16672 23468 16724 23477
rect 19064 23604 19116 23656
rect 18972 23536 19024 23588
rect 19892 23715 19944 23724
rect 19892 23681 19901 23715
rect 19901 23681 19935 23715
rect 19935 23681 19944 23715
rect 22008 23715 22060 23724
rect 19892 23672 19944 23681
rect 22008 23681 22017 23715
rect 22017 23681 22051 23715
rect 22051 23681 22060 23715
rect 22008 23672 22060 23681
rect 22744 23715 22796 23724
rect 22744 23681 22753 23715
rect 22753 23681 22787 23715
rect 22787 23681 22796 23715
rect 22744 23672 22796 23681
rect 24032 23749 24041 23783
rect 24041 23749 24075 23783
rect 24075 23749 24084 23783
rect 24032 23740 24084 23749
rect 24584 23740 24636 23792
rect 23756 23647 23808 23656
rect 23756 23613 23765 23647
rect 23765 23613 23799 23647
rect 23799 23613 23808 23647
rect 23756 23604 23808 23613
rect 19064 23468 19116 23520
rect 21824 23511 21876 23520
rect 21824 23477 21833 23511
rect 21833 23477 21867 23511
rect 21867 23477 21876 23511
rect 21824 23468 21876 23477
rect 22928 23468 22980 23520
rect 26332 23468 26384 23520
rect 5672 23366 5724 23418
rect 5736 23366 5788 23418
rect 5800 23366 5852 23418
rect 5864 23366 5916 23418
rect 5928 23366 5980 23418
rect 15118 23366 15170 23418
rect 15182 23366 15234 23418
rect 15246 23366 15298 23418
rect 15310 23366 15362 23418
rect 15374 23366 15426 23418
rect 24563 23366 24615 23418
rect 24627 23366 24679 23418
rect 24691 23366 24743 23418
rect 24755 23366 24807 23418
rect 24819 23366 24871 23418
rect 10048 23264 10100 23316
rect 10140 23264 10192 23316
rect 11244 23264 11296 23316
rect 13728 23264 13780 23316
rect 14372 23307 14424 23316
rect 14372 23273 14381 23307
rect 14381 23273 14415 23307
rect 14415 23273 14424 23307
rect 14372 23264 14424 23273
rect 18512 23264 18564 23316
rect 20812 23264 20864 23316
rect 22100 23264 22152 23316
rect 22744 23264 22796 23316
rect 23848 23264 23900 23316
rect 24400 23264 24452 23316
rect 3976 23128 4028 23180
rect 11428 23196 11480 23248
rect 18052 23196 18104 23248
rect 18972 23196 19024 23248
rect 23664 23196 23716 23248
rect 3332 23060 3384 23112
rect 3792 23103 3844 23112
rect 3792 23069 3801 23103
rect 3801 23069 3835 23103
rect 3835 23069 3844 23103
rect 3792 23060 3844 23069
rect 3884 23103 3936 23112
rect 3884 23069 3893 23103
rect 3893 23069 3927 23103
rect 3927 23069 3936 23103
rect 3884 23060 3936 23069
rect 4712 23060 4764 23112
rect 3240 22992 3292 23044
rect 1676 22924 1728 22976
rect 4160 22924 4212 22976
rect 4344 22924 4396 22976
rect 4804 22924 4856 22976
rect 5540 22992 5592 23044
rect 7196 22992 7248 23044
rect 7932 23035 7984 23044
rect 7932 23001 7941 23035
rect 7941 23001 7975 23035
rect 7975 23001 7984 23035
rect 7932 22992 7984 23001
rect 9036 22992 9088 23044
rect 10324 23171 10376 23180
rect 10324 23137 10349 23171
rect 10349 23137 10376 23171
rect 10324 23128 10376 23137
rect 11704 23128 11756 23180
rect 9864 22992 9916 23044
rect 10232 23060 10284 23112
rect 11244 23060 11296 23112
rect 13084 23128 13136 23180
rect 15476 23128 15528 23180
rect 18788 23128 18840 23180
rect 20996 23128 21048 23180
rect 23756 23128 23808 23180
rect 15108 23103 15160 23112
rect 11336 23035 11388 23044
rect 8116 22924 8168 22976
rect 8208 22924 8260 22976
rect 10232 22967 10284 22976
rect 10232 22933 10241 22967
rect 10241 22933 10275 22967
rect 10275 22933 10284 22967
rect 11336 23001 11345 23035
rect 11345 23001 11379 23035
rect 11379 23001 11388 23035
rect 11336 22992 11388 23001
rect 11796 22992 11848 23044
rect 12900 23035 12952 23044
rect 12900 23001 12909 23035
rect 12909 23001 12943 23035
rect 12943 23001 12952 23035
rect 12900 22992 12952 23001
rect 10232 22924 10284 22933
rect 11520 22924 11572 22976
rect 13176 22992 13228 23044
rect 15108 23069 15117 23103
rect 15117 23069 15151 23103
rect 15151 23069 15160 23103
rect 15108 23060 15160 23069
rect 15292 23103 15344 23112
rect 15292 23069 15301 23103
rect 15301 23069 15335 23103
rect 15335 23069 15344 23103
rect 15292 23060 15344 23069
rect 18420 23103 18472 23112
rect 18420 23069 18429 23103
rect 18429 23069 18463 23103
rect 18463 23069 18472 23103
rect 18420 23060 18472 23069
rect 16672 22992 16724 23044
rect 16764 22992 16816 23044
rect 17132 23035 17184 23044
rect 17132 23001 17141 23035
rect 17141 23001 17175 23035
rect 17175 23001 17184 23035
rect 17132 22992 17184 23001
rect 18696 23035 18748 23044
rect 18696 23001 18705 23035
rect 18705 23001 18739 23035
rect 18739 23001 18748 23035
rect 18696 22992 18748 23001
rect 21824 22992 21876 23044
rect 22468 23035 22520 23044
rect 22468 23001 22477 23035
rect 22477 23001 22511 23035
rect 22511 23001 22520 23035
rect 22468 22992 22520 23001
rect 22560 22992 22612 23044
rect 23296 23060 23348 23112
rect 19616 22967 19668 22976
rect 19616 22933 19625 22967
rect 19625 22933 19659 22967
rect 19659 22933 19668 22967
rect 19616 22924 19668 22933
rect 19708 22967 19760 22976
rect 19708 22933 19717 22967
rect 19717 22933 19751 22967
rect 19751 22933 19760 22967
rect 19708 22924 19760 22933
rect 23020 22924 23072 22976
rect 23204 22924 23256 22976
rect 26240 22992 26292 23044
rect 23848 22924 23900 22976
rect 24216 22924 24268 22976
rect 10395 22822 10447 22874
rect 10459 22822 10511 22874
rect 10523 22822 10575 22874
rect 10587 22822 10639 22874
rect 10651 22822 10703 22874
rect 19840 22822 19892 22874
rect 19904 22822 19956 22874
rect 19968 22822 20020 22874
rect 20032 22822 20084 22874
rect 20096 22822 20148 22874
rect 3056 22720 3108 22772
rect 2872 22652 2924 22704
rect 4344 22720 4396 22772
rect 4436 22720 4488 22772
rect 7196 22763 7248 22772
rect 7196 22729 7205 22763
rect 7205 22729 7239 22763
rect 7239 22729 7248 22763
rect 7196 22720 7248 22729
rect 7932 22720 7984 22772
rect 9772 22763 9824 22772
rect 9772 22729 9781 22763
rect 9781 22729 9815 22763
rect 9815 22729 9824 22763
rect 9772 22720 9824 22729
rect 9864 22763 9916 22772
rect 9864 22729 9873 22763
rect 9873 22729 9907 22763
rect 9907 22729 9916 22763
rect 9864 22720 9916 22729
rect 4252 22652 4304 22704
rect 1676 22627 1728 22636
rect 1676 22593 1710 22627
rect 1710 22593 1728 22627
rect 1676 22584 1728 22593
rect 3792 22584 3844 22636
rect 3976 22584 4028 22636
rect 4160 22627 4212 22636
rect 4160 22593 4169 22627
rect 4169 22593 4203 22627
rect 4203 22593 4212 22627
rect 7748 22652 7800 22704
rect 4160 22584 4212 22593
rect 3424 22516 3476 22568
rect 8116 22584 8168 22636
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 9588 22695 9640 22704
rect 9588 22661 9597 22695
rect 9597 22661 9631 22695
rect 9631 22661 9640 22695
rect 9588 22652 9640 22661
rect 10416 22652 10468 22704
rect 10876 22652 10928 22704
rect 11336 22627 11388 22636
rect 11336 22593 11345 22627
rect 11345 22593 11379 22627
rect 11379 22593 11388 22627
rect 11336 22584 11388 22593
rect 11520 22627 11572 22636
rect 11520 22593 11529 22627
rect 11529 22593 11563 22627
rect 11563 22593 11572 22627
rect 11520 22584 11572 22593
rect 11612 22584 11664 22636
rect 12440 22652 12492 22704
rect 12624 22652 12676 22704
rect 13176 22584 13228 22636
rect 15660 22720 15712 22772
rect 15292 22652 15344 22704
rect 16856 22652 16908 22704
rect 4436 22448 4488 22500
rect 9680 22448 9732 22500
rect 10692 22448 10744 22500
rect 11704 22516 11756 22568
rect 11612 22491 11664 22500
rect 3056 22423 3108 22432
rect 3056 22389 3065 22423
rect 3065 22389 3099 22423
rect 3099 22389 3108 22423
rect 3056 22380 3108 22389
rect 3884 22423 3936 22432
rect 3884 22389 3893 22423
rect 3893 22389 3927 22423
rect 3927 22389 3936 22423
rect 3884 22380 3936 22389
rect 4252 22423 4304 22432
rect 4252 22389 4261 22423
rect 4261 22389 4295 22423
rect 4295 22389 4304 22423
rect 4252 22380 4304 22389
rect 7932 22380 7984 22432
rect 11060 22380 11112 22432
rect 11612 22457 11621 22491
rect 11621 22457 11655 22491
rect 11655 22457 11664 22491
rect 11612 22448 11664 22457
rect 11796 22448 11848 22500
rect 12532 22448 12584 22500
rect 15108 22584 15160 22636
rect 15476 22584 15528 22636
rect 15844 22627 15896 22636
rect 15844 22593 15853 22627
rect 15853 22593 15887 22627
rect 15887 22593 15896 22627
rect 15844 22584 15896 22593
rect 18696 22652 18748 22704
rect 19708 22720 19760 22772
rect 21732 22720 21784 22772
rect 22008 22720 22060 22772
rect 22652 22720 22704 22772
rect 22836 22720 22888 22772
rect 18972 22627 19024 22636
rect 18972 22593 18981 22627
rect 18981 22593 19015 22627
rect 19015 22593 19024 22627
rect 18972 22584 19024 22593
rect 20904 22652 20956 22704
rect 20720 22627 20772 22636
rect 19064 22559 19116 22568
rect 19064 22525 19073 22559
rect 19073 22525 19107 22559
rect 19107 22525 19116 22559
rect 19064 22516 19116 22525
rect 19248 22448 19300 22500
rect 20720 22593 20738 22627
rect 20738 22593 20772 22627
rect 20720 22584 20772 22593
rect 20996 22627 21048 22636
rect 20996 22593 21005 22627
rect 21005 22593 21039 22627
rect 21039 22593 21048 22627
rect 20996 22584 21048 22593
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 22192 22584 22244 22636
rect 22560 22627 22612 22636
rect 22560 22593 22569 22627
rect 22569 22593 22603 22627
rect 22603 22593 22612 22627
rect 22560 22584 22612 22593
rect 22744 22584 22796 22636
rect 23756 22584 23808 22636
rect 24216 22559 24268 22568
rect 24216 22525 24225 22559
rect 24225 22525 24259 22559
rect 24259 22525 24268 22559
rect 24216 22516 24268 22525
rect 13360 22423 13412 22432
rect 13360 22389 13369 22423
rect 13369 22389 13403 22423
rect 13403 22389 13412 22423
rect 13360 22380 13412 22389
rect 14740 22423 14792 22432
rect 14740 22389 14749 22423
rect 14749 22389 14783 22423
rect 14783 22389 14792 22423
rect 14740 22380 14792 22389
rect 15660 22380 15712 22432
rect 15844 22380 15896 22432
rect 18512 22380 18564 22432
rect 20628 22380 20680 22432
rect 23296 22448 23348 22500
rect 22284 22423 22336 22432
rect 22284 22389 22293 22423
rect 22293 22389 22327 22423
rect 22327 22389 22336 22423
rect 22284 22380 22336 22389
rect 26240 22380 26292 22432
rect 5672 22278 5724 22330
rect 5736 22278 5788 22330
rect 5800 22278 5852 22330
rect 5864 22278 5916 22330
rect 5928 22278 5980 22330
rect 15118 22278 15170 22330
rect 15182 22278 15234 22330
rect 15246 22278 15298 22330
rect 15310 22278 15362 22330
rect 15374 22278 15426 22330
rect 24563 22278 24615 22330
rect 24627 22278 24679 22330
rect 24691 22278 24743 22330
rect 24755 22278 24807 22330
rect 24819 22278 24871 22330
rect 3424 22176 3476 22228
rect 9404 22176 9456 22228
rect 12808 22176 12860 22228
rect 15016 22176 15068 22228
rect 19340 22176 19392 22228
rect 22376 22176 22428 22228
rect 22468 22176 22520 22228
rect 25596 22176 25648 22228
rect 2872 22108 2924 22160
rect 9956 22108 10008 22160
rect 10232 22108 10284 22160
rect 8208 22040 8260 22092
rect 9772 22040 9824 22092
rect 10600 22108 10652 22160
rect 11520 22108 11572 22160
rect 2780 21972 2832 22024
rect 3884 21972 3936 22024
rect 4160 21972 4212 22024
rect 4436 21972 4488 22024
rect 4712 21972 4764 22024
rect 6920 22015 6972 22024
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 6920 21972 6972 21981
rect 8944 21972 8996 22024
rect 9312 22015 9364 22024
rect 9312 21981 9321 22015
rect 9321 21981 9355 22015
rect 9355 21981 9364 22015
rect 9588 22015 9640 22024
rect 9312 21972 9364 21981
rect 9588 21981 9597 22015
rect 9597 21981 9631 22015
rect 9631 21981 9640 22015
rect 9588 21972 9640 21981
rect 15476 22108 15528 22160
rect 16488 22040 16540 22092
rect 18512 22083 18564 22092
rect 18512 22049 18521 22083
rect 18521 22049 18555 22083
rect 18555 22049 18564 22083
rect 18512 22040 18564 22049
rect 5356 21904 5408 21956
rect 4252 21836 4304 21888
rect 4344 21836 4396 21888
rect 6460 21904 6512 21956
rect 7932 21904 7984 21956
rect 6276 21879 6328 21888
rect 6276 21845 6285 21879
rect 6285 21845 6319 21879
rect 6319 21845 6328 21879
rect 6276 21836 6328 21845
rect 10692 22015 10744 22024
rect 10692 21981 10701 22015
rect 10701 21981 10735 22015
rect 10735 21981 10744 22015
rect 10692 21972 10744 21981
rect 10876 21972 10928 22024
rect 11520 21972 11572 22024
rect 13268 21972 13320 22024
rect 15200 21972 15252 22024
rect 18788 22040 18840 22092
rect 19064 22040 19116 22092
rect 20720 22040 20772 22092
rect 20812 22040 20864 22092
rect 10324 21904 10376 21956
rect 11704 21904 11756 21956
rect 12164 21947 12216 21956
rect 12164 21913 12173 21947
rect 12173 21913 12207 21947
rect 12207 21913 12216 21947
rect 12164 21904 12216 21913
rect 14924 21904 14976 21956
rect 15936 21904 15988 21956
rect 16856 21904 16908 21956
rect 19156 21972 19208 22024
rect 19340 21972 19392 22024
rect 18972 21904 19024 21956
rect 19708 21972 19760 22024
rect 8760 21836 8812 21888
rect 12808 21836 12860 21888
rect 12992 21836 13044 21888
rect 13544 21836 13596 21888
rect 16028 21836 16080 21888
rect 17868 21836 17920 21888
rect 17960 21836 18012 21888
rect 18328 21836 18380 21888
rect 19340 21836 19392 21888
rect 22284 21904 22336 21956
rect 22652 22040 22704 22092
rect 22836 21972 22888 22024
rect 23112 22040 23164 22092
rect 23572 22040 23624 22092
rect 24124 22083 24176 22092
rect 24124 22049 24133 22083
rect 24133 22049 24167 22083
rect 24167 22049 24176 22083
rect 24124 22040 24176 22049
rect 23848 22015 23900 22024
rect 23848 21981 23857 22015
rect 23857 21981 23891 22015
rect 23891 21981 23900 22015
rect 23848 21972 23900 21981
rect 23112 21947 23164 21956
rect 22100 21836 22152 21888
rect 22836 21836 22888 21888
rect 23112 21913 23121 21947
rect 23121 21913 23155 21947
rect 23155 21913 23164 21947
rect 23112 21904 23164 21913
rect 25228 21904 25280 21956
rect 23480 21836 23532 21888
rect 24032 21879 24084 21888
rect 24032 21845 24041 21879
rect 24041 21845 24075 21879
rect 24075 21845 24084 21879
rect 24032 21836 24084 21845
rect 10395 21734 10447 21786
rect 10459 21734 10511 21786
rect 10523 21734 10575 21786
rect 10587 21734 10639 21786
rect 10651 21734 10703 21786
rect 19840 21734 19892 21786
rect 19904 21734 19956 21786
rect 19968 21734 20020 21786
rect 20032 21734 20084 21786
rect 20096 21734 20148 21786
rect 3332 21496 3384 21548
rect 3608 21539 3660 21548
rect 3608 21505 3618 21539
rect 3618 21505 3652 21539
rect 3652 21505 3660 21539
rect 3608 21496 3660 21505
rect 3976 21564 4028 21616
rect 4896 21632 4948 21684
rect 4160 21496 4212 21548
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 6460 21632 6512 21684
rect 6276 21564 6328 21616
rect 6920 21632 6972 21684
rect 7748 21632 7800 21684
rect 8944 21632 8996 21684
rect 9864 21632 9916 21684
rect 10784 21632 10836 21684
rect 11244 21632 11296 21684
rect 12256 21632 12308 21684
rect 13544 21632 13596 21684
rect 15200 21632 15252 21684
rect 16396 21632 16448 21684
rect 16856 21675 16908 21684
rect 16856 21641 16865 21675
rect 16865 21641 16899 21675
rect 16899 21641 16908 21675
rect 16856 21632 16908 21641
rect 19432 21675 19484 21684
rect 19432 21641 19441 21675
rect 19441 21641 19475 21675
rect 19475 21641 19484 21675
rect 19432 21632 19484 21641
rect 22192 21632 22244 21684
rect 6368 21539 6420 21548
rect 6368 21505 6377 21539
rect 6377 21505 6411 21539
rect 6411 21505 6420 21539
rect 6368 21496 6420 21505
rect 8300 21564 8352 21616
rect 8760 21564 8812 21616
rect 10140 21564 10192 21616
rect 10324 21564 10376 21616
rect 12164 21607 12216 21616
rect 8024 21496 8076 21548
rect 4160 21360 4212 21412
rect 5448 21360 5500 21412
rect 6736 21403 6788 21412
rect 6736 21369 6745 21403
rect 6745 21369 6779 21403
rect 6779 21369 6788 21403
rect 6736 21360 6788 21369
rect 7840 21428 7892 21480
rect 9588 21496 9640 21548
rect 10784 21539 10836 21548
rect 10784 21505 10793 21539
rect 10793 21505 10827 21539
rect 10827 21505 10836 21539
rect 10784 21496 10836 21505
rect 12164 21573 12173 21607
rect 12173 21573 12207 21607
rect 12207 21573 12216 21607
rect 12164 21564 12216 21573
rect 12992 21564 13044 21616
rect 14740 21564 14792 21616
rect 15476 21564 15528 21616
rect 12808 21496 12860 21548
rect 15844 21496 15896 21548
rect 22836 21564 22888 21616
rect 20904 21539 20956 21548
rect 20904 21505 20913 21539
rect 20913 21505 20947 21539
rect 20947 21505 20956 21539
rect 20904 21496 20956 21505
rect 9956 21471 10008 21480
rect 9956 21437 9982 21471
rect 9982 21437 10008 21471
rect 9956 21428 10008 21437
rect 10692 21471 10744 21480
rect 3884 21292 3936 21344
rect 6092 21335 6144 21344
rect 6092 21301 6101 21335
rect 6101 21301 6135 21335
rect 6135 21301 6144 21335
rect 6092 21292 6144 21301
rect 9220 21360 9272 21412
rect 9312 21360 9364 21412
rect 10692 21437 10701 21471
rect 10701 21437 10735 21471
rect 10735 21437 10744 21471
rect 10692 21428 10744 21437
rect 11520 21428 11572 21480
rect 13728 21471 13780 21480
rect 13728 21437 13737 21471
rect 13737 21437 13771 21471
rect 13771 21437 13780 21471
rect 13728 21428 13780 21437
rect 14924 21428 14976 21480
rect 7840 21335 7892 21344
rect 7840 21301 7849 21335
rect 7849 21301 7883 21335
rect 7883 21301 7892 21335
rect 7840 21292 7892 21301
rect 9404 21292 9456 21344
rect 10876 21360 10928 21412
rect 11428 21360 11480 21412
rect 12348 21360 12400 21412
rect 11520 21335 11572 21344
rect 11520 21301 11529 21335
rect 11529 21301 11563 21335
rect 11563 21301 11572 21335
rect 11520 21292 11572 21301
rect 14096 21292 14148 21344
rect 16120 21360 16172 21412
rect 18052 21360 18104 21412
rect 19248 21360 19300 21412
rect 19432 21360 19484 21412
rect 20536 21360 20588 21412
rect 15476 21292 15528 21344
rect 16212 21292 16264 21344
rect 20904 21292 20956 21344
rect 22008 21496 22060 21548
rect 22284 21539 22336 21548
rect 22284 21505 22333 21539
rect 22333 21505 22336 21539
rect 22284 21496 22336 21505
rect 22744 21539 22796 21548
rect 22376 21360 22428 21412
rect 22468 21360 22520 21412
rect 22744 21505 22753 21539
rect 22753 21505 22787 21539
rect 22787 21505 22796 21539
rect 22744 21496 22796 21505
rect 23848 21632 23900 21684
rect 23572 21607 23624 21616
rect 23572 21573 23581 21607
rect 23581 21573 23615 21607
rect 23615 21573 23624 21607
rect 23572 21564 23624 21573
rect 24032 21564 24084 21616
rect 22652 21428 22704 21480
rect 23112 21360 23164 21412
rect 22836 21335 22888 21344
rect 22836 21301 22845 21335
rect 22845 21301 22879 21335
rect 22879 21301 22888 21335
rect 22836 21292 22888 21301
rect 25228 21292 25280 21344
rect 5672 21190 5724 21242
rect 5736 21190 5788 21242
rect 5800 21190 5852 21242
rect 5864 21190 5916 21242
rect 5928 21190 5980 21242
rect 15118 21190 15170 21242
rect 15182 21190 15234 21242
rect 15246 21190 15298 21242
rect 15310 21190 15362 21242
rect 15374 21190 15426 21242
rect 24563 21190 24615 21242
rect 24627 21190 24679 21242
rect 24691 21190 24743 21242
rect 24755 21190 24807 21242
rect 24819 21190 24871 21242
rect 2872 20995 2924 21004
rect 2872 20961 2881 20995
rect 2881 20961 2915 20995
rect 2915 20961 2924 20995
rect 2872 20952 2924 20961
rect 3608 21088 3660 21140
rect 5356 21131 5408 21140
rect 4068 21020 4120 21072
rect 5356 21097 5365 21131
rect 5365 21097 5399 21131
rect 5399 21097 5408 21131
rect 5356 21088 5408 21097
rect 8944 21088 8996 21140
rect 9036 21088 9088 21140
rect 12440 21088 12492 21140
rect 13820 21131 13872 21140
rect 13820 21097 13829 21131
rect 13829 21097 13863 21131
rect 13863 21097 13872 21131
rect 13820 21088 13872 21097
rect 16948 21088 17000 21140
rect 3332 20927 3384 20936
rect 3332 20893 3341 20927
rect 3341 20893 3375 20927
rect 3375 20893 3384 20927
rect 3332 20884 3384 20893
rect 6092 21020 6144 21072
rect 7840 21020 7892 21072
rect 14924 21020 14976 21072
rect 20812 21088 20864 21140
rect 22008 21088 22060 21140
rect 22468 21088 22520 21140
rect 1860 20816 1912 20868
rect 2964 20859 3016 20868
rect 2964 20825 2973 20859
rect 2973 20825 3007 20859
rect 3007 20825 3016 20859
rect 2964 20816 3016 20825
rect 3240 20816 3292 20868
rect 3976 20884 4028 20936
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 4620 20884 4672 20936
rect 5448 20927 5500 20936
rect 1400 20748 1452 20800
rect 3516 20791 3568 20800
rect 3516 20757 3525 20791
rect 3525 20757 3559 20791
rect 3559 20757 3568 20791
rect 3516 20748 3568 20757
rect 4160 20748 4212 20800
rect 5448 20893 5457 20927
rect 5457 20893 5491 20927
rect 5491 20893 5500 20927
rect 5448 20884 5500 20893
rect 6092 20884 6144 20936
rect 6920 20884 6972 20936
rect 7932 20927 7984 20936
rect 7932 20893 7941 20927
rect 7941 20893 7975 20927
rect 7975 20893 7984 20927
rect 7932 20884 7984 20893
rect 9312 20884 9364 20936
rect 12624 20927 12676 20936
rect 12624 20893 12633 20927
rect 12633 20893 12667 20927
rect 12667 20893 12676 20927
rect 12624 20884 12676 20893
rect 13544 20927 13596 20936
rect 13544 20893 13553 20927
rect 13553 20893 13587 20927
rect 13587 20893 13596 20927
rect 13544 20884 13596 20893
rect 14556 20927 14608 20936
rect 4804 20748 4856 20800
rect 9128 20816 9180 20868
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 15200 20884 15252 20936
rect 15660 20884 15712 20936
rect 17960 20952 18012 21004
rect 7472 20748 7524 20800
rect 8116 20791 8168 20800
rect 8116 20757 8125 20791
rect 8125 20757 8159 20791
rect 8159 20757 8168 20791
rect 8116 20748 8168 20757
rect 14096 20816 14148 20868
rect 16120 20859 16172 20868
rect 16120 20825 16129 20859
rect 16129 20825 16163 20859
rect 16163 20825 16172 20859
rect 16120 20816 16172 20825
rect 18052 20816 18104 20868
rect 19064 20952 19116 21004
rect 18788 20884 18840 20936
rect 19340 20884 19392 20936
rect 19616 20884 19668 20936
rect 20720 20927 20772 20936
rect 20720 20893 20729 20927
rect 20729 20893 20763 20927
rect 20763 20893 20772 20927
rect 20720 20884 20772 20893
rect 20904 20884 20956 20936
rect 11520 20748 11572 20800
rect 12992 20791 13044 20800
rect 12992 20757 13001 20791
rect 13001 20757 13035 20791
rect 13035 20757 13044 20791
rect 12992 20748 13044 20757
rect 13636 20748 13688 20800
rect 15476 20748 15528 20800
rect 15752 20748 15804 20800
rect 16672 20791 16724 20800
rect 16672 20757 16681 20791
rect 16681 20757 16715 20791
rect 16715 20757 16724 20791
rect 16672 20748 16724 20757
rect 17408 20748 17460 20800
rect 20812 20816 20864 20868
rect 22192 20884 22244 20936
rect 22652 20952 22704 21004
rect 23388 21020 23440 21072
rect 24124 21020 24176 21072
rect 23112 20952 23164 21004
rect 23204 20884 23256 20936
rect 23940 20884 23992 20936
rect 25596 20816 25648 20868
rect 20352 20748 20404 20800
rect 22192 20748 22244 20800
rect 23112 20748 23164 20800
rect 10395 20646 10447 20698
rect 10459 20646 10511 20698
rect 10523 20646 10575 20698
rect 10587 20646 10639 20698
rect 10651 20646 10703 20698
rect 19840 20646 19892 20698
rect 19904 20646 19956 20698
rect 19968 20646 20020 20698
rect 20032 20646 20084 20698
rect 20096 20646 20148 20698
rect 2412 20587 2464 20596
rect 2412 20553 2421 20587
rect 2421 20553 2455 20587
rect 2455 20553 2464 20587
rect 2412 20544 2464 20553
rect 3056 20544 3108 20596
rect 3976 20587 4028 20596
rect 3976 20553 3985 20587
rect 3985 20553 4019 20587
rect 4019 20553 4028 20587
rect 3976 20544 4028 20553
rect 6368 20544 6420 20596
rect 6460 20587 6512 20596
rect 6460 20553 6469 20587
rect 6469 20553 6503 20587
rect 6503 20553 6512 20587
rect 6920 20587 6972 20596
rect 6460 20544 6512 20553
rect 6920 20553 6929 20587
rect 6929 20553 6963 20587
rect 6963 20553 6972 20587
rect 6920 20544 6972 20553
rect 17316 20587 17368 20596
rect 17316 20553 17325 20587
rect 17325 20553 17359 20587
rect 17359 20553 17368 20587
rect 17316 20544 17368 20553
rect 20352 20544 20404 20596
rect 20812 20544 20864 20596
rect 21548 20544 21600 20596
rect 1860 20519 1912 20528
rect 1860 20485 1869 20519
rect 1869 20485 1903 20519
rect 1903 20485 1912 20519
rect 1860 20476 1912 20485
rect 2964 20476 3016 20528
rect 3332 20476 3384 20528
rect 2872 20408 2924 20460
rect 4252 20476 4304 20528
rect 7472 20476 7524 20528
rect 8116 20476 8168 20528
rect 3608 20451 3660 20460
rect 3608 20417 3617 20451
rect 3617 20417 3651 20451
rect 3651 20417 3660 20451
rect 3608 20408 3660 20417
rect 4160 20408 4212 20460
rect 5264 20408 5316 20460
rect 6644 20408 6696 20460
rect 6736 20408 6788 20460
rect 10048 20408 10100 20460
rect 10692 20451 10744 20460
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 10968 20408 11020 20460
rect 11244 20451 11296 20460
rect 11244 20417 11253 20451
rect 11253 20417 11287 20451
rect 11287 20417 11296 20451
rect 11244 20408 11296 20417
rect 11612 20408 11664 20460
rect 11980 20451 12032 20460
rect 1400 20204 1452 20256
rect 3056 20340 3108 20392
rect 3240 20340 3292 20392
rect 3516 20383 3568 20392
rect 3516 20349 3525 20383
rect 3525 20349 3559 20383
rect 3559 20349 3568 20383
rect 3516 20340 3568 20349
rect 4712 20383 4764 20392
rect 4712 20349 4721 20383
rect 4721 20349 4755 20383
rect 4755 20349 4764 20383
rect 4712 20340 4764 20349
rect 7472 20340 7524 20392
rect 8116 20340 8168 20392
rect 9680 20383 9732 20392
rect 9128 20315 9180 20324
rect 9128 20281 9137 20315
rect 9137 20281 9171 20315
rect 9171 20281 9180 20315
rect 9128 20272 9180 20281
rect 4344 20247 4396 20256
rect 4344 20213 4353 20247
rect 4353 20213 4387 20247
rect 4387 20213 4396 20247
rect 4344 20204 4396 20213
rect 6644 20247 6696 20256
rect 6644 20213 6653 20247
rect 6653 20213 6687 20247
rect 6687 20213 6696 20247
rect 6644 20204 6696 20213
rect 8392 20204 8444 20256
rect 9680 20349 9689 20383
rect 9689 20349 9723 20383
rect 9723 20349 9732 20383
rect 9680 20340 9732 20349
rect 11980 20417 11989 20451
rect 11989 20417 12023 20451
rect 12023 20417 12032 20451
rect 11980 20408 12032 20417
rect 12164 20451 12216 20460
rect 12164 20417 12173 20451
rect 12173 20417 12207 20451
rect 12207 20417 12216 20451
rect 13912 20476 13964 20528
rect 14832 20476 14884 20528
rect 12164 20408 12216 20417
rect 13084 20408 13136 20460
rect 13360 20408 13412 20460
rect 14096 20451 14148 20460
rect 14096 20417 14105 20451
rect 14105 20417 14139 20451
rect 14139 20417 14148 20451
rect 14096 20408 14148 20417
rect 14188 20408 14240 20460
rect 10784 20315 10836 20324
rect 10784 20281 10793 20315
rect 10793 20281 10827 20315
rect 10827 20281 10836 20315
rect 10784 20272 10836 20281
rect 11152 20272 11204 20324
rect 14372 20340 14424 20392
rect 14648 20340 14700 20392
rect 13636 20272 13688 20324
rect 15200 20408 15252 20460
rect 15660 20451 15712 20460
rect 15660 20417 15669 20451
rect 15669 20417 15703 20451
rect 15703 20417 15712 20451
rect 15660 20408 15712 20417
rect 15752 20408 15804 20460
rect 16028 20408 16080 20460
rect 16304 20451 16356 20460
rect 16304 20417 16313 20451
rect 16313 20417 16347 20451
rect 16347 20417 16356 20451
rect 16304 20408 16356 20417
rect 15936 20383 15988 20392
rect 15936 20349 15945 20383
rect 15945 20349 15979 20383
rect 15979 20349 15988 20383
rect 15936 20340 15988 20349
rect 16764 20451 16816 20460
rect 16764 20417 16773 20451
rect 16773 20417 16807 20451
rect 16807 20417 16816 20451
rect 16764 20408 16816 20417
rect 17500 20408 17552 20460
rect 18420 20408 18472 20460
rect 18696 20408 18748 20460
rect 19248 20408 19300 20460
rect 23388 20544 23440 20596
rect 25596 20587 25648 20596
rect 20536 20476 20588 20528
rect 22100 20476 22152 20528
rect 22376 20476 22428 20528
rect 17960 20340 18012 20392
rect 18972 20340 19024 20392
rect 20444 20408 20496 20460
rect 25596 20553 25605 20587
rect 25605 20553 25639 20587
rect 25639 20553 25648 20587
rect 25596 20544 25648 20553
rect 24124 20519 24176 20528
rect 24124 20485 24133 20519
rect 24133 20485 24167 20519
rect 24167 20485 24176 20519
rect 24124 20476 24176 20485
rect 25136 20476 25188 20528
rect 13452 20204 13504 20256
rect 14556 20204 14608 20256
rect 15292 20272 15344 20324
rect 15660 20272 15712 20324
rect 16120 20272 16172 20324
rect 19064 20315 19116 20324
rect 19064 20281 19073 20315
rect 19073 20281 19107 20315
rect 19107 20281 19116 20315
rect 19064 20272 19116 20281
rect 19616 20272 19668 20324
rect 23296 20340 23348 20392
rect 16304 20204 16356 20256
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 17040 20247 17092 20256
rect 17040 20213 17049 20247
rect 17049 20213 17083 20247
rect 17083 20213 17092 20247
rect 17040 20204 17092 20213
rect 18788 20247 18840 20256
rect 18788 20213 18797 20247
rect 18797 20213 18831 20247
rect 18831 20213 18840 20247
rect 20444 20272 20496 20324
rect 18788 20204 18840 20213
rect 5672 20102 5724 20154
rect 5736 20102 5788 20154
rect 5800 20102 5852 20154
rect 5864 20102 5916 20154
rect 5928 20102 5980 20154
rect 15118 20102 15170 20154
rect 15182 20102 15234 20154
rect 15246 20102 15298 20154
rect 15310 20102 15362 20154
rect 15374 20102 15426 20154
rect 24563 20102 24615 20154
rect 24627 20102 24679 20154
rect 24691 20102 24743 20154
rect 24755 20102 24807 20154
rect 24819 20102 24871 20154
rect 2504 20043 2556 20052
rect 2504 20009 2513 20043
rect 2513 20009 2547 20043
rect 2547 20009 2556 20043
rect 2504 20000 2556 20009
rect 2872 20043 2924 20052
rect 2872 20009 2881 20043
rect 2881 20009 2915 20043
rect 2915 20009 2924 20043
rect 2872 20000 2924 20009
rect 5264 20043 5316 20052
rect 5264 20009 5273 20043
rect 5273 20009 5307 20043
rect 5307 20009 5316 20043
rect 5264 20000 5316 20009
rect 7932 20043 7984 20052
rect 7932 20009 7941 20043
rect 7941 20009 7975 20043
rect 7975 20009 7984 20043
rect 7932 20000 7984 20009
rect 8208 20043 8260 20052
rect 8208 20009 8217 20043
rect 8217 20009 8251 20043
rect 8251 20009 8260 20043
rect 8208 20000 8260 20009
rect 11152 20000 11204 20052
rect 11980 20000 12032 20052
rect 13820 20000 13872 20052
rect 15568 20000 15620 20052
rect 15752 20043 15804 20052
rect 15752 20009 15761 20043
rect 15761 20009 15795 20043
rect 15795 20009 15804 20043
rect 15752 20000 15804 20009
rect 16580 20043 16632 20052
rect 16580 20009 16589 20043
rect 16589 20009 16623 20043
rect 16623 20009 16632 20043
rect 16580 20000 16632 20009
rect 18420 20000 18472 20052
rect 22376 20043 22428 20052
rect 22376 20009 22385 20043
rect 22385 20009 22419 20043
rect 22419 20009 22428 20043
rect 22376 20000 22428 20009
rect 23296 20000 23348 20052
rect 24400 20043 24452 20052
rect 24400 20009 24409 20043
rect 24409 20009 24443 20043
rect 24443 20009 24452 20043
rect 24400 20000 24452 20009
rect 25136 20043 25188 20052
rect 25136 20009 25145 20043
rect 25145 20009 25179 20043
rect 25179 20009 25188 20043
rect 25136 20000 25188 20009
rect 4344 19932 4396 19984
rect 4620 19907 4672 19916
rect 4620 19873 4629 19907
rect 4629 19873 4663 19907
rect 4663 19873 4672 19907
rect 4620 19864 4672 19873
rect 3976 19839 4028 19848
rect 3240 19728 3292 19780
rect 3976 19805 3985 19839
rect 3985 19805 4019 19839
rect 4019 19805 4028 19839
rect 3976 19796 4028 19805
rect 6920 19796 6972 19848
rect 7748 19839 7800 19848
rect 7748 19805 7757 19839
rect 7757 19805 7791 19839
rect 7791 19805 7800 19839
rect 7748 19796 7800 19805
rect 8300 19839 8352 19848
rect 8300 19805 8309 19839
rect 8309 19805 8343 19839
rect 8343 19805 8352 19839
rect 8300 19796 8352 19805
rect 10692 19796 10744 19848
rect 11244 19907 11296 19916
rect 11244 19873 11253 19907
rect 11253 19873 11287 19907
rect 11287 19873 11296 19907
rect 11244 19864 11296 19873
rect 11336 19839 11388 19848
rect 11336 19805 11345 19839
rect 11345 19805 11379 19839
rect 11379 19805 11388 19839
rect 11336 19796 11388 19805
rect 11428 19839 11480 19848
rect 11428 19805 11438 19839
rect 11438 19805 11472 19839
rect 11472 19805 11480 19839
rect 11428 19796 11480 19805
rect 11888 19796 11940 19848
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 5356 19728 5408 19780
rect 6368 19728 6420 19780
rect 6644 19771 6696 19780
rect 6644 19737 6653 19771
rect 6653 19737 6687 19771
rect 6687 19737 6696 19771
rect 6644 19728 6696 19737
rect 7288 19728 7340 19780
rect 12716 19728 12768 19780
rect 13176 19771 13228 19780
rect 13176 19737 13185 19771
rect 13185 19737 13219 19771
rect 13219 19737 13228 19771
rect 13176 19728 13228 19737
rect 17040 19932 17092 19984
rect 22560 19932 22612 19984
rect 25044 19932 25096 19984
rect 13544 19864 13596 19916
rect 14372 19864 14424 19916
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 15568 19839 15620 19848
rect 15568 19805 15577 19839
rect 15577 19805 15611 19839
rect 15611 19805 15620 19839
rect 15568 19796 15620 19805
rect 16120 19796 16172 19848
rect 16764 19796 16816 19848
rect 17868 19864 17920 19916
rect 17960 19839 18012 19848
rect 17960 19805 17969 19839
rect 17969 19805 18003 19839
rect 18003 19805 18012 19839
rect 17960 19796 18012 19805
rect 22192 19839 22244 19848
rect 15476 19728 15528 19780
rect 17776 19728 17828 19780
rect 22192 19805 22201 19839
rect 22201 19805 22235 19839
rect 22235 19805 22244 19839
rect 22192 19796 22244 19805
rect 22560 19796 22612 19848
rect 23204 19864 23256 19916
rect 21548 19728 21600 19780
rect 3056 19703 3108 19712
rect 3056 19669 3065 19703
rect 3065 19669 3099 19703
rect 3099 19669 3108 19703
rect 3056 19660 3108 19669
rect 4896 19703 4948 19712
rect 4896 19669 4905 19703
rect 4905 19669 4939 19703
rect 4939 19669 4948 19703
rect 6276 19703 6328 19712
rect 4896 19660 4948 19669
rect 6276 19669 6285 19703
rect 6285 19669 6319 19703
rect 6319 19669 6328 19703
rect 6276 19660 6328 19669
rect 11244 19660 11296 19712
rect 13636 19660 13688 19712
rect 18604 19660 18656 19712
rect 19708 19660 19760 19712
rect 20260 19703 20312 19712
rect 20260 19669 20269 19703
rect 20269 19669 20303 19703
rect 20303 19669 20312 19703
rect 20260 19660 20312 19669
rect 23204 19728 23256 19780
rect 23940 19839 23992 19848
rect 23940 19805 23954 19839
rect 23954 19805 23988 19839
rect 23988 19805 23992 19839
rect 23940 19796 23992 19805
rect 24676 19796 24728 19848
rect 23020 19660 23072 19712
rect 26516 19728 26568 19780
rect 27528 19728 27580 19780
rect 24032 19660 24084 19712
rect 24400 19660 24452 19712
rect 10395 19558 10447 19610
rect 10459 19558 10511 19610
rect 10523 19558 10575 19610
rect 10587 19558 10639 19610
rect 10651 19558 10703 19610
rect 19840 19558 19892 19610
rect 19904 19558 19956 19610
rect 19968 19558 20020 19610
rect 20032 19558 20084 19610
rect 20096 19558 20148 19610
rect 3608 19456 3660 19508
rect 4344 19499 4396 19508
rect 4344 19465 4353 19499
rect 4353 19465 4387 19499
rect 4387 19465 4396 19499
rect 4344 19456 4396 19465
rect 4252 19388 4304 19440
rect 4436 19363 4488 19372
rect 4436 19329 4445 19363
rect 4445 19329 4479 19363
rect 4479 19329 4488 19363
rect 4436 19320 4488 19329
rect 4896 19320 4948 19372
rect 2596 19252 2648 19304
rect 3056 19295 3108 19304
rect 3056 19261 3065 19295
rect 3065 19261 3099 19295
rect 3099 19261 3108 19295
rect 3056 19252 3108 19261
rect 4528 19252 4580 19304
rect 5356 19363 5408 19372
rect 5356 19329 5365 19363
rect 5365 19329 5399 19363
rect 5399 19329 5408 19363
rect 5356 19320 5408 19329
rect 5540 19363 5592 19372
rect 5540 19329 5549 19363
rect 5549 19329 5583 19363
rect 5583 19329 5592 19363
rect 5540 19320 5592 19329
rect 6368 19363 6420 19372
rect 6368 19329 6377 19363
rect 6377 19329 6411 19363
rect 6411 19329 6420 19363
rect 6368 19320 6420 19329
rect 7748 19320 7800 19372
rect 9680 19456 9732 19508
rect 10600 19388 10652 19440
rect 11336 19456 11388 19508
rect 11980 19499 12032 19508
rect 11980 19465 11989 19499
rect 11989 19465 12023 19499
rect 12023 19465 12032 19499
rect 11980 19456 12032 19465
rect 11244 19388 11296 19440
rect 11060 19363 11112 19372
rect 11060 19329 11069 19363
rect 11069 19329 11103 19363
rect 11103 19329 11112 19363
rect 11060 19320 11112 19329
rect 11152 19363 11204 19372
rect 11152 19329 11161 19363
rect 11161 19329 11195 19363
rect 11195 19329 11204 19363
rect 11612 19388 11664 19440
rect 11704 19388 11756 19440
rect 12256 19388 12308 19440
rect 13728 19456 13780 19508
rect 14004 19456 14056 19508
rect 14372 19456 14424 19508
rect 11152 19320 11204 19329
rect 12072 19320 12124 19372
rect 12716 19320 12768 19372
rect 12808 19320 12860 19372
rect 13084 19320 13136 19372
rect 14648 19320 14700 19372
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 15844 19320 15896 19372
rect 18236 19456 18288 19508
rect 19708 19456 19760 19508
rect 20260 19456 20312 19508
rect 20352 19456 20404 19508
rect 24676 19499 24728 19508
rect 24676 19465 24685 19499
rect 24685 19465 24719 19499
rect 24719 19465 24728 19499
rect 24676 19456 24728 19465
rect 26516 19499 26568 19508
rect 26516 19465 26525 19499
rect 26525 19465 26559 19499
rect 26559 19465 26568 19499
rect 26516 19456 26568 19465
rect 17224 19320 17276 19372
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 17960 19320 18012 19372
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 19248 19320 19300 19372
rect 13360 19252 13412 19304
rect 16212 19252 16264 19304
rect 18788 19295 18840 19304
rect 18788 19261 18797 19295
rect 18797 19261 18831 19295
rect 18831 19261 18840 19295
rect 18788 19252 18840 19261
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 19616 19295 19668 19304
rect 19616 19261 19625 19295
rect 19625 19261 19659 19295
rect 19659 19261 19668 19295
rect 19616 19252 19668 19261
rect 20076 19388 20128 19440
rect 19892 19363 19944 19372
rect 19892 19329 19901 19363
rect 19901 19329 19935 19363
rect 19935 19329 19944 19363
rect 19892 19320 19944 19329
rect 20720 19388 20772 19440
rect 23388 19388 23440 19440
rect 25044 19431 25096 19440
rect 20260 19320 20312 19372
rect 24492 19363 24544 19372
rect 24492 19329 24501 19363
rect 24501 19329 24535 19363
rect 24535 19329 24544 19363
rect 24492 19320 24544 19329
rect 25044 19397 25053 19431
rect 25053 19397 25087 19431
rect 25087 19397 25096 19431
rect 25044 19388 25096 19397
rect 26056 19388 26108 19440
rect 2412 19159 2464 19168
rect 2412 19125 2421 19159
rect 2421 19125 2455 19159
rect 2455 19125 2464 19159
rect 2412 19116 2464 19125
rect 5540 19116 5592 19168
rect 8760 19159 8812 19168
rect 8760 19125 8769 19159
rect 8769 19125 8803 19159
rect 8803 19125 8812 19159
rect 8760 19116 8812 19125
rect 18236 19184 18288 19236
rect 12072 19116 12124 19168
rect 12992 19116 13044 19168
rect 17316 19159 17368 19168
rect 17316 19125 17325 19159
rect 17325 19125 17359 19159
rect 17359 19125 17368 19159
rect 17316 19116 17368 19125
rect 19892 19116 19944 19168
rect 20352 19116 20404 19168
rect 5672 19014 5724 19066
rect 5736 19014 5788 19066
rect 5800 19014 5852 19066
rect 5864 19014 5916 19066
rect 5928 19014 5980 19066
rect 15118 19014 15170 19066
rect 15182 19014 15234 19066
rect 15246 19014 15298 19066
rect 15310 19014 15362 19066
rect 15374 19014 15426 19066
rect 24563 19014 24615 19066
rect 24627 19014 24679 19066
rect 24691 19014 24743 19066
rect 24755 19014 24807 19066
rect 24819 19014 24871 19066
rect 2412 18776 2464 18828
rect 2596 18819 2648 18828
rect 2596 18785 2605 18819
rect 2605 18785 2639 18819
rect 2639 18785 2648 18819
rect 2596 18776 2648 18785
rect 2504 18708 2556 18760
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 4804 18708 4856 18760
rect 7748 18819 7800 18828
rect 7748 18785 7757 18819
rect 7757 18785 7791 18819
rect 7791 18785 7800 18819
rect 7748 18776 7800 18785
rect 8208 18776 8260 18828
rect 7472 18708 7524 18760
rect 2688 18615 2740 18624
rect 2688 18581 2697 18615
rect 2697 18581 2731 18615
rect 2731 18581 2740 18615
rect 5540 18640 5592 18692
rect 7564 18640 7616 18692
rect 8024 18708 8076 18760
rect 8668 18844 8720 18896
rect 10876 18844 10928 18896
rect 8576 18776 8628 18828
rect 9956 18776 10008 18828
rect 11428 18844 11480 18896
rect 8668 18640 8720 18692
rect 2688 18572 2740 18581
rect 6276 18572 6328 18624
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 10324 18708 10376 18760
rect 13084 18912 13136 18964
rect 12072 18844 12124 18896
rect 12532 18844 12584 18896
rect 12900 18887 12952 18896
rect 12900 18853 12909 18887
rect 12909 18853 12943 18887
rect 12943 18853 12952 18887
rect 12900 18844 12952 18853
rect 12440 18776 12492 18828
rect 12532 18751 12584 18760
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 12716 18751 12768 18760
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 12716 18708 12768 18717
rect 11704 18640 11756 18692
rect 12992 18751 13044 18760
rect 12992 18717 13001 18751
rect 13001 18717 13035 18751
rect 13035 18717 13044 18751
rect 12992 18708 13044 18717
rect 13544 18776 13596 18828
rect 19248 18912 19300 18964
rect 19524 18912 19576 18964
rect 20076 18912 20128 18964
rect 20444 18912 20496 18964
rect 18788 18844 18840 18896
rect 22560 18955 22612 18964
rect 22560 18921 22569 18955
rect 22569 18921 22603 18955
rect 22603 18921 22612 18955
rect 22560 18912 22612 18921
rect 22928 18912 22980 18964
rect 13452 18751 13504 18760
rect 13452 18717 13461 18751
rect 13461 18717 13495 18751
rect 13495 18717 13504 18751
rect 13452 18708 13504 18717
rect 13636 18708 13688 18760
rect 14188 18751 14240 18760
rect 14188 18717 14197 18751
rect 14197 18717 14231 18751
rect 14231 18717 14240 18751
rect 14188 18708 14240 18717
rect 14648 18776 14700 18828
rect 14372 18751 14424 18760
rect 14372 18717 14396 18751
rect 14396 18717 14424 18751
rect 14372 18708 14424 18717
rect 14556 18751 14608 18760
rect 14556 18717 14565 18751
rect 14565 18717 14599 18751
rect 14599 18717 14608 18751
rect 14556 18708 14608 18717
rect 15476 18751 15528 18760
rect 10876 18572 10928 18624
rect 12716 18572 12768 18624
rect 13084 18572 13136 18624
rect 14832 18640 14884 18692
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 15660 18751 15712 18760
rect 15660 18717 15669 18751
rect 15669 18717 15703 18751
rect 15703 18717 15712 18751
rect 15660 18708 15712 18717
rect 16488 18819 16540 18828
rect 15936 18708 15988 18760
rect 16488 18785 16497 18819
rect 16497 18785 16531 18819
rect 16531 18785 16540 18819
rect 16488 18776 16540 18785
rect 18236 18776 18288 18828
rect 18972 18776 19024 18828
rect 19708 18776 19760 18828
rect 20444 18819 20496 18828
rect 20444 18785 20453 18819
rect 20453 18785 20487 18819
rect 20487 18785 20496 18819
rect 20444 18776 20496 18785
rect 16120 18751 16172 18760
rect 16120 18717 16129 18751
rect 16129 18717 16163 18751
rect 16163 18717 16172 18751
rect 16304 18751 16356 18760
rect 16120 18708 16172 18717
rect 16304 18717 16313 18751
rect 16313 18717 16347 18751
rect 16347 18717 16356 18751
rect 16304 18708 16356 18717
rect 18788 18708 18840 18760
rect 19524 18708 19576 18760
rect 20720 18776 20772 18828
rect 23480 18844 23532 18896
rect 23756 18955 23808 18964
rect 23756 18921 23765 18955
rect 23765 18921 23799 18955
rect 23799 18921 23808 18955
rect 23756 18912 23808 18921
rect 23940 18912 23992 18964
rect 26056 18912 26108 18964
rect 15292 18615 15344 18624
rect 15292 18581 15301 18615
rect 15301 18581 15335 18615
rect 15335 18581 15344 18615
rect 15292 18572 15344 18581
rect 15568 18572 15620 18624
rect 17316 18640 17368 18692
rect 19432 18640 19484 18692
rect 16212 18572 16264 18624
rect 18420 18572 18472 18624
rect 19892 18640 19944 18692
rect 22744 18751 22796 18760
rect 22744 18717 22753 18751
rect 22753 18717 22787 18751
rect 22787 18717 22796 18751
rect 22744 18708 22796 18717
rect 22928 18708 22980 18760
rect 23756 18776 23808 18828
rect 20720 18640 20772 18692
rect 22376 18640 22428 18692
rect 23112 18683 23164 18692
rect 23112 18649 23121 18683
rect 23121 18649 23155 18683
rect 23155 18649 23164 18683
rect 23112 18640 23164 18649
rect 20260 18572 20312 18624
rect 22652 18572 22704 18624
rect 24492 18708 24544 18760
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 10395 18470 10447 18522
rect 10459 18470 10511 18522
rect 10523 18470 10575 18522
rect 10587 18470 10639 18522
rect 10651 18470 10703 18522
rect 19840 18470 19892 18522
rect 19904 18470 19956 18522
rect 19968 18470 20020 18522
rect 20032 18470 20084 18522
rect 20096 18470 20148 18522
rect 1860 18411 1912 18420
rect 1860 18377 1869 18411
rect 1869 18377 1903 18411
rect 1903 18377 1912 18411
rect 1860 18368 1912 18377
rect 2228 18368 2280 18420
rect 2596 18368 2648 18420
rect 2688 18368 2740 18420
rect 4436 18368 4488 18420
rect 7472 18411 7524 18420
rect 7472 18377 7481 18411
rect 7481 18377 7515 18411
rect 7515 18377 7524 18411
rect 7472 18368 7524 18377
rect 2504 18164 2556 18216
rect 4344 18232 4396 18284
rect 4620 18275 4672 18284
rect 4620 18241 4629 18275
rect 4629 18241 4663 18275
rect 4663 18241 4672 18275
rect 4620 18232 4672 18241
rect 6368 18232 6420 18284
rect 7564 18275 7616 18284
rect 7564 18241 7573 18275
rect 7573 18241 7607 18275
rect 7607 18241 7616 18275
rect 7564 18232 7616 18241
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7748 18232 7800 18241
rect 8208 18368 8260 18420
rect 9220 18368 9272 18420
rect 12348 18368 12400 18420
rect 8576 18300 8628 18352
rect 8760 18300 8812 18352
rect 11244 18300 11296 18352
rect 11704 18300 11756 18352
rect 4068 18207 4120 18216
rect 4068 18173 4077 18207
rect 4077 18173 4111 18207
rect 4111 18173 4120 18207
rect 4068 18164 4120 18173
rect 3240 18096 3292 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 2504 18028 2556 18080
rect 3516 18096 3568 18148
rect 10324 18164 10376 18216
rect 11244 18164 11296 18216
rect 11428 18232 11480 18284
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 12624 18300 12676 18352
rect 14188 18368 14240 18420
rect 16304 18368 16356 18420
rect 4528 18096 4580 18148
rect 7840 18139 7892 18148
rect 7840 18105 7849 18139
rect 7849 18105 7883 18139
rect 7883 18105 7892 18139
rect 7840 18096 7892 18105
rect 10048 18096 10100 18148
rect 12072 18164 12124 18216
rect 13176 18232 13228 18284
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 14372 18232 14424 18284
rect 13360 18164 13412 18216
rect 15476 18300 15528 18352
rect 15292 18232 15344 18284
rect 18420 18300 18472 18352
rect 19432 18300 19484 18352
rect 22928 18368 22980 18420
rect 23112 18368 23164 18420
rect 18788 18232 18840 18284
rect 19616 18232 19668 18284
rect 16764 18207 16816 18216
rect 16764 18173 16773 18207
rect 16773 18173 16807 18207
rect 16807 18173 16816 18207
rect 16764 18164 16816 18173
rect 22652 18275 22704 18284
rect 22652 18241 22661 18275
rect 22661 18241 22695 18275
rect 22695 18241 22704 18275
rect 22652 18232 22704 18241
rect 23388 18300 23440 18352
rect 24952 18300 25004 18352
rect 4160 18028 4212 18080
rect 6092 18028 6144 18080
rect 11336 18028 11388 18080
rect 11428 18028 11480 18080
rect 13176 18096 13228 18148
rect 13820 18096 13872 18148
rect 14648 18096 14700 18148
rect 14832 18139 14884 18148
rect 14832 18105 14841 18139
rect 14841 18105 14875 18139
rect 14875 18105 14884 18139
rect 14832 18096 14884 18105
rect 19340 18139 19392 18148
rect 19340 18105 19349 18139
rect 19349 18105 19383 18139
rect 19383 18105 19392 18139
rect 19340 18096 19392 18105
rect 19708 18096 19760 18148
rect 23480 18164 23532 18216
rect 13360 18028 13412 18080
rect 14924 18028 14976 18080
rect 16580 18028 16632 18080
rect 20260 18028 20312 18080
rect 20720 18028 20772 18080
rect 22744 18071 22796 18080
rect 22744 18037 22753 18071
rect 22753 18037 22787 18071
rect 22787 18037 22796 18071
rect 22744 18028 22796 18037
rect 23204 18028 23256 18080
rect 5672 17926 5724 17978
rect 5736 17926 5788 17978
rect 5800 17926 5852 17978
rect 5864 17926 5916 17978
rect 5928 17926 5980 17978
rect 15118 17926 15170 17978
rect 15182 17926 15234 17978
rect 15246 17926 15298 17978
rect 15310 17926 15362 17978
rect 15374 17926 15426 17978
rect 24563 17926 24615 17978
rect 24627 17926 24679 17978
rect 24691 17926 24743 17978
rect 24755 17926 24807 17978
rect 24819 17926 24871 17978
rect 20 17824 72 17876
rect 7196 17824 7248 17876
rect 9220 17867 9272 17876
rect 9220 17833 9229 17867
rect 9229 17833 9263 17867
rect 9263 17833 9272 17867
rect 9220 17824 9272 17833
rect 6644 17799 6696 17808
rect 6644 17765 6653 17799
rect 6653 17765 6687 17799
rect 6687 17765 6696 17799
rect 6644 17756 6696 17765
rect 11704 17824 11756 17876
rect 11980 17867 12032 17876
rect 11980 17833 11989 17867
rect 11989 17833 12023 17867
rect 12023 17833 12032 17867
rect 11980 17824 12032 17833
rect 12440 17867 12492 17876
rect 12440 17833 12449 17867
rect 12449 17833 12483 17867
rect 12483 17833 12492 17867
rect 12440 17824 12492 17833
rect 11060 17756 11112 17808
rect 12808 17824 12860 17876
rect 13452 17824 13504 17876
rect 14832 17824 14884 17876
rect 16304 17824 16356 17876
rect 17592 17824 17644 17876
rect 14188 17799 14240 17808
rect 14188 17765 14197 17799
rect 14197 17765 14231 17799
rect 14231 17765 14240 17799
rect 14188 17756 14240 17765
rect 1492 17552 1544 17604
rect 4712 17620 4764 17672
rect 3792 17552 3844 17604
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 7380 17688 7432 17740
rect 13544 17731 13596 17740
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 13820 17688 13872 17740
rect 16764 17756 16816 17808
rect 17684 17756 17736 17808
rect 6552 17620 6604 17629
rect 6828 17620 6880 17672
rect 7748 17620 7800 17672
rect 2780 17527 2832 17536
rect 2780 17493 2789 17527
rect 2789 17493 2823 17527
rect 2823 17493 2832 17527
rect 2780 17484 2832 17493
rect 3056 17527 3108 17536
rect 3056 17493 3065 17527
rect 3065 17493 3099 17527
rect 3099 17493 3108 17527
rect 3056 17484 3108 17493
rect 3516 17484 3568 17536
rect 5264 17527 5316 17536
rect 5264 17493 5273 17527
rect 5273 17493 5307 17527
rect 5307 17493 5316 17527
rect 5264 17484 5316 17493
rect 6000 17484 6052 17536
rect 7012 17552 7064 17604
rect 8852 17620 8904 17672
rect 10784 17663 10836 17672
rect 10784 17629 10793 17663
rect 10793 17629 10827 17663
rect 10827 17629 10836 17663
rect 10784 17620 10836 17629
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 8116 17527 8168 17536
rect 8116 17493 8125 17527
rect 8125 17493 8159 17527
rect 8159 17493 8168 17527
rect 8116 17484 8168 17493
rect 9496 17552 9548 17604
rect 10324 17552 10376 17604
rect 11244 17620 11296 17672
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 12072 17620 12124 17672
rect 12808 17620 12860 17672
rect 13084 17620 13136 17672
rect 14004 17620 14056 17672
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 16580 17688 16632 17740
rect 14832 17620 14884 17672
rect 16028 17663 16080 17672
rect 16028 17629 16037 17663
rect 16037 17629 16071 17663
rect 16071 17629 16080 17663
rect 16028 17620 16080 17629
rect 16856 17620 16908 17672
rect 17224 17663 17276 17672
rect 9772 17484 9824 17536
rect 10876 17484 10928 17536
rect 13176 17552 13228 17604
rect 11888 17484 11940 17536
rect 13268 17484 13320 17536
rect 14648 17484 14700 17536
rect 16120 17484 16172 17536
rect 16396 17552 16448 17604
rect 17224 17629 17233 17663
rect 17233 17629 17267 17663
rect 17267 17629 17276 17663
rect 17224 17620 17276 17629
rect 18512 17824 18564 17876
rect 19708 17756 19760 17808
rect 19156 17688 19208 17740
rect 19432 17731 19484 17740
rect 19432 17697 19441 17731
rect 19441 17697 19475 17731
rect 19475 17697 19484 17731
rect 19432 17688 19484 17697
rect 20168 17824 20220 17876
rect 22468 17731 22520 17740
rect 22468 17697 22477 17731
rect 22477 17697 22511 17731
rect 22511 17697 22520 17731
rect 22468 17688 22520 17697
rect 23388 17688 23440 17740
rect 24400 17688 24452 17740
rect 18420 17663 18472 17672
rect 18420 17629 18429 17663
rect 18429 17629 18463 17663
rect 18463 17629 18472 17663
rect 18420 17620 18472 17629
rect 18512 17663 18564 17672
rect 18512 17629 18521 17663
rect 18521 17629 18555 17663
rect 18555 17629 18564 17663
rect 18512 17620 18564 17629
rect 20168 17663 20220 17672
rect 20168 17629 20177 17663
rect 20177 17629 20211 17663
rect 20211 17629 20220 17663
rect 20168 17620 20220 17629
rect 20352 17663 20404 17672
rect 20352 17629 20360 17663
rect 20360 17629 20394 17663
rect 20394 17629 20404 17663
rect 20352 17620 20404 17629
rect 20536 17663 20588 17672
rect 20536 17629 20545 17663
rect 20545 17629 20579 17663
rect 20579 17629 20588 17663
rect 20536 17620 20588 17629
rect 22652 17620 22704 17672
rect 23204 17663 23256 17672
rect 23204 17629 23213 17663
rect 23213 17629 23247 17663
rect 23247 17629 23256 17663
rect 23204 17620 23256 17629
rect 17316 17484 17368 17536
rect 18144 17527 18196 17536
rect 18144 17493 18153 17527
rect 18153 17493 18187 17527
rect 18187 17493 18196 17527
rect 18144 17484 18196 17493
rect 19340 17484 19392 17536
rect 24860 17595 24912 17604
rect 24860 17561 24869 17595
rect 24869 17561 24903 17595
rect 24903 17561 24912 17595
rect 24860 17552 24912 17561
rect 25504 17552 25556 17604
rect 23204 17484 23256 17536
rect 24216 17484 24268 17536
rect 24768 17484 24820 17536
rect 10395 17382 10447 17434
rect 10459 17382 10511 17434
rect 10523 17382 10575 17434
rect 10587 17382 10639 17434
rect 10651 17382 10703 17434
rect 19840 17382 19892 17434
rect 19904 17382 19956 17434
rect 19968 17382 20020 17434
rect 20032 17382 20084 17434
rect 20096 17382 20148 17434
rect 2228 17323 2280 17332
rect 2228 17289 2237 17323
rect 2237 17289 2271 17323
rect 2271 17289 2280 17323
rect 2228 17280 2280 17289
rect 2780 17280 2832 17332
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 7012 17280 7064 17332
rect 7196 17280 7248 17332
rect 7564 17323 7616 17332
rect 7564 17289 7573 17323
rect 7573 17289 7607 17323
rect 7607 17289 7616 17323
rect 7564 17280 7616 17289
rect 7656 17280 7708 17332
rect 8852 17323 8904 17332
rect 3148 17144 3200 17196
rect 5264 17212 5316 17264
rect 6828 17255 6880 17264
rect 6828 17221 6837 17255
rect 6837 17221 6871 17255
rect 6871 17221 6880 17255
rect 6828 17212 6880 17221
rect 4896 17144 4948 17196
rect 5540 17144 5592 17196
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 7104 17144 7156 17196
rect 7196 17187 7248 17196
rect 7196 17153 7205 17187
rect 7205 17153 7239 17187
rect 7239 17153 7248 17187
rect 7472 17187 7524 17196
rect 7196 17144 7248 17153
rect 7472 17153 7495 17187
rect 7495 17153 7524 17187
rect 7472 17144 7524 17153
rect 7840 17187 7892 17196
rect 4252 17119 4304 17128
rect 4252 17085 4261 17119
rect 4261 17085 4295 17119
rect 4295 17085 4304 17119
rect 4252 17076 4304 17085
rect 4436 17119 4488 17128
rect 4436 17085 4445 17119
rect 4445 17085 4479 17119
rect 4479 17085 4488 17119
rect 4436 17076 4488 17085
rect 6920 17076 6972 17128
rect 7840 17153 7849 17187
rect 7849 17153 7883 17187
rect 7883 17153 7892 17187
rect 7840 17144 7892 17153
rect 8852 17289 8861 17323
rect 8861 17289 8895 17323
rect 8895 17289 8904 17323
rect 8852 17280 8904 17289
rect 9220 17280 9272 17332
rect 10784 17323 10836 17332
rect 10784 17289 10793 17323
rect 10793 17289 10827 17323
rect 10827 17289 10836 17323
rect 10784 17280 10836 17289
rect 11244 17280 11296 17332
rect 12072 17280 12124 17332
rect 12348 17280 12400 17332
rect 13544 17280 13596 17332
rect 2964 17008 3016 17060
rect 1308 16940 1360 16992
rect 7380 17008 7432 17060
rect 3792 16983 3844 16992
rect 3792 16949 3801 16983
rect 3801 16949 3835 16983
rect 3835 16949 3844 16983
rect 3792 16940 3844 16949
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 4896 16940 4948 16949
rect 6644 16940 6696 16992
rect 7472 16940 7524 16992
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 8024 17076 8076 17128
rect 9220 17144 9272 17196
rect 10324 17212 10376 17264
rect 14004 17280 14056 17332
rect 15016 17323 15068 17332
rect 15016 17289 15025 17323
rect 15025 17289 15059 17323
rect 15059 17289 15068 17323
rect 15016 17280 15068 17289
rect 9956 17144 10008 17196
rect 10968 17144 11020 17196
rect 11520 17187 11572 17196
rect 11520 17153 11529 17187
rect 11529 17153 11563 17187
rect 11563 17153 11572 17187
rect 11520 17144 11572 17153
rect 12624 17144 12676 17196
rect 13084 17187 13136 17196
rect 8484 17076 8536 17128
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 13360 17187 13412 17196
rect 13360 17153 13369 17187
rect 13369 17153 13403 17187
rect 13403 17153 13412 17187
rect 13360 17144 13412 17153
rect 13544 17187 13596 17196
rect 13544 17153 13553 17187
rect 13553 17153 13587 17187
rect 13587 17153 13596 17187
rect 13544 17144 13596 17153
rect 18052 17280 18104 17332
rect 18788 17280 18840 17332
rect 19708 17280 19760 17332
rect 20352 17280 20404 17332
rect 21180 17280 21232 17332
rect 25504 17323 25556 17332
rect 25504 17289 25513 17323
rect 25513 17289 25547 17323
rect 25547 17289 25556 17323
rect 25504 17280 25556 17289
rect 25688 17280 25740 17332
rect 15936 17212 15988 17264
rect 14648 17144 14700 17196
rect 14740 17076 14792 17128
rect 14648 17008 14700 17060
rect 16212 17144 16264 17196
rect 16764 17212 16816 17264
rect 18144 17212 18196 17264
rect 19156 17212 19208 17264
rect 23848 17212 23900 17264
rect 24216 17212 24268 17264
rect 24768 17255 24820 17264
rect 16580 17144 16632 17196
rect 17224 17144 17276 17196
rect 17960 17187 18012 17196
rect 17960 17153 17969 17187
rect 17969 17153 18003 17187
rect 18003 17153 18012 17187
rect 17960 17144 18012 17153
rect 18236 17187 18288 17196
rect 18236 17153 18245 17187
rect 18245 17153 18279 17187
rect 18279 17153 18288 17187
rect 18236 17144 18288 17153
rect 15660 17076 15712 17128
rect 16856 17076 16908 17128
rect 24768 17221 24777 17255
rect 24777 17221 24811 17255
rect 24811 17221 24820 17255
rect 24768 17212 24820 17221
rect 24952 17187 25004 17196
rect 24952 17153 24955 17187
rect 24955 17153 25004 17187
rect 22652 17119 22704 17128
rect 22652 17085 22661 17119
rect 22661 17085 22695 17119
rect 22695 17085 22704 17119
rect 22652 17076 22704 17085
rect 23480 17076 23532 17128
rect 24400 17119 24452 17128
rect 24400 17085 24409 17119
rect 24409 17085 24443 17119
rect 24443 17085 24452 17119
rect 24400 17076 24452 17085
rect 24952 17144 25004 17153
rect 25320 17187 25372 17196
rect 25320 17153 25329 17187
rect 25329 17153 25363 17187
rect 25363 17153 25372 17187
rect 25320 17144 25372 17153
rect 25688 17076 25740 17128
rect 16580 17008 16632 17060
rect 8576 16940 8628 16992
rect 9312 16940 9364 16992
rect 9772 16940 9824 16992
rect 11796 16940 11848 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 17776 16983 17828 16992
rect 17776 16949 17785 16983
rect 17785 16949 17819 16983
rect 17819 16949 17828 16983
rect 17776 16940 17828 16949
rect 24860 17008 24912 17060
rect 24308 16940 24360 16992
rect 5672 16838 5724 16890
rect 5736 16838 5788 16890
rect 5800 16838 5852 16890
rect 5864 16838 5916 16890
rect 5928 16838 5980 16890
rect 15118 16838 15170 16890
rect 15182 16838 15234 16890
rect 15246 16838 15298 16890
rect 15310 16838 15362 16890
rect 15374 16838 15426 16890
rect 24563 16838 24615 16890
rect 24627 16838 24679 16890
rect 24691 16838 24743 16890
rect 24755 16838 24807 16890
rect 24819 16838 24871 16890
rect 3056 16736 3108 16788
rect 2872 16668 2924 16720
rect 3148 16668 3200 16720
rect 2964 16600 3016 16652
rect 4712 16600 4764 16652
rect 8208 16736 8260 16788
rect 8576 16779 8628 16788
rect 8576 16745 8585 16779
rect 8585 16745 8619 16779
rect 8619 16745 8628 16779
rect 8576 16736 8628 16745
rect 12992 16779 13044 16788
rect 12992 16745 13001 16779
rect 13001 16745 13035 16779
rect 13035 16745 13044 16779
rect 12992 16736 13044 16745
rect 13268 16779 13320 16788
rect 13268 16745 13277 16779
rect 13277 16745 13311 16779
rect 13311 16745 13320 16779
rect 13268 16736 13320 16745
rect 13544 16779 13596 16788
rect 7012 16711 7064 16720
rect 7012 16677 7021 16711
rect 7021 16677 7055 16711
rect 7055 16677 7064 16711
rect 7012 16668 7064 16677
rect 8024 16668 8076 16720
rect 9220 16668 9272 16720
rect 9956 16711 10008 16720
rect 7840 16600 7892 16652
rect 8484 16600 8536 16652
rect 9312 16643 9364 16652
rect 9312 16609 9321 16643
rect 9321 16609 9355 16643
rect 9355 16609 9364 16643
rect 9312 16600 9364 16609
rect 9956 16677 9965 16711
rect 9965 16677 9999 16711
rect 9999 16677 10008 16711
rect 9956 16668 10008 16677
rect 9680 16600 9732 16652
rect 2780 16575 2832 16584
rect 2780 16541 2789 16575
rect 2789 16541 2823 16575
rect 2823 16541 2832 16575
rect 2780 16532 2832 16541
rect 2504 16464 2556 16516
rect 4436 16532 4488 16584
rect 5264 16532 5316 16584
rect 6000 16532 6052 16584
rect 4896 16464 4948 16516
rect 7564 16532 7616 16584
rect 8576 16532 8628 16584
rect 8852 16532 8904 16584
rect 10876 16532 10928 16584
rect 11244 16575 11296 16584
rect 11244 16541 11253 16575
rect 11253 16541 11287 16575
rect 11287 16541 11296 16575
rect 11244 16532 11296 16541
rect 11428 16575 11480 16584
rect 11428 16541 11437 16575
rect 11437 16541 11471 16575
rect 11471 16541 11480 16575
rect 11428 16532 11480 16541
rect 4252 16439 4304 16448
rect 4252 16405 4261 16439
rect 4261 16405 4295 16439
rect 4295 16405 4304 16439
rect 4252 16396 4304 16405
rect 4712 16439 4764 16448
rect 4712 16405 4721 16439
rect 4721 16405 4755 16439
rect 4755 16405 4764 16439
rect 7472 16464 7524 16516
rect 4712 16396 4764 16405
rect 7380 16396 7432 16448
rect 8300 16464 8352 16516
rect 11336 16464 11388 16516
rect 12256 16532 12308 16584
rect 13176 16600 13228 16652
rect 13544 16745 13553 16779
rect 13553 16745 13587 16779
rect 13587 16745 13596 16779
rect 13544 16736 13596 16745
rect 14648 16736 14700 16788
rect 15016 16736 15068 16788
rect 19708 16736 19760 16788
rect 18512 16711 18564 16720
rect 18512 16677 18521 16711
rect 18521 16677 18555 16711
rect 18555 16677 18564 16711
rect 18512 16668 18564 16677
rect 12808 16532 12860 16584
rect 13360 16575 13412 16584
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 12440 16464 12492 16516
rect 13268 16464 13320 16516
rect 13544 16532 13596 16584
rect 15476 16600 15528 16652
rect 18236 16600 18288 16652
rect 14832 16575 14884 16584
rect 14832 16541 14841 16575
rect 14841 16541 14875 16575
rect 14875 16541 14884 16575
rect 14832 16532 14884 16541
rect 17316 16532 17368 16584
rect 17776 16532 17828 16584
rect 20168 16668 20220 16720
rect 20352 16736 20404 16788
rect 22652 16779 22704 16788
rect 22652 16745 22661 16779
rect 22661 16745 22695 16779
rect 22695 16745 22704 16779
rect 22652 16736 22704 16745
rect 23480 16736 23532 16788
rect 23848 16779 23900 16788
rect 23848 16745 23857 16779
rect 23857 16745 23891 16779
rect 23891 16745 23900 16779
rect 23848 16736 23900 16745
rect 25320 16736 25372 16788
rect 20536 16668 20588 16720
rect 20168 16575 20220 16584
rect 14464 16439 14516 16448
rect 14464 16405 14473 16439
rect 14473 16405 14507 16439
rect 14507 16405 14516 16439
rect 14464 16396 14516 16405
rect 15660 16464 15712 16516
rect 16120 16464 16172 16516
rect 20168 16541 20176 16575
rect 20176 16541 20210 16575
rect 20210 16541 20220 16575
rect 20168 16532 20220 16541
rect 22468 16600 22520 16652
rect 16672 16396 16724 16448
rect 17224 16396 17276 16448
rect 20444 16464 20496 16516
rect 18420 16396 18472 16448
rect 19432 16396 19484 16448
rect 23388 16532 23440 16584
rect 23480 16464 23532 16516
rect 23572 16396 23624 16448
rect 24308 16532 24360 16584
rect 24492 16464 24544 16516
rect 24124 16439 24176 16448
rect 24124 16405 24133 16439
rect 24133 16405 24167 16439
rect 24167 16405 24176 16439
rect 24584 16439 24636 16448
rect 24124 16396 24176 16405
rect 24584 16405 24593 16439
rect 24593 16405 24627 16439
rect 24627 16405 24636 16439
rect 24584 16396 24636 16405
rect 26148 16396 26200 16448
rect 10395 16294 10447 16346
rect 10459 16294 10511 16346
rect 10523 16294 10575 16346
rect 10587 16294 10639 16346
rect 10651 16294 10703 16346
rect 19840 16294 19892 16346
rect 19904 16294 19956 16346
rect 19968 16294 20020 16346
rect 20032 16294 20084 16346
rect 20096 16294 20148 16346
rect 4528 16192 4580 16244
rect 4712 16192 4764 16244
rect 5356 16192 5408 16244
rect 2228 16124 2280 16176
rect 2136 16099 2188 16108
rect 2136 16065 2145 16099
rect 2145 16065 2179 16099
rect 2179 16065 2188 16099
rect 2136 16056 2188 16065
rect 2504 15988 2556 16040
rect 2964 15920 3016 15972
rect 3792 16124 3844 16176
rect 3976 16124 4028 16176
rect 3608 16056 3660 16108
rect 4160 16056 4212 16108
rect 4896 16056 4948 16108
rect 5264 16056 5316 16108
rect 7104 16192 7156 16244
rect 7840 16167 7892 16176
rect 7840 16133 7849 16167
rect 7849 16133 7883 16167
rect 7883 16133 7892 16167
rect 8668 16192 8720 16244
rect 9496 16192 9548 16244
rect 16028 16192 16080 16244
rect 18328 16192 18380 16244
rect 18880 16192 18932 16244
rect 19432 16235 19484 16244
rect 19432 16201 19441 16235
rect 19441 16201 19475 16235
rect 19475 16201 19484 16235
rect 19432 16192 19484 16201
rect 7840 16124 7892 16133
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 8392 16056 8444 16108
rect 14648 16124 14700 16176
rect 14740 16167 14792 16176
rect 14740 16133 14749 16167
rect 14749 16133 14783 16167
rect 14783 16133 14792 16167
rect 14740 16124 14792 16133
rect 17592 16124 17644 16176
rect 20536 16192 20588 16244
rect 21180 16192 21232 16244
rect 23204 16192 23256 16244
rect 23388 16192 23440 16244
rect 23572 16192 23624 16244
rect 24216 16192 24268 16244
rect 26148 16192 26200 16244
rect 23664 16124 23716 16176
rect 24124 16124 24176 16176
rect 8760 16056 8812 16108
rect 9496 16099 9548 16108
rect 3516 16031 3568 16040
rect 3516 15997 3525 16031
rect 3525 15997 3559 16031
rect 3559 15997 3568 16031
rect 3516 15988 3568 15997
rect 5448 15988 5500 16040
rect 6092 15988 6144 16040
rect 6736 15988 6788 16040
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 15844 16056 15896 16108
rect 18052 16056 18104 16108
rect 18420 16056 18472 16108
rect 19248 16056 19300 16108
rect 10140 15988 10192 16040
rect 14372 15988 14424 16040
rect 15476 15988 15528 16040
rect 18788 16031 18840 16040
rect 18788 15997 18797 16031
rect 18797 15997 18831 16031
rect 18831 15997 18840 16031
rect 18788 15988 18840 15997
rect 18880 15988 18932 16040
rect 20444 16056 20496 16108
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 24400 16056 24452 16108
rect 25228 16031 25280 16040
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 2320 15852 2372 15904
rect 13360 15920 13412 15972
rect 3884 15852 3936 15904
rect 6552 15852 6604 15904
rect 7656 15895 7708 15904
rect 7656 15861 7665 15895
rect 7665 15861 7699 15895
rect 7699 15861 7708 15895
rect 7656 15852 7708 15861
rect 7748 15852 7800 15904
rect 8024 15852 8076 15904
rect 8484 15852 8536 15904
rect 8760 15895 8812 15904
rect 8760 15861 8769 15895
rect 8769 15861 8803 15895
rect 8803 15861 8812 15895
rect 8760 15852 8812 15861
rect 9680 15895 9732 15904
rect 9680 15861 9689 15895
rect 9689 15861 9723 15895
rect 9723 15861 9732 15895
rect 9680 15852 9732 15861
rect 13268 15895 13320 15904
rect 13268 15861 13277 15895
rect 13277 15861 13311 15895
rect 13311 15861 13320 15895
rect 13268 15852 13320 15861
rect 14924 15852 14976 15904
rect 17960 15852 18012 15904
rect 18788 15852 18840 15904
rect 19156 15852 19208 15904
rect 25228 15997 25237 16031
rect 25237 15997 25271 16031
rect 25271 15997 25280 16031
rect 25228 15988 25280 15997
rect 20444 15920 20496 15972
rect 20352 15852 20404 15904
rect 20628 15895 20680 15904
rect 20628 15861 20637 15895
rect 20637 15861 20671 15895
rect 20671 15861 20680 15895
rect 20628 15852 20680 15861
rect 26792 15852 26844 15904
rect 5672 15750 5724 15802
rect 5736 15750 5788 15802
rect 5800 15750 5852 15802
rect 5864 15750 5916 15802
rect 5928 15750 5980 15802
rect 15118 15750 15170 15802
rect 15182 15750 15234 15802
rect 15246 15750 15298 15802
rect 15310 15750 15362 15802
rect 15374 15750 15426 15802
rect 24563 15750 24615 15802
rect 24627 15750 24679 15802
rect 24691 15750 24743 15802
rect 24755 15750 24807 15802
rect 24819 15750 24871 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 2964 15691 3016 15700
rect 2964 15657 2973 15691
rect 2973 15657 3007 15691
rect 3007 15657 3016 15691
rect 2964 15648 3016 15657
rect 3516 15648 3568 15700
rect 1584 15580 1636 15632
rect 6552 15648 6604 15700
rect 4160 15623 4212 15632
rect 4160 15589 4169 15623
rect 4169 15589 4203 15623
rect 4203 15589 4212 15623
rect 4160 15580 4212 15589
rect 3884 15555 3936 15564
rect 3884 15521 3893 15555
rect 3893 15521 3927 15555
rect 3927 15521 3936 15555
rect 3884 15512 3936 15521
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 2780 15487 2832 15496
rect 2780 15453 2789 15487
rect 2789 15453 2823 15487
rect 2823 15453 2832 15487
rect 2780 15444 2832 15453
rect 4252 15444 4304 15496
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 7104 15580 7156 15632
rect 7288 15555 7340 15564
rect 7288 15521 7297 15555
rect 7297 15521 7331 15555
rect 7331 15521 7340 15555
rect 7288 15512 7340 15521
rect 7104 15444 7156 15496
rect 7380 15487 7432 15496
rect 7380 15453 7390 15487
rect 7390 15453 7424 15487
rect 7424 15453 7432 15487
rect 7380 15444 7432 15453
rect 7748 15487 7800 15496
rect 7472 15376 7524 15428
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 8300 15648 8352 15700
rect 10048 15648 10100 15700
rect 10968 15648 11020 15700
rect 11060 15648 11112 15700
rect 11612 15648 11664 15700
rect 12624 15648 12676 15700
rect 14648 15691 14700 15700
rect 14648 15657 14657 15691
rect 14657 15657 14691 15691
rect 14691 15657 14700 15691
rect 14648 15648 14700 15657
rect 17592 15648 17644 15700
rect 17868 15648 17920 15700
rect 18880 15648 18932 15700
rect 20536 15648 20588 15700
rect 24492 15648 24544 15700
rect 25228 15648 25280 15700
rect 8024 15580 8076 15632
rect 8116 15512 8168 15564
rect 8024 15487 8076 15496
rect 8024 15453 8033 15487
rect 8033 15453 8067 15487
rect 8067 15453 8076 15487
rect 10968 15555 11020 15564
rect 10968 15521 10977 15555
rect 10977 15521 11011 15555
rect 11011 15521 11020 15555
rect 10968 15512 11020 15521
rect 11336 15512 11388 15564
rect 17132 15512 17184 15564
rect 8024 15444 8076 15453
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 8668 15444 8720 15496
rect 14924 15444 14976 15496
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 18144 15512 18196 15564
rect 19248 15512 19300 15564
rect 9404 15376 9456 15428
rect 10324 15376 10376 15428
rect 11704 15376 11756 15428
rect 12532 15376 12584 15428
rect 17316 15376 17368 15428
rect 17960 15376 18012 15428
rect 18420 15444 18472 15496
rect 20628 15444 20680 15496
rect 21640 15487 21692 15496
rect 21640 15453 21649 15487
rect 21649 15453 21683 15487
rect 21683 15453 21692 15487
rect 21640 15444 21692 15453
rect 23572 15487 23624 15496
rect 23572 15453 23581 15487
rect 23581 15453 23615 15487
rect 23615 15453 23624 15487
rect 23572 15444 23624 15453
rect 24032 15580 24084 15632
rect 25044 15580 25096 15632
rect 26516 15512 26568 15564
rect 18604 15376 18656 15428
rect 22008 15419 22060 15428
rect 22008 15385 22042 15419
rect 22042 15385 22060 15419
rect 22008 15376 22060 15385
rect 23204 15376 23256 15428
rect 24308 15444 24360 15496
rect 24860 15444 24912 15496
rect 26792 15444 26844 15496
rect 4988 15308 5040 15360
rect 8576 15308 8628 15360
rect 17132 15308 17184 15360
rect 18328 15351 18380 15360
rect 18328 15317 18337 15351
rect 18337 15317 18371 15351
rect 18371 15317 18380 15351
rect 18328 15308 18380 15317
rect 22284 15308 22336 15360
rect 24216 15308 24268 15360
rect 25136 15308 25188 15360
rect 25412 15308 25464 15360
rect 10395 15206 10447 15258
rect 10459 15206 10511 15258
rect 10523 15206 10575 15258
rect 10587 15206 10639 15258
rect 10651 15206 10703 15258
rect 19840 15206 19892 15258
rect 19904 15206 19956 15258
rect 19968 15206 20020 15258
rect 20032 15206 20084 15258
rect 20096 15206 20148 15258
rect 3240 15104 3292 15156
rect 7380 15104 7432 15156
rect 7840 15104 7892 15156
rect 8024 15104 8076 15156
rect 8300 15104 8352 15156
rect 10324 15104 10376 15156
rect 11704 15147 11756 15156
rect 11704 15113 11713 15147
rect 11713 15113 11747 15147
rect 11747 15113 11756 15147
rect 11704 15104 11756 15113
rect 12624 15104 12676 15156
rect 1768 15036 1820 15088
rect 4160 15036 4212 15088
rect 6920 15036 6972 15088
rect 4988 15011 5040 15020
rect 4988 14977 4997 15011
rect 4997 14977 5031 15011
rect 5031 14977 5040 15011
rect 4988 14968 5040 14977
rect 7840 15011 7892 15020
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 3424 14943 3476 14952
rect 3424 14909 3433 14943
rect 3433 14909 3467 14943
rect 3467 14909 3476 14943
rect 3424 14900 3476 14909
rect 2964 14875 3016 14884
rect 2964 14841 2973 14875
rect 2973 14841 3007 14875
rect 3007 14841 3016 14875
rect 2964 14832 3016 14841
rect 4436 14900 4488 14952
rect 4620 14832 4672 14884
rect 3976 14807 4028 14816
rect 3976 14773 3985 14807
rect 3985 14773 4019 14807
rect 4019 14773 4028 14807
rect 3976 14764 4028 14773
rect 7840 14977 7849 15011
rect 7849 14977 7883 15011
rect 7883 14977 7892 15011
rect 7840 14968 7892 14977
rect 9312 15011 9364 15020
rect 7288 14943 7340 14952
rect 7288 14909 7297 14943
rect 7297 14909 7331 14943
rect 7331 14909 7340 14943
rect 7288 14900 7340 14909
rect 9312 14977 9321 15011
rect 9321 14977 9355 15011
rect 9355 14977 9364 15011
rect 13268 15036 13320 15088
rect 9312 14968 9364 14977
rect 10048 15011 10100 15020
rect 10048 14977 10057 15011
rect 10057 14977 10091 15011
rect 10091 14977 10100 15011
rect 10048 14968 10100 14977
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 10876 14968 10928 15020
rect 8668 14832 8720 14884
rect 9496 14832 9548 14884
rect 11980 14968 12032 15020
rect 12532 14968 12584 15020
rect 12808 15011 12860 15020
rect 12808 14977 12822 15011
rect 12822 14977 12856 15011
rect 12856 14977 12860 15011
rect 12808 14968 12860 14977
rect 7104 14764 7156 14816
rect 8300 14764 8352 14816
rect 9036 14764 9088 14816
rect 11428 14764 11480 14816
rect 12624 14764 12676 14816
rect 13268 14900 13320 14952
rect 14924 14968 14976 15020
rect 15568 15011 15620 15020
rect 15568 14977 15577 15011
rect 15577 14977 15611 15011
rect 15611 14977 15620 15011
rect 15568 14968 15620 14977
rect 17316 15147 17368 15156
rect 17316 15113 17325 15147
rect 17325 15113 17359 15147
rect 17359 15113 17368 15147
rect 17316 15104 17368 15113
rect 18604 15104 18656 15156
rect 19248 15147 19300 15156
rect 19248 15113 19257 15147
rect 19257 15113 19291 15147
rect 19291 15113 19300 15147
rect 19248 15104 19300 15113
rect 19340 15104 19392 15156
rect 22376 15104 22428 15156
rect 23940 15104 23992 15156
rect 24032 15104 24084 15156
rect 16120 15036 16172 15088
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 17592 14968 17644 15020
rect 18328 15036 18380 15088
rect 25044 15079 25096 15088
rect 17960 14968 18012 15020
rect 18972 14968 19024 15020
rect 16948 14943 17000 14952
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 21180 14943 21232 14952
rect 21180 14909 21189 14943
rect 21189 14909 21223 14943
rect 21223 14909 21232 14943
rect 21180 14900 21232 14909
rect 21640 14900 21692 14952
rect 22560 14968 22612 15020
rect 24492 15011 24544 15020
rect 24492 14977 24501 15011
rect 24501 14977 24535 15011
rect 24535 14977 24544 15011
rect 24492 14968 24544 14977
rect 25044 15045 25053 15079
rect 25053 15045 25087 15079
rect 25087 15045 25096 15079
rect 25044 15036 25096 15045
rect 25596 15036 25648 15088
rect 16672 14764 16724 14816
rect 17132 14764 17184 14816
rect 25412 14764 25464 14816
rect 26516 14807 26568 14816
rect 26516 14773 26525 14807
rect 26525 14773 26559 14807
rect 26559 14773 26568 14807
rect 26516 14764 26568 14773
rect 5672 14662 5724 14714
rect 5736 14662 5788 14714
rect 5800 14662 5852 14714
rect 5864 14662 5916 14714
rect 5928 14662 5980 14714
rect 15118 14662 15170 14714
rect 15182 14662 15234 14714
rect 15246 14662 15298 14714
rect 15310 14662 15362 14714
rect 15374 14662 15426 14714
rect 24563 14662 24615 14714
rect 24627 14662 24679 14714
rect 24691 14662 24743 14714
rect 24755 14662 24807 14714
rect 24819 14662 24871 14714
rect 3424 14560 3476 14612
rect 4160 14560 4212 14612
rect 5540 14560 5592 14612
rect 10784 14603 10836 14612
rect 4068 14492 4120 14544
rect 6184 14492 6236 14544
rect 4620 14424 4672 14476
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 3148 14356 3200 14408
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 5264 14356 5316 14408
rect 6920 14356 6972 14408
rect 7748 14356 7800 14408
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 5080 14288 5132 14340
rect 9680 14356 9732 14408
rect 10784 14569 10793 14603
rect 10793 14569 10827 14603
rect 10827 14569 10836 14603
rect 10784 14560 10836 14569
rect 11612 14492 11664 14544
rect 10784 14356 10836 14408
rect 11612 14356 11664 14408
rect 5632 14220 5684 14272
rect 7012 14263 7064 14272
rect 7012 14229 7021 14263
rect 7021 14229 7055 14263
rect 7055 14229 7064 14263
rect 7012 14220 7064 14229
rect 7196 14220 7248 14272
rect 7748 14220 7800 14272
rect 11428 14288 11480 14340
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 10876 14220 10928 14272
rect 11796 14263 11848 14272
rect 11796 14229 11805 14263
rect 11805 14229 11839 14263
rect 11839 14229 11848 14263
rect 11796 14220 11848 14229
rect 13176 14424 13228 14476
rect 13268 14424 13320 14476
rect 17040 14560 17092 14612
rect 18972 14603 19024 14612
rect 18972 14569 18981 14603
rect 18981 14569 19015 14603
rect 19015 14569 19024 14603
rect 18972 14560 19024 14569
rect 19616 14560 19668 14612
rect 22008 14603 22060 14612
rect 14280 14492 14332 14544
rect 16580 14492 16632 14544
rect 16948 14492 17000 14544
rect 18144 14492 18196 14544
rect 17684 14424 17736 14476
rect 13820 14399 13872 14408
rect 13820 14365 13829 14399
rect 13829 14365 13863 14399
rect 13863 14365 13872 14399
rect 13820 14356 13872 14365
rect 15568 14356 15620 14408
rect 16580 14399 16632 14408
rect 12532 14220 12584 14272
rect 12992 14288 13044 14340
rect 13728 14288 13780 14340
rect 16212 14288 16264 14340
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 16580 14356 16632 14365
rect 17224 14356 17276 14408
rect 17776 14356 17828 14408
rect 18052 14356 18104 14408
rect 18328 14399 18380 14408
rect 18328 14365 18337 14399
rect 18337 14365 18371 14399
rect 18371 14365 18380 14399
rect 18328 14356 18380 14365
rect 16856 14288 16908 14340
rect 18604 14288 18656 14340
rect 19064 14356 19116 14408
rect 19156 14356 19208 14408
rect 19340 14356 19392 14408
rect 22008 14569 22017 14603
rect 22017 14569 22051 14603
rect 22051 14569 22060 14603
rect 22008 14560 22060 14569
rect 25596 14603 25648 14612
rect 25596 14569 25605 14603
rect 25605 14569 25639 14603
rect 25639 14569 25648 14603
rect 25596 14560 25648 14569
rect 21640 14492 21692 14544
rect 22376 14535 22428 14544
rect 22376 14501 22385 14535
rect 22385 14501 22419 14535
rect 22419 14501 22428 14535
rect 22376 14492 22428 14501
rect 20168 14467 20220 14476
rect 20168 14433 20177 14467
rect 20177 14433 20211 14467
rect 20211 14433 20220 14467
rect 20168 14424 20220 14433
rect 26700 14424 26752 14476
rect 21548 14356 21600 14408
rect 21824 14399 21876 14408
rect 21824 14365 21838 14399
rect 21838 14365 21872 14399
rect 21872 14365 21876 14399
rect 25412 14399 25464 14408
rect 21824 14356 21876 14365
rect 25412 14365 25421 14399
rect 25421 14365 25455 14399
rect 25455 14365 25464 14399
rect 25412 14356 25464 14365
rect 14924 14263 14976 14272
rect 14924 14229 14933 14263
rect 14933 14229 14967 14263
rect 14967 14229 14976 14263
rect 14924 14220 14976 14229
rect 17592 14263 17644 14272
rect 17592 14229 17601 14263
rect 17601 14229 17635 14263
rect 17635 14229 17644 14263
rect 17592 14220 17644 14229
rect 17684 14263 17736 14272
rect 17684 14229 17693 14263
rect 17693 14229 17727 14263
rect 17727 14229 17736 14263
rect 18144 14263 18196 14272
rect 17684 14220 17736 14229
rect 18144 14229 18153 14263
rect 18153 14229 18187 14263
rect 18187 14229 18196 14263
rect 18144 14220 18196 14229
rect 18328 14220 18380 14272
rect 19156 14220 19208 14272
rect 20904 14288 20956 14340
rect 21640 14331 21692 14340
rect 21640 14297 21649 14331
rect 21649 14297 21683 14331
rect 21683 14297 21692 14331
rect 21640 14288 21692 14297
rect 22284 14263 22336 14272
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 10395 14118 10447 14170
rect 10459 14118 10511 14170
rect 10523 14118 10575 14170
rect 10587 14118 10639 14170
rect 10651 14118 10703 14170
rect 19840 14118 19892 14170
rect 19904 14118 19956 14170
rect 19968 14118 20020 14170
rect 20032 14118 20084 14170
rect 20096 14118 20148 14170
rect 2504 14016 2556 14068
rect 5080 14016 5132 14068
rect 5632 14016 5684 14068
rect 7196 14016 7248 14068
rect 2596 13880 2648 13932
rect 3148 13948 3200 14000
rect 2872 13923 2924 13932
rect 2872 13889 2881 13923
rect 2881 13889 2915 13923
rect 2915 13889 2924 13923
rect 2872 13880 2924 13889
rect 3976 13948 4028 14000
rect 7656 14016 7708 14068
rect 8300 14016 8352 14068
rect 9312 14059 9364 14068
rect 9312 14025 9321 14059
rect 9321 14025 9355 14059
rect 9355 14025 9364 14059
rect 9312 14016 9364 14025
rect 5540 13923 5592 13932
rect 5540 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 6276 13880 6328 13932
rect 8208 13991 8260 14000
rect 8208 13957 8242 13991
rect 8242 13957 8260 13991
rect 8208 13948 8260 13957
rect 10140 14059 10192 14068
rect 10140 14025 10149 14059
rect 10149 14025 10183 14059
rect 10183 14025 10192 14059
rect 10784 14059 10836 14068
rect 10140 14016 10192 14025
rect 10784 14025 10793 14059
rect 10793 14025 10827 14059
rect 10827 14025 10836 14059
rect 10784 14016 10836 14025
rect 11796 14016 11848 14068
rect 12072 14016 12124 14068
rect 12992 14016 13044 14068
rect 13820 14016 13872 14068
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 7104 13923 7156 13932
rect 7104 13889 7114 13923
rect 7114 13889 7148 13923
rect 7148 13889 7156 13923
rect 7104 13880 7156 13889
rect 7472 13880 7524 13932
rect 1400 13812 1452 13864
rect 5264 13855 5316 13864
rect 5264 13821 5273 13855
rect 5273 13821 5307 13855
rect 5307 13821 5316 13855
rect 5264 13812 5316 13821
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 10140 13880 10192 13932
rect 11888 13880 11940 13932
rect 12716 13948 12768 14000
rect 13176 13948 13228 14000
rect 15476 14016 15528 14068
rect 18696 14059 18748 14068
rect 18696 14025 18705 14059
rect 18705 14025 18739 14059
rect 18739 14025 18748 14059
rect 18696 14016 18748 14025
rect 19616 14016 19668 14068
rect 22008 14016 22060 14068
rect 23020 14016 23072 14068
rect 12072 13923 12124 13932
rect 12072 13889 12081 13923
rect 12081 13889 12115 13923
rect 12115 13889 12124 13923
rect 12072 13880 12124 13889
rect 12808 13880 12860 13932
rect 13820 13880 13872 13932
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 20904 13991 20956 14000
rect 20904 13957 20922 13991
rect 20922 13957 20956 13991
rect 20904 13948 20956 13957
rect 15568 13880 15620 13932
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 17224 13880 17276 13932
rect 6736 13744 6788 13796
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 10416 13719 10468 13728
rect 10416 13685 10425 13719
rect 10425 13685 10459 13719
rect 10459 13685 10468 13719
rect 10416 13676 10468 13685
rect 11980 13744 12032 13796
rect 14924 13812 14976 13864
rect 16212 13812 16264 13864
rect 13820 13787 13872 13796
rect 13820 13753 13829 13787
rect 13829 13753 13863 13787
rect 13863 13753 13872 13787
rect 13820 13744 13872 13753
rect 14280 13744 14332 13796
rect 16672 13719 16724 13728
rect 16672 13685 16681 13719
rect 16681 13685 16715 13719
rect 16715 13685 16724 13719
rect 16672 13676 16724 13685
rect 21640 13880 21692 13932
rect 21180 13855 21232 13864
rect 18604 13744 18656 13796
rect 18788 13744 18840 13796
rect 21180 13821 21189 13855
rect 21189 13821 21223 13855
rect 21223 13821 21232 13855
rect 22100 13923 22152 13932
rect 22100 13889 22134 13923
rect 22134 13889 22152 13923
rect 22100 13880 22152 13889
rect 23664 13923 23716 13932
rect 23664 13889 23698 13923
rect 23698 13889 23716 13923
rect 23664 13880 23716 13889
rect 25044 13880 25096 13932
rect 21180 13812 21232 13821
rect 23388 13855 23440 13864
rect 23388 13821 23397 13855
rect 23397 13821 23431 13855
rect 23431 13821 23440 13855
rect 23388 13812 23440 13821
rect 18512 13719 18564 13728
rect 18512 13685 18521 13719
rect 18521 13685 18555 13719
rect 18555 13685 18564 13719
rect 18512 13676 18564 13685
rect 22744 13676 22796 13728
rect 23296 13676 23348 13728
rect 24124 13676 24176 13728
rect 25136 13676 25188 13728
rect 5672 13574 5724 13626
rect 5736 13574 5788 13626
rect 5800 13574 5852 13626
rect 5864 13574 5916 13626
rect 5928 13574 5980 13626
rect 15118 13574 15170 13626
rect 15182 13574 15234 13626
rect 15246 13574 15298 13626
rect 15310 13574 15362 13626
rect 15374 13574 15426 13626
rect 24563 13574 24615 13626
rect 24627 13574 24679 13626
rect 24691 13574 24743 13626
rect 24755 13574 24807 13626
rect 24819 13574 24871 13626
rect 2780 13472 2832 13524
rect 5356 13472 5408 13524
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 14372 13472 14424 13524
rect 2320 13336 2372 13388
rect 4620 13336 4672 13388
rect 6736 13336 6788 13388
rect 5448 13268 5500 13320
rect 6092 13268 6144 13320
rect 7196 13311 7248 13320
rect 7196 13277 7230 13311
rect 7230 13277 7248 13311
rect 7196 13268 7248 13277
rect 2596 13175 2648 13184
rect 2596 13141 2605 13175
rect 2605 13141 2639 13175
rect 2639 13141 2648 13175
rect 2596 13132 2648 13141
rect 6644 13132 6696 13184
rect 11980 13404 12032 13456
rect 12532 13404 12584 13456
rect 12992 13404 13044 13456
rect 15568 13447 15620 13456
rect 15568 13413 15577 13447
rect 15577 13413 15611 13447
rect 15611 13413 15620 13447
rect 15568 13404 15620 13413
rect 10968 13336 11020 13388
rect 11796 13336 11848 13388
rect 12072 13268 12124 13320
rect 13544 13336 13596 13388
rect 16672 13336 16724 13388
rect 12808 13268 12860 13320
rect 14832 13311 14884 13320
rect 14832 13277 14841 13311
rect 14841 13277 14875 13311
rect 14875 13277 14884 13311
rect 14832 13268 14884 13277
rect 10416 13200 10468 13252
rect 11888 13200 11940 13252
rect 12256 13200 12308 13252
rect 12532 13132 12584 13184
rect 15476 13268 15528 13320
rect 16580 13268 16632 13320
rect 19708 13472 19760 13524
rect 21180 13472 21232 13524
rect 22100 13472 22152 13524
rect 22560 13472 22612 13524
rect 23664 13472 23716 13524
rect 17224 13404 17276 13456
rect 18512 13404 18564 13456
rect 17684 13379 17736 13388
rect 17684 13345 17693 13379
rect 17693 13345 17727 13379
rect 17727 13345 17736 13379
rect 17684 13336 17736 13345
rect 17592 13268 17644 13320
rect 18052 13311 18104 13320
rect 18052 13277 18061 13311
rect 18061 13277 18095 13311
rect 18095 13277 18104 13311
rect 18052 13268 18104 13277
rect 21640 13336 21692 13388
rect 21824 13404 21876 13456
rect 22744 13404 22796 13456
rect 24492 13472 24544 13524
rect 25044 13472 25096 13524
rect 24032 13404 24084 13456
rect 22376 13336 22428 13388
rect 21824 13311 21876 13320
rect 21824 13277 21833 13311
rect 21833 13277 21867 13311
rect 21867 13277 21876 13311
rect 21824 13268 21876 13277
rect 22008 13311 22060 13320
rect 22008 13277 22017 13311
rect 22017 13277 22051 13311
rect 22051 13277 22060 13311
rect 22008 13268 22060 13277
rect 22192 13311 22244 13320
rect 22192 13277 22206 13311
rect 22206 13277 22240 13311
rect 22240 13277 22244 13311
rect 22192 13268 22244 13277
rect 20260 13200 20312 13252
rect 20996 13200 21048 13252
rect 14556 13132 14608 13184
rect 14648 13175 14700 13184
rect 14648 13141 14657 13175
rect 14657 13141 14691 13175
rect 14691 13141 14700 13175
rect 14648 13132 14700 13141
rect 15476 13132 15528 13184
rect 17132 13132 17184 13184
rect 17960 13132 18012 13184
rect 19248 13132 19300 13184
rect 19340 13132 19392 13184
rect 23940 13268 23992 13320
rect 24492 13268 24544 13320
rect 24584 13243 24636 13252
rect 22744 13175 22796 13184
rect 22744 13141 22753 13175
rect 22753 13141 22787 13175
rect 22787 13141 22796 13175
rect 22744 13132 22796 13141
rect 23296 13132 23348 13184
rect 24032 13132 24084 13184
rect 24584 13209 24593 13243
rect 24593 13209 24627 13243
rect 24627 13209 24636 13243
rect 24584 13200 24636 13209
rect 24676 13243 24728 13252
rect 24676 13209 24685 13243
rect 24685 13209 24719 13243
rect 24719 13209 24728 13243
rect 25136 13243 25188 13252
rect 24676 13200 24728 13209
rect 25136 13209 25145 13243
rect 25145 13209 25179 13243
rect 25179 13209 25188 13243
rect 25136 13200 25188 13209
rect 24492 13132 24544 13184
rect 10395 13030 10447 13082
rect 10459 13030 10511 13082
rect 10523 13030 10575 13082
rect 10587 13030 10639 13082
rect 10651 13030 10703 13082
rect 19840 13030 19892 13082
rect 19904 13030 19956 13082
rect 19968 13030 20020 13082
rect 20032 13030 20084 13082
rect 20096 13030 20148 13082
rect 3608 12928 3660 12980
rect 4068 12928 4120 12980
rect 8668 12971 8720 12980
rect 8668 12937 8677 12971
rect 8677 12937 8711 12971
rect 8711 12937 8720 12971
rect 8668 12928 8720 12937
rect 3056 12860 3108 12912
rect 3884 12860 3936 12912
rect 5540 12860 5592 12912
rect 6736 12903 6788 12912
rect 6736 12869 6745 12903
rect 6745 12869 6779 12903
rect 6779 12869 6788 12903
rect 6736 12860 6788 12869
rect 8852 12860 8904 12912
rect 9496 12860 9548 12912
rect 10048 12860 10100 12912
rect 12348 12928 12400 12980
rect 12532 12971 12584 12980
rect 12532 12937 12541 12971
rect 12541 12937 12575 12971
rect 12575 12937 12584 12971
rect 12532 12928 12584 12937
rect 13268 12928 13320 12980
rect 13544 12928 13596 12980
rect 17500 12928 17552 12980
rect 18328 12928 18380 12980
rect 19708 12928 19760 12980
rect 20260 12971 20312 12980
rect 20260 12937 20269 12971
rect 20269 12937 20303 12971
rect 20303 12937 20312 12971
rect 20260 12928 20312 12937
rect 20996 12928 21048 12980
rect 22284 12971 22336 12980
rect 22284 12937 22293 12971
rect 22293 12937 22327 12971
rect 22327 12937 22336 12971
rect 22284 12928 22336 12937
rect 23572 12928 23624 12980
rect 23940 12928 23992 12980
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 6644 12835 6696 12844
rect 6644 12801 6653 12835
rect 6653 12801 6687 12835
rect 6687 12801 6696 12835
rect 6644 12792 6696 12801
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 4160 12724 4212 12776
rect 4436 12724 4488 12776
rect 8760 12792 8812 12844
rect 10968 12860 11020 12912
rect 11796 12835 11848 12844
rect 11796 12801 11800 12835
rect 11800 12801 11834 12835
rect 11834 12801 11848 12835
rect 11796 12792 11848 12801
rect 8392 12724 8444 12776
rect 2780 12656 2832 12708
rect 7932 12699 7984 12708
rect 7932 12665 7941 12699
rect 7941 12665 7975 12699
rect 7975 12665 7984 12699
rect 7932 12656 7984 12665
rect 2964 12588 3016 12640
rect 4436 12631 4488 12640
rect 4436 12597 4445 12631
rect 4445 12597 4479 12631
rect 4479 12597 4488 12631
rect 4436 12588 4488 12597
rect 6368 12588 6420 12640
rect 8668 12588 8720 12640
rect 12072 12792 12124 12844
rect 12256 12835 12308 12844
rect 12256 12801 12265 12835
rect 12265 12801 12299 12835
rect 12299 12801 12308 12835
rect 12900 12860 12952 12912
rect 14556 12860 14608 12912
rect 19340 12860 19392 12912
rect 19524 12860 19576 12912
rect 22100 12903 22152 12912
rect 22100 12869 22109 12903
rect 22109 12869 22143 12903
rect 22143 12869 22152 12903
rect 22100 12860 22152 12869
rect 23296 12860 23348 12912
rect 24124 12903 24176 12912
rect 24124 12869 24133 12903
rect 24133 12869 24167 12903
rect 24167 12869 24176 12903
rect 24124 12860 24176 12869
rect 12256 12792 12308 12801
rect 14004 12792 14056 12844
rect 14280 12792 14332 12844
rect 17040 12792 17092 12844
rect 21088 12792 21140 12844
rect 22468 12792 22520 12844
rect 23940 12835 23992 12844
rect 23940 12801 23949 12835
rect 23949 12801 23983 12835
rect 23983 12801 23992 12835
rect 23940 12792 23992 12801
rect 24492 12792 24544 12844
rect 25412 12792 25464 12844
rect 25688 12792 25740 12844
rect 12348 12724 12400 12776
rect 12992 12724 13044 12776
rect 18420 12724 18472 12776
rect 20076 12724 20128 12776
rect 23664 12656 23716 12708
rect 24676 12699 24728 12708
rect 24676 12665 24685 12699
rect 24685 12665 24719 12699
rect 24719 12665 24728 12699
rect 24676 12656 24728 12665
rect 14556 12631 14608 12640
rect 14556 12597 14565 12631
rect 14565 12597 14599 12631
rect 14599 12597 14608 12631
rect 14556 12588 14608 12597
rect 20444 12588 20496 12640
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 24492 12631 24544 12640
rect 24492 12597 24501 12631
rect 24501 12597 24535 12631
rect 24535 12597 24544 12631
rect 24492 12588 24544 12597
rect 5672 12486 5724 12538
rect 5736 12486 5788 12538
rect 5800 12486 5852 12538
rect 5864 12486 5916 12538
rect 5928 12486 5980 12538
rect 15118 12486 15170 12538
rect 15182 12486 15234 12538
rect 15246 12486 15298 12538
rect 15310 12486 15362 12538
rect 15374 12486 15426 12538
rect 24563 12486 24615 12538
rect 24627 12486 24679 12538
rect 24691 12486 24743 12538
rect 24755 12486 24807 12538
rect 24819 12486 24871 12538
rect 2596 12384 2648 12436
rect 5264 12427 5316 12436
rect 5264 12393 5273 12427
rect 5273 12393 5307 12427
rect 5307 12393 5316 12427
rect 5264 12384 5316 12393
rect 6184 12384 6236 12436
rect 7656 12384 7708 12436
rect 8760 12384 8812 12436
rect 9496 12427 9548 12436
rect 9496 12393 9505 12427
rect 9505 12393 9539 12427
rect 9539 12393 9548 12427
rect 9496 12384 9548 12393
rect 12808 12427 12860 12436
rect 3424 12359 3476 12368
rect 3424 12325 3433 12359
rect 3433 12325 3467 12359
rect 3467 12325 3476 12359
rect 3424 12316 3476 12325
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 3056 12291 3108 12300
rect 3056 12257 3065 12291
rect 3065 12257 3099 12291
rect 3099 12257 3108 12291
rect 3056 12248 3108 12257
rect 5540 12248 5592 12300
rect 9680 12316 9732 12368
rect 10140 12316 10192 12368
rect 5264 12180 5316 12232
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 6736 12180 6788 12232
rect 7932 12180 7984 12232
rect 1952 12112 2004 12164
rect 4436 12112 4488 12164
rect 11152 12248 11204 12300
rect 11336 12248 11388 12300
rect 9496 12180 9548 12232
rect 3792 12044 3844 12096
rect 3976 12044 4028 12096
rect 4988 12044 5040 12096
rect 6184 12044 6236 12096
rect 6460 12044 6512 12096
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11428 12223 11480 12232
rect 9680 12044 9732 12096
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 12072 12248 12124 12300
rect 12808 12393 12817 12427
rect 12817 12393 12851 12427
rect 12851 12393 12860 12427
rect 12808 12384 12860 12393
rect 14004 12384 14056 12436
rect 17684 12384 17736 12436
rect 15660 12316 15712 12368
rect 17592 12316 17644 12368
rect 18052 12316 18104 12368
rect 12440 12180 12492 12232
rect 14556 12180 14608 12232
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 15476 12248 15528 12300
rect 19524 12384 19576 12436
rect 21548 12384 21600 12436
rect 22100 12384 22152 12436
rect 18328 12316 18380 12368
rect 15200 12223 15252 12232
rect 15200 12189 15209 12223
rect 15209 12189 15243 12223
rect 15243 12189 15252 12223
rect 15200 12180 15252 12189
rect 15660 12223 15712 12232
rect 12992 12155 13044 12164
rect 11612 12087 11664 12096
rect 11612 12053 11621 12087
rect 11621 12053 11655 12087
rect 11655 12053 11664 12087
rect 11612 12044 11664 12053
rect 12992 12121 13001 12155
rect 13001 12121 13035 12155
rect 13035 12121 13044 12155
rect 12992 12112 13044 12121
rect 12624 12044 12676 12096
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 17776 12223 17828 12232
rect 17776 12189 17785 12223
rect 17785 12189 17819 12223
rect 17819 12189 17828 12223
rect 17776 12180 17828 12189
rect 17868 12180 17920 12232
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 19248 12248 19300 12300
rect 19340 12248 19392 12300
rect 20076 12248 20128 12300
rect 22744 12180 22796 12232
rect 23388 12248 23440 12300
rect 22928 12180 22980 12232
rect 23572 12223 23624 12232
rect 23572 12189 23581 12223
rect 23581 12189 23615 12223
rect 23615 12189 23624 12223
rect 23572 12180 23624 12189
rect 23848 12223 23900 12232
rect 23848 12189 23857 12223
rect 23857 12189 23891 12223
rect 23891 12189 23900 12223
rect 23848 12180 23900 12189
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 17500 12044 17552 12096
rect 17868 12044 17920 12096
rect 18604 12112 18656 12164
rect 20444 12112 20496 12164
rect 22376 12112 22428 12164
rect 23664 12112 23716 12164
rect 24400 12180 24452 12232
rect 18144 12044 18196 12096
rect 18236 12044 18288 12096
rect 20996 12044 21048 12096
rect 21180 12087 21232 12096
rect 21180 12053 21189 12087
rect 21189 12053 21223 12087
rect 21223 12053 21232 12087
rect 21180 12044 21232 12053
rect 22192 12044 22244 12096
rect 24032 12044 24084 12096
rect 10395 11942 10447 11994
rect 10459 11942 10511 11994
rect 10523 11942 10575 11994
rect 10587 11942 10639 11994
rect 10651 11942 10703 11994
rect 19840 11942 19892 11994
rect 19904 11942 19956 11994
rect 19968 11942 20020 11994
rect 20032 11942 20084 11994
rect 20096 11942 20148 11994
rect 1952 11883 2004 11892
rect 1952 11849 1961 11883
rect 1961 11849 1995 11883
rect 1995 11849 2004 11883
rect 1952 11840 2004 11849
rect 4068 11840 4120 11892
rect 4988 11815 5040 11824
rect 2780 11704 2832 11756
rect 2964 11747 3016 11756
rect 2964 11713 2973 11747
rect 2973 11713 3007 11747
rect 3007 11713 3016 11747
rect 2964 11704 3016 11713
rect 3792 11747 3844 11756
rect 3792 11713 3801 11747
rect 3801 11713 3835 11747
rect 3835 11713 3844 11747
rect 3792 11704 3844 11713
rect 4988 11781 4997 11815
rect 4997 11781 5031 11815
rect 5031 11781 5040 11815
rect 4988 11772 5040 11781
rect 4620 11747 4672 11756
rect 4620 11713 4629 11747
rect 4629 11713 4663 11747
rect 4663 11713 4672 11747
rect 6000 11840 6052 11892
rect 8760 11840 8812 11892
rect 4620 11704 4672 11713
rect 4160 11636 4212 11688
rect 5540 11636 5592 11688
rect 6736 11772 6788 11824
rect 8852 11815 8904 11824
rect 8852 11781 8861 11815
rect 8861 11781 8895 11815
rect 8895 11781 8904 11815
rect 8852 11772 8904 11781
rect 9220 11840 9272 11892
rect 15016 11840 15068 11892
rect 15200 11840 15252 11892
rect 6460 11704 6512 11756
rect 7748 11704 7800 11756
rect 10140 11704 10192 11756
rect 3424 11568 3476 11620
rect 3884 11500 3936 11552
rect 5172 11500 5224 11552
rect 7748 11543 7800 11552
rect 7748 11509 7757 11543
rect 7757 11509 7791 11543
rect 7791 11509 7800 11543
rect 7748 11500 7800 11509
rect 10416 11500 10468 11552
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 10784 11543 10836 11552
rect 10784 11509 10793 11543
rect 10793 11509 10827 11543
rect 10827 11509 10836 11543
rect 10784 11500 10836 11509
rect 11612 11772 11664 11824
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 11980 11704 12032 11756
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12808 11772 12860 11824
rect 13912 11772 13964 11824
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 14832 11704 14884 11756
rect 15476 11772 15528 11824
rect 11244 11500 11296 11552
rect 11612 11500 11664 11552
rect 13820 11636 13872 11688
rect 17316 11840 17368 11892
rect 17776 11840 17828 11892
rect 18236 11840 18288 11892
rect 19432 11883 19484 11892
rect 19432 11849 19441 11883
rect 19441 11849 19475 11883
rect 19475 11849 19484 11883
rect 19432 11840 19484 11849
rect 21548 11883 21600 11892
rect 21548 11849 21557 11883
rect 21557 11849 21591 11883
rect 21591 11849 21600 11883
rect 21548 11840 21600 11849
rect 24492 11840 24544 11892
rect 16396 11772 16448 11824
rect 17132 11704 17184 11756
rect 21824 11747 21876 11756
rect 15568 11636 15620 11688
rect 16672 11636 16724 11688
rect 17868 11679 17920 11688
rect 17868 11645 17877 11679
rect 17877 11645 17911 11679
rect 17911 11645 17920 11679
rect 17868 11636 17920 11645
rect 18420 11636 18472 11688
rect 19892 11679 19944 11688
rect 12992 11500 13044 11552
rect 13176 11500 13228 11552
rect 14556 11500 14608 11552
rect 15936 11500 15988 11552
rect 16120 11568 16172 11620
rect 17776 11568 17828 11620
rect 19892 11645 19901 11679
rect 19901 11645 19935 11679
rect 19935 11645 19944 11679
rect 19892 11636 19944 11645
rect 18328 11543 18380 11552
rect 18328 11509 18337 11543
rect 18337 11509 18371 11543
rect 18371 11509 18380 11543
rect 18328 11500 18380 11509
rect 21824 11713 21833 11747
rect 21833 11713 21867 11747
rect 21867 11713 21876 11747
rect 21824 11704 21876 11713
rect 22192 11747 22244 11756
rect 22192 11713 22206 11747
rect 22206 11713 22240 11747
rect 22240 11713 22244 11747
rect 22192 11704 22244 11713
rect 22652 11704 22704 11756
rect 23204 11704 23256 11756
rect 23388 11704 23440 11756
rect 22376 11611 22428 11620
rect 22376 11577 22385 11611
rect 22385 11577 22419 11611
rect 22419 11577 22428 11611
rect 22376 11568 22428 11577
rect 21364 11543 21416 11552
rect 21364 11509 21373 11543
rect 21373 11509 21407 11543
rect 21407 11509 21416 11543
rect 21364 11500 21416 11509
rect 23940 11543 23992 11552
rect 23940 11509 23949 11543
rect 23949 11509 23983 11543
rect 23983 11509 23992 11543
rect 23940 11500 23992 11509
rect 25412 11500 25464 11552
rect 25872 11543 25924 11552
rect 25872 11509 25881 11543
rect 25881 11509 25915 11543
rect 25915 11509 25924 11543
rect 25872 11500 25924 11509
rect 5672 11398 5724 11450
rect 5736 11398 5788 11450
rect 5800 11398 5852 11450
rect 5864 11398 5916 11450
rect 5928 11398 5980 11450
rect 15118 11398 15170 11450
rect 15182 11398 15234 11450
rect 15246 11398 15298 11450
rect 15310 11398 15362 11450
rect 15374 11398 15426 11450
rect 24563 11398 24615 11450
rect 24627 11398 24679 11450
rect 24691 11398 24743 11450
rect 24755 11398 24807 11450
rect 24819 11398 24871 11450
rect 2688 11296 2740 11348
rect 4804 11296 4856 11348
rect 6368 11296 6420 11348
rect 7288 11296 7340 11348
rect 10784 11296 10836 11348
rect 11980 11296 12032 11348
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 6644 11228 6696 11280
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 6000 11160 6052 11212
rect 6368 11092 6420 11144
rect 7748 11160 7800 11212
rect 9680 11228 9732 11280
rect 11244 11228 11296 11280
rect 10048 11160 10100 11212
rect 10416 11160 10468 11212
rect 1400 11024 1452 11076
rect 2412 11067 2464 11076
rect 2412 11033 2421 11067
rect 2421 11033 2455 11067
rect 2455 11033 2464 11067
rect 2412 11024 2464 11033
rect 9588 11092 9640 11144
rect 10140 11024 10192 11076
rect 10600 11024 10652 11076
rect 11612 11160 11664 11212
rect 12348 11228 12400 11280
rect 16120 11296 16172 11348
rect 17132 11339 17184 11348
rect 17132 11305 17141 11339
rect 17141 11305 17175 11339
rect 17175 11305 17184 11339
rect 17132 11296 17184 11305
rect 13912 11160 13964 11212
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 15476 11228 15528 11280
rect 15568 11160 15620 11212
rect 15660 11160 15712 11212
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 14832 11092 14884 11144
rect 17684 11228 17736 11280
rect 17592 11203 17644 11212
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 19892 11296 19944 11348
rect 21180 11296 21232 11348
rect 26240 11296 26292 11348
rect 17592 11160 17644 11169
rect 19248 11203 19300 11212
rect 19248 11169 19257 11203
rect 19257 11169 19291 11203
rect 19291 11169 19300 11203
rect 19248 11160 19300 11169
rect 4252 10956 4304 11008
rect 5724 10999 5776 11008
rect 5724 10965 5733 10999
rect 5733 10965 5767 10999
rect 5767 10965 5776 10999
rect 5724 10956 5776 10965
rect 9128 10956 9180 11008
rect 12992 10999 13044 11008
rect 12992 10965 13001 10999
rect 13001 10965 13035 10999
rect 13035 10965 13044 10999
rect 12992 10956 13044 10965
rect 14556 10956 14608 11008
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 15936 11024 15988 11076
rect 17408 11092 17460 11144
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 18144 11135 18196 11144
rect 18144 11101 18153 11135
rect 18153 11101 18187 11135
rect 18187 11101 18196 11135
rect 18144 11092 18196 11101
rect 18328 11135 18380 11144
rect 18328 11101 18336 11135
rect 18336 11101 18370 11135
rect 18370 11101 18380 11135
rect 18328 11092 18380 11101
rect 19892 11092 19944 11144
rect 16396 10956 16448 11008
rect 17960 10999 18012 11008
rect 17960 10965 17969 10999
rect 17969 10965 18003 10999
rect 18003 10965 18012 10999
rect 17960 10956 18012 10965
rect 10395 10854 10447 10906
rect 10459 10854 10511 10906
rect 10523 10854 10575 10906
rect 10587 10854 10639 10906
rect 10651 10854 10703 10906
rect 19840 10854 19892 10906
rect 19904 10854 19956 10906
rect 19968 10854 20020 10906
rect 20032 10854 20084 10906
rect 20096 10854 20148 10906
rect 2412 10752 2464 10804
rect 3240 10752 3292 10804
rect 3976 10752 4028 10804
rect 5724 10752 5776 10804
rect 12348 10752 12400 10804
rect 16396 10795 16448 10804
rect 16396 10761 16405 10795
rect 16405 10761 16439 10795
rect 16439 10761 16448 10795
rect 16396 10752 16448 10761
rect 17868 10752 17920 10804
rect 22468 10752 22520 10804
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 2320 10616 2372 10668
rect 3976 10659 4028 10668
rect 3976 10625 3994 10659
rect 3994 10625 4028 10659
rect 3976 10616 4028 10625
rect 4620 10659 4672 10668
rect 4620 10625 4629 10659
rect 4629 10625 4663 10659
rect 4663 10625 4672 10659
rect 4620 10616 4672 10625
rect 9128 10684 9180 10736
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 6736 10616 6788 10668
rect 9680 10659 9732 10668
rect 9680 10625 9729 10659
rect 9729 10625 9732 10659
rect 9680 10616 9732 10625
rect 2596 10548 2648 10600
rect 4528 10591 4580 10600
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 4528 10557 4537 10591
rect 4537 10557 4571 10591
rect 4571 10557 4580 10591
rect 4528 10548 4580 10557
rect 1676 10412 1728 10421
rect 5540 10412 5592 10464
rect 6000 10455 6052 10464
rect 6000 10421 6009 10455
rect 6009 10421 6043 10455
rect 6043 10421 6052 10455
rect 6000 10412 6052 10421
rect 6920 10412 6972 10464
rect 9404 10412 9456 10464
rect 11060 10616 11112 10668
rect 12440 10616 12492 10668
rect 14280 10616 14332 10668
rect 15568 10616 15620 10668
rect 17960 10684 18012 10736
rect 19340 10616 19392 10668
rect 22100 10659 22152 10668
rect 22100 10625 22109 10659
rect 22109 10625 22143 10659
rect 22143 10625 22152 10659
rect 22100 10616 22152 10625
rect 22284 10616 22336 10668
rect 10324 10412 10376 10464
rect 17132 10548 17184 10600
rect 22652 10616 22704 10668
rect 22928 10659 22980 10668
rect 22928 10625 22937 10659
rect 22937 10625 22971 10659
rect 22971 10625 22980 10659
rect 22928 10616 22980 10625
rect 23112 10659 23164 10668
rect 23112 10625 23121 10659
rect 23121 10625 23155 10659
rect 23155 10625 23164 10659
rect 23112 10616 23164 10625
rect 22468 10591 22520 10600
rect 22468 10557 22477 10591
rect 22477 10557 22511 10591
rect 22511 10557 22520 10591
rect 23204 10591 23256 10600
rect 22468 10548 22520 10557
rect 23204 10557 23213 10591
rect 23213 10557 23247 10591
rect 23247 10557 23256 10591
rect 23204 10548 23256 10557
rect 23480 10548 23532 10600
rect 23020 10480 23072 10532
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 24952 10659 25004 10668
rect 23940 10616 23992 10625
rect 24952 10625 24961 10659
rect 24961 10625 24995 10659
rect 24995 10625 25004 10659
rect 24952 10616 25004 10625
rect 25504 10616 25556 10668
rect 24492 10548 24544 10600
rect 12164 10412 12216 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12716 10455 12768 10464
rect 12440 10412 12492 10421
rect 12716 10421 12725 10455
rect 12725 10421 12759 10455
rect 12759 10421 12768 10455
rect 12716 10412 12768 10421
rect 13636 10412 13688 10464
rect 16580 10412 16632 10464
rect 17408 10412 17460 10464
rect 22192 10412 22244 10464
rect 23296 10412 23348 10464
rect 23756 10412 23808 10464
rect 25044 10412 25096 10464
rect 5672 10310 5724 10362
rect 5736 10310 5788 10362
rect 5800 10310 5852 10362
rect 5864 10310 5916 10362
rect 5928 10310 5980 10362
rect 15118 10310 15170 10362
rect 15182 10310 15234 10362
rect 15246 10310 15298 10362
rect 15310 10310 15362 10362
rect 15374 10310 15426 10362
rect 24563 10310 24615 10362
rect 24627 10310 24679 10362
rect 24691 10310 24743 10362
rect 24755 10310 24807 10362
rect 24819 10310 24871 10362
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 3976 10208 4028 10260
rect 4068 10208 4120 10260
rect 13820 10208 13872 10260
rect 14096 10208 14148 10260
rect 4528 10140 4580 10192
rect 2596 10072 2648 10124
rect 2872 10072 2924 10124
rect 4252 10115 4304 10124
rect 2780 10004 2832 10056
rect 4252 10081 4261 10115
rect 4261 10081 4295 10115
rect 4295 10081 4304 10115
rect 4252 10072 4304 10081
rect 2964 9936 3016 9988
rect 3332 9868 3384 9920
rect 4160 9911 4212 9920
rect 4160 9877 4169 9911
rect 4169 9877 4203 9911
rect 4203 9877 4212 9911
rect 4160 9868 4212 9877
rect 5540 10072 5592 10124
rect 12256 10072 12308 10124
rect 14464 10115 14516 10124
rect 14464 10081 14473 10115
rect 14473 10081 14507 10115
rect 14507 10081 14516 10115
rect 14464 10072 14516 10081
rect 14648 10115 14700 10124
rect 14648 10081 14657 10115
rect 14657 10081 14691 10115
rect 14691 10081 14700 10115
rect 14648 10072 14700 10081
rect 16304 10208 16356 10260
rect 19708 10208 19760 10260
rect 22100 10208 22152 10260
rect 22376 10208 22428 10260
rect 23112 10208 23164 10260
rect 24952 10208 25004 10260
rect 15476 10072 15528 10124
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 15844 10004 15896 10056
rect 6000 9936 6052 9988
rect 11060 9936 11112 9988
rect 4988 9868 5040 9920
rect 7196 9911 7248 9920
rect 7196 9877 7205 9911
rect 7205 9877 7239 9911
rect 7239 9877 7248 9911
rect 7196 9868 7248 9877
rect 8944 9911 8996 9920
rect 8944 9877 8953 9911
rect 8953 9877 8987 9911
rect 8987 9877 8996 9911
rect 8944 9868 8996 9877
rect 11980 9868 12032 9920
rect 13176 9936 13228 9988
rect 13360 9936 13412 9988
rect 15200 9936 15252 9988
rect 22192 10140 22244 10192
rect 23204 10140 23256 10192
rect 22652 10072 22704 10124
rect 22100 10004 22152 10056
rect 22468 10004 22520 10056
rect 23204 10047 23256 10056
rect 22928 9868 22980 9920
rect 23204 10013 23213 10047
rect 23213 10013 23247 10047
rect 23247 10013 23256 10047
rect 23204 10004 23256 10013
rect 23388 10047 23440 10056
rect 23388 10013 23397 10047
rect 23397 10013 23431 10047
rect 23431 10013 23440 10047
rect 23388 10004 23440 10013
rect 23848 10140 23900 10192
rect 24952 10072 25004 10124
rect 23940 10004 23992 10056
rect 23112 9979 23164 9988
rect 23112 9945 23121 9979
rect 23121 9945 23155 9979
rect 23155 9945 23164 9979
rect 23112 9936 23164 9945
rect 23756 9936 23808 9988
rect 23572 9868 23624 9920
rect 24768 9911 24820 9920
rect 24768 9877 24777 9911
rect 24777 9877 24811 9911
rect 24811 9877 24820 9911
rect 24768 9868 24820 9877
rect 25136 9936 25188 9988
rect 25504 9868 25556 9920
rect 25596 9868 25648 9920
rect 10395 9766 10447 9818
rect 10459 9766 10511 9818
rect 10523 9766 10575 9818
rect 10587 9766 10639 9818
rect 10651 9766 10703 9818
rect 19840 9766 19892 9818
rect 19904 9766 19956 9818
rect 19968 9766 20020 9818
rect 20032 9766 20084 9818
rect 20096 9766 20148 9818
rect 2780 9707 2832 9716
rect 2780 9673 2789 9707
rect 2789 9673 2823 9707
rect 2823 9673 2832 9707
rect 2780 9664 2832 9673
rect 4620 9664 4672 9716
rect 6368 9664 6420 9716
rect 1676 9639 1728 9648
rect 1676 9605 1710 9639
rect 1710 9605 1728 9639
rect 1676 9596 1728 9605
rect 2688 9596 2740 9648
rect 2872 9596 2924 9648
rect 2964 9596 3016 9648
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 2780 9460 2832 9512
rect 3148 9460 3200 9512
rect 3792 9503 3844 9512
rect 3792 9469 3801 9503
rect 3801 9469 3835 9503
rect 3835 9469 3844 9503
rect 3792 9460 3844 9469
rect 4160 9528 4212 9580
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 6092 9596 6144 9648
rect 4620 9460 4672 9512
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 5080 9460 5132 9512
rect 6092 9460 6144 9512
rect 8944 9596 8996 9648
rect 9680 9596 9732 9648
rect 9772 9596 9824 9648
rect 7196 9528 7248 9580
rect 7288 9528 7340 9580
rect 4344 9367 4396 9376
rect 4344 9333 4353 9367
rect 4353 9333 4387 9367
rect 4387 9333 4396 9367
rect 4344 9324 4396 9333
rect 6920 9324 6972 9376
rect 7104 9324 7156 9376
rect 7932 9367 7984 9376
rect 7932 9333 7941 9367
rect 7941 9333 7975 9367
rect 7975 9333 7984 9367
rect 7932 9324 7984 9333
rect 9772 9324 9824 9376
rect 10324 9528 10376 9580
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 10876 9392 10928 9444
rect 10968 9392 11020 9444
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11888 9596 11940 9648
rect 12716 9664 12768 9716
rect 13176 9664 13228 9716
rect 13728 9664 13780 9716
rect 14372 9664 14424 9716
rect 14924 9664 14976 9716
rect 19156 9707 19208 9716
rect 11520 9528 11572 9537
rect 11888 9460 11940 9512
rect 12348 9571 12400 9580
rect 12348 9537 12357 9571
rect 12357 9537 12391 9571
rect 12391 9537 12400 9571
rect 12348 9528 12400 9537
rect 12532 9528 12584 9580
rect 13636 9571 13688 9580
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 15200 9639 15252 9648
rect 15200 9605 15209 9639
rect 15209 9605 15243 9639
rect 15243 9605 15252 9639
rect 15200 9596 15252 9605
rect 19156 9673 19165 9707
rect 19165 9673 19199 9707
rect 19199 9673 19208 9707
rect 19156 9664 19208 9673
rect 18972 9596 19024 9648
rect 15108 9571 15160 9580
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15108 9528 15160 9537
rect 15844 9571 15896 9580
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 13912 9460 13964 9512
rect 15016 9460 15068 9512
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 18236 9528 18288 9580
rect 19708 9596 19760 9648
rect 23480 9664 23532 9716
rect 25504 9707 25556 9716
rect 25504 9673 25513 9707
rect 25513 9673 25547 9707
rect 25547 9673 25556 9707
rect 25504 9664 25556 9673
rect 21180 9596 21232 9648
rect 22284 9596 22336 9648
rect 23296 9596 23348 9648
rect 20628 9528 20680 9580
rect 17132 9460 17184 9512
rect 12532 9392 12584 9444
rect 13360 9392 13412 9444
rect 11060 9324 11112 9376
rect 11244 9367 11296 9376
rect 11244 9333 11253 9367
rect 11253 9333 11287 9367
rect 11287 9333 11296 9367
rect 11244 9324 11296 9333
rect 11796 9367 11848 9376
rect 11796 9333 11805 9367
rect 11805 9333 11839 9367
rect 11839 9333 11848 9367
rect 11796 9324 11848 9333
rect 14648 9367 14700 9376
rect 14648 9333 14657 9367
rect 14657 9333 14691 9367
rect 14691 9333 14700 9367
rect 14648 9324 14700 9333
rect 17316 9324 17368 9376
rect 19064 9392 19116 9444
rect 20996 9392 21048 9444
rect 23204 9528 23256 9580
rect 24768 9571 24820 9580
rect 22744 9460 22796 9512
rect 23020 9392 23072 9444
rect 24768 9537 24777 9571
rect 24777 9537 24811 9571
rect 24811 9537 24820 9571
rect 24768 9528 24820 9537
rect 25044 9571 25096 9580
rect 25044 9537 25053 9571
rect 25053 9537 25087 9571
rect 25087 9537 25096 9571
rect 25044 9528 25096 9537
rect 25596 9571 25648 9580
rect 25136 9460 25188 9512
rect 25596 9537 25605 9571
rect 25605 9537 25639 9571
rect 25639 9537 25648 9571
rect 25596 9528 25648 9537
rect 25504 9460 25556 9512
rect 24492 9392 24544 9444
rect 18880 9367 18932 9376
rect 18880 9333 18889 9367
rect 18889 9333 18923 9367
rect 18923 9333 18932 9367
rect 19708 9367 19760 9376
rect 18880 9324 18932 9333
rect 19708 9333 19717 9367
rect 19717 9333 19751 9367
rect 19751 9333 19760 9367
rect 19708 9324 19760 9333
rect 20352 9324 20404 9376
rect 22376 9324 22428 9376
rect 23388 9324 23440 9376
rect 5672 9222 5724 9274
rect 5736 9222 5788 9274
rect 5800 9222 5852 9274
rect 5864 9222 5916 9274
rect 5928 9222 5980 9274
rect 15118 9222 15170 9274
rect 15182 9222 15234 9274
rect 15246 9222 15298 9274
rect 15310 9222 15362 9274
rect 15374 9222 15426 9274
rect 24563 9222 24615 9274
rect 24627 9222 24679 9274
rect 24691 9222 24743 9274
rect 24755 9222 24807 9274
rect 24819 9222 24871 9274
rect 4160 9120 4212 9172
rect 4712 9120 4764 9172
rect 7288 9120 7340 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 11520 9120 11572 9172
rect 12992 9120 13044 9172
rect 12164 9052 12216 9104
rect 14004 9120 14056 9172
rect 15016 9163 15068 9172
rect 15016 9129 15025 9163
rect 15025 9129 15059 9163
rect 15059 9129 15068 9163
rect 15016 9120 15068 9129
rect 18236 9163 18288 9172
rect 18236 9129 18245 9163
rect 18245 9129 18279 9163
rect 18279 9129 18288 9163
rect 18236 9120 18288 9129
rect 22284 9163 22336 9172
rect 22284 9129 22293 9163
rect 22293 9129 22327 9163
rect 22327 9129 22336 9163
rect 22284 9120 22336 9129
rect 22928 9120 22980 9172
rect 25504 9120 25556 9172
rect 15384 9052 15436 9104
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 3240 8916 3292 8968
rect 5080 8959 5132 8968
rect 5080 8925 5089 8959
rect 5089 8925 5123 8959
rect 5123 8925 5132 8959
rect 5080 8916 5132 8925
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 8300 8916 8352 8968
rect 8760 8916 8812 8968
rect 10692 8984 10744 9036
rect 11244 8984 11296 9036
rect 17776 8984 17828 9036
rect 21548 9052 21600 9104
rect 22744 9095 22796 9104
rect 22744 9061 22753 9095
rect 22753 9061 22787 9095
rect 22787 9061 22796 9095
rect 22744 9052 22796 9061
rect 12256 8916 12308 8968
rect 13728 8959 13780 8968
rect 13728 8925 13737 8959
rect 13737 8925 13771 8959
rect 13771 8925 13780 8959
rect 13728 8916 13780 8925
rect 17132 8916 17184 8968
rect 19340 8959 19392 8968
rect 19340 8925 19349 8959
rect 19349 8925 19383 8959
rect 19383 8925 19392 8959
rect 19340 8916 19392 8925
rect 20996 9027 21048 9036
rect 20996 8993 21005 9027
rect 21005 8993 21039 9027
rect 21039 8993 21048 9027
rect 20996 8984 21048 8993
rect 20352 8959 20404 8968
rect 3608 8848 3660 8900
rect 4068 8848 4120 8900
rect 6828 8823 6880 8832
rect 6828 8789 6837 8823
rect 6837 8789 6871 8823
rect 6871 8789 6880 8823
rect 6828 8780 6880 8789
rect 7564 8848 7616 8900
rect 11796 8848 11848 8900
rect 12348 8848 12400 8900
rect 14004 8848 14056 8900
rect 10968 8780 11020 8832
rect 13820 8780 13872 8832
rect 15200 8780 15252 8832
rect 15844 8823 15896 8832
rect 15844 8789 15853 8823
rect 15853 8789 15887 8823
rect 15887 8789 15896 8823
rect 15844 8780 15896 8789
rect 16856 8780 16908 8832
rect 20352 8925 20361 8959
rect 20361 8925 20395 8959
rect 20395 8925 20404 8959
rect 20352 8916 20404 8925
rect 20628 8916 20680 8968
rect 21180 8916 21232 8968
rect 21272 8848 21324 8900
rect 18052 8780 18104 8832
rect 18604 8823 18656 8832
rect 18604 8789 18613 8823
rect 18613 8789 18647 8823
rect 18647 8789 18656 8823
rect 18604 8780 18656 8789
rect 18696 8823 18748 8832
rect 18696 8789 18705 8823
rect 18705 8789 18739 8823
rect 18739 8789 18748 8823
rect 18696 8780 18748 8789
rect 18880 8780 18932 8832
rect 20352 8780 20404 8832
rect 21088 8780 21140 8832
rect 21824 8984 21876 9036
rect 21640 8959 21692 8968
rect 21640 8925 21649 8959
rect 21649 8925 21683 8959
rect 21683 8925 21692 8959
rect 21640 8916 21692 8925
rect 22284 8848 22336 8900
rect 23020 8916 23072 8968
rect 23296 8959 23348 8968
rect 23296 8925 23305 8959
rect 23305 8925 23339 8959
rect 23339 8925 23348 8959
rect 23296 8916 23348 8925
rect 23848 8959 23900 8968
rect 23848 8925 23857 8959
rect 23857 8925 23891 8959
rect 23891 8925 23900 8959
rect 23848 8916 23900 8925
rect 24032 8959 24084 8968
rect 24032 8925 24041 8959
rect 24041 8925 24075 8959
rect 24075 8925 24084 8959
rect 24032 8916 24084 8925
rect 23756 8848 23808 8900
rect 23112 8780 23164 8832
rect 24124 8780 24176 8832
rect 24952 8848 25004 8900
rect 10395 8678 10447 8730
rect 10459 8678 10511 8730
rect 10523 8678 10575 8730
rect 10587 8678 10639 8730
rect 10651 8678 10703 8730
rect 19840 8678 19892 8730
rect 19904 8678 19956 8730
rect 19968 8678 20020 8730
rect 20032 8678 20084 8730
rect 20096 8678 20148 8730
rect 5080 8576 5132 8628
rect 6092 8619 6144 8628
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 7564 8619 7616 8628
rect 7564 8585 7573 8619
rect 7573 8585 7607 8619
rect 7607 8585 7616 8619
rect 7564 8576 7616 8585
rect 2228 8440 2280 8492
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 6460 8508 6512 8560
rect 9220 8551 9272 8560
rect 9220 8517 9229 8551
rect 9229 8517 9263 8551
rect 9263 8517 9272 8551
rect 9220 8508 9272 8517
rect 5448 8372 5500 8424
rect 5540 8372 5592 8424
rect 6828 8440 6880 8492
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 9680 8483 9732 8492
rect 9680 8449 9684 8483
rect 9684 8449 9718 8483
rect 9718 8449 9732 8483
rect 9680 8440 9732 8449
rect 9956 8508 10008 8560
rect 12256 8576 12308 8628
rect 12164 8508 12216 8560
rect 12348 8551 12400 8560
rect 12348 8517 12357 8551
rect 12357 8517 12391 8551
rect 12391 8517 12400 8551
rect 12348 8508 12400 8517
rect 2136 8279 2188 8288
rect 2136 8245 2145 8279
rect 2145 8245 2179 8279
rect 2179 8245 2188 8279
rect 2136 8236 2188 8245
rect 4160 8236 4212 8288
rect 6920 8372 6972 8424
rect 7104 8372 7156 8424
rect 8116 8372 8168 8424
rect 9312 8304 9364 8356
rect 10232 8372 10284 8424
rect 10508 8304 10560 8356
rect 6276 8236 6328 8288
rect 9128 8236 9180 8288
rect 9588 8236 9640 8288
rect 10324 8236 10376 8288
rect 10692 8440 10744 8492
rect 10876 8483 10928 8492
rect 10876 8449 10885 8483
rect 10885 8449 10919 8483
rect 10919 8449 10928 8483
rect 10876 8440 10928 8449
rect 12532 8483 12584 8492
rect 12532 8449 12535 8483
rect 12535 8449 12584 8483
rect 12532 8440 12584 8449
rect 14924 8576 14976 8628
rect 16212 8576 16264 8628
rect 19156 8619 19208 8628
rect 13820 8508 13872 8560
rect 15200 8551 15252 8560
rect 15200 8517 15209 8551
rect 15209 8517 15243 8551
rect 15243 8517 15252 8551
rect 15200 8508 15252 8517
rect 14648 8440 14700 8492
rect 12348 8372 12400 8424
rect 12716 8372 12768 8424
rect 13084 8415 13136 8424
rect 13084 8381 13093 8415
rect 13093 8381 13127 8415
rect 13127 8381 13136 8415
rect 13084 8372 13136 8381
rect 14832 8372 14884 8424
rect 15384 8440 15436 8492
rect 15660 8440 15712 8492
rect 17132 8508 17184 8560
rect 18236 8508 18288 8560
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 17960 8483 18012 8492
rect 17960 8449 17969 8483
rect 17969 8449 18003 8483
rect 18003 8449 18012 8483
rect 17960 8440 18012 8449
rect 19156 8585 19165 8619
rect 19165 8585 19199 8619
rect 19199 8585 19208 8619
rect 19156 8576 19208 8585
rect 19340 8619 19392 8628
rect 19340 8585 19349 8619
rect 19349 8585 19383 8619
rect 19383 8585 19392 8619
rect 19340 8576 19392 8585
rect 23020 8576 23072 8628
rect 24032 8619 24084 8628
rect 24032 8585 24041 8619
rect 24041 8585 24075 8619
rect 24075 8585 24084 8619
rect 24032 8576 24084 8585
rect 16948 8372 17000 8424
rect 17316 8415 17368 8424
rect 17316 8381 17325 8415
rect 17325 8381 17359 8415
rect 17359 8381 17368 8415
rect 17316 8372 17368 8381
rect 11336 8347 11388 8356
rect 11336 8313 11345 8347
rect 11345 8313 11379 8347
rect 11379 8313 11388 8347
rect 11336 8304 11388 8313
rect 15936 8304 15988 8356
rect 16212 8304 16264 8356
rect 11888 8236 11940 8288
rect 12624 8279 12676 8288
rect 12624 8245 12633 8279
rect 12633 8245 12667 8279
rect 12667 8245 12676 8279
rect 12624 8236 12676 8245
rect 14924 8236 14976 8288
rect 15476 8236 15528 8288
rect 18512 8415 18564 8424
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 19432 8440 19484 8492
rect 20352 8508 20404 8560
rect 21364 8508 21416 8560
rect 19708 8440 19760 8492
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 21456 8440 21508 8449
rect 21916 8440 21968 8492
rect 22100 8440 22152 8492
rect 22284 8483 22336 8492
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 24124 8483 24176 8492
rect 22284 8440 22336 8449
rect 24124 8449 24133 8483
rect 24133 8449 24167 8483
rect 24167 8449 24176 8483
rect 24124 8440 24176 8449
rect 24492 8440 24544 8492
rect 18604 8347 18656 8356
rect 18604 8313 18613 8347
rect 18613 8313 18647 8347
rect 18647 8313 18656 8347
rect 18604 8304 18656 8313
rect 21640 8415 21692 8424
rect 21640 8381 21649 8415
rect 21649 8381 21683 8415
rect 21683 8381 21692 8415
rect 21640 8372 21692 8381
rect 19340 8304 19392 8356
rect 19708 8304 19760 8356
rect 21548 8304 21600 8356
rect 22008 8304 22060 8356
rect 23112 8304 23164 8356
rect 17684 8236 17736 8288
rect 18880 8236 18932 8288
rect 20996 8236 21048 8288
rect 23204 8236 23256 8288
rect 5672 8134 5724 8186
rect 5736 8134 5788 8186
rect 5800 8134 5852 8186
rect 5864 8134 5916 8186
rect 5928 8134 5980 8186
rect 15118 8134 15170 8186
rect 15182 8134 15234 8186
rect 15246 8134 15298 8186
rect 15310 8134 15362 8186
rect 15374 8134 15426 8186
rect 24563 8134 24615 8186
rect 24627 8134 24679 8186
rect 24691 8134 24743 8186
rect 24755 8134 24807 8186
rect 24819 8134 24871 8186
rect 6460 8032 6512 8084
rect 9220 8032 9272 8084
rect 13084 8032 13136 8084
rect 13728 8075 13780 8084
rect 13728 8041 13737 8075
rect 13737 8041 13771 8075
rect 13771 8041 13780 8075
rect 13728 8032 13780 8041
rect 15016 8075 15068 8084
rect 15016 8041 15025 8075
rect 15025 8041 15059 8075
rect 15059 8041 15068 8075
rect 15016 8032 15068 8041
rect 15660 8032 15712 8084
rect 17960 8032 18012 8084
rect 20536 8032 20588 8084
rect 21180 8032 21232 8084
rect 21272 8032 21324 8084
rect 5540 7964 5592 8016
rect 6092 7964 6144 8016
rect 12532 7964 12584 8016
rect 13176 8007 13228 8016
rect 13176 7973 13185 8007
rect 13185 7973 13219 8007
rect 13219 7973 13228 8007
rect 13176 7964 13228 7973
rect 1400 7828 1452 7880
rect 8300 7896 8352 7948
rect 11060 7896 11112 7948
rect 14832 7964 14884 8016
rect 15384 7964 15436 8016
rect 1768 7803 1820 7812
rect 1768 7769 1802 7803
rect 1802 7769 1820 7803
rect 1768 7760 1820 7769
rect 4344 7760 4396 7812
rect 3516 7692 3568 7744
rect 3976 7692 4028 7744
rect 5264 7735 5316 7744
rect 5264 7701 5273 7735
rect 5273 7701 5307 7735
rect 5307 7701 5316 7735
rect 5540 7828 5592 7880
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 6828 7828 6880 7880
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 12348 7828 12400 7880
rect 6184 7760 6236 7812
rect 9312 7760 9364 7812
rect 10324 7803 10376 7812
rect 10324 7769 10333 7803
rect 10333 7769 10367 7803
rect 10367 7769 10376 7803
rect 10324 7760 10376 7769
rect 11336 7760 11388 7812
rect 11888 7760 11940 7812
rect 13360 7896 13412 7948
rect 14280 7896 14332 7948
rect 17040 7964 17092 8016
rect 17776 8007 17828 8016
rect 17776 7973 17785 8007
rect 17785 7973 17819 8007
rect 17819 7973 17828 8007
rect 17776 7964 17828 7973
rect 21824 8032 21876 8084
rect 21916 7964 21968 8016
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 13176 7828 13228 7880
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 14924 7828 14976 7837
rect 15476 7828 15528 7880
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 15936 7828 15988 7837
rect 16856 7828 16908 7880
rect 17224 7896 17276 7948
rect 25872 8032 25924 8084
rect 23020 7939 23072 7948
rect 23020 7905 23029 7939
rect 23029 7905 23063 7939
rect 23063 7905 23072 7939
rect 23020 7896 23072 7905
rect 17868 7828 17920 7880
rect 18236 7828 18288 7880
rect 19064 7828 19116 7880
rect 21180 7871 21232 7880
rect 21180 7837 21189 7871
rect 21189 7837 21223 7871
rect 21223 7837 21232 7871
rect 21180 7828 21232 7837
rect 24492 7896 24544 7948
rect 24676 7828 24728 7880
rect 15384 7803 15436 7812
rect 5264 7692 5316 7701
rect 7288 7692 7340 7744
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 10232 7692 10284 7744
rect 15384 7769 15393 7803
rect 15393 7769 15427 7803
rect 15427 7769 15436 7803
rect 15384 7760 15436 7769
rect 13360 7692 13412 7744
rect 13544 7692 13596 7744
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 16396 7735 16448 7744
rect 16396 7701 16405 7735
rect 16405 7701 16439 7735
rect 16439 7701 16448 7735
rect 16396 7692 16448 7701
rect 18512 7760 18564 7812
rect 17316 7692 17368 7744
rect 18696 7692 18748 7744
rect 24952 7760 25004 7812
rect 20996 7692 21048 7744
rect 23388 7735 23440 7744
rect 23388 7701 23397 7735
rect 23397 7701 23431 7735
rect 23431 7701 23440 7735
rect 23388 7692 23440 7701
rect 24768 7735 24820 7744
rect 24768 7701 24777 7735
rect 24777 7701 24811 7735
rect 24811 7701 24820 7735
rect 24768 7692 24820 7701
rect 10395 7590 10447 7642
rect 10459 7590 10511 7642
rect 10523 7590 10575 7642
rect 10587 7590 10639 7642
rect 10651 7590 10703 7642
rect 19840 7590 19892 7642
rect 19904 7590 19956 7642
rect 19968 7590 20020 7642
rect 20032 7590 20084 7642
rect 20096 7590 20148 7642
rect 1768 7531 1820 7540
rect 1768 7497 1777 7531
rect 1777 7497 1811 7531
rect 1811 7497 1820 7531
rect 1768 7488 1820 7497
rect 2136 7488 2188 7540
rect 3792 7531 3844 7540
rect 3792 7497 3801 7531
rect 3801 7497 3835 7531
rect 3835 7497 3844 7531
rect 3792 7488 3844 7497
rect 3608 7420 3660 7472
rect 4252 7463 4304 7472
rect 4252 7429 4261 7463
rect 4261 7429 4295 7463
rect 4295 7429 4304 7463
rect 6644 7488 6696 7540
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 7288 7531 7340 7540
rect 7288 7497 7297 7531
rect 7297 7497 7331 7531
rect 7331 7497 7340 7531
rect 7288 7488 7340 7497
rect 11152 7488 11204 7540
rect 11428 7488 11480 7540
rect 14740 7488 14792 7540
rect 4252 7420 4304 7429
rect 3516 7395 3568 7404
rect 2688 7284 2740 7336
rect 2412 7216 2464 7268
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 3608 7327 3660 7336
rect 3608 7293 3617 7327
rect 3617 7293 3651 7327
rect 3651 7293 3660 7327
rect 3608 7284 3660 7293
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 6000 7395 6052 7404
rect 6000 7361 6009 7395
rect 6009 7361 6043 7395
rect 6043 7361 6052 7395
rect 6000 7352 6052 7361
rect 8944 7420 8996 7472
rect 9312 7420 9364 7472
rect 12624 7420 12676 7472
rect 13544 7420 13596 7472
rect 4528 7216 4580 7268
rect 4068 7148 4120 7200
rect 4344 7191 4396 7200
rect 4344 7157 4353 7191
rect 4353 7157 4387 7191
rect 4387 7157 4396 7191
rect 4344 7148 4396 7157
rect 4896 7148 4948 7200
rect 16396 7352 16448 7404
rect 17684 7463 17736 7472
rect 17684 7429 17693 7463
rect 17693 7429 17727 7463
rect 17727 7429 17736 7463
rect 17684 7420 17736 7429
rect 17960 7488 18012 7540
rect 21180 7488 21232 7540
rect 24768 7531 24820 7540
rect 24768 7497 24777 7531
rect 24777 7497 24811 7531
rect 24811 7497 24820 7531
rect 24768 7488 24820 7497
rect 7104 7327 7156 7336
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 7104 7284 7156 7293
rect 9588 7327 9640 7336
rect 9588 7293 9597 7327
rect 9597 7293 9631 7327
rect 9631 7293 9640 7327
rect 9588 7284 9640 7293
rect 12256 7327 12308 7336
rect 12256 7293 12265 7327
rect 12265 7293 12299 7327
rect 12299 7293 12308 7327
rect 12256 7284 12308 7293
rect 17960 7352 18012 7404
rect 18236 7395 18288 7404
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 18512 7352 18564 7404
rect 18972 7420 19024 7472
rect 18788 7352 18840 7404
rect 21364 7420 21416 7472
rect 21824 7420 21876 7472
rect 19708 7352 19760 7404
rect 19800 7284 19852 7336
rect 20260 7327 20312 7336
rect 17868 7259 17920 7268
rect 17868 7225 17877 7259
rect 17877 7225 17911 7259
rect 17911 7225 17920 7259
rect 17868 7216 17920 7225
rect 17960 7216 18012 7268
rect 20260 7293 20269 7327
rect 20269 7293 20303 7327
rect 20303 7293 20312 7327
rect 20260 7284 20312 7293
rect 20444 7352 20496 7404
rect 21088 7395 21140 7404
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 23020 7352 23072 7404
rect 23204 7395 23256 7404
rect 23204 7361 23213 7395
rect 23213 7361 23247 7395
rect 23247 7361 23256 7395
rect 23204 7352 23256 7361
rect 23388 7395 23440 7404
rect 23388 7361 23397 7395
rect 23397 7361 23431 7395
rect 23431 7361 23440 7395
rect 23388 7352 23440 7361
rect 21272 7327 21324 7336
rect 21272 7293 21281 7327
rect 21281 7293 21315 7327
rect 21315 7293 21324 7327
rect 21272 7284 21324 7293
rect 22652 7284 22704 7336
rect 23480 7327 23532 7336
rect 23480 7293 23489 7327
rect 23489 7293 23523 7327
rect 23523 7293 23532 7327
rect 23480 7284 23532 7293
rect 21640 7216 21692 7268
rect 22192 7259 22244 7268
rect 22192 7225 22201 7259
rect 22201 7225 22235 7259
rect 22235 7225 22244 7259
rect 22192 7216 22244 7225
rect 22284 7216 22336 7268
rect 23388 7216 23440 7268
rect 23940 7352 23992 7404
rect 24676 7420 24728 7472
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 25780 7395 25832 7404
rect 25780 7361 25789 7395
rect 25789 7361 25823 7395
rect 25823 7361 25832 7395
rect 25780 7352 25832 7361
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 14004 7191 14056 7200
rect 14004 7157 14013 7191
rect 14013 7157 14047 7191
rect 14047 7157 14056 7191
rect 14004 7148 14056 7157
rect 14740 7148 14792 7200
rect 18052 7148 18104 7200
rect 18696 7191 18748 7200
rect 18696 7157 18705 7191
rect 18705 7157 18739 7191
rect 18739 7157 18748 7191
rect 18696 7148 18748 7157
rect 25964 7191 26016 7200
rect 25964 7157 25973 7191
rect 25973 7157 26007 7191
rect 26007 7157 26016 7191
rect 25964 7148 26016 7157
rect 5672 7046 5724 7098
rect 5736 7046 5788 7098
rect 5800 7046 5852 7098
rect 5864 7046 5916 7098
rect 5928 7046 5980 7098
rect 15118 7046 15170 7098
rect 15182 7046 15234 7098
rect 15246 7046 15298 7098
rect 15310 7046 15362 7098
rect 15374 7046 15426 7098
rect 24563 7046 24615 7098
rect 24627 7046 24679 7098
rect 24691 7046 24743 7098
rect 24755 7046 24807 7098
rect 24819 7046 24871 7098
rect 2688 6987 2740 6996
rect 2688 6953 2697 6987
rect 2697 6953 2731 6987
rect 2731 6953 2740 6987
rect 2688 6944 2740 6953
rect 6000 6944 6052 6996
rect 10324 6944 10376 6996
rect 11980 6944 12032 6996
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 18052 6944 18104 6996
rect 18604 6987 18656 6996
rect 18604 6953 18613 6987
rect 18613 6953 18647 6987
rect 18647 6953 18656 6987
rect 18604 6944 18656 6953
rect 18972 6944 19024 6996
rect 20260 6987 20312 6996
rect 20260 6953 20269 6987
rect 20269 6953 20303 6987
rect 20303 6953 20312 6987
rect 20260 6944 20312 6953
rect 22100 6944 22152 6996
rect 25780 6987 25832 6996
rect 2228 6808 2280 6860
rect 4528 6876 4580 6928
rect 19708 6876 19760 6928
rect 20076 6876 20128 6928
rect 21088 6876 21140 6928
rect 12072 6808 12124 6860
rect 13912 6808 13964 6860
rect 17776 6851 17828 6860
rect 2412 6740 2464 6792
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 4620 6740 4672 6792
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 5540 6740 5592 6792
rect 4160 6672 4212 6724
rect 4252 6672 4304 6724
rect 6000 6672 6052 6724
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 7104 6740 7156 6792
rect 7748 6740 7800 6792
rect 8392 6740 8444 6792
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 3240 6604 3292 6656
rect 8852 6672 8904 6724
rect 9220 6604 9272 6656
rect 11888 6740 11940 6792
rect 16948 6740 17000 6792
rect 17132 6740 17184 6792
rect 11244 6604 11296 6656
rect 17776 6817 17785 6851
rect 17785 6817 17819 6851
rect 17819 6817 17828 6851
rect 17776 6808 17828 6817
rect 19800 6808 19852 6860
rect 20444 6808 20496 6860
rect 20536 6808 20588 6860
rect 21272 6808 21324 6860
rect 21364 6851 21416 6860
rect 21364 6817 21373 6851
rect 21373 6817 21407 6851
rect 21407 6817 21416 6851
rect 21364 6808 21416 6817
rect 22100 6808 22152 6860
rect 17960 6740 18012 6792
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 18880 6740 18932 6792
rect 21548 6783 21600 6792
rect 12256 6604 12308 6656
rect 14464 6647 14516 6656
rect 14464 6613 14473 6647
rect 14473 6613 14507 6647
rect 14507 6613 14516 6647
rect 14464 6604 14516 6613
rect 14832 6647 14884 6656
rect 14832 6613 14841 6647
rect 14841 6613 14875 6647
rect 14875 6613 14884 6647
rect 14832 6604 14884 6613
rect 14924 6647 14976 6656
rect 14924 6613 14933 6647
rect 14933 6613 14967 6647
rect 14967 6613 14976 6647
rect 20076 6672 20128 6724
rect 14924 6604 14976 6613
rect 17960 6604 18012 6656
rect 18236 6604 18288 6656
rect 20260 6604 20312 6656
rect 20536 6604 20588 6656
rect 21548 6749 21557 6783
rect 21557 6749 21591 6783
rect 21591 6749 21600 6783
rect 21548 6740 21600 6749
rect 25780 6953 25789 6987
rect 25789 6953 25823 6987
rect 25823 6953 25832 6987
rect 25780 6944 25832 6953
rect 22652 6876 22704 6928
rect 23388 6876 23440 6928
rect 22284 6740 22336 6792
rect 22928 6808 22980 6860
rect 23204 6783 23256 6792
rect 22468 6672 22520 6724
rect 21548 6604 21600 6656
rect 23204 6749 23213 6783
rect 23213 6749 23247 6783
rect 23247 6749 23256 6783
rect 23204 6740 23256 6749
rect 24860 6876 24912 6928
rect 25044 6740 25096 6792
rect 25320 6783 25372 6792
rect 25320 6749 25329 6783
rect 25329 6749 25363 6783
rect 25363 6749 25372 6783
rect 25320 6740 25372 6749
rect 24952 6672 25004 6724
rect 25504 6715 25556 6724
rect 25504 6681 25513 6715
rect 25513 6681 25547 6715
rect 25547 6681 25556 6715
rect 25504 6672 25556 6681
rect 25688 6715 25740 6724
rect 25688 6681 25697 6715
rect 25697 6681 25731 6715
rect 25731 6681 25740 6715
rect 25688 6672 25740 6681
rect 24860 6604 24912 6656
rect 25136 6604 25188 6656
rect 27712 6604 27764 6656
rect 10395 6502 10447 6554
rect 10459 6502 10511 6554
rect 10523 6502 10575 6554
rect 10587 6502 10639 6554
rect 10651 6502 10703 6554
rect 19840 6502 19892 6554
rect 19904 6502 19956 6554
rect 19968 6502 20020 6554
rect 20032 6502 20084 6554
rect 20096 6502 20148 6554
rect 4344 6400 4396 6452
rect 4620 6400 4672 6452
rect 4068 6332 4120 6384
rect 10232 6400 10284 6452
rect 12072 6400 12124 6452
rect 12256 6443 12308 6452
rect 12256 6409 12265 6443
rect 12265 6409 12299 6443
rect 12299 6409 12308 6443
rect 12256 6400 12308 6409
rect 14924 6400 14976 6452
rect 20352 6400 20404 6452
rect 22468 6443 22520 6452
rect 6000 6375 6052 6384
rect 6000 6341 6009 6375
rect 6009 6341 6043 6375
rect 6043 6341 6052 6375
rect 6000 6332 6052 6341
rect 2228 6264 2280 6316
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 4252 6264 4304 6316
rect 4620 6264 4672 6316
rect 4896 6264 4948 6316
rect 6184 6264 6236 6316
rect 1492 6239 1544 6248
rect 1492 6205 1501 6239
rect 1501 6205 1535 6239
rect 1535 6205 1544 6239
rect 1492 6196 1544 6205
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 8852 6307 8904 6316
rect 6368 6264 6420 6273
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 11060 6332 11112 6384
rect 11888 6332 11940 6384
rect 14464 6375 14516 6384
rect 9404 6307 9456 6316
rect 9404 6273 9438 6307
rect 9438 6273 9456 6307
rect 9404 6264 9456 6273
rect 11704 6264 11756 6316
rect 4804 6128 4856 6180
rect 5448 6128 5500 6180
rect 3332 6060 3384 6112
rect 5264 6060 5316 6112
rect 6000 6128 6052 6180
rect 12164 6307 12216 6316
rect 12164 6273 12173 6307
rect 12173 6273 12207 6307
rect 12207 6273 12216 6307
rect 12164 6264 12216 6273
rect 12900 6307 12952 6316
rect 12900 6273 12934 6307
rect 12934 6273 12952 6307
rect 14464 6341 14498 6375
rect 14498 6341 14516 6375
rect 14464 6332 14516 6341
rect 12900 6264 12952 6273
rect 12348 6196 12400 6248
rect 15476 6264 15528 6316
rect 18696 6332 18748 6384
rect 20076 6332 20128 6384
rect 22468 6409 22477 6443
rect 22477 6409 22511 6443
rect 22511 6409 22520 6443
rect 22468 6400 22520 6409
rect 22652 6400 22704 6452
rect 22928 6443 22980 6452
rect 22928 6409 22937 6443
rect 22937 6409 22971 6443
rect 22971 6409 22980 6443
rect 22928 6400 22980 6409
rect 24768 6443 24820 6452
rect 24768 6409 24777 6443
rect 24777 6409 24811 6443
rect 24811 6409 24820 6443
rect 24768 6400 24820 6409
rect 25136 6443 25188 6452
rect 25136 6409 25145 6443
rect 25145 6409 25179 6443
rect 25179 6409 25188 6443
rect 25136 6400 25188 6409
rect 25320 6400 25372 6452
rect 25964 6400 26016 6452
rect 21548 6332 21600 6384
rect 16948 6264 17000 6316
rect 17960 6307 18012 6316
rect 17960 6273 17969 6307
rect 17969 6273 18003 6307
rect 18003 6273 18012 6307
rect 17960 6264 18012 6273
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 19892 6307 19944 6316
rect 18604 6264 18656 6273
rect 19892 6273 19901 6307
rect 19901 6273 19935 6307
rect 19935 6273 19944 6307
rect 19892 6264 19944 6273
rect 20812 6307 20864 6316
rect 20812 6273 20821 6307
rect 20821 6273 20855 6307
rect 20855 6273 20864 6307
rect 20812 6264 20864 6273
rect 26240 6332 26292 6384
rect 9772 6060 9824 6112
rect 11152 6060 11204 6112
rect 11704 6060 11756 6112
rect 12164 6060 12216 6112
rect 18052 6196 18104 6248
rect 23204 6264 23256 6316
rect 24860 6264 24912 6316
rect 25504 6264 25556 6316
rect 14372 6060 14424 6112
rect 14556 6060 14608 6112
rect 19340 6128 19392 6180
rect 23388 6239 23440 6248
rect 23388 6205 23397 6239
rect 23397 6205 23431 6239
rect 23431 6205 23440 6239
rect 23388 6196 23440 6205
rect 24492 6239 24544 6248
rect 23020 6128 23072 6180
rect 24492 6205 24501 6239
rect 24501 6205 24535 6239
rect 24535 6205 24544 6239
rect 24492 6196 24544 6205
rect 25964 6239 26016 6248
rect 24124 6128 24176 6180
rect 25964 6205 25973 6239
rect 25973 6205 26007 6239
rect 26007 6205 26016 6239
rect 25964 6196 26016 6205
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 18788 6060 18840 6112
rect 19708 6103 19760 6112
rect 19708 6069 19717 6103
rect 19717 6069 19751 6103
rect 19751 6069 19760 6103
rect 19708 6060 19760 6069
rect 22192 6060 22244 6112
rect 24400 6060 24452 6112
rect 5672 5958 5724 6010
rect 5736 5958 5788 6010
rect 5800 5958 5852 6010
rect 5864 5958 5916 6010
rect 5928 5958 5980 6010
rect 15118 5958 15170 6010
rect 15182 5958 15234 6010
rect 15246 5958 15298 6010
rect 15310 5958 15362 6010
rect 15374 5958 15426 6010
rect 24563 5958 24615 6010
rect 24627 5958 24679 6010
rect 24691 5958 24743 6010
rect 24755 5958 24807 6010
rect 24819 5958 24871 6010
rect 2228 5899 2280 5908
rect 2228 5865 2237 5899
rect 2237 5865 2271 5899
rect 2271 5865 2280 5899
rect 2228 5856 2280 5865
rect 4896 5899 4948 5908
rect 4896 5865 4905 5899
rect 4905 5865 4939 5899
rect 4939 5865 4948 5899
rect 4896 5856 4948 5865
rect 6092 5856 6144 5908
rect 6368 5856 6420 5908
rect 9404 5856 9456 5908
rect 14832 5856 14884 5908
rect 18696 5899 18748 5908
rect 18696 5865 18705 5899
rect 18705 5865 18739 5899
rect 18739 5865 18748 5899
rect 18696 5856 18748 5865
rect 2596 5788 2648 5840
rect 4160 5788 4212 5840
rect 5816 5788 5868 5840
rect 6184 5788 6236 5840
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 3148 5559 3200 5568
rect 2688 5516 2740 5525
rect 3148 5525 3157 5559
rect 3157 5525 3191 5559
rect 3191 5525 3200 5559
rect 3148 5516 3200 5525
rect 4712 5720 4764 5772
rect 6276 5720 6328 5772
rect 9772 5763 9824 5772
rect 4252 5652 4304 5704
rect 5264 5695 5316 5704
rect 4620 5627 4672 5636
rect 4620 5593 4629 5627
rect 4629 5593 4663 5627
rect 4663 5593 4672 5627
rect 4620 5584 4672 5593
rect 4804 5627 4856 5636
rect 4804 5593 4813 5627
rect 4813 5593 4847 5627
rect 4847 5593 4856 5627
rect 4804 5584 4856 5593
rect 4068 5516 4120 5568
rect 4896 5516 4948 5568
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 5908 5652 5960 5704
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 9772 5729 9781 5763
rect 9781 5729 9815 5763
rect 9815 5729 9824 5763
rect 9772 5720 9824 5729
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 6184 5652 6236 5661
rect 8484 5652 8536 5704
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 13820 5652 13872 5704
rect 14556 5652 14608 5704
rect 15292 5788 15344 5840
rect 15568 5788 15620 5840
rect 19616 5831 19668 5840
rect 15200 5695 15252 5704
rect 15200 5661 15209 5695
rect 15209 5661 15243 5695
rect 15243 5661 15252 5695
rect 15200 5652 15252 5661
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 18420 5652 18472 5704
rect 19616 5797 19625 5831
rect 19625 5797 19659 5831
rect 19659 5797 19668 5831
rect 19616 5788 19668 5797
rect 19892 5856 19944 5908
rect 20812 5856 20864 5908
rect 21088 5899 21140 5908
rect 20076 5788 20128 5840
rect 19432 5720 19484 5772
rect 18696 5695 18748 5704
rect 18696 5661 18705 5695
rect 18705 5661 18739 5695
rect 18739 5661 18748 5695
rect 18696 5652 18748 5661
rect 6000 5627 6052 5636
rect 6000 5593 6009 5627
rect 6009 5593 6043 5627
rect 6043 5593 6052 5627
rect 6000 5584 6052 5593
rect 8300 5627 8352 5636
rect 8300 5593 8318 5627
rect 8318 5593 8352 5627
rect 8300 5584 8352 5593
rect 12072 5584 12124 5636
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 9496 5516 9548 5568
rect 12624 5516 12676 5568
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 13268 5516 13320 5568
rect 17684 5559 17736 5568
rect 17684 5525 17693 5559
rect 17693 5525 17727 5559
rect 17727 5525 17736 5559
rect 17684 5516 17736 5525
rect 18052 5516 18104 5568
rect 19524 5695 19576 5704
rect 19524 5661 19533 5695
rect 19533 5661 19567 5695
rect 19567 5661 19576 5695
rect 19524 5652 19576 5661
rect 20076 5695 20128 5704
rect 20076 5661 20085 5695
rect 20085 5661 20119 5695
rect 20119 5661 20128 5695
rect 20076 5652 20128 5661
rect 20260 5695 20312 5704
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 21088 5865 21097 5899
rect 21097 5865 21131 5899
rect 21131 5865 21140 5899
rect 21088 5856 21140 5865
rect 21640 5899 21692 5908
rect 21640 5865 21649 5899
rect 21649 5865 21683 5899
rect 21683 5865 21692 5899
rect 21640 5856 21692 5865
rect 22376 5856 22428 5908
rect 23296 5856 23348 5908
rect 24124 5899 24176 5908
rect 20996 5788 21048 5840
rect 22008 5788 22060 5840
rect 23388 5788 23440 5840
rect 24124 5865 24133 5899
rect 24133 5865 24167 5899
rect 24167 5865 24176 5899
rect 24124 5856 24176 5865
rect 24400 5856 24452 5908
rect 24768 5788 24820 5840
rect 20628 5584 20680 5636
rect 24308 5720 24360 5772
rect 22008 5652 22060 5704
rect 22652 5695 22704 5704
rect 20996 5516 21048 5568
rect 21456 5516 21508 5568
rect 22008 5516 22060 5568
rect 22652 5661 22661 5695
rect 22661 5661 22695 5695
rect 22695 5661 22704 5695
rect 22652 5652 22704 5661
rect 24124 5695 24176 5704
rect 24124 5661 24133 5695
rect 24133 5661 24167 5695
rect 24167 5661 24176 5695
rect 24400 5695 24452 5704
rect 24124 5652 24176 5661
rect 24400 5661 24409 5695
rect 24409 5661 24443 5695
rect 24443 5661 24452 5695
rect 24400 5652 24452 5661
rect 25688 5720 25740 5772
rect 25596 5652 25648 5704
rect 26424 5584 26476 5636
rect 23756 5559 23808 5568
rect 23756 5525 23765 5559
rect 23765 5525 23799 5559
rect 23799 5525 23808 5559
rect 23756 5516 23808 5525
rect 10395 5414 10447 5466
rect 10459 5414 10511 5466
rect 10523 5414 10575 5466
rect 10587 5414 10639 5466
rect 10651 5414 10703 5466
rect 19840 5414 19892 5466
rect 19904 5414 19956 5466
rect 19968 5414 20020 5466
rect 20032 5414 20084 5466
rect 20096 5414 20148 5466
rect 2688 5312 2740 5364
rect 4252 5355 4304 5364
rect 4252 5321 4261 5355
rect 4261 5321 4295 5355
rect 4295 5321 4304 5355
rect 4252 5312 4304 5321
rect 5816 5287 5868 5296
rect 5816 5253 5825 5287
rect 5825 5253 5859 5287
rect 5859 5253 5868 5287
rect 5816 5244 5868 5253
rect 6092 5244 6144 5296
rect 6276 5244 6328 5296
rect 11428 5312 11480 5364
rect 11704 5355 11756 5364
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 12900 5312 12952 5364
rect 13176 5312 13228 5364
rect 15200 5312 15252 5364
rect 3148 5176 3200 5228
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 4068 5108 4120 5160
rect 3976 5040 4028 5092
rect 12624 5287 12676 5296
rect 7012 5176 7064 5228
rect 7104 5108 7156 5160
rect 9220 5108 9272 5160
rect 10600 5176 10652 5228
rect 10876 5219 10928 5228
rect 10876 5185 10885 5219
rect 10885 5185 10919 5219
rect 10919 5185 10928 5219
rect 10876 5176 10928 5185
rect 11060 5219 11112 5228
rect 11060 5185 11069 5219
rect 11069 5185 11103 5219
rect 11103 5185 11112 5219
rect 11060 5176 11112 5185
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 11428 5176 11480 5228
rect 12072 5219 12124 5228
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 12624 5253 12633 5287
rect 12633 5253 12667 5287
rect 12667 5253 12676 5287
rect 12624 5244 12676 5253
rect 13820 5287 13872 5296
rect 13820 5253 13829 5287
rect 13829 5253 13863 5287
rect 13863 5253 13872 5287
rect 13820 5244 13872 5253
rect 14372 5244 14424 5296
rect 12716 5219 12768 5228
rect 10692 5151 10744 5160
rect 10692 5117 10701 5151
rect 10701 5117 10735 5151
rect 10735 5117 10744 5151
rect 11520 5151 11572 5160
rect 10692 5108 10744 5117
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 12716 5185 12725 5219
rect 12725 5185 12759 5219
rect 12759 5185 12768 5219
rect 12716 5176 12768 5185
rect 13268 5176 13320 5228
rect 14556 5176 14608 5228
rect 15016 5219 15068 5228
rect 13820 5108 13872 5160
rect 14372 5151 14424 5160
rect 14372 5117 14381 5151
rect 14381 5117 14415 5151
rect 14415 5117 14424 5151
rect 14372 5108 14424 5117
rect 14464 5151 14516 5160
rect 14464 5117 14473 5151
rect 14473 5117 14507 5151
rect 14507 5117 14516 5151
rect 14464 5108 14516 5117
rect 8300 5040 8352 5092
rect 9496 5083 9548 5092
rect 9496 5049 9505 5083
rect 9505 5049 9539 5083
rect 9539 5049 9548 5083
rect 9496 5040 9548 5049
rect 13544 5040 13596 5092
rect 15016 5185 15025 5219
rect 15025 5185 15059 5219
rect 15059 5185 15068 5219
rect 15016 5176 15068 5185
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 17684 5312 17736 5364
rect 19708 5312 19760 5364
rect 20628 5355 20680 5364
rect 17592 5244 17644 5296
rect 17776 5244 17828 5296
rect 19524 5244 19576 5296
rect 20628 5321 20637 5355
rect 20637 5321 20671 5355
rect 20671 5321 20680 5355
rect 20628 5312 20680 5321
rect 19708 5176 19760 5228
rect 22284 5244 22336 5296
rect 20812 5219 20864 5228
rect 20812 5185 20821 5219
rect 20821 5185 20855 5219
rect 20855 5185 20864 5219
rect 20812 5176 20864 5185
rect 21916 5219 21968 5228
rect 21916 5185 21925 5219
rect 21925 5185 21959 5219
rect 21959 5185 21968 5219
rect 21916 5176 21968 5185
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22376 5219 22428 5228
rect 22100 5176 22152 5185
rect 22376 5185 22385 5219
rect 22385 5185 22419 5219
rect 22419 5185 22428 5219
rect 22376 5176 22428 5185
rect 15844 5108 15896 5160
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 19248 5108 19300 5160
rect 19432 5108 19484 5160
rect 21364 5108 21416 5160
rect 3884 5015 3936 5024
rect 3884 4981 3893 5015
rect 3893 4981 3927 5015
rect 3927 4981 3936 5015
rect 3884 4972 3936 4981
rect 8760 4972 8812 5024
rect 13360 4972 13412 5024
rect 18420 5040 18472 5092
rect 21456 5040 21508 5092
rect 17408 4972 17460 5024
rect 20260 4972 20312 5024
rect 23388 5176 23440 5228
rect 23756 5219 23808 5228
rect 23756 5185 23765 5219
rect 23765 5185 23799 5219
rect 23799 5185 23808 5219
rect 23756 5176 23808 5185
rect 24400 5312 24452 5364
rect 24124 5244 24176 5296
rect 24768 5219 24820 5228
rect 24768 5185 24777 5219
rect 24777 5185 24811 5219
rect 24811 5185 24820 5219
rect 24768 5176 24820 5185
rect 22836 5108 22888 5160
rect 23020 5040 23072 5092
rect 22928 4972 22980 5024
rect 23572 5015 23624 5024
rect 23572 4981 23581 5015
rect 23581 4981 23615 5015
rect 23615 4981 23624 5015
rect 23572 4972 23624 4981
rect 25044 5219 25096 5228
rect 25044 5185 25053 5219
rect 25053 5185 25087 5219
rect 25087 5185 25096 5219
rect 25044 5176 25096 5185
rect 27252 5312 27304 5364
rect 25596 5176 25648 5228
rect 26424 5219 26476 5228
rect 26424 5185 26433 5219
rect 26433 5185 26467 5219
rect 26467 5185 26476 5219
rect 26424 5176 26476 5185
rect 27436 5219 27488 5228
rect 27436 5185 27459 5219
rect 27459 5185 27488 5219
rect 27436 5176 27488 5185
rect 27712 5219 27764 5228
rect 27712 5185 27721 5219
rect 27721 5185 27755 5219
rect 27755 5185 27764 5219
rect 27712 5176 27764 5185
rect 24492 5040 24544 5092
rect 27528 5108 27580 5160
rect 27344 5040 27396 5092
rect 26884 4972 26936 5024
rect 5672 4870 5724 4922
rect 5736 4870 5788 4922
rect 5800 4870 5852 4922
rect 5864 4870 5916 4922
rect 5928 4870 5980 4922
rect 15118 4870 15170 4922
rect 15182 4870 15234 4922
rect 15246 4870 15298 4922
rect 15310 4870 15362 4922
rect 15374 4870 15426 4922
rect 24563 4870 24615 4922
rect 24627 4870 24679 4922
rect 24691 4870 24743 4922
rect 24755 4870 24807 4922
rect 24819 4870 24871 4922
rect 4804 4768 4856 4820
rect 10600 4811 10652 4820
rect 10600 4777 10609 4811
rect 10609 4777 10643 4811
rect 10643 4777 10652 4811
rect 10600 4768 10652 4777
rect 10876 4700 10928 4752
rect 12992 4768 13044 4820
rect 15476 4768 15528 4820
rect 15844 4811 15896 4820
rect 15844 4777 15853 4811
rect 15853 4777 15887 4811
rect 15887 4777 15896 4811
rect 15844 4768 15896 4777
rect 14556 4743 14608 4752
rect 1492 4632 1544 4684
rect 1584 4564 1636 4616
rect 8484 4632 8536 4684
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 3884 4564 3936 4616
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 8760 4564 8812 4616
rect 10692 4607 10744 4616
rect 10692 4573 10702 4607
rect 10702 4573 10736 4607
rect 10736 4573 10744 4607
rect 10692 4564 10744 4573
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 8944 4496 8996 4548
rect 11060 4496 11112 4548
rect 12716 4632 12768 4684
rect 14556 4709 14565 4743
rect 14565 4709 14599 4743
rect 14599 4709 14608 4743
rect 14556 4700 14608 4709
rect 14740 4700 14792 4752
rect 19340 4700 19392 4752
rect 22468 4768 22520 4820
rect 22836 4811 22888 4820
rect 22836 4777 22845 4811
rect 22845 4777 22879 4811
rect 22879 4777 22888 4811
rect 22836 4768 22888 4777
rect 22928 4768 22980 4820
rect 25044 4768 25096 4820
rect 25596 4811 25648 4820
rect 25596 4777 25605 4811
rect 25605 4777 25639 4811
rect 25639 4777 25648 4811
rect 25596 4768 25648 4777
rect 25964 4768 26016 4820
rect 13176 4564 13228 4616
rect 13360 4564 13412 4616
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 15016 4632 15068 4684
rect 19708 4675 19760 4684
rect 19708 4641 19717 4675
rect 19717 4641 19751 4675
rect 19751 4641 19760 4675
rect 19708 4632 19760 4641
rect 26240 4700 26292 4752
rect 27344 4743 27396 4752
rect 14464 4564 14516 4616
rect 1400 4471 1452 4480
rect 1400 4437 1409 4471
rect 1409 4437 1443 4471
rect 1443 4437 1452 4471
rect 1400 4428 1452 4437
rect 6920 4428 6972 4480
rect 7012 4471 7064 4480
rect 7012 4437 7021 4471
rect 7021 4437 7055 4471
rect 7055 4437 7064 4471
rect 7012 4428 7064 4437
rect 9404 4428 9456 4480
rect 11152 4428 11204 4480
rect 12440 4539 12492 4548
rect 12440 4505 12449 4539
rect 12449 4505 12483 4539
rect 12483 4505 12492 4539
rect 14372 4539 14424 4548
rect 12440 4496 12492 4505
rect 14372 4505 14381 4539
rect 14381 4505 14415 4539
rect 14415 4505 14424 4539
rect 16672 4564 16724 4616
rect 17132 4564 17184 4616
rect 17776 4607 17828 4616
rect 17776 4573 17785 4607
rect 17785 4573 17819 4607
rect 17819 4573 17828 4607
rect 17776 4564 17828 4573
rect 19616 4607 19668 4616
rect 19616 4573 19625 4607
rect 19625 4573 19659 4607
rect 19659 4573 19668 4607
rect 19616 4564 19668 4573
rect 21364 4607 21416 4616
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 22008 4564 22060 4616
rect 22376 4564 22428 4616
rect 23572 4675 23624 4684
rect 14372 4496 14424 4505
rect 15476 4496 15528 4548
rect 17408 4496 17460 4548
rect 21916 4539 21968 4548
rect 21916 4505 21925 4539
rect 21925 4505 21959 4539
rect 21959 4505 21968 4539
rect 21916 4496 21968 4505
rect 22284 4496 22336 4548
rect 23572 4641 23581 4675
rect 23581 4641 23615 4675
rect 23615 4641 23624 4675
rect 23572 4632 23624 4641
rect 23480 4564 23532 4616
rect 24400 4632 24452 4684
rect 25872 4632 25924 4684
rect 26884 4675 26936 4684
rect 26884 4641 26893 4675
rect 26893 4641 26927 4675
rect 26927 4641 26936 4675
rect 26884 4632 26936 4641
rect 27344 4709 27353 4743
rect 27353 4709 27387 4743
rect 27387 4709 27396 4743
rect 27344 4700 27396 4709
rect 24124 4564 24176 4616
rect 27436 4632 27488 4684
rect 27252 4607 27304 4616
rect 27252 4573 27261 4607
rect 27261 4573 27295 4607
rect 27295 4573 27304 4607
rect 27528 4607 27580 4616
rect 27252 4564 27304 4573
rect 27528 4573 27537 4607
rect 27537 4573 27571 4607
rect 27571 4573 27580 4607
rect 27528 4564 27580 4573
rect 24492 4496 24544 4548
rect 13268 4428 13320 4480
rect 17960 4428 18012 4480
rect 19064 4428 19116 4480
rect 19524 4428 19576 4480
rect 20996 4471 21048 4480
rect 20996 4437 21005 4471
rect 21005 4437 21039 4471
rect 21039 4437 21048 4471
rect 20996 4428 21048 4437
rect 22468 4471 22520 4480
rect 22468 4437 22477 4471
rect 22477 4437 22511 4471
rect 22511 4437 22520 4471
rect 22468 4428 22520 4437
rect 23388 4428 23440 4480
rect 23480 4428 23532 4480
rect 24124 4428 24176 4480
rect 25136 4471 25188 4480
rect 25136 4437 25145 4471
rect 25145 4437 25179 4471
rect 25179 4437 25188 4471
rect 25136 4428 25188 4437
rect 26240 4428 26292 4480
rect 10395 4326 10447 4378
rect 10459 4326 10511 4378
rect 10523 4326 10575 4378
rect 10587 4326 10639 4378
rect 10651 4326 10703 4378
rect 19840 4326 19892 4378
rect 19904 4326 19956 4378
rect 19968 4326 20020 4378
rect 20032 4326 20084 4378
rect 20096 4326 20148 4378
rect 6920 4224 6972 4276
rect 8944 4267 8996 4276
rect 8944 4233 8953 4267
rect 8953 4233 8987 4267
rect 8987 4233 8996 4267
rect 8944 4224 8996 4233
rect 9404 4267 9456 4276
rect 9404 4233 9413 4267
rect 9413 4233 9447 4267
rect 9447 4233 9456 4267
rect 9404 4224 9456 4233
rect 13544 4224 13596 4276
rect 3792 4156 3844 4208
rect 5908 4131 5960 4140
rect 5908 4097 5926 4131
rect 5926 4097 5960 4131
rect 5908 4088 5960 4097
rect 9496 4156 9548 4208
rect 11244 4199 11296 4208
rect 11244 4165 11253 4199
rect 11253 4165 11287 4199
rect 11287 4165 11296 4199
rect 11244 4156 11296 4165
rect 12440 4156 12492 4208
rect 15660 4156 15712 4208
rect 17960 4156 18012 4208
rect 18420 4199 18472 4208
rect 18420 4165 18429 4199
rect 18429 4165 18463 4199
rect 18463 4165 18472 4199
rect 18420 4156 18472 4165
rect 18512 4156 18564 4208
rect 19708 4224 19760 4276
rect 21916 4224 21968 4276
rect 22376 4224 22428 4276
rect 23480 4224 23532 4276
rect 23572 4224 23624 4276
rect 26240 4224 26292 4276
rect 27252 4267 27304 4276
rect 27252 4233 27261 4267
rect 27261 4233 27295 4267
rect 27295 4233 27304 4267
rect 27252 4224 27304 4233
rect 19064 4156 19116 4208
rect 6644 4020 6696 4072
rect 7012 4063 7064 4072
rect 7012 4029 7021 4063
rect 7021 4029 7055 4063
rect 7055 4029 7064 4063
rect 9864 4088 9916 4140
rect 10140 4088 10192 4140
rect 11152 4088 11204 4140
rect 13176 4088 13228 4140
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 13728 4131 13780 4140
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 15568 4088 15620 4140
rect 15752 4088 15804 4140
rect 16948 4131 17000 4140
rect 16948 4097 16957 4131
rect 16957 4097 16991 4131
rect 16991 4097 17000 4131
rect 16948 4088 17000 4097
rect 17592 4131 17644 4140
rect 17592 4097 17601 4131
rect 17601 4097 17635 4131
rect 17635 4097 17644 4131
rect 17592 4088 17644 4097
rect 7012 4020 7064 4029
rect 6736 3952 6788 4004
rect 9588 4020 9640 4072
rect 14648 4020 14700 4072
rect 16580 4020 16632 4072
rect 12808 3952 12860 4004
rect 18144 3952 18196 4004
rect 20720 4131 20772 4140
rect 20720 4097 20729 4131
rect 20729 4097 20763 4131
rect 20763 4097 20772 4131
rect 20720 4088 20772 4097
rect 25136 4156 25188 4208
rect 27528 4156 27580 4208
rect 21272 4088 21324 4140
rect 23940 4088 23992 4140
rect 26516 4088 26568 4140
rect 21548 4020 21600 4072
rect 22468 3952 22520 4004
rect 5448 3884 5500 3936
rect 6000 3884 6052 3936
rect 6460 3884 6512 3936
rect 11060 3884 11112 3936
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 12164 3884 12216 3893
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 15016 3884 15068 3936
rect 18420 3884 18472 3936
rect 19064 3884 19116 3936
rect 22744 3884 22796 3936
rect 29828 4088 29880 4140
rect 24952 3884 25004 3936
rect 5672 3782 5724 3834
rect 5736 3782 5788 3834
rect 5800 3782 5852 3834
rect 5864 3782 5916 3834
rect 5928 3782 5980 3834
rect 15118 3782 15170 3834
rect 15182 3782 15234 3834
rect 15246 3782 15298 3834
rect 15310 3782 15362 3834
rect 15374 3782 15426 3834
rect 24563 3782 24615 3834
rect 24627 3782 24679 3834
rect 24691 3782 24743 3834
rect 24755 3782 24807 3834
rect 24819 3782 24871 3834
rect 6644 3723 6696 3732
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 9220 3680 9272 3732
rect 9404 3680 9456 3732
rect 4160 3612 4212 3664
rect 9588 3612 9640 3664
rect 1768 3544 1820 3596
rect 6368 3544 6420 3596
rect 6644 3544 6696 3596
rect 8116 3544 8168 3596
rect 12716 3680 12768 3732
rect 13176 3723 13228 3732
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 5448 3408 5500 3460
rect 7932 3408 7984 3460
rect 9036 3408 9088 3460
rect 11060 3612 11112 3664
rect 11244 3544 11296 3596
rect 13176 3689 13185 3723
rect 13185 3689 13219 3723
rect 13219 3689 13228 3723
rect 13176 3680 13228 3689
rect 15476 3680 15528 3732
rect 17592 3723 17644 3732
rect 13544 3612 13596 3664
rect 15844 3612 15896 3664
rect 17592 3689 17601 3723
rect 17601 3689 17635 3723
rect 17635 3689 17644 3723
rect 17592 3680 17644 3689
rect 21272 3723 21324 3732
rect 21272 3689 21281 3723
rect 21281 3689 21315 3723
rect 21315 3689 21324 3723
rect 21272 3680 21324 3689
rect 21548 3680 21600 3732
rect 22468 3723 22520 3732
rect 13360 3544 13412 3596
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11520 3519 11572 3528
rect 11060 3476 11112 3485
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 13268 3519 13320 3528
rect 13268 3485 13278 3519
rect 13278 3485 13312 3519
rect 13312 3485 13320 3519
rect 13728 3587 13780 3596
rect 13728 3553 13737 3587
rect 13737 3553 13771 3587
rect 13771 3553 13780 3587
rect 13728 3544 13780 3553
rect 13268 3476 13320 3485
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 15660 3544 15712 3596
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15068 3519
rect 15016 3476 15068 3485
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 15568 3476 15620 3528
rect 16580 3544 16632 3596
rect 17132 3587 17184 3596
rect 17132 3553 17141 3587
rect 17141 3553 17175 3587
rect 17175 3553 17184 3587
rect 17132 3544 17184 3553
rect 18052 3612 18104 3664
rect 20720 3612 20772 3664
rect 21824 3612 21876 3664
rect 11796 3451 11848 3460
rect 11796 3417 11830 3451
rect 11830 3417 11848 3451
rect 11796 3408 11848 3417
rect 13820 3408 13872 3460
rect 9956 3340 10008 3392
rect 11520 3340 11572 3392
rect 12348 3340 12400 3392
rect 13268 3340 13320 3392
rect 14464 3408 14516 3460
rect 16028 3451 16080 3460
rect 16028 3417 16037 3451
rect 16037 3417 16071 3451
rect 16071 3417 16080 3451
rect 16028 3408 16080 3417
rect 17316 3519 17368 3528
rect 17316 3485 17325 3519
rect 17325 3485 17359 3519
rect 17359 3485 17368 3519
rect 17316 3476 17368 3485
rect 18420 3587 18472 3596
rect 18420 3553 18429 3587
rect 18429 3553 18463 3587
rect 18463 3553 18472 3587
rect 18420 3544 18472 3553
rect 18052 3476 18104 3528
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 19524 3451 19576 3460
rect 19524 3417 19558 3451
rect 19558 3417 19576 3451
rect 19524 3408 19576 3417
rect 19708 3408 19760 3460
rect 21272 3408 21324 3460
rect 22468 3689 22477 3723
rect 22477 3689 22511 3723
rect 22511 3689 22520 3723
rect 22468 3680 22520 3689
rect 23204 3723 23256 3732
rect 23204 3689 23213 3723
rect 23213 3689 23247 3723
rect 23247 3689 23256 3723
rect 23204 3680 23256 3689
rect 26792 3680 26844 3732
rect 27344 3680 27396 3732
rect 25872 3544 25924 3596
rect 21548 3519 21600 3528
rect 21548 3485 21557 3519
rect 21557 3485 21591 3519
rect 21591 3485 21600 3519
rect 21548 3476 21600 3485
rect 22008 3519 22060 3528
rect 22008 3485 22017 3519
rect 22017 3485 22051 3519
rect 22051 3485 22060 3519
rect 22008 3476 22060 3485
rect 23572 3476 23624 3528
rect 23848 3476 23900 3528
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 16948 3383 17000 3392
rect 16948 3349 16957 3383
rect 16957 3349 16991 3383
rect 16991 3349 17000 3383
rect 16948 3340 17000 3349
rect 18880 3383 18932 3392
rect 18880 3349 18889 3383
rect 18889 3349 18923 3383
rect 18923 3349 18932 3383
rect 18880 3340 18932 3349
rect 22008 3340 22060 3392
rect 23756 3408 23808 3460
rect 23664 3383 23716 3392
rect 23664 3349 23673 3383
rect 23673 3349 23707 3383
rect 23707 3349 23716 3383
rect 23664 3340 23716 3349
rect 10395 3238 10447 3290
rect 10459 3238 10511 3290
rect 10523 3238 10575 3290
rect 10587 3238 10639 3290
rect 10651 3238 10703 3290
rect 19840 3238 19892 3290
rect 19904 3238 19956 3290
rect 19968 3238 20020 3290
rect 20032 3238 20084 3290
rect 20096 3238 20148 3290
rect 11060 3136 11112 3188
rect 11796 3136 11848 3188
rect 12164 3136 12216 3188
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 11520 3068 11572 3120
rect 9588 3043 9640 3052
rect 9588 3009 9622 3043
rect 9622 3009 9640 3043
rect 9588 3000 9640 3009
rect 10140 3000 10192 3052
rect 2964 2975 3016 2984
rect 2964 2941 2973 2975
rect 2973 2941 3007 2975
rect 3007 2941 3016 2975
rect 2964 2932 3016 2941
rect 7840 2975 7892 2984
rect 7840 2941 7849 2975
rect 7849 2941 7883 2975
rect 7883 2941 7892 2975
rect 7840 2932 7892 2941
rect 13268 3136 13320 3188
rect 15292 3136 15344 3188
rect 12348 3000 12400 3052
rect 12716 3043 12768 3052
rect 12716 3009 12725 3043
rect 12725 3009 12759 3043
rect 12759 3009 12768 3043
rect 12716 3000 12768 3009
rect 13636 3000 13688 3052
rect 15568 3111 15620 3120
rect 15568 3077 15577 3111
rect 15577 3077 15611 3111
rect 15611 3077 15620 3111
rect 15568 3068 15620 3077
rect 15752 3111 15804 3120
rect 15752 3077 15761 3111
rect 15761 3077 15795 3111
rect 15795 3077 15804 3111
rect 15752 3068 15804 3077
rect 16028 3136 16080 3188
rect 17132 3136 17184 3188
rect 17408 3136 17460 3188
rect 21272 3179 21324 3188
rect 21272 3145 21281 3179
rect 21281 3145 21315 3179
rect 21315 3145 21324 3179
rect 21272 3136 21324 3145
rect 23572 3179 23624 3188
rect 23572 3145 23581 3179
rect 23581 3145 23615 3179
rect 23615 3145 23624 3179
rect 23572 3136 23624 3145
rect 23940 3136 23992 3188
rect 16948 3111 17000 3120
rect 16948 3077 16982 3111
rect 16982 3077 17000 3111
rect 16948 3068 17000 3077
rect 18880 3068 18932 3120
rect 13820 3000 13872 3052
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 19708 3043 19760 3052
rect 14924 2932 14976 2984
rect 18052 2907 18104 2916
rect 18052 2873 18061 2907
rect 18061 2873 18095 2907
rect 18095 2873 18104 2907
rect 18052 2864 18104 2873
rect 10048 2796 10100 2848
rect 15476 2796 15528 2848
rect 18328 2796 18380 2848
rect 19708 3009 19717 3043
rect 19717 3009 19751 3043
rect 19751 3009 19760 3043
rect 19708 3000 19760 3009
rect 20996 3000 21048 3052
rect 22192 3043 22244 3052
rect 22192 3009 22226 3043
rect 22226 3009 22244 3043
rect 22192 3000 22244 3009
rect 23572 3000 23624 3052
rect 24952 3068 25004 3120
rect 24124 3043 24176 3052
rect 24124 3009 24158 3043
rect 24158 3009 24176 3043
rect 24124 3000 24176 3009
rect 25780 3043 25832 3052
rect 25780 3009 25789 3043
rect 25789 3009 25823 3043
rect 25823 3009 25832 3043
rect 25780 3000 25832 3009
rect 26056 3000 26108 3052
rect 26792 3043 26844 3052
rect 26792 3009 26801 3043
rect 26801 3009 26835 3043
rect 26835 3009 26844 3043
rect 26792 3000 26844 3009
rect 25872 2932 25924 2984
rect 26148 2932 26200 2984
rect 23848 2864 23900 2916
rect 26332 2864 26384 2916
rect 25228 2839 25280 2848
rect 25228 2805 25237 2839
rect 25237 2805 25271 2839
rect 25271 2805 25280 2839
rect 25228 2796 25280 2805
rect 5672 2694 5724 2746
rect 5736 2694 5788 2746
rect 5800 2694 5852 2746
rect 5864 2694 5916 2746
rect 5928 2694 5980 2746
rect 15118 2694 15170 2746
rect 15182 2694 15234 2746
rect 15246 2694 15298 2746
rect 15310 2694 15362 2746
rect 15374 2694 15426 2746
rect 24563 2694 24615 2746
rect 24627 2694 24679 2746
rect 24691 2694 24743 2746
rect 24755 2694 24807 2746
rect 24819 2694 24871 2746
rect 3056 2592 3108 2644
rect 9404 2592 9456 2644
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 12716 2592 12768 2644
rect 13360 2635 13412 2644
rect 13360 2601 13369 2635
rect 13369 2601 13403 2635
rect 13403 2601 13412 2635
rect 13360 2592 13412 2601
rect 14280 2592 14332 2644
rect 17316 2592 17368 2644
rect 25780 2592 25832 2644
rect 26516 2592 26568 2644
rect 10048 2499 10100 2508
rect 10048 2465 10057 2499
rect 10057 2465 10091 2499
rect 10091 2465 10100 2499
rect 10048 2456 10100 2465
rect 10140 2499 10192 2508
rect 10140 2465 10149 2499
rect 10149 2465 10183 2499
rect 10183 2465 10192 2499
rect 10140 2456 10192 2465
rect 23480 2524 23532 2576
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 12072 2388 12124 2440
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 14464 2388 14516 2397
rect 17408 2388 17460 2440
rect 21824 2431 21876 2440
rect 21824 2397 21833 2431
rect 21833 2397 21867 2431
rect 21867 2397 21876 2431
rect 21824 2388 21876 2397
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 23848 2456 23900 2508
rect 23756 2431 23808 2440
rect 23756 2397 23765 2431
rect 23765 2397 23799 2431
rect 23799 2397 23808 2431
rect 23756 2388 23808 2397
rect 23572 2320 23624 2372
rect 25228 2524 25280 2576
rect 26056 2524 26108 2576
rect 26148 2320 26200 2372
rect 23664 2252 23716 2304
rect 10395 2150 10447 2202
rect 10459 2150 10511 2202
rect 10523 2150 10575 2202
rect 10587 2150 10639 2202
rect 10651 2150 10703 2202
rect 19840 2150 19892 2202
rect 19904 2150 19956 2202
rect 19968 2150 20020 2202
rect 20032 2150 20084 2202
rect 20096 2150 20148 2202
rect 3332 1300 3384 1352
rect 6552 1300 6604 1352
rect 8576 1300 8628 1352
rect 26240 1300 26292 1352
<< metal2 >>
rect 32 31878 612 31906
rect 662 31889 718 32689
rect 32 17882 60 31878
rect 584 31770 612 31878
rect 676 31770 704 31889
rect 584 31742 704 31770
rect 1596 31878 1900 31906
rect 1950 31889 2006 32689
rect 3238 31889 3294 32689
rect 3974 32056 4030 32065
rect 3974 31991 4030 32000
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1412 24274 1440 25842
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1400 20800 1452 20806
rect 1400 20742 1452 20748
rect 1412 20262 1440 20742
rect 1400 20256 1452 20262
rect 1400 20198 1452 20204
rect 20 17876 72 17882
rect 20 17818 72 17824
rect 1308 16992 1360 16998
rect 1308 16934 1360 16940
rect 1320 3534 1348 16934
rect 1412 16574 1440 20198
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17610 1532 18022
rect 1492 17604 1544 17610
rect 1492 17546 1544 17552
rect 1412 16546 1532 16574
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 13870 1440 14894
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 12306 1440 13806
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1412 10674 1440 11018
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 7886 1440 9454
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 6338 1440 7822
rect 1504 6914 1532 16546
rect 1596 15638 1624 31878
rect 1872 31770 1900 31878
rect 1964 31770 1992 31889
rect 1872 31742 1992 31770
rect 3252 29714 3280 31889
rect 3988 30394 4016 31991
rect 4618 31889 4674 32689
rect 5906 31889 5962 32689
rect 4066 30696 4122 30705
rect 4066 30631 4122 30640
rect 4080 30598 4108 30631
rect 4068 30592 4120 30598
rect 4068 30534 4120 30540
rect 3976 30388 4028 30394
rect 3976 30330 4028 30336
rect 4068 29844 4120 29850
rect 4068 29786 4120 29792
rect 3240 29708 3292 29714
rect 3240 29650 3292 29656
rect 4080 29345 4108 29786
rect 4632 29714 4660 31889
rect 5920 31770 5948 31889
rect 6012 31878 6224 31906
rect 7286 31889 7342 32689
rect 8574 31889 8630 32689
rect 6012 31770 6040 31878
rect 5920 31742 6040 31770
rect 5672 29948 5980 29968
rect 5672 29946 5678 29948
rect 5734 29946 5758 29948
rect 5814 29946 5838 29948
rect 5894 29946 5918 29948
rect 5974 29946 5980 29948
rect 5734 29894 5736 29946
rect 5916 29894 5918 29946
rect 5672 29892 5678 29894
rect 5734 29892 5758 29894
rect 5814 29892 5838 29894
rect 5894 29892 5918 29894
rect 5974 29892 5980 29894
rect 5672 29872 5980 29892
rect 4620 29708 4672 29714
rect 4620 29650 4672 29656
rect 5172 29640 5224 29646
rect 5172 29582 5224 29588
rect 4066 29336 4122 29345
rect 4066 29271 4122 29280
rect 5184 29238 5212 29582
rect 5632 29572 5684 29578
rect 5632 29514 5684 29520
rect 5644 29306 5672 29514
rect 5632 29300 5684 29306
rect 5632 29242 5684 29248
rect 5172 29232 5224 29238
rect 5172 29174 5224 29180
rect 3976 29164 4028 29170
rect 3976 29106 4028 29112
rect 3988 28762 4016 29106
rect 4160 28960 4212 28966
rect 4160 28902 4212 28908
rect 3976 28756 4028 28762
rect 3976 28698 4028 28704
rect 4172 28558 4200 28902
rect 4344 28756 4396 28762
rect 4344 28698 4396 28704
rect 4160 28552 4212 28558
rect 4160 28494 4212 28500
rect 4252 28552 4304 28558
rect 4252 28494 4304 28500
rect 4264 28098 4292 28494
rect 4172 28070 4292 28098
rect 4066 27976 4122 27985
rect 4066 27911 4122 27920
rect 4080 27674 4108 27911
rect 4068 27668 4120 27674
rect 4068 27610 4120 27616
rect 4172 27470 4200 28070
rect 4252 28008 4304 28014
rect 4252 27950 4304 27956
rect 4264 27538 4292 27950
rect 4356 27606 4384 28698
rect 5184 28626 5212 29174
rect 5908 29164 5960 29170
rect 5960 29124 6040 29152
rect 5908 29106 5960 29112
rect 5672 28860 5980 28880
rect 5672 28858 5678 28860
rect 5734 28858 5758 28860
rect 5814 28858 5838 28860
rect 5894 28858 5918 28860
rect 5974 28858 5980 28860
rect 5734 28806 5736 28858
rect 5916 28806 5918 28858
rect 5672 28804 5678 28806
rect 5734 28804 5758 28806
rect 5814 28804 5838 28806
rect 5894 28804 5918 28806
rect 5974 28804 5980 28806
rect 5672 28784 5980 28804
rect 5172 28620 5224 28626
rect 5172 28562 5224 28568
rect 4528 28552 4580 28558
rect 4528 28494 4580 28500
rect 4540 28218 4568 28494
rect 4528 28212 4580 28218
rect 4528 28154 4580 28160
rect 4344 27600 4396 27606
rect 4344 27542 4396 27548
rect 4252 27532 4304 27538
rect 4252 27474 4304 27480
rect 4160 27464 4212 27470
rect 4160 27406 4212 27412
rect 3884 27328 3936 27334
rect 3884 27270 3936 27276
rect 3896 27062 3924 27270
rect 3884 27056 3936 27062
rect 3884 26998 3936 27004
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 2688 26920 2740 26926
rect 2688 26862 2740 26868
rect 2700 25974 2728 26862
rect 3344 26382 3372 26930
rect 4068 26852 4120 26858
rect 4068 26794 4120 26800
rect 4080 26625 4108 26794
rect 4066 26616 4122 26625
rect 4172 26586 4200 27406
rect 4264 27130 4292 27474
rect 4252 27124 4304 27130
rect 4252 27066 4304 27072
rect 4356 26790 4384 27542
rect 4436 27464 4488 27470
rect 4436 27406 4488 27412
rect 4448 27130 4476 27406
rect 4436 27124 4488 27130
rect 4436 27066 4488 27072
rect 4988 26988 5040 26994
rect 4988 26930 5040 26936
rect 4344 26784 4396 26790
rect 4344 26726 4396 26732
rect 4066 26551 4122 26560
rect 4160 26580 4212 26586
rect 4160 26522 4212 26528
rect 2780 26376 2832 26382
rect 2780 26318 2832 26324
rect 3332 26376 3384 26382
rect 3332 26318 3384 26324
rect 2688 25968 2740 25974
rect 2688 25910 2740 25916
rect 2596 25900 2648 25906
rect 2596 25842 2648 25848
rect 2608 25498 2636 25842
rect 2792 25702 2820 26318
rect 3056 26240 3108 26246
rect 3056 26182 3108 26188
rect 2780 25696 2832 25702
rect 2780 25638 2832 25644
rect 2596 25492 2648 25498
rect 2596 25434 2648 25440
rect 2792 25294 2820 25638
rect 3068 25498 3096 26182
rect 3056 25492 3108 25498
rect 3056 25434 3108 25440
rect 2780 25288 2832 25294
rect 2780 25230 2832 25236
rect 2792 24886 2820 25230
rect 2780 24880 2832 24886
rect 2780 24822 2832 24828
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 1952 24132 2004 24138
rect 1952 24074 2004 24080
rect 1964 23798 1992 24074
rect 2608 23866 2636 24550
rect 2596 23860 2648 23866
rect 2596 23802 2648 23808
rect 1952 23792 2004 23798
rect 1952 23734 2004 23740
rect 2792 23730 2820 24822
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 2884 24410 2912 24754
rect 3240 24744 3292 24750
rect 3240 24686 3292 24692
rect 2872 24404 2924 24410
rect 2872 24346 2924 24352
rect 2884 23798 2912 24346
rect 3056 24268 3108 24274
rect 3056 24210 3108 24216
rect 2872 23792 2924 23798
rect 2872 23734 2924 23740
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 3068 23662 3096 24210
rect 3252 24206 3280 24686
rect 3344 24290 3372 26318
rect 3884 25900 3936 25906
rect 3884 25842 3936 25848
rect 3896 25498 3924 25842
rect 3976 25696 4028 25702
rect 3976 25638 4028 25644
rect 3884 25492 3936 25498
rect 3884 25434 3936 25440
rect 3988 25158 4016 25638
rect 4172 25362 4200 26522
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4908 25906 4936 26318
rect 4896 25900 4948 25906
rect 4896 25842 4948 25848
rect 4160 25356 4212 25362
rect 4160 25298 4212 25304
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4436 25288 4488 25294
rect 4436 25230 4488 25236
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3344 24262 3464 24290
rect 3436 24206 3464 24262
rect 3240 24200 3292 24206
rect 3240 24142 3292 24148
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3148 24132 3200 24138
rect 3148 24074 3200 24080
rect 3160 23798 3188 24074
rect 3252 23866 3280 24142
rect 3332 24064 3384 24070
rect 3332 24006 3384 24012
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3148 23792 3200 23798
rect 3148 23734 3200 23740
rect 3056 23656 3108 23662
rect 3056 23598 3108 23604
rect 2780 23588 2832 23594
rect 2780 23530 2832 23536
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1688 22642 1716 22918
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 2792 22030 2820 23530
rect 3160 22794 3188 23734
rect 3344 23118 3372 24006
rect 3332 23112 3384 23118
rect 3332 23054 3384 23060
rect 3240 23044 3292 23050
rect 3240 22986 3292 22992
rect 3068 22778 3188 22794
rect 3056 22772 3188 22778
rect 3108 22766 3188 22772
rect 3056 22714 3108 22720
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 2884 22166 2912 22646
rect 3056 22432 3108 22438
rect 3056 22374 3108 22380
rect 2872 22160 2924 22166
rect 2872 22102 2924 22108
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 1860 20868 1912 20874
rect 1860 20810 1912 20816
rect 1872 20534 1900 20810
rect 2412 20596 2464 20602
rect 2792 20584 2820 21966
rect 2884 21010 2912 22102
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 2464 20556 2820 20584
rect 2412 20538 2464 20544
rect 1860 20528 1912 20534
rect 1860 20470 1912 20476
rect 2516 20058 2544 20556
rect 2976 20534 3004 20810
rect 3068 20602 3096 22374
rect 3252 22094 3280 22986
rect 3436 22574 3464 24142
rect 3608 24132 3660 24138
rect 3608 24074 3660 24080
rect 3620 23866 3648 24074
rect 3608 23860 3660 23866
rect 3608 23802 3660 23808
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3804 23118 3832 23666
rect 3884 23656 3936 23662
rect 3884 23598 3936 23604
rect 3896 23118 3924 23598
rect 3988 23186 4016 25094
rect 4080 24682 4108 25230
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 4344 24608 4396 24614
rect 4344 24550 4396 24556
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4066 23896 4122 23905
rect 4066 23831 4122 23840
rect 4080 23594 4108 23831
rect 4264 23730 4292 24210
rect 4356 24206 4384 24550
rect 4344 24200 4396 24206
rect 4344 24142 4396 24148
rect 4356 23866 4384 24142
rect 4344 23860 4396 23866
rect 4344 23802 4396 23808
rect 4252 23724 4304 23730
rect 4252 23666 4304 23672
rect 4068 23588 4120 23594
rect 4068 23530 4120 23536
rect 3976 23180 4028 23186
rect 3976 23122 4028 23128
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 3884 23112 3936 23118
rect 3884 23054 3936 23060
rect 3804 22642 3832 23054
rect 3792 22636 3844 22642
rect 3792 22578 3844 22584
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3436 22234 3464 22510
rect 3896 22438 3924 23054
rect 3988 22642 4016 23122
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4344 22976 4396 22982
rect 4344 22918 4396 22924
rect 4172 22642 4200 22918
rect 4356 22778 4384 22918
rect 4448 22778 4476 25230
rect 4908 24818 4936 25842
rect 5000 25430 5028 26930
rect 5184 26450 5212 28562
rect 6012 28422 6040 29124
rect 6092 29028 6144 29034
rect 6092 28970 6144 28976
rect 6104 28762 6132 28970
rect 6092 28756 6144 28762
rect 6092 28698 6144 28704
rect 6000 28416 6052 28422
rect 6000 28358 6052 28364
rect 5672 27772 5980 27792
rect 5672 27770 5678 27772
rect 5734 27770 5758 27772
rect 5814 27770 5838 27772
rect 5894 27770 5918 27772
rect 5974 27770 5980 27772
rect 5734 27718 5736 27770
rect 5916 27718 5918 27770
rect 5672 27716 5678 27718
rect 5734 27716 5758 27718
rect 5814 27716 5838 27718
rect 5894 27716 5918 27718
rect 5974 27716 5980 27718
rect 5672 27696 5980 27716
rect 6012 26994 6040 28358
rect 6000 26988 6052 26994
rect 6000 26930 6052 26936
rect 5540 26784 5592 26790
rect 5540 26726 5592 26732
rect 5172 26444 5224 26450
rect 5172 26386 5224 26392
rect 5184 26042 5212 26386
rect 5552 26382 5580 26726
rect 5672 26684 5980 26704
rect 5672 26682 5678 26684
rect 5734 26682 5758 26684
rect 5814 26682 5838 26684
rect 5894 26682 5918 26684
rect 5974 26682 5980 26684
rect 5734 26630 5736 26682
rect 5916 26630 5918 26682
rect 5672 26628 5678 26630
rect 5734 26628 5758 26630
rect 5814 26628 5838 26630
rect 5894 26628 5918 26630
rect 5974 26628 5980 26630
rect 5672 26608 5980 26628
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 6012 26042 6040 26930
rect 6092 26784 6144 26790
rect 6092 26726 6144 26732
rect 5172 26036 5224 26042
rect 5172 25978 5224 25984
rect 6000 26036 6052 26042
rect 6000 25978 6052 25984
rect 4988 25424 5040 25430
rect 4988 25366 5040 25372
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4724 24410 4752 24754
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 4908 24206 4936 24754
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 4344 22772 4396 22778
rect 4344 22714 4396 22720
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4252 22704 4304 22710
rect 4252 22646 4304 22652
rect 3976 22636 4028 22642
rect 3976 22578 4028 22584
rect 4160 22636 4212 22642
rect 4160 22578 4212 22584
rect 4264 22438 4292 22646
rect 4436 22500 4488 22506
rect 4436 22442 4488 22448
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 3160 22066 3280 22094
rect 3056 20596 3108 20602
rect 3056 20538 3108 20544
rect 2964 20528 3016 20534
rect 2964 20470 3016 20476
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2884 20058 2912 20402
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2424 18834 2452 19110
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2516 18766 2544 19994
rect 3068 19718 3096 20334
rect 3160 19825 3188 22066
rect 3884 22024 3936 22030
rect 3884 21966 3936 21972
rect 4160 22024 4212 22030
rect 4160 21966 4212 21972
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3344 20942 3372 21490
rect 3620 21146 3648 21490
rect 3896 21350 3924 21966
rect 4172 21706 4200 21966
rect 4264 21894 4292 22374
rect 4448 22030 4476 22442
rect 4724 22030 4752 23054
rect 4816 22982 4844 23666
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4436 22024 4488 22030
rect 4436 21966 4488 21972
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 3988 21678 4200 21706
rect 3988 21622 4016 21678
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4172 21418 4200 21490
rect 4160 21412 4212 21418
rect 4160 21354 4212 21360
rect 3884 21344 3936 21350
rect 3884 21286 3936 21292
rect 3608 21140 3660 21146
rect 3608 21082 3660 21088
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 3240 20868 3292 20874
rect 3240 20810 3292 20816
rect 3252 20398 3280 20810
rect 3344 20534 3372 20878
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3332 20528 3384 20534
rect 3332 20470 3384 20476
rect 3528 20398 3556 20742
rect 3896 20482 3924 21286
rect 4066 21176 4122 21185
rect 4066 21111 4122 21120
rect 4080 21078 4108 21111
rect 4068 21072 4120 21078
rect 4068 21014 4120 21020
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3988 20602 4016 20878
rect 4172 20806 4200 21354
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3608 20460 3660 20466
rect 3896 20454 4016 20482
rect 4172 20466 4200 20742
rect 4264 20534 4292 21830
rect 4356 20942 4384 21830
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 3608 20402 3660 20408
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 3146 19816 3202 19825
rect 3146 19751 3202 19760
rect 3240 19780 3292 19786
rect 3240 19722 3292 19728
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 3068 19310 3096 19654
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2608 18834 2636 19246
rect 2596 18828 2648 18834
rect 2596 18770 2648 18776
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1872 18426 1900 18634
rect 2608 18426 2636 18770
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2700 18426 2728 18566
rect 1860 18420 1912 18426
rect 1860 18362 1912 18368
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2240 17338 2268 18362
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2516 18086 2544 18158
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2240 16182 2268 17274
rect 2516 16522 2544 18022
rect 2504 16516 2556 16522
rect 2504 16458 2556 16464
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1584 15632 1636 15638
rect 1584 15574 1636 15580
rect 1780 15094 1808 15846
rect 2148 15706 2176 16050
rect 2516 16046 2544 16458
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2332 15502 2360 15846
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 1768 15088 1820 15094
rect 1768 15030 1820 15036
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2516 14074 2544 14350
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13394 2360 13670
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2608 13190 2636 13874
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2608 12442 2636 13126
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 1964 11898 1992 12106
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 2700 11354 2728 18362
rect 3252 18154 3280 19722
rect 3528 18154 3556 20334
rect 3620 19514 3648 20402
rect 3988 19854 4016 20454
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4356 20346 4384 20878
rect 4264 20318 4384 20346
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3608 19508 3660 19514
rect 3608 19450 3660 19456
rect 3698 18456 3754 18465
rect 3698 18391 3754 18400
rect 3240 18148 3292 18154
rect 3240 18090 3292 18096
rect 3516 18148 3568 18154
rect 3516 18090 3568 18096
rect 2780 17536 2832 17542
rect 2780 17478 2832 17484
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 2792 17338 2820 17478
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2792 16590 2820 17274
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2792 13530 2820 15438
rect 2884 13938 2912 16662
rect 2976 16658 3004 17002
rect 3068 16794 3096 17478
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 3160 16726 3188 17138
rect 3528 17105 3556 17478
rect 3712 17105 3740 18391
rect 3792 17604 3844 17610
rect 3792 17546 3844 17552
rect 3514 17096 3570 17105
rect 3514 17031 3570 17040
rect 3698 17096 3754 17105
rect 3698 17031 3754 17040
rect 3804 16998 3832 17546
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 3988 16182 4016 19790
rect 4264 19446 4292 20318
rect 4344 20256 4396 20262
rect 4344 20198 4396 20204
rect 4356 19990 4384 20198
rect 4344 19984 4396 19990
rect 4344 19926 4396 19932
rect 4356 19514 4384 19926
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4252 19440 4304 19446
rect 4252 19382 4304 19388
rect 4264 18408 4292 19382
rect 4448 19378 4476 21966
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 4632 19922 4660 20878
rect 4724 20398 4752 21966
rect 4908 21690 4936 24142
rect 5000 23730 5028 25366
rect 5184 25362 5212 25978
rect 6104 25770 6132 26726
rect 6092 25764 6144 25770
rect 6092 25706 6144 25712
rect 5672 25596 5980 25616
rect 5672 25594 5678 25596
rect 5734 25594 5758 25596
rect 5814 25594 5838 25596
rect 5894 25594 5918 25596
rect 5974 25594 5980 25596
rect 5734 25542 5736 25594
rect 5916 25542 5918 25594
rect 5672 25540 5678 25542
rect 5734 25540 5758 25542
rect 5814 25540 5838 25542
rect 5894 25540 5918 25542
rect 5974 25540 5980 25542
rect 5672 25520 5980 25540
rect 5172 25356 5224 25362
rect 5172 25298 5224 25304
rect 5184 24750 5212 25298
rect 5172 24744 5224 24750
rect 5172 24686 5224 24692
rect 5184 24206 5212 24686
rect 6104 24682 6132 25706
rect 6092 24676 6144 24682
rect 6092 24618 6144 24624
rect 5672 24508 5980 24528
rect 5672 24506 5678 24508
rect 5734 24506 5758 24508
rect 5814 24506 5838 24508
rect 5894 24506 5918 24508
rect 5974 24506 5980 24508
rect 5734 24454 5736 24506
rect 5916 24454 5918 24506
rect 5672 24452 5678 24454
rect 5734 24452 5758 24454
rect 5814 24452 5838 24454
rect 5894 24452 5918 24454
rect 5974 24452 5980 24454
rect 5672 24432 5980 24452
rect 5172 24200 5224 24206
rect 5172 24142 5224 24148
rect 5540 24132 5592 24138
rect 5540 24074 5592 24080
rect 5552 23866 5580 24074
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 4988 23724 5040 23730
rect 4988 23666 5040 23672
rect 5000 23526 5028 23666
rect 6104 23526 6132 24618
rect 4988 23520 5040 23526
rect 4988 23462 5040 23468
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 6092 23520 6144 23526
rect 6092 23462 6144 23468
rect 5552 23050 5580 23462
rect 5672 23420 5980 23440
rect 5672 23418 5678 23420
rect 5734 23418 5758 23420
rect 5814 23418 5838 23420
rect 5894 23418 5918 23420
rect 5974 23418 5980 23420
rect 5734 23366 5736 23418
rect 5916 23366 5918 23418
rect 5672 23364 5678 23366
rect 5734 23364 5758 23366
rect 5814 23364 5838 23366
rect 5894 23364 5918 23366
rect 5974 23364 5980 23366
rect 5672 23344 5980 23364
rect 5540 23044 5592 23050
rect 5540 22986 5592 22992
rect 5672 22332 5980 22352
rect 5672 22330 5678 22332
rect 5734 22330 5758 22332
rect 5814 22330 5838 22332
rect 5894 22330 5918 22332
rect 5974 22330 5980 22332
rect 5734 22278 5736 22330
rect 5916 22278 5918 22330
rect 5672 22276 5678 22278
rect 5734 22276 5758 22278
rect 5814 22276 5838 22278
rect 5894 22276 5918 22278
rect 5974 22276 5980 22278
rect 5672 22256 5980 22276
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 4896 21684 4948 21690
rect 4896 21626 4948 21632
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4816 20806 4844 21490
rect 5368 21146 5396 21898
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 5460 20942 5488 21354
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 5672 21244 5980 21264
rect 5672 21242 5678 21244
rect 5734 21242 5758 21244
rect 5814 21242 5838 21244
rect 5894 21242 5918 21244
rect 5974 21242 5980 21244
rect 5734 21190 5736 21242
rect 5916 21190 5918 21242
rect 5672 21188 5678 21190
rect 5734 21188 5758 21190
rect 5814 21188 5838 21190
rect 5894 21188 5918 21190
rect 5974 21188 5980 21190
rect 5672 21168 5980 21188
rect 6104 21078 6132 21286
rect 6092 21072 6144 21078
rect 6092 21014 6144 21020
rect 6104 20942 6132 21014
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 6092 20936 6144 20942
rect 6092 20878 6144 20884
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4620 19916 4672 19922
rect 4620 19858 4672 19864
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4448 18426 4476 19314
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4436 18420 4488 18426
rect 4264 18380 4384 18408
rect 4356 18290 4384 18380
rect 4436 18362 4488 18368
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4068 18216 4120 18222
rect 4120 18176 4292 18204
rect 4068 18158 4120 18164
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4172 17338 4200 18022
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4264 17134 4292 18176
rect 4540 18154 4568 19246
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4528 18148 4580 18154
rect 4528 18090 4580 18096
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4264 16454 4292 17070
rect 4448 16590 4476 17070
rect 4632 16776 4660 18226
rect 4724 17678 4752 20334
rect 5276 20058 5304 20402
rect 5672 20156 5980 20176
rect 5672 20154 5678 20156
rect 5734 20154 5758 20156
rect 5814 20154 5838 20156
rect 5894 20154 5918 20156
rect 5974 20154 5980 20156
rect 5734 20102 5736 20154
rect 5916 20102 5918 20154
rect 5672 20100 5678 20102
rect 5734 20100 5758 20102
rect 5814 20100 5838 20102
rect 5894 20100 5918 20102
rect 5974 20100 5980 20102
rect 5672 20080 5980 20100
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4908 19378 4936 19654
rect 5368 19378 5396 19722
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4540 16748 4660 16776
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 3792 16176 3844 16182
rect 3976 16176 4028 16182
rect 3844 16124 3924 16130
rect 3792 16118 3924 16124
rect 3976 16118 4028 16124
rect 3608 16108 3660 16114
rect 3804 16102 3924 16118
rect 3608 16050 3660 16056
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2976 15706 3004 15914
rect 3528 15706 3556 15982
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 2976 14890 3004 15642
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 2964 14884 3016 14890
rect 2964 14826 3016 14832
rect 3252 14414 3280 15098
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3436 14618 3464 14894
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3160 14006 3188 14350
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2792 12714 2820 13466
rect 3620 12986 3648 16050
rect 3896 15910 3924 16102
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15570 3924 15846
rect 4172 15638 4200 16050
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 11762 2820 12650
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2976 11762 3004 12582
rect 3068 12306 3096 12854
rect 3620 12434 3648 12922
rect 3896 12918 3924 15506
rect 4172 15094 4200 15574
rect 4264 15502 4292 16390
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3988 14006 4016 14758
rect 4172 14618 4200 15030
rect 4448 14958 4476 16526
rect 4540 16250 4568 16748
rect 4632 16658 4752 16674
rect 4632 16652 4764 16658
rect 4632 16646 4712 16652
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 4080 14385 4108 14486
rect 4066 14376 4122 14385
rect 4066 14311 4122 14320
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 4066 13016 4122 13025
rect 4066 12951 4068 12960
rect 4120 12951 4122 12960
rect 4068 12922 4120 12928
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3436 12406 3648 12434
rect 3436 12374 3464 12406
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 3436 11626 3464 12310
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3804 11762 3832 12038
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3988 11665 4016 12038
rect 4080 11898 4108 12786
rect 4448 12782 4476 14894
rect 4632 14890 4660 16646
rect 4712 16594 4764 16600
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4724 16250 4752 16390
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4620 14884 4672 14890
rect 4620 14826 4672 14832
rect 4632 14482 4660 14826
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4632 13394 4660 14418
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4172 11694 4200 12718
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4448 12170 4476 12582
rect 4436 12164 4488 12170
rect 4436 12106 4488 12112
rect 4632 11762 4660 13330
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4160 11688 4212 11694
rect 3974 11656 4030 11665
rect 3424 11620 3476 11626
rect 4160 11630 4212 11636
rect 3974 11591 4030 11600
rect 3424 11562 3476 11568
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 2688 11348 2740 11354
rect 2608 11308 2688 11336
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2424 10810 2452 11018
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 9654 1716 10406
rect 2332 10266 2360 10610
rect 2608 10606 2636 11308
rect 2688 11290 2740 11296
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2608 10130 2636 10542
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2792 9722 2820 9998
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2136 8288 2188 8294
rect 2136 8230 2188 8236
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1780 7546 1808 7754
rect 2148 7546 2176 8230
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1504 6886 1624 6914
rect 1412 6310 1532 6338
rect 1504 6254 1532 6310
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1504 4690 1532 6190
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1596 4622 1624 6886
rect 2240 6866 2268 8434
rect 2700 7342 2728 9590
rect 2792 9518 2820 9658
rect 2884 9654 2912 10066
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2976 9654 3004 9930
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 3252 9586 3280 10746
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3344 9586 3372 9862
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3160 8974 3188 9454
rect 3252 8974 3280 9522
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3608 8900 3660 8906
rect 3608 8842 3660 8848
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7410 3556 7686
rect 3620 7478 3648 8842
rect 3804 7546 3832 9454
rect 3896 7585 3924 11494
rect 4632 11336 4660 11698
rect 4816 11354 4844 18702
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 5276 17270 5304 17478
rect 5264 17264 5316 17270
rect 5264 17206 5316 17212
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4908 16998 4936 17138
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4908 16522 4936 16934
rect 5276 16590 5304 17206
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4908 16114 4936 16458
rect 5276 16114 5304 16526
rect 5368 16250 5396 19314
rect 5552 19174 5580 19314
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5552 18698 5580 19110
rect 5672 19068 5980 19088
rect 5672 19066 5678 19068
rect 5734 19066 5758 19068
rect 5814 19066 5838 19068
rect 5894 19066 5918 19068
rect 5974 19066 5980 19068
rect 5734 19014 5736 19066
rect 5916 19014 5918 19066
rect 5672 19012 5678 19014
rect 5734 19012 5758 19014
rect 5814 19012 5838 19014
rect 5894 19012 5918 19014
rect 5974 19012 5980 19014
rect 5672 18992 5980 19012
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 5672 17980 5980 18000
rect 5672 17978 5678 17980
rect 5734 17978 5758 17980
rect 5814 17978 5838 17980
rect 5894 17978 5918 17980
rect 5974 17978 5980 17980
rect 5734 17926 5736 17978
rect 5916 17926 5918 17978
rect 5672 17924 5678 17926
rect 5734 17924 5758 17926
rect 5814 17924 5838 17926
rect 5894 17924 5918 17926
rect 5974 17924 5980 17926
rect 5672 17904 5980 17924
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5448 16040 5500 16046
rect 5552 16028 5580 17138
rect 5672 16892 5980 16912
rect 5672 16890 5678 16892
rect 5734 16890 5758 16892
rect 5814 16890 5838 16892
rect 5894 16890 5918 16892
rect 5974 16890 5980 16892
rect 5734 16838 5736 16890
rect 5916 16838 5918 16890
rect 5672 16836 5678 16838
rect 5734 16836 5758 16838
rect 5814 16836 5838 16838
rect 5894 16836 5918 16838
rect 5974 16836 5980 16838
rect 5672 16816 5980 16836
rect 6012 16590 6040 17478
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 6104 16046 6132 18022
rect 5500 16000 5580 16028
rect 5448 15982 5500 15988
rect 5354 15736 5410 15745
rect 5354 15671 5410 15680
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 5000 15026 5028 15302
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 5092 14074 5120 14282
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 5276 13870 5304 14350
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5276 12442 5304 13806
rect 5368 13530 5396 15671
rect 5552 14618 5580 16000
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 5672 15804 5980 15824
rect 5672 15802 5678 15804
rect 5734 15802 5758 15804
rect 5814 15802 5838 15804
rect 5894 15802 5918 15804
rect 5974 15802 5980 15804
rect 5734 15750 5736 15802
rect 5916 15750 5918 15802
rect 5672 15748 5678 15750
rect 5734 15748 5758 15750
rect 5814 15748 5838 15750
rect 5894 15748 5918 15750
rect 5974 15748 5980 15750
rect 5672 15728 5980 15748
rect 5672 14716 5980 14736
rect 5672 14714 5678 14716
rect 5734 14714 5758 14716
rect 5814 14714 5838 14716
rect 5894 14714 5918 14716
rect 5974 14714 5980 14716
rect 5734 14662 5736 14714
rect 5916 14662 5918 14714
rect 5672 14660 5678 14662
rect 5734 14660 5758 14662
rect 5814 14660 5838 14662
rect 5894 14660 5918 14662
rect 5974 14660 5980 14662
rect 5672 14640 5980 14660
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5552 13938 5580 14554
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5644 14074 5672 14214
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5672 13628 5980 13648
rect 5672 13626 5678 13628
rect 5734 13626 5758 13628
rect 5814 13626 5838 13628
rect 5894 13626 5918 13628
rect 5974 13626 5980 13628
rect 5734 13574 5736 13626
rect 5916 13574 5918 13626
rect 5672 13572 5678 13574
rect 5734 13572 5758 13574
rect 5814 13572 5838 13574
rect 5894 13572 5918 13574
rect 5974 13572 5980 13574
rect 5672 13552 5980 13572
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 6104 13326 6132 15982
rect 6196 14550 6224 31878
rect 7104 29708 7156 29714
rect 7104 29650 7156 29656
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6932 29238 6960 29446
rect 6920 29232 6972 29238
rect 6920 29174 6972 29180
rect 7116 29102 7144 29650
rect 7104 29096 7156 29102
rect 7104 29038 7156 29044
rect 7012 28552 7064 28558
rect 7012 28494 7064 28500
rect 7024 28218 7052 28494
rect 7012 28212 7064 28218
rect 7012 28154 7064 28160
rect 7116 28014 7144 29038
rect 7104 28008 7156 28014
rect 7104 27950 7156 27956
rect 6552 27872 6604 27878
rect 6552 27814 6604 27820
rect 6564 26994 6592 27814
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 7116 26926 7144 27950
rect 6644 26920 6696 26926
rect 6644 26862 6696 26868
rect 7104 26920 7156 26926
rect 7104 26862 7156 26868
rect 6460 26784 6512 26790
rect 6460 26726 6512 26732
rect 6472 25906 6500 26726
rect 6656 26586 6684 26862
rect 6644 26580 6696 26586
rect 6644 26522 6696 26528
rect 6460 25900 6512 25906
rect 6460 25842 6512 25848
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 6748 25498 6776 25842
rect 6920 25696 6972 25702
rect 6920 25638 6972 25644
rect 6736 25492 6788 25498
rect 6736 25434 6788 25440
rect 6932 25294 6960 25638
rect 7300 25378 7328 31889
rect 8588 31770 8616 31889
rect 8680 31878 8892 31906
rect 9954 31889 10010 32689
rect 11242 31889 11298 32689
rect 12530 31889 12586 32689
rect 13910 31889 13966 32689
rect 15198 31889 15254 32689
rect 8680 31770 8708 31878
rect 8588 31742 8708 31770
rect 7380 29504 7432 29510
rect 7380 29446 7432 29452
rect 7392 28626 7420 29446
rect 7380 28620 7432 28626
rect 7380 28562 7432 28568
rect 8576 28552 8628 28558
rect 8576 28494 8628 28500
rect 8392 28416 8444 28422
rect 8392 28358 8444 28364
rect 8404 28150 8432 28358
rect 8392 28144 8444 28150
rect 8392 28086 8444 28092
rect 8588 27606 8616 28494
rect 8576 27600 8628 27606
rect 8576 27542 8628 27548
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 8300 27464 8352 27470
rect 8300 27406 8352 27412
rect 7564 26852 7616 26858
rect 7564 26794 7616 26800
rect 7116 25350 7328 25378
rect 7576 25362 7604 26794
rect 7852 26246 7880 27406
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 8220 27062 8248 27270
rect 8208 27056 8260 27062
rect 8208 26998 8260 27004
rect 8312 26586 8340 27406
rect 8300 26580 8352 26586
rect 8300 26522 8352 26528
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 7840 26240 7892 26246
rect 7840 26182 7892 26188
rect 7748 25696 7800 25702
rect 7748 25638 7800 25644
rect 7564 25356 7616 25362
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6828 25152 6880 25158
rect 6828 25094 6880 25100
rect 6460 24064 6512 24070
rect 6460 24006 6512 24012
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6472 23798 6500 24006
rect 6748 23866 6776 24006
rect 6736 23860 6788 23866
rect 6736 23802 6788 23808
rect 6460 23792 6512 23798
rect 6460 23734 6512 23740
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6564 22094 6592 23666
rect 6840 23662 6868 25094
rect 6920 24676 6972 24682
rect 6920 24618 6972 24624
rect 6932 24274 6960 24618
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 6828 23656 6880 23662
rect 6828 23598 6880 23604
rect 6472 22066 6592 22094
rect 6472 21962 6500 22066
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6460 21956 6512 21962
rect 6460 21898 6512 21904
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6288 21622 6316 21830
rect 6932 21690 6960 21966
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 6276 21616 6328 21622
rect 6276 21558 6328 21564
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6380 20602 6408 21490
rect 6472 20602 6500 21626
rect 6736 21412 6788 21418
rect 6736 21354 6788 21360
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6748 20466 6776 21354
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 6932 20602 6960 20878
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6656 20262 6684 20402
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6656 19786 6684 20198
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6644 19780 6696 19786
rect 6644 19722 6696 19728
rect 6276 19712 6328 19718
rect 6276 19654 6328 19660
rect 6288 18630 6316 19654
rect 6380 19378 6408 19722
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 6276 18624 6328 18630
rect 6276 18566 6328 18572
rect 6380 18290 6408 19314
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6564 17202 6592 17614
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6656 16998 6684 17750
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6748 16046 6776 20402
rect 6932 19854 6960 20538
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6840 17270 6868 17614
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 7024 17490 7052 17546
rect 6932 17462 7052 17490
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6932 17134 6960 17462
rect 7116 17377 7144 25350
rect 7564 25298 7616 25304
rect 7380 25220 7432 25226
rect 7380 25162 7432 25168
rect 7472 25220 7524 25226
rect 7472 25162 7524 25168
rect 7392 24818 7420 25162
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7484 24750 7512 25162
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7300 24138 7328 24550
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 7288 24132 7340 24138
rect 7288 24074 7340 24080
rect 7208 23866 7236 24074
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 7472 23724 7524 23730
rect 7576 23712 7604 25298
rect 7760 24886 7788 25638
rect 7852 25294 7880 26182
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 7748 24880 7800 24886
rect 7748 24822 7800 24828
rect 7524 23684 7604 23712
rect 7472 23666 7524 23672
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 7932 23044 7984 23050
rect 7932 22986 7984 22992
rect 7208 22778 7236 22986
rect 7944 22778 7972 22986
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7932 22772 7984 22778
rect 7932 22714 7984 22720
rect 7748 22704 7800 22710
rect 7748 22646 7800 22652
rect 7760 21690 7788 22646
rect 7932 22432 7984 22438
rect 7932 22374 7984 22380
rect 7944 21962 7972 22374
rect 7932 21956 7984 21962
rect 7932 21898 7984 21904
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7484 20534 7512 20742
rect 7472 20528 7524 20534
rect 7472 20470 7524 20476
rect 7472 20392 7524 20398
rect 7472 20334 7524 20340
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7102 17368 7158 17377
rect 7012 17332 7064 17338
rect 7208 17338 7236 17818
rect 7102 17303 7158 17312
rect 7196 17332 7248 17338
rect 7012 17274 7064 17280
rect 7196 17274 7248 17280
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6564 15706 6592 15846
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6184 14544 6236 14550
rect 6184 14486 6236 14492
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 5448 13320 5500 13326
rect 6092 13320 6144 13326
rect 5500 13280 5580 13308
rect 5448 13262 5500 13268
rect 5552 12918 5580 13280
rect 6092 13262 6144 13268
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5276 12238 5304 12378
rect 5552 12306 5580 12854
rect 5672 12540 5980 12560
rect 5672 12538 5678 12540
rect 5734 12538 5758 12540
rect 5814 12538 5838 12540
rect 5894 12538 5918 12540
rect 5974 12538 5980 12540
rect 5734 12486 5736 12538
rect 5916 12486 5918 12538
rect 5672 12484 5678 12486
rect 5734 12484 5758 12486
rect 5814 12484 5838 12486
rect 5894 12484 5918 12486
rect 5974 12484 5980 12486
rect 5672 12464 5980 12484
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 6196 12238 6224 12378
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6196 12102 6224 12174
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 5000 11830 5028 12038
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 4540 11308 4660 11336
rect 4804 11348 4856 11354
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3988 10810 4016 11086
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3988 10266 4016 10610
rect 4066 10296 4122 10305
rect 3976 10260 4028 10266
rect 4066 10231 4068 10240
rect 3976 10202 4028 10208
rect 4120 10231 4122 10240
rect 4068 10202 4120 10208
rect 4264 10130 4292 10950
rect 4540 10606 4568 11308
rect 4804 11290 4856 11296
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4540 10198 4568 10542
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4172 9586 4200 9862
rect 4632 9722 4660 10610
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4172 9178 4200 9522
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4066 8936 4122 8945
rect 4066 8871 4068 8880
rect 4120 8871 4122 8880
rect 4068 8842 4120 8848
rect 4160 8288 4212 8294
rect 4080 8248 4160 8276
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3882 7576 3938 7585
rect 3792 7540 3844 7546
rect 3882 7511 3938 7520
rect 3792 7482 3844 7488
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3620 7342 3648 7414
rect 3988 7410 4016 7686
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2424 6798 2452 7210
rect 2700 7002 2728 7278
rect 4080 7206 4108 8248
rect 4160 8230 4212 8236
rect 4356 7818 4384 9318
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4252 7472 4304 7478
rect 4304 7432 4384 7460
rect 4252 7414 4304 7420
rect 4356 7206 4384 7432
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 2688 6996 2740 7002
rect 2608 6956 2688 6984
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2240 5914 2268 6258
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2608 5846 2636 6956
rect 2688 6938 2740 6944
rect 4356 6798 4384 7142
rect 4540 6934 4568 7210
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 4632 6798 4660 9454
rect 4724 9178 4752 9522
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 6322 3280 6598
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 4080 6225 4108 6326
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 3344 5710 3372 6054
rect 4172 5846 4200 6666
rect 4264 6322 4292 6666
rect 4356 6458 4384 6734
rect 4632 6458 4660 6734
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4816 6338 4844 11290
rect 5184 11150 5212 11494
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5552 10470 5580 11630
rect 5672 11452 5980 11472
rect 5672 11450 5678 11452
rect 5734 11450 5758 11452
rect 5814 11450 5838 11452
rect 5894 11450 5918 11452
rect 5974 11450 5980 11452
rect 5734 11398 5736 11450
rect 5916 11398 5918 11450
rect 5672 11396 5678 11398
rect 5734 11396 5758 11398
rect 5814 11396 5838 11398
rect 5894 11396 5918 11398
rect 5974 11396 5980 11398
rect 5672 11376 5980 11396
rect 6012 11218 6040 11834
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10810 5764 10950
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 6012 10554 6040 11154
rect 6012 10526 6132 10554
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5552 10130 5580 10406
rect 5672 10364 5980 10384
rect 5672 10362 5678 10364
rect 5734 10362 5758 10364
rect 5814 10362 5838 10364
rect 5894 10362 5918 10364
rect 5974 10362 5980 10364
rect 5734 10310 5736 10362
rect 5916 10310 5918 10362
rect 5672 10308 5678 10310
rect 5734 10308 5758 10310
rect 5814 10308 5838 10310
rect 5894 10308 5918 10310
rect 5974 10308 5980 10310
rect 5672 10288 5980 10308
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 6012 9994 6040 10406
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 5000 9518 5028 9862
rect 6104 9654 6132 10526
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6196 9466 6224 12038
rect 6288 9602 6316 13874
rect 6748 13802 6776 15438
rect 6932 15094 6960 17070
rect 7024 16726 7052 17274
rect 7208 17202 7236 17274
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 7116 16250 7144 17138
rect 7300 17082 7328 19722
rect 7484 18766 7512 20334
rect 7760 19854 7788 21626
rect 8036 21554 8064 26318
rect 8392 25152 8444 25158
rect 8392 25094 8444 25100
rect 8760 25152 8812 25158
rect 8760 25094 8812 25100
rect 8404 24954 8432 25094
rect 8392 24948 8444 24954
rect 8392 24890 8444 24896
rect 8772 24886 8800 25094
rect 8760 24880 8812 24886
rect 8760 24822 8812 24828
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8772 23730 8800 24006
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 8128 22642 8156 22918
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 8220 22098 8248 22918
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 7840 21480 7892 21486
rect 7840 21422 7892 21428
rect 7852 21350 7880 21422
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7852 21078 7880 21286
rect 7840 21072 7892 21078
rect 7840 21014 7892 21020
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 7944 20058 7972 20878
rect 8116 20800 8168 20806
rect 8116 20742 8168 20748
rect 8128 20534 8156 20742
rect 8116 20528 8168 20534
rect 8116 20470 8168 20476
rect 8116 20392 8168 20398
rect 8220 20346 8248 22034
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8772 21622 8800 21830
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 8760 21616 8812 21622
rect 8760 21558 8812 21564
rect 8168 20340 8248 20346
rect 8116 20334 8248 20340
rect 8128 20318 8248 20334
rect 8220 20058 8248 20318
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8312 19854 8340 21558
rect 8864 21026 8892 31878
rect 9312 29572 9364 29578
rect 9312 29514 9364 29520
rect 9324 29306 9352 29514
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9772 28416 9824 28422
rect 9772 28358 9824 28364
rect 9784 28150 9812 28358
rect 9772 28144 9824 28150
rect 9772 28086 9824 28092
rect 9036 28008 9088 28014
rect 9036 27950 9088 27956
rect 9312 28008 9364 28014
rect 9312 27950 9364 27956
rect 8944 27872 8996 27878
rect 8944 27814 8996 27820
rect 8956 27538 8984 27814
rect 9048 27606 9076 27950
rect 9036 27600 9088 27606
rect 9036 27542 9088 27548
rect 9324 27538 9352 27950
rect 8944 27532 8996 27538
rect 8944 27474 8996 27480
rect 9312 27532 9364 27538
rect 9312 27474 9364 27480
rect 9324 26994 9352 27474
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 9416 26994 9444 27406
rect 9312 26988 9364 26994
rect 9312 26930 9364 26936
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9220 25968 9272 25974
rect 9220 25910 9272 25916
rect 9232 24954 9260 25910
rect 9600 25838 9628 26318
rect 9404 25832 9456 25838
rect 9404 25774 9456 25780
rect 9588 25832 9640 25838
rect 9588 25774 9640 25780
rect 9416 25498 9444 25774
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 9220 24948 9272 24954
rect 9220 24890 9272 24896
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9508 24274 9536 24550
rect 9496 24268 9548 24274
rect 9496 24210 9548 24216
rect 9600 24206 9628 25774
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9784 23730 9812 24754
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9036 23044 9088 23050
rect 9036 22986 9088 22992
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8956 21690 8984 21966
rect 8944 21684 8996 21690
rect 8944 21626 8996 21632
rect 8956 21146 8984 21626
rect 9048 21146 9076 22986
rect 9784 22778 9812 23666
rect 9876 23050 9904 24006
rect 9864 23044 9916 23050
rect 9864 22986 9916 22992
rect 9876 22953 9904 22986
rect 9862 22944 9918 22953
rect 9862 22879 9918 22888
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9588 22704 9640 22710
rect 9508 22664 9588 22692
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9416 22234 9444 22578
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9312 22024 9364 22030
rect 9508 21978 9536 22664
rect 9588 22646 9640 22652
rect 9680 22500 9732 22506
rect 9680 22442 9732 22448
rect 9692 22094 9720 22442
rect 9600 22066 9720 22094
rect 9600 22030 9628 22066
rect 9364 21972 9536 21978
rect 9312 21966 9536 21972
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9324 21950 9536 21966
rect 9324 21418 9352 21950
rect 9588 21548 9640 21554
rect 9692 21536 9720 22066
rect 9770 22128 9826 22137
rect 9770 22063 9772 22072
rect 9824 22063 9826 22072
rect 9772 22034 9824 22040
rect 9876 21690 9904 22714
rect 9968 22166 9996 31889
rect 10395 30492 10703 30512
rect 10395 30490 10401 30492
rect 10457 30490 10481 30492
rect 10537 30490 10561 30492
rect 10617 30490 10641 30492
rect 10697 30490 10703 30492
rect 10457 30438 10459 30490
rect 10639 30438 10641 30490
rect 10395 30436 10401 30438
rect 10457 30436 10481 30438
rect 10537 30436 10561 30438
rect 10617 30436 10641 30438
rect 10697 30436 10703 30438
rect 10395 30416 10703 30436
rect 11152 30252 11204 30258
rect 11152 30194 11204 30200
rect 11164 29646 11192 30194
rect 11152 29640 11204 29646
rect 11152 29582 11204 29588
rect 10324 29572 10376 29578
rect 10324 29514 10376 29520
rect 10336 29306 10364 29514
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10968 29504 11020 29510
rect 10968 29446 11020 29452
rect 10395 29404 10703 29424
rect 10395 29402 10401 29404
rect 10457 29402 10481 29404
rect 10537 29402 10561 29404
rect 10617 29402 10641 29404
rect 10697 29402 10703 29404
rect 10457 29350 10459 29402
rect 10639 29350 10641 29402
rect 10395 29348 10401 29350
rect 10457 29348 10481 29350
rect 10537 29348 10561 29350
rect 10617 29348 10641 29350
rect 10697 29348 10703 29350
rect 10395 29328 10703 29348
rect 10324 29300 10376 29306
rect 10324 29242 10376 29248
rect 10796 29238 10824 29446
rect 10784 29232 10836 29238
rect 10784 29174 10836 29180
rect 10980 29170 11008 29446
rect 10968 29164 11020 29170
rect 10968 29106 11020 29112
rect 10140 29096 10192 29102
rect 10140 29038 10192 29044
rect 10876 29096 10928 29102
rect 10876 29038 10928 29044
rect 10048 28212 10100 28218
rect 10048 28154 10100 28160
rect 10060 27334 10088 28154
rect 10048 27328 10100 27334
rect 10048 27270 10100 27276
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 10060 26353 10088 26726
rect 10046 26344 10102 26353
rect 10046 26279 10102 26288
rect 10152 26042 10180 29038
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10244 27674 10272 28494
rect 10395 28316 10703 28336
rect 10395 28314 10401 28316
rect 10457 28314 10481 28316
rect 10537 28314 10561 28316
rect 10617 28314 10641 28316
rect 10697 28314 10703 28316
rect 10457 28262 10459 28314
rect 10639 28262 10641 28314
rect 10395 28260 10401 28262
rect 10457 28260 10481 28262
rect 10537 28260 10561 28262
rect 10617 28260 10641 28262
rect 10697 28260 10703 28262
rect 10395 28240 10703 28260
rect 10232 27668 10284 27674
rect 10232 27610 10284 27616
rect 10784 27532 10836 27538
rect 10784 27474 10836 27480
rect 10395 27228 10703 27248
rect 10395 27226 10401 27228
rect 10457 27226 10481 27228
rect 10537 27226 10561 27228
rect 10617 27226 10641 27228
rect 10697 27226 10703 27228
rect 10457 27174 10459 27226
rect 10639 27174 10641 27226
rect 10395 27172 10401 27174
rect 10457 27172 10481 27174
rect 10537 27172 10561 27174
rect 10617 27172 10641 27174
rect 10697 27172 10703 27174
rect 10395 27152 10703 27172
rect 10324 26988 10376 26994
rect 10324 26930 10376 26936
rect 10336 26586 10364 26930
rect 10796 26586 10824 27474
rect 10888 27402 10916 29038
rect 11164 28626 11192 29582
rect 11256 28626 11284 31889
rect 12256 30048 12308 30054
rect 12256 29990 12308 29996
rect 12268 29578 12296 29990
rect 12544 29714 12572 31889
rect 12532 29708 12584 29714
rect 12532 29650 12584 29656
rect 12256 29572 12308 29578
rect 12256 29514 12308 29520
rect 11612 29504 11664 29510
rect 11612 29446 11664 29452
rect 11624 29170 11652 29446
rect 12544 29306 12572 29650
rect 13636 29640 13688 29646
rect 13636 29582 13688 29588
rect 12992 29572 13044 29578
rect 12992 29514 13044 29520
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 13004 29238 13032 29514
rect 12992 29232 13044 29238
rect 12992 29174 13044 29180
rect 11612 29164 11664 29170
rect 11612 29106 11664 29112
rect 12532 29164 12584 29170
rect 12532 29106 12584 29112
rect 12900 29164 12952 29170
rect 12900 29106 12952 29112
rect 13268 29164 13320 29170
rect 13268 29106 13320 29112
rect 12164 29096 12216 29102
rect 12164 29038 12216 29044
rect 11152 28620 11204 28626
rect 11152 28562 11204 28568
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 11980 28620 12032 28626
rect 11980 28562 12032 28568
rect 11164 28506 11192 28562
rect 11164 28478 11284 28506
rect 11152 28416 11204 28422
rect 11152 28358 11204 28364
rect 11164 28150 11192 28358
rect 11152 28144 11204 28150
rect 11152 28086 11204 28092
rect 11256 27538 11284 28478
rect 11336 27600 11388 27606
rect 11336 27542 11388 27548
rect 11244 27532 11296 27538
rect 11244 27474 11296 27480
rect 10876 27396 10928 27402
rect 10876 27338 10928 27344
rect 10888 26994 10916 27338
rect 11256 27130 11284 27474
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 10968 27056 11020 27062
rect 10968 26998 11020 27004
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10980 26586 11008 26998
rect 11060 26988 11112 26994
rect 11060 26930 11112 26936
rect 10324 26580 10376 26586
rect 10324 26522 10376 26528
rect 10784 26580 10836 26586
rect 10784 26522 10836 26528
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 11072 26450 11100 26930
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 10968 26308 11020 26314
rect 10968 26250 11020 26256
rect 10395 26140 10703 26160
rect 10395 26138 10401 26140
rect 10457 26138 10481 26140
rect 10537 26138 10561 26140
rect 10617 26138 10641 26140
rect 10697 26138 10703 26140
rect 10457 26086 10459 26138
rect 10639 26086 10641 26138
rect 10395 26084 10401 26086
rect 10457 26084 10481 26086
rect 10537 26084 10561 26086
rect 10617 26084 10641 26086
rect 10697 26084 10703 26086
rect 10395 26064 10703 26084
rect 10140 26036 10192 26042
rect 10140 25978 10192 25984
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10140 25832 10192 25838
rect 10140 25774 10192 25780
rect 10152 24750 10180 25774
rect 10888 25226 10916 25842
rect 10980 25838 11008 26250
rect 10968 25832 11020 25838
rect 10968 25774 11020 25780
rect 10980 25362 11008 25774
rect 11348 25770 11376 27542
rect 11612 27328 11664 27334
rect 11612 27270 11664 27276
rect 11624 27062 11652 27270
rect 11612 27056 11664 27062
rect 11612 26998 11664 27004
rect 11428 26240 11480 26246
rect 11428 26182 11480 26188
rect 11336 25764 11388 25770
rect 11336 25706 11388 25712
rect 10968 25356 11020 25362
rect 10968 25298 11020 25304
rect 10876 25220 10928 25226
rect 10876 25162 10928 25168
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10140 24744 10192 24750
rect 10140 24686 10192 24692
rect 10152 23322 10180 24686
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10048 23316 10100 23322
rect 10048 23258 10100 23264
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10060 22794 10088 23258
rect 10244 23118 10272 23462
rect 10336 23186 10364 25094
rect 10395 25052 10703 25072
rect 10395 25050 10401 25052
rect 10457 25050 10481 25052
rect 10537 25050 10561 25052
rect 10617 25050 10641 25052
rect 10697 25050 10703 25052
rect 10457 24998 10459 25050
rect 10639 24998 10641 25050
rect 10395 24996 10401 24998
rect 10457 24996 10481 24998
rect 10537 24996 10561 24998
rect 10617 24996 10641 24998
rect 10697 24996 10703 24998
rect 10395 24976 10703 24996
rect 10416 24880 10468 24886
rect 10600 24880 10652 24886
rect 10468 24840 10600 24868
rect 10416 24822 10468 24828
rect 10600 24822 10652 24828
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 10428 24274 10456 24550
rect 10796 24410 10824 24754
rect 10784 24404 10836 24410
rect 10784 24346 10836 24352
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 10395 23964 10703 23984
rect 10395 23962 10401 23964
rect 10457 23962 10481 23964
rect 10537 23962 10561 23964
rect 10617 23962 10641 23964
rect 10697 23962 10703 23964
rect 10457 23910 10459 23962
rect 10639 23910 10641 23962
rect 10395 23908 10401 23910
rect 10457 23908 10481 23910
rect 10537 23908 10561 23910
rect 10617 23908 10641 23910
rect 10697 23908 10703 23910
rect 10395 23888 10703 23908
rect 10888 23866 10916 25162
rect 10980 24750 11008 25298
rect 10968 24744 11020 24750
rect 10968 24686 11020 24692
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10232 23112 10284 23118
rect 10284 23060 10364 23066
rect 10232 23054 10364 23060
rect 10244 23038 10364 23054
rect 10232 22976 10284 22982
rect 10232 22918 10284 22924
rect 10244 22794 10272 22918
rect 10060 22766 10272 22794
rect 9956 22160 10008 22166
rect 9956 22102 10008 22108
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9640 21508 9720 21536
rect 9588 21490 9640 21496
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 9220 21412 9272 21418
rect 9220 21354 9272 21360
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 8864 20998 9076 21026
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 7760 19378 7788 19790
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 8208 18828 8260 18834
rect 8260 18788 8340 18816
rect 8208 18770 8260 18776
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7484 18426 7512 18702
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7576 18290 7604 18634
rect 7760 18290 7788 18770
rect 8024 18760 8076 18766
rect 8076 18720 8156 18748
rect 8024 18702 8076 18708
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7208 17054 7328 17082
rect 7392 17066 7420 17682
rect 7576 17490 7604 18226
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7484 17462 7696 17490
rect 7484 17202 7512 17462
rect 7668 17338 7696 17462
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7380 17060 7432 17066
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7116 15638 7144 16186
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 7116 14822 7144 15438
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6932 13870 6960 14350
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 13938 7052 14214
rect 7116 13938 7144 14758
rect 7208 14278 7236 17054
rect 7380 17002 7432 17008
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7484 16522 7512 16934
rect 7576 16590 7604 17274
rect 7654 17232 7710 17241
rect 7654 17167 7710 17176
rect 7668 16946 7696 17167
rect 7760 17134 7788 17614
rect 7852 17202 7880 18090
rect 8128 17542 8156 18720
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 7668 16918 7788 16946
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7472 16516 7524 16522
rect 7472 16458 7524 16464
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7392 16114 7420 16390
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7760 15910 7788 16918
rect 8036 16726 8064 17070
rect 8024 16720 8076 16726
rect 8024 16662 8076 16668
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7852 16182 7880 16594
rect 7840 16176 7892 16182
rect 7840 16118 7892 16124
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7300 14958 7328 15506
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7392 15162 7420 15438
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6748 13394 6776 13738
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6656 12850 6684 13126
rect 6748 12918 6776 13330
rect 7208 13326 7236 14010
rect 7484 13938 7512 15370
rect 7668 14074 7696 15846
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7760 14414 7788 15438
rect 7852 15162 7880 16118
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 8036 15638 8064 15846
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 8128 15570 8156 17478
rect 8220 16794 8248 18362
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8312 16522 8340 18788
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 8312 15706 8340 16458
rect 8404 16114 8432 20198
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8588 18358 8616 18770
rect 8680 18698 8708 18838
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8772 18358 8800 19110
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8760 18352 8812 18358
rect 8760 18294 8812 18300
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8864 17338 8892 17614
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8496 16658 8524 17070
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8588 16794 8616 16934
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8864 16590 8892 17274
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8036 15162 8064 15438
rect 8312 15162 8340 15438
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 7852 15026 7880 15098
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8312 14414 8340 14758
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 12238 6408 12582
rect 6748 12238 6776 12854
rect 7484 12850 7512 13874
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6380 11354 6408 12174
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6472 11762 6500 12038
rect 6748 11830 6776 12174
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6380 10674 6408 11086
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6380 9722 6408 10610
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6288 9574 6592 9602
rect 5092 8974 5120 9454
rect 5672 9276 5980 9296
rect 5672 9274 5678 9276
rect 5734 9274 5758 9276
rect 5814 9274 5838 9276
rect 5894 9274 5918 9276
rect 5974 9274 5980 9276
rect 5734 9222 5736 9274
rect 5916 9222 5918 9274
rect 5672 9220 5678 9222
rect 5734 9220 5758 9222
rect 5814 9220 5838 9222
rect 5894 9220 5918 9222
rect 5974 9220 5980 9222
rect 5672 9200 5980 9220
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5092 8634 5120 8910
rect 6104 8634 6132 9454
rect 6196 9438 6408 9466
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5276 7750 5304 8434
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5460 7834 5488 8366
rect 5552 8022 5580 8366
rect 6104 8242 6132 8570
rect 6276 8288 6328 8294
rect 6104 8214 6224 8242
rect 6276 8230 6328 8236
rect 5672 8188 5980 8208
rect 5672 8186 5678 8188
rect 5734 8186 5758 8188
rect 5814 8186 5838 8188
rect 5894 8186 5918 8188
rect 5974 8186 5980 8188
rect 5734 8134 5736 8186
rect 5916 8134 5918 8186
rect 5672 8132 5678 8134
rect 5734 8132 5758 8134
rect 5814 8132 5838 8134
rect 5894 8132 5918 8134
rect 5974 8132 5980 8134
rect 5672 8112 5980 8132
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6104 7886 6132 7958
rect 5540 7880 5592 7886
rect 5460 7828 5540 7834
rect 5460 7822 5592 7828
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5460 7806 5580 7822
rect 6196 7818 6224 8214
rect 6288 7886 6316 8230
rect 6380 7970 6408 9438
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6472 8566 6500 8910
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6472 8090 6500 8502
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6380 7942 6500 7970
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 6798 4936 7142
rect 5552 6798 5580 7806
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5672 7100 5980 7120
rect 5672 7098 5678 7100
rect 5734 7098 5758 7100
rect 5814 7098 5838 7100
rect 5894 7098 5918 7100
rect 5974 7098 5980 7100
rect 5734 7046 5736 7098
rect 5916 7046 5918 7098
rect 5672 7044 5678 7046
rect 5734 7044 5758 7046
rect 5814 7044 5838 7046
rect 5894 7044 5918 7046
rect 5974 7044 5980 7046
rect 5672 7024 5980 7044
rect 6012 7002 6040 7346
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 5540 6792 5592 6798
rect 6184 6792 6236 6798
rect 5540 6734 5592 6740
rect 6104 6752 6184 6780
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 6012 6390 6040 6666
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4724 6310 4844 6338
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 4896 6316 4948 6322
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 2700 5370 2728 5510
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 3160 5234 3188 5510
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 4080 5166 4108 5510
rect 4264 5370 4292 5646
rect 4632 5642 4660 6258
rect 4724 5778 4752 6310
rect 4896 6258 4948 6264
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4816 5642 4844 6122
rect 4908 5914 4936 6258
rect 6104 6202 6132 6752
rect 6184 6734 6236 6740
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6012 6186 6132 6202
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 6000 6180 6132 6186
rect 6052 6174 6132 6180
rect 6000 6122 6052 6128
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5276 5710 5304 6054
rect 5460 5710 5488 6122
rect 5672 6012 5980 6032
rect 5672 6010 5678 6012
rect 5734 6010 5758 6012
rect 5814 6010 5838 6012
rect 5894 6010 5918 6012
rect 5974 6010 5980 6012
rect 5734 5958 5736 6010
rect 5916 5958 5918 6010
rect 5672 5956 5678 5958
rect 5734 5956 5758 5958
rect 5814 5956 5838 5958
rect 5894 5956 5918 5958
rect 5974 5956 5980 5958
rect 5672 5936 5980 5956
rect 5816 5840 5868 5846
rect 6012 5828 6040 6122
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5816 5782 5868 5788
rect 5920 5800 6040 5828
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4622 3924 4966
rect 3988 4865 4016 5034
rect 3974 4856 4030 4865
rect 4816 4826 4844 5578
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4908 5234 4936 5510
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 3974 4791 4030 4800
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 1400 4480 1452 4486
rect 1400 4422 1452 4428
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1412 3505 1440 4422
rect 3804 4214 3832 4558
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 5460 3942 5488 5646
rect 5828 5302 5856 5782
rect 5920 5710 5948 5800
rect 6104 5710 6132 5850
rect 6196 5846 6224 6258
rect 6380 5914 6408 6258
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6184 5840 6236 5846
rect 6472 5794 6500 7942
rect 6184 5782 6236 5788
rect 6196 5710 6224 5782
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6380 5766 6500 5794
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5672 4924 5980 4944
rect 5672 4922 5678 4924
rect 5734 4922 5758 4924
rect 5814 4922 5838 4924
rect 5894 4922 5918 4924
rect 5974 4922 5980 4924
rect 5734 4870 5736 4922
rect 5916 4870 5918 4922
rect 5672 4868 5678 4870
rect 5734 4868 5758 4870
rect 5814 4868 5838 4870
rect 5894 4868 5918 4870
rect 5974 4868 5980 4870
rect 5672 4848 5980 4868
rect 6012 4622 6040 5578
rect 6092 5296 6144 5302
rect 6196 5284 6224 5646
rect 6288 5302 6316 5714
rect 6144 5256 6224 5284
rect 6276 5296 6328 5302
rect 6092 5238 6144 5244
rect 6276 5238 6328 5244
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5448 3936 5500 3942
rect 5920 3924 5948 4082
rect 6000 3936 6052 3942
rect 5920 3896 6000 3924
rect 5448 3878 5500 3884
rect 6000 3878 6052 3884
rect 5672 3836 5980 3856
rect 5672 3834 5678 3836
rect 5734 3834 5758 3836
rect 5814 3834 5838 3836
rect 5894 3834 5918 3836
rect 5974 3834 5980 3836
rect 5734 3782 5736 3834
rect 5916 3782 5918 3834
rect 5672 3780 5678 3782
rect 5734 3780 5758 3782
rect 5814 3780 5838 3782
rect 5894 3780 5918 3782
rect 5974 3780 5980 3782
rect 5672 3760 5980 3780
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1308 3470 1360 3476
rect 1398 3496 1454 3505
rect 584 800 612 3470
rect 1398 3431 1454 3440
rect 1780 800 1808 3538
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2976 800 3004 2926
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3068 2145 3096 2586
rect 3054 2136 3110 2145
rect 3054 2071 3110 2080
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 570 0 626 800
rect 1766 0 1822 800
rect 2962 0 3018 800
rect 3344 785 3372 1294
rect 4172 800 4200 3606
rect 6380 3602 6408 5766
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6472 3534 6500 3878
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5460 800 5488 3402
rect 5672 2748 5980 2768
rect 5672 2746 5678 2748
rect 5734 2746 5758 2748
rect 5814 2746 5838 2748
rect 5894 2746 5918 2748
rect 5974 2746 5980 2748
rect 5734 2694 5736 2746
rect 5916 2694 5918 2746
rect 5672 2692 5678 2694
rect 5734 2692 5758 2694
rect 5814 2692 5838 2694
rect 5894 2692 5918 2694
rect 5974 2692 5980 2694
rect 5672 2672 5980 2692
rect 6564 1358 6592 9574
rect 6656 9042 6684 11222
rect 6748 10674 6776 11766
rect 7300 11354 7328 12786
rect 7656 12436 7708 12442
rect 7760 12434 7788 14214
rect 8220 14006 8248 14214
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8312 13530 8340 14010
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8404 12782 8432 16050
rect 8484 15904 8536 15910
rect 8588 15892 8616 16526
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8536 15864 8616 15892
rect 8484 15846 8536 15852
rect 8588 15366 8616 15864
rect 8680 15502 8708 16186
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8772 15910 8800 16050
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7708 12406 7788 12434
rect 7656 12378 7708 12384
rect 7760 11762 7788 12406
rect 7944 12238 7972 12650
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7760 11218 7788 11494
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6932 9382 6960 10406
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9586 7236 9862
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6656 7546 6684 8978
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6840 8498 6868 8774
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6932 8430 6960 9318
rect 7116 8634 7144 9318
rect 7300 9178 7328 9522
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7576 8634 7604 8842
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7546 6868 7822
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6656 5234 6684 7482
rect 7116 7342 7144 8366
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7546 7328 7686
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7116 6798 7144 7278
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7760 6798 7788 7142
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7024 5234 7052 5510
rect 6644 5228 6696 5234
rect 7012 5228 7064 5234
rect 6696 5188 6776 5216
rect 6644 5170 6696 5176
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6656 3738 6684 4014
rect 6748 4010 6776 5188
rect 7012 5170 7064 5176
rect 7116 5166 7144 6734
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 7012 4480 7064 4486
rect 7116 4468 7144 5102
rect 7064 4440 7144 4468
rect 7012 4422 7064 4428
rect 6932 4282 6960 4422
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 7024 4078 7052 4422
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6552 1352 6604 1358
rect 6552 1294 6604 1300
rect 6656 800 6684 3538
rect 7944 3466 7972 9318
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8128 7206 8156 8366
rect 8312 7954 8340 8910
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 3602 8156 7142
rect 8312 6780 8340 7890
rect 8392 6792 8444 6798
rect 8312 6752 8392 6780
rect 8444 6752 8524 6780
rect 8392 6734 8444 6740
rect 8496 5710 8524 6752
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8312 5098 8340 5578
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8496 4690 8524 5646
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7852 800 7880 2926
rect 8588 1358 8616 15302
rect 8680 14890 8708 15438
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8680 12646 8708 12922
rect 8772 12850 8800 15846
rect 9048 14822 9076 20998
rect 9232 20924 9260 21354
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 9312 20936 9364 20942
rect 9232 20896 9312 20924
rect 9312 20878 9364 20884
rect 9128 20868 9180 20874
rect 9128 20810 9180 20816
rect 9140 20330 9168 20810
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9232 17882 9260 18362
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9232 17338 9260 17818
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9232 16726 9260 17138
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9324 16658 9352 16934
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9416 15434 9444 21286
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9692 19514 9720 20334
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9968 18834 9996 21422
rect 10060 20466 10088 22766
rect 10336 22692 10364 23038
rect 10395 22876 10703 22896
rect 10395 22874 10401 22876
rect 10457 22874 10481 22876
rect 10537 22874 10561 22876
rect 10617 22874 10641 22876
rect 10697 22874 10703 22876
rect 10457 22822 10459 22874
rect 10639 22822 10641 22874
rect 10395 22820 10401 22822
rect 10457 22820 10481 22822
rect 10537 22820 10561 22822
rect 10617 22820 10641 22822
rect 10697 22820 10703 22822
rect 10395 22800 10703 22820
rect 10796 22760 10824 23666
rect 10612 22732 10824 22760
rect 10152 22664 10364 22692
rect 10416 22704 10468 22710
rect 10414 22672 10416 22681
rect 10468 22672 10470 22681
rect 10152 21622 10180 22664
rect 10414 22607 10470 22616
rect 10612 22166 10640 22732
rect 10876 22704 10928 22710
rect 10876 22646 10928 22652
rect 10692 22500 10744 22506
rect 10692 22442 10744 22448
rect 10232 22160 10284 22166
rect 10232 22102 10284 22108
rect 10600 22160 10652 22166
rect 10600 22102 10652 22108
rect 10140 21616 10192 21622
rect 10140 21558 10192 21564
rect 10244 21434 10272 22102
rect 10704 22030 10732 22442
rect 10888 22030 10916 22646
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10324 21956 10376 21962
rect 10324 21898 10376 21904
rect 10336 21622 10364 21898
rect 10395 21788 10703 21808
rect 10395 21786 10401 21788
rect 10457 21786 10481 21788
rect 10537 21786 10561 21788
rect 10617 21786 10641 21788
rect 10697 21786 10703 21788
rect 10457 21734 10459 21786
rect 10639 21734 10641 21786
rect 10395 21732 10401 21734
rect 10457 21732 10481 21734
rect 10537 21732 10561 21734
rect 10617 21732 10641 21734
rect 10697 21732 10703 21734
rect 10395 21712 10703 21732
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10324 21616 10376 21622
rect 10324 21558 10376 21564
rect 10796 21554 10824 21626
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10152 21406 10272 21434
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10060 18154 10088 18702
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9508 16250 9536 17546
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9784 16998 9812 17478
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9968 16726 9996 17138
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9404 15428 9456 15434
rect 9404 15370 9456 15376
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9324 14074 9352 14962
rect 9508 14890 9536 16050
rect 9692 15910 9720 16594
rect 10152 16046 10180 21406
rect 10704 20890 10732 21422
rect 10888 21418 10916 21966
rect 10876 21412 10928 21418
rect 10876 21354 10928 21360
rect 10704 20862 10824 20890
rect 10395 20700 10703 20720
rect 10395 20698 10401 20700
rect 10457 20698 10481 20700
rect 10537 20698 10561 20700
rect 10617 20698 10641 20700
rect 10697 20698 10703 20700
rect 10457 20646 10459 20698
rect 10639 20646 10641 20698
rect 10395 20644 10401 20646
rect 10457 20644 10481 20646
rect 10537 20644 10561 20646
rect 10617 20644 10641 20646
rect 10697 20644 10703 20646
rect 10395 20624 10703 20644
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10704 19854 10732 20402
rect 10796 20330 10824 20862
rect 10980 20466 11008 24686
rect 11348 24274 11376 25706
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 11060 24132 11112 24138
rect 11060 24074 11112 24080
rect 11072 22438 11100 24074
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 11164 20330 11192 24142
rect 11440 23526 11468 26182
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 11704 25832 11756 25838
rect 11702 25800 11704 25809
rect 11756 25800 11758 25809
rect 11624 25758 11702 25786
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11532 24614 11560 24686
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 11532 24410 11560 24550
rect 11520 24404 11572 24410
rect 11520 24346 11572 24352
rect 11428 23520 11480 23526
rect 11428 23462 11480 23468
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11256 23118 11284 23258
rect 11440 23254 11468 23462
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11256 21690 11284 23054
rect 11336 23044 11388 23050
rect 11336 22986 11388 22992
rect 11348 22642 11376 22986
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11440 21418 11468 23190
rect 11520 22976 11572 22982
rect 11520 22918 11572 22924
rect 11532 22642 11560 22918
rect 11624 22642 11652 25758
rect 11702 25735 11758 25744
rect 11808 25498 11836 25842
rect 11796 25492 11848 25498
rect 11796 25434 11848 25440
rect 11796 25152 11848 25158
rect 11796 25094 11848 25100
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11716 23186 11744 23598
rect 11808 23526 11836 25094
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11808 23050 11836 23462
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 11520 22636 11572 22642
rect 11520 22578 11572 22584
rect 11612 22636 11664 22642
rect 11612 22578 11664 22584
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 11612 22500 11664 22506
rect 11612 22442 11664 22448
rect 11520 22160 11572 22166
rect 11518 22128 11520 22137
rect 11572 22128 11574 22137
rect 11518 22063 11574 22072
rect 11532 22030 11560 22063
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11532 21486 11560 21966
rect 11520 21480 11572 21486
rect 11520 21422 11572 21428
rect 11428 21412 11480 21418
rect 11428 21354 11480 21360
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11532 20806 11560 21286
rect 11520 20800 11572 20806
rect 11520 20742 11572 20748
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 10784 20324 10836 20330
rect 10784 20266 10836 20272
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10395 19612 10703 19632
rect 10395 19610 10401 19612
rect 10457 19610 10481 19612
rect 10537 19610 10561 19612
rect 10617 19610 10641 19612
rect 10697 19610 10703 19612
rect 10457 19558 10459 19610
rect 10639 19558 10641 19610
rect 10395 19556 10401 19558
rect 10457 19556 10481 19558
rect 10537 19556 10561 19558
rect 10617 19556 10641 19558
rect 10697 19556 10703 19558
rect 10395 19536 10703 19556
rect 10600 19440 10652 19446
rect 10966 19408 11022 19417
rect 10652 19388 10966 19394
rect 10600 19382 10966 19388
rect 10612 19366 10966 19382
rect 11164 19378 11192 19994
rect 11256 19922 11284 20402
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11256 19446 11284 19654
rect 11348 19514 11376 19790
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 11244 19440 11296 19446
rect 11244 19382 11296 19388
rect 10966 19343 11022 19352
rect 11060 19372 11112 19378
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10336 18222 10364 18702
rect 10888 18630 10916 18838
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10395 18524 10703 18544
rect 10395 18522 10401 18524
rect 10457 18522 10481 18524
rect 10537 18522 10561 18524
rect 10617 18522 10641 18524
rect 10697 18522 10703 18524
rect 10457 18470 10459 18522
rect 10639 18470 10641 18522
rect 10395 18468 10401 18470
rect 10457 18468 10481 18470
rect 10537 18468 10561 18470
rect 10617 18468 10641 18470
rect 10697 18468 10703 18470
rect 10395 18448 10703 18468
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10888 17678 10916 18566
rect 10784 17672 10836 17678
rect 10876 17672 10928 17678
rect 10784 17614 10836 17620
rect 10874 17640 10876 17649
rect 10928 17640 10930 17649
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10336 17270 10364 17546
rect 10395 17436 10703 17456
rect 10395 17434 10401 17436
rect 10457 17434 10481 17436
rect 10537 17434 10561 17436
rect 10617 17434 10641 17436
rect 10697 17434 10703 17436
rect 10457 17382 10459 17434
rect 10639 17382 10641 17434
rect 10395 17380 10401 17382
rect 10457 17380 10481 17382
rect 10537 17380 10561 17382
rect 10617 17380 10641 17382
rect 10697 17380 10703 17382
rect 10395 17360 10703 17380
rect 10796 17338 10824 17614
rect 10874 17575 10930 17584
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 10888 16590 10916 17478
rect 10980 17320 11008 19343
rect 11060 19314 11112 19320
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11072 17814 11100 19314
rect 11256 18358 11284 19382
rect 11244 18352 11296 18358
rect 11244 18294 11296 18300
rect 11348 18306 11376 19450
rect 11440 18902 11468 19790
rect 11532 19334 11560 20742
rect 11624 20466 11652 22442
rect 11716 21962 11744 22510
rect 11808 22506 11836 22986
rect 11796 22500 11848 22506
rect 11796 22442 11848 22448
rect 11992 22094 12020 28562
rect 12176 26994 12204 29038
rect 12440 28076 12492 28082
rect 12440 28018 12492 28024
rect 12348 27600 12400 27606
rect 12452 27554 12480 28018
rect 12400 27548 12480 27554
rect 12348 27542 12480 27548
rect 12360 27526 12480 27542
rect 12164 26988 12216 26994
rect 12164 26930 12216 26936
rect 12544 26790 12572 29106
rect 12912 28558 12940 29106
rect 13280 28558 13308 29106
rect 13648 29102 13676 29582
rect 13636 29096 13688 29102
rect 13636 29038 13688 29044
rect 13924 29084 13952 31889
rect 15212 31770 15240 31889
rect 15304 31878 15516 31906
rect 16578 31889 16634 32689
rect 17866 31889 17922 32689
rect 19246 31889 19302 32689
rect 20534 31889 20590 32689
rect 21822 31889 21878 32689
rect 23202 31889 23258 32689
rect 24490 31889 24546 32689
rect 25870 31889 25926 32689
rect 27158 31889 27214 32689
rect 28538 31889 28594 32689
rect 29826 31889 29882 32689
rect 15304 31770 15332 31878
rect 15212 31742 15332 31770
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 14648 30048 14700 30054
rect 14648 29990 14700 29996
rect 14660 29578 14688 29990
rect 14648 29572 14700 29578
rect 14648 29514 14700 29520
rect 14372 29504 14424 29510
rect 14372 29446 14424 29452
rect 14384 29238 14412 29446
rect 14372 29232 14424 29238
rect 14372 29174 14424 29180
rect 14096 29096 14148 29102
rect 13924 29056 14096 29084
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 13268 28552 13320 28558
rect 13268 28494 13320 28500
rect 12624 27872 12676 27878
rect 12624 27814 12676 27820
rect 12636 27402 12664 27814
rect 12716 27532 12768 27538
rect 12716 27474 12768 27480
rect 12624 27396 12676 27402
rect 12624 27338 12676 27344
rect 12622 27160 12678 27169
rect 12622 27095 12624 27104
rect 12676 27095 12678 27104
rect 12624 27066 12676 27072
rect 12728 26994 12756 27474
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 12164 26240 12216 26246
rect 12164 26182 12216 26188
rect 12176 25974 12204 26182
rect 12164 25968 12216 25974
rect 12164 25910 12216 25916
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12544 25702 12572 25842
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 12256 25696 12308 25702
rect 12532 25696 12584 25702
rect 12256 25638 12308 25644
rect 12530 25664 12532 25673
rect 12584 25664 12586 25673
rect 12084 25294 12112 25638
rect 12268 25498 12296 25638
rect 12530 25599 12586 25608
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12532 24880 12584 24886
rect 12532 24822 12584 24828
rect 12164 24812 12216 24818
rect 12164 24754 12216 24760
rect 12176 23866 12204 24754
rect 12440 24608 12492 24614
rect 12544 24562 12572 24822
rect 12636 24682 12664 25094
rect 12728 24818 12756 25230
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12820 24750 12848 25094
rect 12808 24744 12860 24750
rect 12808 24686 12860 24692
rect 12912 24682 12940 28494
rect 12992 27328 13044 27334
rect 12992 27270 13044 27276
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 13004 27130 13032 27270
rect 12992 27124 13044 27130
rect 12992 27066 13044 27072
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 13004 25430 13032 25638
rect 12992 25424 13044 25430
rect 12992 25366 13044 25372
rect 12624 24676 12676 24682
rect 12624 24618 12676 24624
rect 12900 24676 12952 24682
rect 12900 24618 12952 24624
rect 12912 24562 12940 24618
rect 13004 24614 13032 25366
rect 13096 24750 13124 27270
rect 13176 26580 13228 26586
rect 13176 26522 13228 26528
rect 13188 26382 13216 26522
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 13174 25800 13230 25809
rect 13174 25735 13176 25744
rect 13228 25735 13230 25744
rect 13176 25706 13228 25712
rect 13280 25294 13308 28494
rect 13648 27470 13676 29038
rect 13728 28960 13780 28966
rect 13728 28902 13780 28908
rect 13740 28762 13768 28902
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 13924 28490 13952 29056
rect 14096 29038 14148 29044
rect 14936 28762 14964 30194
rect 15118 29948 15426 29968
rect 15118 29946 15124 29948
rect 15180 29946 15204 29948
rect 15260 29946 15284 29948
rect 15340 29946 15364 29948
rect 15420 29946 15426 29948
rect 15180 29894 15182 29946
rect 15362 29894 15364 29946
rect 15118 29892 15124 29894
rect 15180 29892 15204 29894
rect 15260 29892 15284 29894
rect 15340 29892 15364 29894
rect 15420 29892 15426 29894
rect 15118 29872 15426 29892
rect 15384 29572 15436 29578
rect 15384 29514 15436 29520
rect 15396 29306 15424 29514
rect 15384 29300 15436 29306
rect 15384 29242 15436 29248
rect 15118 28860 15426 28880
rect 15118 28858 15124 28860
rect 15180 28858 15204 28860
rect 15260 28858 15284 28860
rect 15340 28858 15364 28860
rect 15420 28858 15426 28860
rect 15180 28806 15182 28858
rect 15362 28806 15364 28858
rect 15118 28804 15124 28806
rect 15180 28804 15204 28806
rect 15260 28804 15284 28806
rect 15340 28804 15364 28806
rect 15420 28804 15426 28806
rect 15118 28784 15426 28804
rect 14924 28756 14976 28762
rect 14924 28698 14976 28704
rect 15488 28694 15516 31878
rect 15660 29708 15712 29714
rect 15660 29650 15712 29656
rect 15672 29102 15700 29650
rect 15844 29504 15896 29510
rect 15844 29446 15896 29452
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 15476 28688 15528 28694
rect 15476 28630 15528 28636
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 13912 28484 13964 28490
rect 13912 28426 13964 28432
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13636 27464 13688 27470
rect 13636 27406 13688 27412
rect 13360 27396 13412 27402
rect 13360 27338 13412 27344
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 13372 27062 13400 27338
rect 13740 27146 13768 27338
rect 13648 27118 13768 27146
rect 13360 27056 13412 27062
rect 13360 26998 13412 27004
rect 13544 26988 13596 26994
rect 13544 26930 13596 26936
rect 13556 26450 13584 26930
rect 13544 26444 13596 26450
rect 13544 26386 13596 26392
rect 13452 25424 13504 25430
rect 13452 25366 13504 25372
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13280 24886 13308 25230
rect 13464 24886 13492 25366
rect 13556 25276 13584 26386
rect 13648 25702 13676 27118
rect 13832 25770 13860 28086
rect 14016 26246 14044 28358
rect 14096 28076 14148 28082
rect 14096 28018 14148 28024
rect 14108 27470 14136 28018
rect 14556 27940 14608 27946
rect 14556 27882 14608 27888
rect 14464 27872 14516 27878
rect 14464 27814 14516 27820
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14108 26994 14136 27406
rect 14476 27130 14504 27814
rect 14568 27470 14596 27882
rect 15118 27772 15426 27792
rect 15118 27770 15124 27772
rect 15180 27770 15204 27772
rect 15260 27770 15284 27772
rect 15340 27770 15364 27772
rect 15420 27770 15426 27772
rect 15180 27718 15182 27770
rect 15362 27718 15364 27770
rect 15118 27716 15124 27718
rect 15180 27716 15204 27718
rect 15260 27716 15284 27718
rect 15340 27716 15364 27718
rect 15420 27716 15426 27718
rect 15118 27696 15426 27716
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14568 27130 14596 27406
rect 15198 27160 15254 27169
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14924 27124 14976 27130
rect 15198 27095 15254 27104
rect 14924 27066 14976 27072
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14096 26852 14148 26858
rect 14096 26794 14148 26800
rect 14004 26240 14056 26246
rect 14004 26182 14056 26188
rect 13820 25764 13872 25770
rect 13820 25706 13872 25712
rect 13636 25696 13688 25702
rect 13636 25638 13688 25644
rect 13636 25288 13688 25294
rect 13556 25248 13636 25276
rect 13636 25230 13688 25236
rect 13268 24880 13320 24886
rect 13268 24822 13320 24828
rect 13452 24880 13504 24886
rect 13452 24822 13504 24828
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 12492 24556 12572 24562
rect 12440 24550 12572 24556
rect 12452 24534 12572 24550
rect 12164 23860 12216 23866
rect 12164 23802 12216 23808
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 11992 22066 12112 22094
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11624 19446 11652 20402
rect 11716 19446 11744 21898
rect 11794 21040 11850 21049
rect 11794 20975 11850 20984
rect 11612 19440 11664 19446
rect 11612 19382 11664 19388
rect 11704 19440 11756 19446
rect 11704 19382 11756 19388
rect 11532 19306 11652 19334
rect 11428 18896 11480 18902
rect 11480 18856 11560 18884
rect 11428 18838 11480 18844
rect 11348 18290 11468 18306
rect 11348 18284 11480 18290
rect 11348 18278 11428 18284
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 11256 17678 11284 18158
rect 11348 18086 11376 18278
rect 11428 18226 11480 18232
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11244 17332 11296 17338
rect 10980 17292 11192 17320
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10395 16348 10703 16368
rect 10395 16346 10401 16348
rect 10457 16346 10481 16348
rect 10537 16346 10561 16348
rect 10617 16346 10641 16348
rect 10697 16346 10703 16348
rect 10457 16294 10459 16346
rect 10639 16294 10641 16346
rect 10395 16292 10401 16294
rect 10457 16292 10481 16294
rect 10537 16292 10561 16294
rect 10617 16292 10641 16294
rect 10697 16292 10703 16294
rect 10395 16272 10703 16292
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9692 14414 9720 15846
rect 10980 15706 11008 17138
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10060 15026 10088 15642
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 10336 15162 10364 15370
rect 10395 15260 10703 15280
rect 10395 15258 10401 15260
rect 10457 15258 10481 15260
rect 10537 15258 10561 15260
rect 10617 15258 10641 15260
rect 10697 15258 10703 15260
rect 10457 15206 10459 15258
rect 10639 15206 10641 15258
rect 10395 15204 10401 15206
rect 10457 15204 10481 15206
rect 10537 15204 10561 15206
rect 10617 15204 10641 15206
rect 10697 15204 10703 15206
rect 10395 15184 10703 15204
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10796 14618 10824 14962
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10395 14172 10703 14192
rect 10395 14170 10401 14172
rect 10457 14170 10481 14172
rect 10537 14170 10561 14172
rect 10617 14170 10641 14172
rect 10697 14170 10703 14172
rect 10457 14118 10459 14170
rect 10639 14118 10641 14170
rect 10395 14116 10401 14118
rect 10457 14116 10481 14118
rect 10537 14116 10561 14118
rect 10617 14116 10641 14118
rect 10697 14116 10703 14118
rect 10395 14096 10703 14116
rect 10796 14074 10824 14350
rect 10888 14278 10916 14962
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10152 13938 10180 14010
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8772 12442 8800 12786
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8772 11898 8800 12378
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8864 11830 8892 12854
rect 9508 12442 9536 12854
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9496 12232 9548 12238
rect 9692 12220 9720 12310
rect 9548 12192 9720 12220
rect 9496 12174 9548 12180
rect 9680 12096 9732 12102
rect 9600 12056 9680 12084
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9140 10742 9168 10950
rect 9128 10736 9180 10742
rect 9128 10678 9180 10684
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8956 9654 8984 9862
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 9140 9178 9168 9998
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8772 8498 8800 8910
rect 9232 8566 9260 11834
rect 9600 11150 9628 12056
rect 9680 12038 9732 12044
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9692 10674 9720 11222
rect 10060 11218 10088 12854
rect 10152 12374 10180 13874
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10428 13258 10456 13670
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10395 13084 10703 13104
rect 10395 13082 10401 13084
rect 10457 13082 10481 13084
rect 10537 13082 10561 13084
rect 10617 13082 10641 13084
rect 10697 13082 10703 13084
rect 10457 13030 10459 13082
rect 10639 13030 10641 13082
rect 10395 13028 10401 13030
rect 10457 13028 10481 13030
rect 10537 13028 10561 13030
rect 10617 13028 10641 13030
rect 10697 13028 10703 13030
rect 10395 13008 10703 13028
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 10152 11762 10180 12310
rect 10395 11996 10703 12016
rect 10395 11994 10401 11996
rect 10457 11994 10481 11996
rect 10537 11994 10561 11996
rect 10617 11994 10641 11996
rect 10697 11994 10703 11996
rect 10457 11942 10459 11994
rect 10639 11942 10641 11994
rect 10395 11940 10401 11942
rect 10457 11940 10481 11942
rect 10537 11940 10561 11942
rect 10617 11940 10641 11942
rect 10697 11940 10703 11942
rect 10395 11920 10703 11940
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10152 11082 10180 11698
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10428 11218 10456 11494
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10612 11082 10640 11494
rect 10796 11354 10824 11494
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10395 10908 10703 10928
rect 10395 10906 10401 10908
rect 10457 10906 10481 10908
rect 10537 10906 10561 10908
rect 10617 10906 10641 10908
rect 10697 10906 10703 10908
rect 10457 10854 10459 10906
rect 10639 10854 10641 10906
rect 10395 10852 10401 10854
rect 10457 10852 10481 10854
rect 10537 10852 10561 10854
rect 10617 10852 10641 10854
rect 10697 10852 10703 10854
rect 10395 10832 10703 10852
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 7886 9168 8230
rect 9232 8090 9260 8502
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9324 7818 9352 8298
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 7478 8984 7686
rect 9324 7478 9352 7754
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9416 7324 9444 10406
rect 9692 9654 9720 10610
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9692 8514 9720 9590
rect 9784 9382 9812 9590
rect 10336 9586 10364 10406
rect 10395 9820 10703 9840
rect 10395 9818 10401 9820
rect 10457 9818 10481 9820
rect 10537 9818 10561 9820
rect 10617 9818 10641 9820
rect 10697 9818 10703 9820
rect 10457 9766 10459 9818
rect 10639 9766 10641 9818
rect 10395 9764 10401 9766
rect 10457 9764 10481 9766
rect 10537 9764 10561 9766
rect 10617 9764 10641 9766
rect 10697 9764 10703 9766
rect 10395 9744 10703 9764
rect 10888 9704 10916 14214
rect 10980 13394 11008 15506
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10980 12918 11008 13330
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 11072 12322 11100 15642
rect 10980 12294 11100 12322
rect 11164 12306 11192 17292
rect 11244 17274 11296 17280
rect 11256 16590 11284 17274
rect 11440 16590 11468 18022
rect 11532 17202 11560 18856
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11428 16584 11480 16590
rect 11480 16544 11560 16572
rect 11428 16526 11480 16532
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 11348 15570 11376 16458
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11440 14346 11468 14758
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11532 12434 11560 16544
rect 11624 15706 11652 19306
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11716 18358 11744 18634
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11808 18170 11836 20975
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11992 20058 12020 20402
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11716 18142 11836 18170
rect 11716 17882 11744 18142
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11900 17542 11928 19790
rect 12084 19666 12112 22066
rect 12164 21956 12216 21962
rect 12164 21898 12216 21904
rect 12176 21622 12204 21898
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12176 20369 12204 20402
rect 12162 20360 12218 20369
rect 12162 20295 12218 20304
rect 12268 19972 12296 21626
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12360 20074 12388 21354
rect 12452 21146 12480 22646
rect 12544 22506 12572 24534
rect 12820 24534 12940 24562
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12716 24132 12768 24138
rect 12716 24074 12768 24080
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12636 23730 12664 24006
rect 12728 23866 12756 24074
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12636 22710 12664 23666
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12532 22500 12584 22506
rect 12532 22442 12584 22448
rect 12820 22234 12848 24534
rect 13096 24274 13124 24686
rect 13084 24268 13136 24274
rect 13084 24210 13136 24216
rect 13096 23662 13124 24210
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 13084 23656 13136 23662
rect 13084 23598 13136 23604
rect 13084 23180 13136 23186
rect 13084 23122 13136 23128
rect 12900 23044 12952 23050
rect 12900 22986 12952 22992
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 12820 21894 12848 22170
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12360 20046 12572 20074
rect 12268 19944 12480 19972
rect 12084 19638 12204 19666
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11992 17882 12020 19450
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 12084 19174 12112 19314
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 12084 18902 12112 19110
rect 12072 18896 12124 18902
rect 12072 18838 12124 18844
rect 12084 18222 12112 18838
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11980 17672 12032 17678
rect 11978 17640 11980 17649
rect 12072 17672 12124 17678
rect 12032 17640 12034 17649
rect 12072 17614 12124 17620
rect 11978 17575 12034 17584
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 12084 17338 12112 17614
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12176 17241 12204 19638
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12268 17921 12296 19382
rect 12452 18834 12480 19944
rect 12544 18902 12572 20046
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12360 18290 12388 18362
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12254 17912 12310 17921
rect 12254 17847 12310 17856
rect 12360 17338 12388 18226
rect 12452 17882 12480 18770
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12348 17332 12400 17338
rect 12268 17292 12348 17320
rect 12162 17232 12218 17241
rect 12162 17167 12218 17176
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11716 15162 11744 15370
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11624 14414 11652 14486
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11440 12406 11560 12434
rect 11152 12300 11204 12306
rect 10980 10554 11008 12294
rect 11152 12242 11204 12248
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11072 10674 11100 12174
rect 11348 11762 11376 12242
rect 11440 12238 11468 12406
rect 11428 12232 11480 12238
rect 11624 12186 11652 14350
rect 11808 14278 11836 16934
rect 12268 16590 12296 17292
rect 12348 17274 12400 17280
rect 12544 16708 12572 18702
rect 12636 18358 12664 20878
rect 12716 19780 12768 19786
rect 12716 19722 12768 19728
rect 12728 19378 12756 19722
rect 12820 19378 12848 21490
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12728 18630 12756 18702
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12636 17202 12664 18294
rect 12820 17882 12848 19314
rect 12912 18902 12940 22986
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 13004 21622 13032 21830
rect 12992 21616 13044 21622
rect 12992 21558 13044 21564
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 13004 19854 13032 20742
rect 13096 20466 13124 23122
rect 13188 23050 13216 23666
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 13188 22642 13216 22986
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 13372 22094 13400 22374
rect 13280 22066 13400 22094
rect 13648 22094 13676 25230
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13740 23322 13768 23598
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13648 22066 13860 22094
rect 13280 22030 13308 22066
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13556 21690 13584 21830
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 13556 20942 13584 21626
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13084 20460 13136 20466
rect 13360 20460 13412 20466
rect 13136 20420 13308 20448
rect 13084 20402 13136 20408
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13176 19780 13228 19786
rect 13176 19722 13228 19728
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 13004 18766 13032 19110
rect 13096 18970 13124 19314
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12806 17776 12862 17785
rect 12806 17711 12862 17720
rect 12820 17678 12848 17711
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12452 16680 12572 16708
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12452 16522 12480 16680
rect 12636 16574 12664 17138
rect 13004 16794 13032 18702
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13096 17678 13124 18566
rect 13188 18290 13216 19722
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13188 18154 13216 18226
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 13280 17785 13308 20420
rect 13360 20402 13412 20408
rect 13372 19310 13400 20402
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13372 18222 13400 19246
rect 13464 18766 13492 20198
rect 13556 19922 13584 20878
rect 13636 20800 13688 20806
rect 13636 20742 13688 20748
rect 13648 20330 13676 20742
rect 13636 20324 13688 20330
rect 13636 20266 13688 20272
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13648 19718 13676 20266
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13556 18612 13584 18770
rect 13648 18766 13676 19654
rect 13740 19514 13768 21422
rect 13832 21146 13860 22066
rect 14016 21298 14044 26182
rect 14108 25838 14136 26794
rect 14476 26790 14504 26930
rect 14464 26784 14516 26790
rect 14464 26726 14516 26732
rect 14568 26586 14596 27066
rect 14936 26858 14964 27066
rect 15212 26994 15240 27095
rect 15200 26988 15252 26994
rect 15200 26930 15252 26936
rect 14924 26852 14976 26858
rect 14924 26794 14976 26800
rect 15488 26790 15516 28494
rect 15672 27470 15700 29038
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 15660 27464 15712 27470
rect 15660 27406 15712 27412
rect 14832 26784 14884 26790
rect 14832 26726 14884 26732
rect 15476 26784 15528 26790
rect 15476 26726 15528 26732
rect 14556 26580 14608 26586
rect 14556 26522 14608 26528
rect 14568 26314 14596 26522
rect 14844 26382 14872 26726
rect 15118 26684 15426 26704
rect 15118 26682 15124 26684
rect 15180 26682 15204 26684
rect 15260 26682 15284 26684
rect 15340 26682 15364 26684
rect 15420 26682 15426 26684
rect 15180 26630 15182 26682
rect 15362 26630 15364 26682
rect 15118 26628 15124 26630
rect 15180 26628 15204 26630
rect 15260 26628 15284 26630
rect 15340 26628 15364 26630
rect 15420 26628 15426 26630
rect 15118 26608 15426 26628
rect 14924 26512 14976 26518
rect 14924 26454 14976 26460
rect 15016 26512 15068 26518
rect 15016 26454 15068 26460
rect 14832 26376 14884 26382
rect 14832 26318 14884 26324
rect 14556 26308 14608 26314
rect 14556 26250 14608 26256
rect 14464 26240 14516 26246
rect 14464 26182 14516 26188
rect 14476 25906 14504 26182
rect 14464 25900 14516 25906
rect 14464 25842 14516 25848
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 14568 25770 14596 26250
rect 14740 26240 14792 26246
rect 14740 26182 14792 26188
rect 14752 25906 14780 26182
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 14832 25832 14884 25838
rect 14832 25774 14884 25780
rect 14556 25764 14608 25770
rect 14556 25706 14608 25712
rect 14372 25696 14424 25702
rect 14372 25638 14424 25644
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14292 24562 14320 25230
rect 14384 24886 14412 25638
rect 14740 25492 14792 25498
rect 14844 25480 14872 25774
rect 14936 25498 14964 26454
rect 15028 25906 15056 26454
rect 15488 26382 15516 26726
rect 15476 26376 15528 26382
rect 15476 26318 15528 26324
rect 15566 26344 15622 26353
rect 15672 26314 15700 27406
rect 15764 27062 15792 27814
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 15752 26852 15804 26858
rect 15752 26794 15804 26800
rect 15764 26586 15792 26794
rect 15752 26580 15804 26586
rect 15752 26522 15804 26528
rect 15566 26279 15622 26288
rect 15660 26308 15712 26314
rect 15580 26042 15608 26279
rect 15660 26250 15712 26256
rect 15764 26058 15792 26522
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 15672 26030 15792 26058
rect 15476 25968 15528 25974
rect 15672 25922 15700 26030
rect 15528 25916 15700 25922
rect 15476 25910 15700 25916
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 15108 25900 15160 25906
rect 15488 25894 15700 25910
rect 15752 25900 15804 25906
rect 15108 25842 15160 25848
rect 15752 25842 15804 25848
rect 15120 25786 15148 25842
rect 15028 25770 15148 25786
rect 15016 25764 15148 25770
rect 15068 25758 15148 25764
rect 15016 25706 15068 25712
rect 14792 25452 14872 25480
rect 14740 25434 14792 25440
rect 14844 25158 14872 25452
rect 14924 25492 14976 25498
rect 15028 25480 15056 25706
rect 15118 25596 15426 25616
rect 15118 25594 15124 25596
rect 15180 25594 15204 25596
rect 15260 25594 15284 25596
rect 15340 25594 15364 25596
rect 15420 25594 15426 25596
rect 15180 25542 15182 25594
rect 15362 25542 15364 25594
rect 15118 25540 15124 25542
rect 15180 25540 15204 25542
rect 15260 25540 15284 25542
rect 15340 25540 15364 25542
rect 15420 25540 15426 25542
rect 15118 25520 15426 25540
rect 15028 25452 15148 25480
rect 14924 25434 14976 25440
rect 15120 25226 15148 25452
rect 15568 25288 15620 25294
rect 15566 25256 15568 25265
rect 15620 25256 15622 25265
rect 15108 25220 15160 25226
rect 15764 25226 15792 25842
rect 15856 25265 15884 29446
rect 15936 29164 15988 29170
rect 15936 29106 15988 29112
rect 15948 28762 15976 29106
rect 15936 28756 15988 28762
rect 15936 28698 15988 28704
rect 16212 28688 16264 28694
rect 16212 28630 16264 28636
rect 15936 28416 15988 28422
rect 15936 28358 15988 28364
rect 15948 28150 15976 28358
rect 15936 28144 15988 28150
rect 15936 28086 15988 28092
rect 16028 26988 16080 26994
rect 16028 26930 16080 26936
rect 15842 25256 15898 25265
rect 15566 25191 15622 25200
rect 15752 25220 15804 25226
rect 15108 25162 15160 25168
rect 14648 25152 14700 25158
rect 14648 25094 14700 25100
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 15120 25106 15148 25162
rect 14660 24886 14688 25094
rect 14372 24880 14424 24886
rect 14372 24822 14424 24828
rect 14648 24880 14700 24886
rect 14648 24822 14700 24828
rect 14844 24818 14872 25094
rect 15120 25078 15332 25106
rect 15304 24886 15332 25078
rect 15292 24880 15344 24886
rect 15292 24822 15344 24828
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14372 24608 14424 24614
rect 14292 24556 14372 24562
rect 14292 24550 14424 24556
rect 14292 24534 14412 24550
rect 14096 21344 14148 21350
rect 14016 21292 14096 21298
rect 14016 21286 14148 21292
rect 14016 21270 14136 21286
rect 13820 21140 13872 21146
rect 13872 21100 13952 21128
rect 13820 21082 13872 21088
rect 13924 20534 13952 21100
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 14016 20346 14044 21270
rect 14096 20868 14148 20874
rect 14096 20810 14148 20816
rect 14108 20466 14136 20810
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 13924 20318 14044 20346
rect 14094 20360 14150 20369
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13832 19417 13860 19994
rect 13818 19408 13874 19417
rect 13818 19343 13874 19352
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13556 18584 13676 18612
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13266 17776 13322 17785
rect 13266 17711 13322 17720
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 13082 17368 13138 17377
rect 13082 17303 13138 17312
rect 13096 17202 13124 17303
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 13188 16658 13216 17546
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 16794 13308 17478
rect 13372 17202 13400 18022
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 12808 16584 12860 16590
rect 12636 16546 12808 16574
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 14074 11836 14214
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11808 12850 11836 13330
rect 11900 13258 11928 13874
rect 11992 13802 12020 14962
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12084 13938 12112 14010
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11992 13462 12020 13738
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11808 12434 11836 12786
rect 11428 12174 11480 12180
rect 11532 12158 11652 12186
rect 11716 12406 11836 12434
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11256 11286 11284 11494
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10980 10526 11192 10554
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 10796 9676 10916 9704
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9956 8560 10008 8566
rect 9692 8508 9956 8514
rect 9692 8502 10008 8508
rect 9692 8498 9996 8502
rect 9680 8492 9996 8498
rect 9732 8486 9996 8492
rect 10336 8480 10364 9522
rect 10796 9058 10824 9676
rect 11072 9602 11100 9930
rect 10888 9586 11100 9602
rect 10876 9580 11100 9586
rect 10928 9574 11100 9580
rect 10876 9522 10928 9528
rect 10888 9450 10916 9522
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10704 9042 10824 9058
rect 10692 9036 10824 9042
rect 10744 9030 10824 9036
rect 10692 8978 10744 8984
rect 10395 8732 10703 8752
rect 10395 8730 10401 8732
rect 10457 8730 10481 8732
rect 10537 8730 10561 8732
rect 10617 8730 10641 8732
rect 10697 8730 10703 8732
rect 10457 8678 10459 8730
rect 10639 8678 10641 8730
rect 10395 8676 10401 8678
rect 10457 8676 10481 8678
rect 10537 8676 10561 8678
rect 10617 8676 10641 8678
rect 10697 8676 10703 8678
rect 10395 8656 10703 8676
rect 10692 8492 10744 8498
rect 10336 8452 10692 8480
rect 9680 8434 9732 8440
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9600 7342 9628 8230
rect 10244 7750 10272 8366
rect 10520 8362 10548 8452
rect 10796 8480 10824 9030
rect 10980 8838 11008 9386
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10876 8492 10928 8498
rect 10796 8452 10876 8480
rect 10692 8434 10744 8440
rect 10876 8434 10928 8440
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10336 7818 10364 8230
rect 11072 7954 11100 9318
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 9324 7296 9444 7324
rect 9588 7336 9640 7342
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8864 6322 8892 6666
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 9232 5166 9260 6598
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8772 4622 8800 4966
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8944 4548 8996 4554
rect 8944 4490 8996 4496
rect 8956 4282 8984 4490
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 9232 3738 9260 5102
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 9048 3058 9076 3402
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 9048 870 9168 898
rect 9048 800 9076 870
rect 3330 776 3386 785
rect 3330 711 3386 720
rect 4158 0 4214 800
rect 5446 0 5502 800
rect 6642 0 6698 800
rect 7838 0 7894 800
rect 9034 0 9090 800
rect 9140 762 9168 870
rect 9324 762 9352 7296
rect 9588 7278 9640 7284
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9416 5914 9444 6258
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9508 5574 9536 6734
rect 10244 6458 10272 7686
rect 10395 7644 10703 7664
rect 10395 7642 10401 7644
rect 10457 7642 10481 7644
rect 10537 7642 10561 7644
rect 10617 7642 10641 7644
rect 10697 7642 10703 7644
rect 10457 7590 10459 7642
rect 10639 7590 10641 7642
rect 10395 7588 10401 7590
rect 10457 7588 10481 7590
rect 10537 7588 10561 7590
rect 10617 7588 10641 7590
rect 10697 7588 10703 7590
rect 10395 7568 10703 7588
rect 11072 7206 11100 7890
rect 11164 7546 11192 10526
rect 11532 9586 11560 12158
rect 11612 12096 11664 12102
rect 11716 12084 11744 12406
rect 11664 12056 11744 12084
rect 11612 12038 11664 12044
rect 11624 11830 11652 12038
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11992 11762 12020 13398
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12084 12850 12112 13262
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12268 12850 12296 13194
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12084 12306 12112 12786
rect 12360 12782 12388 12922
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12452 12238 12480 16458
rect 12636 15706 12664 16546
rect 12808 16526 12860 16532
rect 13360 16584 13412 16590
rect 13464 16574 13492 17818
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13556 17338 13584 17682
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13556 16794 13584 17138
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13544 16584 13596 16590
rect 13412 16546 13544 16574
rect 13360 16526 13412 16532
rect 13544 16526 13596 16532
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13280 15910 13308 16458
rect 13372 15978 13400 16526
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12544 15026 12572 15370
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12544 14634 12572 14962
rect 12636 14822 12664 15098
rect 13280 15094 13308 15846
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12544 14606 12664 14634
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12544 13462 12572 14214
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12544 12986 12572 13126
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 11218 11652 11494
rect 11992 11354 12020 11698
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12360 11286 12388 11698
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 9042 11284 9318
rect 11532 9178 11560 9522
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 7818 11376 8298
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5778 9812 6054
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9416 4282 9444 4422
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9508 4214 9536 5034
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9876 4146 9904 5714
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9416 2650 9444 3674
rect 9600 3670 9628 4014
rect 9588 3664 9640 3670
rect 9588 3606 9640 3612
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9600 2650 9628 2994
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9968 2446 9996 3334
rect 10152 3058 10180 4082
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2514 10088 2790
rect 10152 2514 10180 2994
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10336 800 10364 6938
rect 10395 6556 10703 6576
rect 10395 6554 10401 6556
rect 10457 6554 10481 6556
rect 10537 6554 10561 6556
rect 10617 6554 10641 6556
rect 10697 6554 10703 6556
rect 10457 6502 10459 6554
rect 10639 6502 10641 6554
rect 10395 6500 10401 6502
rect 10457 6500 10481 6502
rect 10537 6500 10561 6502
rect 10617 6500 10641 6502
rect 10697 6500 10703 6502
rect 10395 6480 10703 6500
rect 11072 6390 11100 7142
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 10395 5468 10703 5488
rect 10395 5466 10401 5468
rect 10457 5466 10481 5468
rect 10537 5466 10561 5468
rect 10617 5466 10641 5468
rect 10697 5466 10703 5468
rect 10457 5414 10459 5466
rect 10639 5414 10641 5466
rect 10395 5412 10401 5414
rect 10457 5412 10481 5414
rect 10537 5412 10561 5414
rect 10617 5412 10641 5414
rect 10697 5412 10703 5414
rect 10395 5392 10703 5412
rect 11164 5234 11192 6054
rect 11256 5710 11284 6598
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11256 5284 11284 5646
rect 11440 5370 11468 7482
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11256 5256 11376 5284
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11152 5228 11204 5234
rect 11348 5216 11376 5256
rect 11428 5228 11480 5234
rect 11204 5188 11284 5216
rect 11152 5170 11204 5176
rect 10612 4826 10640 5170
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10704 4622 10732 5102
rect 10888 4758 10916 5170
rect 10876 4752 10928 4758
rect 10876 4694 10928 4700
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 11072 4554 11100 5170
rect 11256 4622 11284 5188
rect 11348 5188 11428 5216
rect 11348 4690 11376 5188
rect 11428 5170 11480 5176
rect 11532 5166 11560 5646
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10395 4380 10703 4400
rect 10395 4378 10401 4380
rect 10457 4378 10481 4380
rect 10537 4378 10561 4380
rect 10617 4378 10641 4380
rect 10697 4378 10703 4380
rect 10457 4326 10459 4378
rect 10639 4326 10641 4378
rect 10395 4324 10401 4326
rect 10457 4324 10481 4326
rect 10537 4324 10561 4326
rect 10617 4324 10641 4326
rect 10697 4324 10703 4326
rect 10395 4304 10703 4324
rect 11072 3942 11100 4490
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4146 11192 4422
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11072 3670 11100 3878
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 11060 3528 11112 3534
rect 11164 3482 11192 4082
rect 11256 3602 11284 4150
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11112 3476 11192 3482
rect 11060 3470 11192 3476
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11072 3454 11192 3470
rect 10395 3292 10703 3312
rect 10395 3290 10401 3292
rect 10457 3290 10481 3292
rect 10537 3290 10561 3292
rect 10617 3290 10641 3292
rect 10697 3290 10703 3292
rect 10457 3238 10459 3290
rect 10639 3238 10641 3290
rect 10395 3236 10401 3238
rect 10457 3236 10481 3238
rect 10537 3236 10561 3238
rect 10617 3236 10641 3238
rect 10697 3236 10703 3238
rect 10395 3216 10703 3236
rect 11072 3194 11100 3454
rect 11532 3398 11560 3470
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11532 3126 11560 3334
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 11624 2774 11652 11154
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12360 10810 12388 11086
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12452 10674 12480 12174
rect 12636 12102 12664 14606
rect 12714 14104 12770 14113
rect 12714 14039 12770 14048
rect 12728 14006 12756 14039
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12820 13938 12848 14962
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13280 14482 13308 14894
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 13004 14074 13032 14282
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13188 14006 13216 14418
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12820 13326 12848 13874
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12820 12442 12848 13262
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12820 11830 12848 12378
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12912 11762 12940 12854
rect 13004 12782 13032 13398
rect 13280 12986 13308 14418
rect 13648 13988 13676 18584
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13832 17746 13860 18090
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13740 14113 13768 14282
rect 13726 14104 13782 14113
rect 13832 14074 13860 14350
rect 13726 14039 13782 14048
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13648 13960 13768 13988
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13556 12986 13584 13330
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 12990 12200 13046 12209
rect 12990 12135 12992 12144
rect 13044 12135 13046 12144
rect 12992 12106 13044 12112
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 13188 11558 13216 12038
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13004 11014 13032 11494
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11900 9518 11928 9590
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11796 9376 11848 9382
rect 11992 9353 12020 9862
rect 12176 9489 12204 10406
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12162 9480 12218 9489
rect 12162 9415 12218 9424
rect 11796 9318 11848 9324
rect 11978 9344 12034 9353
rect 11808 8906 11836 9318
rect 11978 9279 12034 9288
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11900 7818 11928 8230
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11992 7002 12020 9279
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12176 8566 12204 9046
rect 12268 8974 12296 10066
rect 12452 9674 12480 10406
rect 12728 9722 12756 10406
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13188 9722 13216 9930
rect 12716 9716 12768 9722
rect 12452 9646 12572 9674
rect 12716 9658 12768 9664
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 12544 9586 12572 9646
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12360 9353 12388 9522
rect 12544 9450 12572 9522
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12346 9344 12402 9353
rect 12346 9279 12402 9288
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12268 8634 12296 8910
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12268 7342 12296 8570
rect 12360 8566 12388 8842
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12544 8498 12572 9386
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12360 7886 12388 8366
rect 12544 8022 12572 8434
rect 12728 8430 12756 9658
rect 12900 9512 12952 9518
rect 12898 9480 12900 9489
rect 12952 9480 12954 9489
rect 13372 9450 13400 9930
rect 13648 9586 13676 10406
rect 13740 9722 13768 13960
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13832 13802 13860 13874
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13924 11914 13952 20318
rect 14094 20295 14150 20304
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14016 18290 14044 19450
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 14016 17338 14044 17614
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14016 12442 14044 12786
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 13924 11886 14044 11914
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13832 10266 13860 11630
rect 13924 11354 13952 11766
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13924 9518 13952 11154
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 12898 9415 12954 9424
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 14016 9178 14044 11886
rect 14108 10266 14136 20295
rect 14200 18766 14228 20402
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14200 18426 14228 18702
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14186 17912 14242 17921
rect 14186 17847 14242 17856
rect 14200 17814 14228 17847
rect 14188 17808 14240 17814
rect 14188 17750 14240 17756
rect 14292 17218 14320 24534
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 14384 23322 14412 24142
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14568 23798 14596 24006
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14752 21622 14780 22374
rect 14740 21616 14792 21622
rect 14740 21558 14792 21564
rect 14556 20936 14608 20942
rect 14476 20896 14556 20924
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14384 19922 14412 20334
rect 14372 19916 14424 19922
rect 14372 19858 14424 19864
rect 14384 19514 14412 19858
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14476 18748 14504 20896
rect 14556 20878 14608 20884
rect 14844 20534 14872 24754
rect 15118 24508 15426 24528
rect 15118 24506 15124 24508
rect 15180 24506 15204 24508
rect 15260 24506 15284 24508
rect 15340 24506 15364 24508
rect 15420 24506 15426 24508
rect 15180 24454 15182 24506
rect 15362 24454 15364 24506
rect 15118 24452 15124 24454
rect 15180 24452 15204 24454
rect 15260 24452 15284 24454
rect 15340 24452 15364 24454
rect 15420 24452 15426 24454
rect 15118 24432 15426 24452
rect 15580 24410 15608 25191
rect 15842 25191 15898 25200
rect 15752 25162 15804 25168
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15856 24410 15884 24550
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15118 23420 15426 23440
rect 15118 23418 15124 23420
rect 15180 23418 15204 23420
rect 15260 23418 15284 23420
rect 15340 23418 15364 23420
rect 15420 23418 15426 23420
rect 15180 23366 15182 23418
rect 15362 23366 15364 23418
rect 15118 23364 15124 23366
rect 15180 23364 15204 23366
rect 15260 23364 15284 23366
rect 15340 23364 15364 23366
rect 15420 23364 15426 23366
rect 15118 23344 15426 23364
rect 15488 23186 15516 23462
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 15120 22642 15148 23054
rect 15304 22710 15332 23054
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15118 22332 15426 22352
rect 15118 22330 15124 22332
rect 15180 22330 15204 22332
rect 15260 22330 15284 22332
rect 15340 22330 15364 22332
rect 15420 22330 15426 22332
rect 15180 22278 15182 22330
rect 15362 22278 15364 22330
rect 15118 22276 15124 22278
rect 15180 22276 15204 22278
rect 15260 22276 15284 22278
rect 15340 22276 15364 22278
rect 15420 22276 15426 22278
rect 15118 22256 15426 22276
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 14924 21956 14976 21962
rect 14924 21898 14976 21904
rect 14936 21486 14964 21898
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 14936 21078 14964 21422
rect 14924 21072 14976 21078
rect 14924 21014 14976 21020
rect 14832 20528 14884 20534
rect 14832 20470 14884 20476
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14556 20256 14608 20262
rect 14556 20198 14608 20204
rect 14568 19854 14596 20198
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14660 19378 14688 20334
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14660 18834 14688 19314
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14556 18760 14608 18766
rect 14476 18720 14556 18748
rect 14384 18290 14412 18702
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14200 17190 14320 17218
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12636 7478 12664 8230
rect 13004 7886 13032 9114
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 13096 8090 13124 8366
rect 13740 8090 13768 8910
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13832 8566 13860 8774
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 13188 7886 13216 7958
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13372 7750 13400 7890
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 7478 13584 7686
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 14016 7206 14044 8842
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11900 6390 11928 6734
rect 12084 6458 12112 6802
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12268 6458 12296 6598
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 11716 6118 11744 6258
rect 12176 6118 12204 6258
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 11716 5370 11744 6054
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 12084 5234 12112 5578
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11808 3194 11836 3402
rect 12176 3194 12204 3878
rect 12360 3398 12388 6190
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 5302 12664 5510
rect 12912 5370 12940 6258
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12728 4690 12756 5170
rect 13004 4826 13032 5646
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13188 5370 13216 5510
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13280 5234 13308 5510
rect 13832 5302 13860 5646
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13268 5228 13320 5234
rect 13188 5188 13268 5216
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 13188 4622 13216 5188
rect 13268 5170 13320 5176
rect 13820 5160 13872 5166
rect 13924 5114 13952 6802
rect 13872 5108 13952 5114
rect 13820 5102 13952 5108
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13832 5086 13952 5102
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13372 4622 13400 4966
rect 13556 4622 13584 5034
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12452 4214 12480 4490
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12728 3738 12756 3878
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12176 2774 12204 3130
rect 12360 3058 12388 3334
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 11532 2746 11652 2774
rect 12084 2746 12204 2774
rect 10395 2204 10703 2224
rect 10395 2202 10401 2204
rect 10457 2202 10481 2204
rect 10537 2202 10561 2204
rect 10617 2202 10641 2204
rect 10697 2202 10703 2204
rect 10457 2150 10459 2202
rect 10639 2150 10641 2202
rect 10395 2148 10401 2150
rect 10457 2148 10481 2150
rect 10537 2148 10561 2150
rect 10617 2148 10641 2150
rect 10697 2148 10703 2150
rect 10395 2128 10703 2148
rect 11532 800 11560 2746
rect 12084 2446 12112 2746
rect 12728 2650 12756 2994
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12820 1986 12848 3946
rect 13188 3738 13216 4082
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13280 3534 13308 4422
rect 13372 3602 13400 4558
rect 13556 4282 13584 4558
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13556 3670 13584 4082
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13740 3602 13768 4082
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13280 3194 13308 3334
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13372 2650 13400 3538
rect 13832 3466 13860 5086
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 13832 3058 13860 3402
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13648 2446 13676 2994
rect 14200 2774 14228 17190
rect 14476 16454 14504 18720
rect 14556 18702 14608 18708
rect 14660 18154 14688 18770
rect 14844 18698 14872 19314
rect 14832 18692 14884 18698
rect 14832 18634 14884 18640
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 14844 17882 14872 18090
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14660 17202 14688 17478
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14648 17060 14700 17066
rect 14648 17002 14700 17008
rect 14660 16794 14688 17002
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 14292 13938 14320 14486
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14292 12850 14320 13738
rect 14384 13530 14412 15982
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14292 11150 14320 12786
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14292 10674 14320 11086
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14476 10130 14504 16390
rect 14752 16182 14780 17070
rect 14844 16590 14872 17614
rect 14936 17377 14964 18022
rect 14922 17368 14978 17377
rect 15028 17338 15056 22170
rect 15488 22166 15516 22578
rect 15476 22160 15528 22166
rect 15476 22102 15528 22108
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15212 21690 15240 21966
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15476 21616 15528 21622
rect 15476 21558 15528 21564
rect 15488 21350 15516 21558
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15118 21244 15426 21264
rect 15118 21242 15124 21244
rect 15180 21242 15204 21244
rect 15260 21242 15284 21244
rect 15340 21242 15364 21244
rect 15420 21242 15426 21244
rect 15180 21190 15182 21242
rect 15362 21190 15364 21242
rect 15118 21188 15124 21190
rect 15180 21188 15204 21190
rect 15260 21188 15284 21190
rect 15340 21188 15364 21190
rect 15420 21188 15426 21190
rect 15118 21168 15426 21188
rect 15488 21128 15516 21286
rect 15304 21100 15516 21128
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15212 20466 15240 20878
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15304 20330 15332 21100
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15118 20156 15426 20176
rect 15118 20154 15124 20156
rect 15180 20154 15204 20156
rect 15260 20154 15284 20156
rect 15340 20154 15364 20156
rect 15420 20154 15426 20156
rect 15180 20102 15182 20154
rect 15362 20102 15364 20154
rect 15118 20100 15124 20102
rect 15180 20100 15204 20102
rect 15260 20100 15284 20102
rect 15340 20100 15364 20102
rect 15420 20100 15426 20102
rect 15118 20080 15426 20100
rect 15488 19786 15516 20742
rect 15580 20058 15608 23666
rect 15752 23656 15804 23662
rect 15752 23598 15804 23604
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15672 22438 15700 22714
rect 15660 22432 15712 22438
rect 15660 22374 15712 22380
rect 15672 21049 15700 22374
rect 15658 21040 15714 21049
rect 15658 20975 15714 20984
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15672 20466 15700 20878
rect 15764 20806 15792 23598
rect 15856 22642 15884 23666
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15856 21554 15884 22374
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15660 20324 15712 20330
rect 15660 20266 15712 20272
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15672 19938 15700 20266
rect 15764 20058 15792 20402
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15672 19910 15792 19938
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15118 19068 15426 19088
rect 15118 19066 15124 19068
rect 15180 19066 15204 19068
rect 15260 19066 15284 19068
rect 15340 19066 15364 19068
rect 15420 19066 15426 19068
rect 15180 19014 15182 19066
rect 15362 19014 15364 19066
rect 15118 19012 15124 19014
rect 15180 19012 15204 19014
rect 15260 19012 15284 19014
rect 15340 19012 15364 19014
rect 15420 19012 15426 19014
rect 15118 18992 15426 19012
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 15304 18290 15332 18566
rect 15488 18358 15516 18702
rect 15580 18630 15608 19790
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15476 18352 15528 18358
rect 15476 18294 15528 18300
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15118 17980 15426 18000
rect 15118 17978 15124 17980
rect 15180 17978 15204 17980
rect 15260 17978 15284 17980
rect 15340 17978 15364 17980
rect 15420 17978 15426 17980
rect 15180 17926 15182 17978
rect 15362 17926 15364 17978
rect 15118 17924 15124 17926
rect 15180 17924 15204 17926
rect 15260 17924 15284 17926
rect 15340 17924 15364 17926
rect 15420 17924 15426 17926
rect 15118 17904 15426 17924
rect 15672 17746 15700 18702
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15764 17626 15792 19910
rect 15856 19378 15884 21490
rect 15948 20398 15976 21898
rect 16040 21894 16068 26930
rect 16120 24880 16172 24886
rect 16120 24822 16172 24828
rect 16028 21888 16080 21894
rect 16028 21830 16080 21836
rect 16132 21418 16160 24822
rect 16120 21412 16172 21418
rect 16120 21354 16172 21360
rect 16132 21026 16160 21354
rect 16224 21350 16252 28630
rect 16396 28076 16448 28082
rect 16396 28018 16448 28024
rect 16304 27668 16356 27674
rect 16304 27610 16356 27616
rect 16316 27130 16344 27610
rect 16304 27124 16356 27130
rect 16304 27066 16356 27072
rect 16408 26586 16436 28018
rect 16592 28014 16620 31889
rect 17040 29844 17092 29850
rect 17040 29786 17092 29792
rect 17052 28762 17080 29786
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17040 28756 17092 28762
rect 17040 28698 17092 28704
rect 17420 28694 17448 29106
rect 17408 28688 17460 28694
rect 17880 28642 17908 31889
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 17960 29708 18012 29714
rect 17960 29650 18012 29656
rect 17408 28630 17460 28636
rect 17788 28614 17908 28642
rect 16580 28008 16632 28014
rect 16580 27950 16632 27956
rect 17592 28008 17644 28014
rect 17592 27950 17644 27956
rect 17224 27668 17276 27674
rect 17224 27610 17276 27616
rect 16672 27396 16724 27402
rect 16672 27338 16724 27344
rect 16684 26994 16712 27338
rect 16856 27328 16908 27334
rect 16856 27270 16908 27276
rect 16672 26988 16724 26994
rect 16672 26930 16724 26936
rect 16764 26988 16816 26994
rect 16868 26976 16896 27270
rect 17236 26994 17264 27610
rect 17406 27024 17462 27033
rect 16816 26948 16896 26976
rect 16764 26930 16816 26936
rect 16488 26784 16540 26790
rect 16488 26726 16540 26732
rect 16396 26580 16448 26586
rect 16396 26522 16448 26528
rect 16500 26450 16528 26726
rect 16868 26450 16896 26948
rect 17224 26988 17276 26994
rect 17406 26959 17408 26968
rect 17224 26930 17276 26936
rect 17460 26959 17462 26968
rect 17408 26930 17460 26936
rect 17040 26920 17092 26926
rect 17040 26862 17092 26868
rect 17132 26920 17184 26926
rect 17132 26862 17184 26868
rect 16488 26444 16540 26450
rect 16488 26386 16540 26392
rect 16856 26444 16908 26450
rect 16856 26386 16908 26392
rect 17052 25974 17080 26862
rect 17144 26042 17172 26862
rect 17224 26444 17276 26450
rect 17224 26386 17276 26392
rect 17132 26036 17184 26042
rect 17132 25978 17184 25984
rect 17040 25968 17092 25974
rect 17040 25910 17092 25916
rect 16764 25696 16816 25702
rect 16764 25638 16816 25644
rect 16776 25362 16804 25638
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 17132 25356 17184 25362
rect 17236 25344 17264 26386
rect 17316 26376 17368 26382
rect 17316 26318 17368 26324
rect 17184 25316 17264 25344
rect 17132 25298 17184 25304
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 16316 24614 16344 25230
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 16304 24608 16356 24614
rect 16304 24550 16356 24556
rect 16316 23730 16344 24550
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16304 23724 16356 23730
rect 16304 23666 16356 23672
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 16684 23050 16712 23462
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16488 22092 16540 22098
rect 16488 22034 16540 22040
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 16132 20998 16252 21026
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15580 17598 15792 17626
rect 14922 17303 14978 17312
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 15028 16794 15056 17274
rect 15118 16892 15426 16912
rect 15118 16890 15124 16892
rect 15180 16890 15204 16892
rect 15260 16890 15284 16892
rect 15340 16890 15364 16892
rect 15420 16890 15426 16892
rect 15180 16838 15182 16890
rect 15362 16838 15364 16890
rect 15118 16836 15124 16838
rect 15180 16836 15204 16838
rect 15260 16836 15284 16838
rect 15340 16836 15364 16838
rect 15420 16836 15426 16838
rect 15118 16816 15426 16836
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14648 16176 14700 16182
rect 14648 16118 14700 16124
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 14660 15706 14688 16118
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14936 15502 14964 15846
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14936 14906 14964 14962
rect 14752 14878 14964 14906
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14648 13184 14700 13190
rect 14752 13172 14780 14878
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 13870 14964 14214
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14832 13320 14884 13326
rect 14936 13308 14964 13806
rect 14884 13280 14964 13308
rect 14832 13262 14884 13268
rect 14752 13144 14872 13172
rect 14648 13126 14700 13132
rect 14568 12918 14596 13126
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14568 12238 14596 12582
rect 14660 12434 14688 13126
rect 14660 12406 14780 12434
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14568 11014 14596 11494
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14384 9722 14412 9998
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14278 7984 14334 7993
rect 14278 7919 14280 7928
rect 14332 7919 14334 7928
rect 14280 7890 14332 7896
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14476 6390 14504 6598
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 14568 6118 14596 10950
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14660 9382 14688 10066
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14660 8498 14688 9318
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14752 7970 14780 12406
rect 14844 12238 14872 13144
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14844 11762 14872 12174
rect 15028 11898 15056 16730
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 16046 15516 16594
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15118 15804 15426 15824
rect 15118 15802 15124 15804
rect 15180 15802 15204 15804
rect 15260 15802 15284 15804
rect 15340 15802 15364 15804
rect 15420 15802 15426 15804
rect 15180 15750 15182 15802
rect 15362 15750 15364 15802
rect 15118 15748 15124 15750
rect 15180 15748 15204 15750
rect 15260 15748 15284 15750
rect 15340 15748 15364 15750
rect 15420 15748 15426 15750
rect 15118 15728 15426 15748
rect 15580 15026 15608 17598
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15672 16522 15700 17070
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15856 16114 15884 19314
rect 15936 18760 15988 18766
rect 16040 18748 16068 20402
rect 16132 20330 16160 20810
rect 16120 20324 16172 20330
rect 16120 20266 16172 20272
rect 16132 19854 16160 20266
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16224 19310 16252 20998
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16316 20262 16344 20402
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 15988 18720 16068 18748
rect 16120 18760 16172 18766
rect 15936 18702 15988 18708
rect 16120 18702 16172 18708
rect 15948 17270 15976 18702
rect 16132 17796 16160 18702
rect 16224 18630 16252 19246
rect 16316 18766 16344 20198
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16316 17882 16344 18362
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16132 17768 16252 17796
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 16040 16250 16068 17614
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16132 16522 16160 17478
rect 16224 17377 16252 17768
rect 16210 17368 16266 17377
rect 16210 17303 16266 17312
rect 16224 17202 16252 17303
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16120 16516 16172 16522
rect 16120 16458 16172 16464
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16132 15094 16160 15438
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15118 14716 15426 14736
rect 15118 14714 15124 14716
rect 15180 14714 15204 14716
rect 15260 14714 15284 14716
rect 15340 14714 15364 14716
rect 15420 14714 15426 14716
rect 15180 14662 15182 14714
rect 15362 14662 15364 14714
rect 15118 14660 15124 14662
rect 15180 14660 15204 14662
rect 15260 14660 15284 14662
rect 15340 14660 15364 14662
rect 15420 14660 15426 14662
rect 15118 14640 15426 14660
rect 15580 14414 15608 14962
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15118 13628 15426 13648
rect 15118 13626 15124 13628
rect 15180 13626 15204 13628
rect 15260 13626 15284 13628
rect 15340 13626 15364 13628
rect 15420 13626 15426 13628
rect 15180 13574 15182 13626
rect 15362 13574 15364 13626
rect 15118 13572 15124 13574
rect 15180 13572 15204 13574
rect 15260 13572 15284 13574
rect 15340 13572 15364 13574
rect 15420 13572 15426 13574
rect 15118 13552 15426 13572
rect 15488 13326 15516 14010
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15580 13462 15608 13874
rect 16224 13870 16252 14282
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15118 12540 15426 12560
rect 15118 12538 15124 12540
rect 15180 12538 15204 12540
rect 15260 12538 15284 12540
rect 15340 12538 15364 12540
rect 15420 12538 15426 12540
rect 15180 12486 15182 12538
rect 15362 12486 15364 12538
rect 15118 12484 15124 12486
rect 15180 12484 15204 12486
rect 15260 12484 15284 12486
rect 15340 12484 15364 12486
rect 15420 12484 15426 12486
rect 15118 12464 15426 12484
rect 15488 12306 15516 13126
rect 15660 12368 15712 12374
rect 15658 12336 15660 12345
rect 15712 12336 15714 12345
rect 15476 12300 15528 12306
rect 15658 12271 15714 12280
rect 15476 12242 15528 12248
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15212 11898 15240 12174
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15488 11830 15516 12242
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14844 11150 14872 11698
rect 15118 11452 15426 11472
rect 15118 11450 15124 11452
rect 15180 11450 15204 11452
rect 15260 11450 15284 11452
rect 15340 11450 15364 11452
rect 15420 11450 15426 11452
rect 15180 11398 15182 11450
rect 15362 11398 15364 11450
rect 15118 11396 15124 11398
rect 15180 11396 15204 11398
rect 15260 11396 15284 11398
rect 15340 11396 15364 11398
rect 15420 11396 15426 11398
rect 15118 11376 15426 11396
rect 15488 11286 15516 11766
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15580 11218 15608 11630
rect 15672 11218 15700 12174
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 15948 11082 15976 11494
rect 16132 11354 16160 11562
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10674 15608 10950
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15118 10364 15426 10384
rect 15118 10362 15124 10364
rect 15180 10362 15204 10364
rect 15260 10362 15284 10364
rect 15340 10362 15364 10364
rect 15420 10362 15426 10364
rect 15180 10310 15182 10362
rect 15362 10310 15364 10362
rect 15118 10308 15124 10310
rect 15180 10308 15204 10310
rect 15260 10308 15284 10310
rect 15340 10308 15364 10310
rect 15420 10308 15426 10310
rect 15118 10288 15426 10308
rect 16316 10266 16344 17818
rect 16408 17610 16436 21626
rect 16500 18834 16528 22034
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16684 20262 16712 20742
rect 16776 20466 16804 22986
rect 16868 22710 16896 24142
rect 16856 22704 16908 22710
rect 16856 22646 16908 22652
rect 16856 21956 16908 21962
rect 16856 21898 16908 21904
rect 16868 21690 16896 21898
rect 16856 21684 16908 21690
rect 16856 21626 16908 21632
rect 16960 21146 16988 25094
rect 17052 24818 17080 25094
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 17144 23050 17172 25298
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 17328 20602 17356 26318
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17316 20596 17368 20602
rect 17316 20538 17368 20544
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16592 18086 16620 19994
rect 16776 19854 16804 20402
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17052 19990 17080 20198
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17236 18578 17264 19314
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17328 18698 17356 19110
rect 17316 18692 17368 18698
rect 17316 18634 17368 18640
rect 17236 18550 17356 18578
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16592 17746 16620 18022
rect 16776 17814 16804 18158
rect 16764 17808 16816 17814
rect 16764 17750 16816 17756
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16396 17604 16448 17610
rect 16396 17546 16448 17552
rect 16592 17202 16620 17682
rect 16776 17270 16804 17750
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16868 17134 16896 17614
rect 17236 17202 17264 17614
rect 17328 17542 17356 18550
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16592 14550 16620 17002
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16454 16712 16934
rect 17328 16590 17356 17478
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 17144 15366 17172 15506
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 16684 14822 16712 14962
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16960 14550 16988 14894
rect 17052 14618 17080 14962
rect 17144 14822 17172 15302
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 17236 14414 17264 16390
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17328 15162 17356 15370
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 16592 13326 16620 14350
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16868 13938 16896 14282
rect 17420 14090 17448 20742
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17328 14062 17448 14090
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16684 13394 16712 13670
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16396 11824 16448 11830
rect 16396 11766 16448 11772
rect 16408 11014 16436 11766
rect 16684 11694 16712 13330
rect 17144 13190 17172 13874
rect 17236 13462 17264 13874
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17052 12102 17080 12786
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17328 11898 17356 14062
rect 17512 12986 17540 20402
rect 17604 17882 17632 27950
rect 17788 27674 17816 28614
rect 17868 28552 17920 28558
rect 17972 28540 18000 29650
rect 18144 29504 18196 29510
rect 18144 29446 18196 29452
rect 18052 28756 18104 28762
rect 18052 28698 18104 28704
rect 18064 28558 18092 28698
rect 17920 28512 18000 28540
rect 18052 28552 18104 28558
rect 17868 28494 17920 28500
rect 18052 28494 18104 28500
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 17776 27668 17828 27674
rect 17776 27610 17828 27616
rect 17866 27432 17922 27441
rect 17866 27367 17868 27376
rect 17920 27367 17922 27376
rect 17868 27338 17920 27344
rect 17868 26240 17920 26246
rect 17868 26182 17920 26188
rect 17880 25498 17908 26182
rect 17868 25492 17920 25498
rect 17868 25434 17920 25440
rect 17868 24404 17920 24410
rect 17868 24346 17920 24352
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17788 23866 17816 24074
rect 17776 23860 17828 23866
rect 17776 23802 17828 23808
rect 17880 23730 17908 24346
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17972 21894 18000 28018
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 18064 24750 18092 27406
rect 18156 27334 18184 29446
rect 18616 29306 18644 30194
rect 18696 30184 18748 30190
rect 18696 30126 18748 30132
rect 18708 29782 18736 30126
rect 19064 30116 19116 30122
rect 19064 30058 19116 30064
rect 18696 29776 18748 29782
rect 18696 29718 18748 29724
rect 18604 29300 18656 29306
rect 18604 29242 18656 29248
rect 18236 29028 18288 29034
rect 18236 28970 18288 28976
rect 18248 28490 18276 28970
rect 18236 28484 18288 28490
rect 18236 28426 18288 28432
rect 18144 27328 18196 27334
rect 18144 27270 18196 27276
rect 18248 27146 18276 28426
rect 18328 28008 18380 28014
rect 18328 27950 18380 27956
rect 18340 27538 18368 27950
rect 18328 27532 18380 27538
rect 18328 27474 18380 27480
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 18156 27118 18276 27146
rect 18156 26382 18184 27118
rect 18432 26382 18460 27406
rect 18512 27056 18564 27062
rect 18512 26998 18564 27004
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 18156 25838 18184 26182
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 18156 24206 18184 25774
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 18064 23254 18092 23666
rect 18052 23248 18104 23254
rect 18052 23190 18104 23196
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17880 21706 17908 21830
rect 17880 21678 18000 21706
rect 17972 21010 18000 21678
rect 18052 21412 18104 21418
rect 18052 21354 18104 21360
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17972 20398 18000 20946
rect 18064 20874 18092 21354
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17972 19938 18000 20334
rect 17880 19922 18000 19938
rect 17868 19916 18000 19922
rect 17920 19910 18000 19916
rect 17868 19858 17920 19864
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17776 19780 17828 19786
rect 17776 19722 17828 19728
rect 17788 19378 17816 19722
rect 17972 19378 18000 19790
rect 18248 19514 18276 25094
rect 18328 24744 18380 24750
rect 18328 24686 18380 24692
rect 18340 24410 18368 24686
rect 18328 24404 18380 24410
rect 18328 24346 18380 24352
rect 18328 23724 18380 23730
rect 18328 23666 18380 23672
rect 18340 23594 18368 23666
rect 18328 23588 18380 23594
rect 18328 23530 18380 23536
rect 18432 23118 18460 26318
rect 18524 23322 18552 26998
rect 18616 26926 18644 29242
rect 18708 28626 18736 29718
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 18696 28620 18748 28626
rect 18696 28562 18748 28568
rect 18708 27606 18736 28562
rect 18984 28558 19012 29582
rect 19076 29578 19104 30058
rect 19064 29572 19116 29578
rect 19064 29514 19116 29520
rect 18972 28552 19024 28558
rect 18972 28494 19024 28500
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 18696 27464 18748 27470
rect 18696 27406 18748 27412
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 18604 26920 18656 26926
rect 18604 26862 18656 26868
rect 18708 26858 18736 27406
rect 18788 27056 18840 27062
rect 18786 27024 18788 27033
rect 18840 27024 18842 27033
rect 18786 26959 18842 26968
rect 18696 26852 18748 26858
rect 18696 26794 18748 26800
rect 18880 26852 18932 26858
rect 18880 26794 18932 26800
rect 18708 26518 18736 26794
rect 18696 26512 18748 26518
rect 18696 26454 18748 26460
rect 18788 26512 18840 26518
rect 18788 26454 18840 26460
rect 18604 26444 18656 26450
rect 18604 26386 18656 26392
rect 18616 23730 18644 26386
rect 18696 26308 18748 26314
rect 18696 26250 18748 26256
rect 18708 24342 18736 26250
rect 18800 26042 18828 26454
rect 18892 26246 18920 26794
rect 18984 26450 19012 27406
rect 19076 27334 19104 29514
rect 19260 28966 19288 31889
rect 19616 30592 19668 30598
rect 19616 30534 19668 30540
rect 19628 30054 19656 30534
rect 19840 30492 20148 30512
rect 19840 30490 19846 30492
rect 19902 30490 19926 30492
rect 19982 30490 20006 30492
rect 20062 30490 20086 30492
rect 20142 30490 20148 30492
rect 19902 30438 19904 30490
rect 20084 30438 20086 30490
rect 19840 30436 19846 30438
rect 19902 30436 19926 30438
rect 19982 30436 20006 30438
rect 20062 30436 20086 30438
rect 20142 30436 20148 30438
rect 19840 30416 20148 30436
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19616 30048 19668 30054
rect 19616 29990 19668 29996
rect 19352 29170 19380 29990
rect 19628 29782 19656 29990
rect 19616 29776 19668 29782
rect 19616 29718 19668 29724
rect 20364 29714 20392 30194
rect 20548 30138 20576 31889
rect 20720 30252 20772 30258
rect 20720 30194 20772 30200
rect 20456 30110 20576 30138
rect 20352 29708 20404 29714
rect 20352 29650 20404 29656
rect 19840 29404 20148 29424
rect 19840 29402 19846 29404
rect 19902 29402 19926 29404
rect 19982 29402 20006 29404
rect 20062 29402 20086 29404
rect 20142 29402 20148 29404
rect 19902 29350 19904 29402
rect 20084 29350 20086 29402
rect 19840 29348 19846 29350
rect 19902 29348 19926 29350
rect 19982 29348 20006 29350
rect 20062 29348 20086 29350
rect 20142 29348 20148 29350
rect 19840 29328 20148 29348
rect 20364 29170 20392 29650
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 20260 29164 20312 29170
rect 20260 29106 20312 29112
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 19248 28960 19300 28966
rect 19248 28902 19300 28908
rect 19840 28316 20148 28336
rect 19840 28314 19846 28316
rect 19902 28314 19926 28316
rect 19982 28314 20006 28316
rect 20062 28314 20086 28316
rect 20142 28314 20148 28316
rect 19902 28262 19904 28314
rect 20084 28262 20086 28314
rect 19840 28260 19846 28262
rect 19902 28260 19926 28262
rect 19982 28260 20006 28262
rect 20062 28260 20086 28262
rect 20142 28260 20148 28262
rect 19840 28240 20148 28260
rect 19248 28212 19300 28218
rect 19248 28154 19300 28160
rect 19260 27470 19288 28154
rect 20272 28082 20300 29106
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 19444 27674 19472 28018
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 19708 27600 19760 27606
rect 19708 27542 19760 27548
rect 19248 27464 19300 27470
rect 19720 27441 19748 27542
rect 19248 27406 19300 27412
rect 19706 27432 19762 27441
rect 19706 27367 19762 27376
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 20168 27328 20220 27334
rect 20168 27270 20220 27276
rect 19352 27062 19380 27270
rect 19840 27228 20148 27248
rect 19840 27226 19846 27228
rect 19902 27226 19926 27228
rect 19982 27226 20006 27228
rect 20062 27226 20086 27228
rect 20142 27226 20148 27228
rect 19902 27174 19904 27226
rect 20084 27174 20086 27226
rect 19840 27172 19846 27174
rect 19902 27172 19926 27174
rect 19982 27172 20006 27174
rect 20062 27172 20086 27174
rect 20142 27172 20148 27174
rect 19840 27152 20148 27172
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 19064 26920 19116 26926
rect 19064 26862 19116 26868
rect 18972 26444 19024 26450
rect 18972 26386 19024 26392
rect 18880 26240 18932 26246
rect 18880 26182 18932 26188
rect 18788 26036 18840 26042
rect 18788 25978 18840 25984
rect 18800 25838 18828 25978
rect 18892 25838 18920 26182
rect 18788 25832 18840 25838
rect 18788 25774 18840 25780
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 19076 25650 19104 26862
rect 19168 26450 19196 26930
rect 19248 26920 19300 26926
rect 19248 26862 19300 26868
rect 19260 26518 19288 26862
rect 19248 26512 19300 26518
rect 19248 26454 19300 26460
rect 19156 26444 19208 26450
rect 19156 26386 19208 26392
rect 19352 25770 19380 26998
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 19536 26790 19564 26930
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19340 25764 19392 25770
rect 19340 25706 19392 25712
rect 18984 25622 19104 25650
rect 18984 24954 19012 25622
rect 19064 25492 19116 25498
rect 19064 25434 19116 25440
rect 18972 24948 19024 24954
rect 18972 24890 19024 24896
rect 18880 24880 18932 24886
rect 18880 24822 18932 24828
rect 18788 24744 18840 24750
rect 18788 24686 18840 24692
rect 18696 24336 18748 24342
rect 18696 24278 18748 24284
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18512 23316 18564 23322
rect 18512 23258 18564 23264
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17682 17912 17738 17921
rect 17592 17876 17644 17882
rect 17682 17847 17738 17856
rect 17592 17818 17644 17824
rect 17696 17814 17724 17847
rect 17684 17808 17736 17814
rect 17684 17750 17736 17756
rect 17592 16176 17644 16182
rect 17592 16118 17644 16124
rect 17604 15706 17632 16118
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17604 15026 17632 15642
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17696 14482 17724 17750
rect 17972 17202 18000 19314
rect 18236 19236 18288 19242
rect 18236 19178 18288 19184
rect 18248 18834 18276 19178
rect 18236 18828 18288 18834
rect 18236 18770 18288 18776
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17788 16590 17816 16934
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17684 14476 17736 14482
rect 17684 14418 17736 14424
rect 17788 14414 17816 16526
rect 18064 16114 18092 17274
rect 18156 17270 18184 17478
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18248 17202 18276 18770
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18248 16658 18276 17138
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 18340 16250 18368 21830
rect 18432 20466 18460 23054
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18524 22098 18552 22374
rect 18512 22092 18564 22098
rect 18512 22034 18564 22040
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18616 20448 18644 23666
rect 18800 23186 18828 24686
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 18694 23080 18750 23089
rect 18694 23015 18696 23024
rect 18748 23015 18750 23024
rect 18696 22986 18748 22992
rect 18708 22710 18736 22986
rect 18696 22704 18748 22710
rect 18696 22646 18748 22652
rect 18800 22098 18828 23122
rect 18788 22092 18840 22098
rect 18788 22034 18840 22040
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18696 20460 18748 20466
rect 18616 20420 18696 20448
rect 18432 20058 18460 20402
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18616 19718 18644 20420
rect 18696 20402 18748 20408
rect 18800 20262 18828 20878
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18432 18358 18460 18566
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18524 17678 18552 17818
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18432 16454 18460 17614
rect 18524 16726 18552 17614
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17604 13326 17632 14214
rect 17696 13394 17724 14214
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17604 12374 17632 13262
rect 17696 12442 17724 13330
rect 17880 13172 17908 15642
rect 17972 15434 18000 15846
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17972 15144 18000 15370
rect 17972 15116 18092 15144
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17972 13190 18000 14962
rect 18064 14414 18092 15116
rect 18156 14550 18184 15506
rect 18432 15502 18460 16050
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18340 15094 18368 15302
rect 18616 15162 18644 15370
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18328 14408 18380 14414
rect 18328 14350 18380 14356
rect 18064 13326 18092 14350
rect 18340 14278 18368 14350
rect 18616 14346 18644 15098
rect 18604 14340 18656 14346
rect 18604 14282 18656 14288
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17788 13144 17908 13172
rect 17960 13184 18012 13190
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 17144 11354 17172 11698
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16408 10810 16436 10950
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14936 9722 14964 9998
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 15212 9654 15240 9930
rect 15200 9648 15252 9654
rect 14936 9586 15148 9602
rect 15200 9590 15252 9596
rect 14936 9580 15160 9586
rect 14936 9574 15108 9580
rect 14936 8634 14964 9574
rect 15108 9522 15160 9528
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15028 9178 15056 9454
rect 15118 9276 15426 9296
rect 15118 9274 15124 9276
rect 15180 9274 15204 9276
rect 15260 9274 15284 9276
rect 15340 9274 15364 9276
rect 15420 9274 15426 9276
rect 15180 9222 15182 9274
rect 15362 9222 15364 9274
rect 15118 9220 15124 9222
rect 15180 9220 15204 9222
rect 15260 9220 15284 9222
rect 15340 9220 15364 9222
rect 15420 9220 15426 9222
rect 15118 9200 15426 9220
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14844 8022 14872 8366
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14660 7942 14780 7970
rect 14832 8016 14884 8022
rect 14832 7958 14884 7964
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14384 5302 14412 6054
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14384 5166 14412 5238
rect 14568 5234 14596 5646
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14384 4554 14412 5102
rect 14476 4622 14504 5102
rect 14568 4758 14596 5170
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14660 4078 14688 7942
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14844 7698 14872 7958
rect 14936 7886 14964 8230
rect 15028 8090 15056 9114
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15212 8566 15240 8774
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15396 8498 15424 9046
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15488 8294 15516 10066
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15856 9586 15884 9998
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15856 8838 15884 9522
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15118 8188 15426 8208
rect 15118 8186 15124 8188
rect 15180 8186 15204 8188
rect 15260 8186 15284 8188
rect 15340 8186 15364 8188
rect 15420 8186 15426 8188
rect 15180 8134 15182 8186
rect 15362 8134 15364 8186
rect 15118 8132 15124 8134
rect 15180 8132 15204 8134
rect 15260 8132 15284 8134
rect 15340 8132 15364 8134
rect 15420 8132 15426 8134
rect 15118 8112 15426 8132
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15396 7818 15424 7958
rect 15488 7886 15516 8230
rect 15672 8090 15700 8434
rect 16224 8362 16252 8570
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 14752 7546 14780 7686
rect 14844 7670 15056 7698
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 4758 14780 7142
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14844 5914 14872 6598
rect 14936 6458 14964 6598
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 15028 6338 15056 7670
rect 15118 7100 15426 7120
rect 15118 7098 15124 7100
rect 15180 7098 15204 7100
rect 15260 7098 15284 7100
rect 15340 7098 15364 7100
rect 15420 7098 15426 7100
rect 15180 7046 15182 7098
rect 15362 7046 15364 7098
rect 15118 7044 15124 7046
rect 15180 7044 15204 7046
rect 15260 7044 15284 7046
rect 15340 7044 15364 7046
rect 15420 7044 15426 7046
rect 15118 7024 15426 7044
rect 15672 7002 15700 8026
rect 15948 7886 15976 8298
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16408 7410 16436 7686
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 14936 6310 15056 6338
rect 15476 6316 15528 6322
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14016 2746 14228 2774
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 12728 1958 12848 1986
rect 12728 800 12756 1958
rect 14016 800 14044 2746
rect 14292 2650 14320 3470
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14476 2446 14504 3402
rect 14936 2990 14964 6310
rect 15476 6258 15528 6264
rect 15118 6012 15426 6032
rect 15118 6010 15124 6012
rect 15180 6010 15204 6012
rect 15260 6010 15284 6012
rect 15340 6010 15364 6012
rect 15420 6010 15426 6012
rect 15180 5958 15182 6010
rect 15362 5958 15364 6010
rect 15118 5956 15124 5958
rect 15180 5956 15204 5958
rect 15260 5956 15284 5958
rect 15340 5956 15364 5958
rect 15420 5956 15426 5958
rect 15118 5936 15426 5956
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15212 5370 15240 5646
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15304 5234 15332 5782
rect 15488 5710 15516 6258
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5846 15608 6054
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 15292 5228 15344 5234
rect 15344 5188 15516 5216
rect 15292 5170 15344 5176
rect 15028 4690 15056 5170
rect 15118 4924 15426 4944
rect 15118 4922 15124 4924
rect 15180 4922 15204 4924
rect 15260 4922 15284 4924
rect 15340 4922 15364 4924
rect 15420 4922 15426 4924
rect 15180 4870 15182 4922
rect 15362 4870 15364 4922
rect 15118 4868 15124 4870
rect 15180 4868 15204 4870
rect 15260 4868 15284 4870
rect 15340 4868 15364 4870
rect 15420 4868 15426 4870
rect 15118 4848 15426 4868
rect 15488 4826 15516 5188
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15856 4826 15884 5102
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 15028 3534 15056 3878
rect 15118 3836 15426 3856
rect 15118 3834 15124 3836
rect 15180 3834 15204 3836
rect 15260 3834 15284 3836
rect 15340 3834 15364 3836
rect 15420 3834 15426 3836
rect 15180 3782 15182 3834
rect 15362 3782 15364 3834
rect 15118 3780 15124 3782
rect 15180 3780 15204 3782
rect 15260 3780 15284 3782
rect 15340 3780 15364 3782
rect 15420 3780 15426 3782
rect 15118 3760 15426 3780
rect 15488 3738 15516 4490
rect 15660 4208 15712 4214
rect 16592 4162 16620 10406
rect 17144 9518 17172 10542
rect 17420 10470 17448 11086
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17144 8974 17172 9454
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16868 7886 16896 8774
rect 17144 8566 17172 8910
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16960 6798 16988 8366
rect 17052 8022 17080 8434
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17144 6798 17172 8502
rect 17328 8430 17356 9318
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17222 7984 17278 7993
rect 17222 7919 17224 7928
rect 17276 7919 17278 7928
rect 17224 7890 17276 7896
rect 17328 7750 17356 8366
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 16960 6322 16988 6734
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 15660 4150 15712 4156
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15580 3534 15608 4082
rect 15672 3602 15700 4150
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 16500 4134 16620 4162
rect 15764 3618 15792 4082
rect 15844 3664 15896 3670
rect 15764 3612 15844 3618
rect 15764 3606 15896 3612
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15764 3590 15884 3606
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15304 3194 15332 3470
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15580 3126 15608 3470
rect 15764 3126 15792 3590
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 16040 3194 16068 3402
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15118 2748 15426 2768
rect 15118 2746 15124 2748
rect 15180 2746 15204 2748
rect 15260 2746 15284 2748
rect 15340 2746 15364 2748
rect 15420 2746 15426 2748
rect 15180 2694 15182 2746
rect 15362 2694 15364 2746
rect 15118 2692 15124 2694
rect 15180 2692 15204 2694
rect 15260 2692 15284 2694
rect 15340 2692 15364 2694
rect 15420 2692 15426 2694
rect 15118 2672 15426 2692
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 15212 870 15332 898
rect 15212 800 15240 870
rect 9140 734 9352 762
rect 10322 0 10378 800
rect 11518 0 11574 800
rect 12714 0 12770 800
rect 14002 0 14058 800
rect 15198 0 15254 800
rect 15304 762 15332 870
rect 15488 762 15516 2790
rect 16500 2774 16528 4134
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16592 3602 16620 4014
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16684 3058 16712 4558
rect 16960 4146 16988 6258
rect 17144 4622 17172 6734
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17420 4554 17448 4966
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16960 3126 16988 3334
rect 17144 3194 17172 3538
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 16948 3120 17000 3126
rect 16948 3062 17000 3068
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16408 2746 16528 2774
rect 16408 800 16436 2746
rect 17328 2650 17356 3470
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17420 2446 17448 3130
rect 17512 2774 17540 12038
rect 17604 11218 17632 12310
rect 17696 11286 17724 12378
rect 17788 12238 17816 13144
rect 17960 13126 18012 13132
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 18064 12238 18092 12310
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18156 12186 18184 14214
rect 18708 14074 18736 19314
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18800 18902 18828 19246
rect 18788 18896 18840 18902
rect 18788 18838 18840 18844
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18800 18290 18828 18702
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18800 17338 18828 18226
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18892 16250 18920 24822
rect 18984 23798 19012 24890
rect 19076 24614 19104 25434
rect 19352 25226 19380 25706
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19444 25362 19472 25638
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19536 25294 19564 26726
rect 20180 26518 20208 27270
rect 20168 26512 20220 26518
rect 20168 26454 20220 26460
rect 19616 26308 19668 26314
rect 19616 26250 19668 26256
rect 19628 26042 19656 26250
rect 19840 26140 20148 26160
rect 19840 26138 19846 26140
rect 19902 26138 19926 26140
rect 19982 26138 20006 26140
rect 20062 26138 20086 26140
rect 20142 26138 20148 26140
rect 19902 26086 19904 26138
rect 20084 26086 20086 26138
rect 19840 26084 19846 26086
rect 19902 26084 19926 26086
rect 19982 26084 20006 26086
rect 20062 26084 20086 26086
rect 20142 26084 20148 26086
rect 19840 26064 20148 26084
rect 19616 26036 19668 26042
rect 19616 25978 19668 25984
rect 20272 25974 20300 28018
rect 20352 27328 20404 27334
rect 20352 27270 20404 27276
rect 20260 25968 20312 25974
rect 20260 25910 20312 25916
rect 20272 25362 20300 25910
rect 20260 25356 20312 25362
rect 20260 25298 20312 25304
rect 20364 25294 20392 27270
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 20352 25288 20404 25294
rect 20352 25230 20404 25236
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 19524 25152 19576 25158
rect 19708 25152 19760 25158
rect 19524 25094 19576 25100
rect 19706 25120 19708 25129
rect 19760 25120 19762 25129
rect 19156 24676 19208 24682
rect 19156 24618 19208 24624
rect 19248 24676 19300 24682
rect 19248 24618 19300 24624
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 19168 23866 19196 24618
rect 19260 24342 19288 24618
rect 19248 24336 19300 24342
rect 19248 24278 19300 24284
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 18972 23792 19024 23798
rect 18972 23734 19024 23740
rect 19156 23724 19208 23730
rect 19208 23684 19288 23712
rect 19156 23666 19208 23672
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 18972 23588 19024 23594
rect 18972 23530 19024 23536
rect 18984 23254 19012 23530
rect 19076 23526 19104 23598
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 18972 23248 19024 23254
rect 18972 23190 19024 23196
rect 18984 22642 19012 23190
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18984 21962 19012 22578
rect 19076 22574 19104 23462
rect 19260 22624 19288 23684
rect 19168 22596 19288 22624
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 19076 22098 19104 22510
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 19168 22030 19196 22596
rect 19248 22500 19300 22506
rect 19248 22442 19300 22448
rect 19156 22024 19208 22030
rect 19156 21966 19208 21972
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 19260 21418 19288 22442
rect 19352 22234 19380 24006
rect 19340 22228 19392 22234
rect 19392 22188 19472 22216
rect 19340 22170 19392 22176
rect 19340 22024 19392 22030
rect 19338 21992 19340 22001
rect 19392 21992 19394 22001
rect 19338 21927 19394 21936
rect 19352 21894 19380 21927
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19444 21690 19472 22188
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 19432 21412 19484 21418
rect 19432 21354 19484 21360
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18984 19310 19012 20334
rect 19076 20330 19104 20946
rect 19260 20466 19288 21354
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19064 20324 19116 20330
rect 19064 20266 19116 20272
rect 19260 19378 19288 20402
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18984 18834 19012 19246
rect 19260 18970 19288 19314
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 19352 18154 19380 20878
rect 19444 18698 19472 21354
rect 19536 18970 19564 25094
rect 19706 25055 19762 25064
rect 19840 25052 20148 25072
rect 19840 25050 19846 25052
rect 19902 25050 19926 25052
rect 19982 25050 20006 25052
rect 20062 25050 20086 25052
rect 20142 25050 20148 25052
rect 19902 24998 19904 25050
rect 20084 24998 20086 25050
rect 19840 24996 19846 24998
rect 19902 24996 19926 24998
rect 19982 24996 20006 24998
rect 20062 24996 20086 24998
rect 20142 24996 20148 24998
rect 19840 24976 20148 24996
rect 20260 24880 20312 24886
rect 20260 24822 20312 24828
rect 19708 24744 19760 24750
rect 19708 24686 19760 24692
rect 19720 24410 19748 24686
rect 19708 24404 19760 24410
rect 19708 24346 19760 24352
rect 19720 23848 19748 24346
rect 20168 24132 20220 24138
rect 20168 24074 20220 24080
rect 19840 23964 20148 23984
rect 19840 23962 19846 23964
rect 19902 23962 19926 23964
rect 19982 23962 20006 23964
rect 20062 23962 20086 23964
rect 20142 23962 20148 23964
rect 19902 23910 19904 23962
rect 20084 23910 20086 23962
rect 19840 23908 19846 23910
rect 19902 23908 19926 23910
rect 19982 23908 20006 23910
rect 20062 23908 20086 23910
rect 20142 23908 20148 23910
rect 19840 23888 20148 23908
rect 20180 23866 20208 24074
rect 20168 23860 20220 23866
rect 19720 23820 19932 23848
rect 19904 23730 19932 23820
rect 20168 23802 20220 23808
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19616 22976 19668 22982
rect 19616 22918 19668 22924
rect 19708 22976 19760 22982
rect 19708 22918 19760 22924
rect 19628 20942 19656 22918
rect 19720 22778 19748 22918
rect 19840 22876 20148 22896
rect 19840 22874 19846 22876
rect 19902 22874 19926 22876
rect 19982 22874 20006 22876
rect 20062 22874 20086 22876
rect 20142 22874 20148 22876
rect 19902 22822 19904 22874
rect 20084 22822 20086 22874
rect 19840 22820 19846 22822
rect 19902 22820 19926 22822
rect 19982 22820 20006 22822
rect 20062 22820 20086 22822
rect 20142 22820 20148 22822
rect 19840 22800 20148 22820
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19720 22030 19748 22714
rect 20272 22094 20300 24822
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20364 23866 20392 24142
rect 20352 23860 20404 23866
rect 20352 23802 20404 23808
rect 20180 22066 20300 22094
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19840 21788 20148 21808
rect 19840 21786 19846 21788
rect 19902 21786 19926 21788
rect 19982 21786 20006 21788
rect 20062 21786 20086 21788
rect 20142 21786 20148 21788
rect 19902 21734 19904 21786
rect 20084 21734 20086 21786
rect 19840 21732 19846 21734
rect 19902 21732 19926 21734
rect 19982 21732 20006 21734
rect 20062 21732 20086 21734
rect 20142 21732 20148 21734
rect 19840 21712 20148 21732
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 19840 20700 20148 20720
rect 19840 20698 19846 20700
rect 19902 20698 19926 20700
rect 19982 20698 20006 20700
rect 20062 20698 20086 20700
rect 20142 20698 20148 20700
rect 19902 20646 19904 20698
rect 20084 20646 20086 20698
rect 19840 20644 19846 20646
rect 19902 20644 19926 20646
rect 19982 20644 20006 20646
rect 20062 20644 20086 20646
rect 20142 20644 20148 20646
rect 19840 20624 20148 20644
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19628 19310 19656 20266
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19720 19514 19748 19654
rect 19840 19612 20148 19632
rect 19840 19610 19846 19612
rect 19902 19610 19926 19612
rect 19982 19610 20006 19612
rect 20062 19610 20086 19612
rect 20142 19610 20148 19612
rect 19902 19558 19904 19610
rect 20084 19558 20086 19610
rect 19840 19556 19846 19558
rect 19902 19556 19926 19558
rect 19982 19556 20006 19558
rect 20062 19556 20086 19558
rect 20142 19556 20148 19558
rect 19840 19536 20148 19556
rect 19708 19508 19760 19514
rect 19708 19450 19760 19456
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19628 18850 19656 19246
rect 19904 19174 19932 19314
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19628 18834 19748 18850
rect 19628 18828 19760 18834
rect 19628 18822 19708 18828
rect 19708 18770 19760 18776
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19444 17746 19472 18294
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19168 17270 19196 17682
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18880 16040 18932 16046
rect 18880 15982 18932 15988
rect 18800 15910 18828 15982
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18800 13802 18828 15846
rect 18892 15706 18920 15982
rect 19168 15910 19196 17206
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 19260 15570 19288 16050
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19260 15162 19288 15506
rect 19352 15162 19380 17478
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19444 16250 19472 16390
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19536 15586 19564 18702
rect 19904 18698 19932 19110
rect 20088 18970 20116 19382
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 19892 18692 19944 18698
rect 19892 18634 19944 18640
rect 19840 18524 20148 18544
rect 19840 18522 19846 18524
rect 19902 18522 19926 18524
rect 19982 18522 20006 18524
rect 20062 18522 20086 18524
rect 20142 18522 20148 18524
rect 19902 18470 19904 18522
rect 20084 18470 20086 18522
rect 19840 18468 19846 18470
rect 19902 18468 19926 18470
rect 19982 18468 20006 18470
rect 20062 18468 20086 18470
rect 20142 18468 20148 18470
rect 19840 18448 20148 18468
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19444 15558 19564 15586
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18984 14618 19012 14962
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 19352 14498 19380 15098
rect 19076 14470 19380 14498
rect 19076 14414 19104 14470
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19156 14408 19208 14414
rect 19340 14408 19392 14414
rect 19156 14350 19208 14356
rect 19338 14376 19340 14385
rect 19392 14376 19394 14385
rect 19168 14278 19196 14350
rect 19338 14311 19394 14320
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18524 13462 18552 13670
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18340 12374 18368 12922
rect 18420 12776 18472 12782
rect 18616 12764 18644 13738
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 18472 12736 18644 12764
rect 18420 12718 18472 12724
rect 18328 12368 18380 12374
rect 18328 12310 18380 12316
rect 17880 12102 17908 12174
rect 18156 12158 18368 12186
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17788 11626 17816 11834
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17696 11150 17724 11222
rect 17880 11150 17908 11630
rect 18156 11150 18184 12038
rect 18248 11898 18276 12038
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18340 11642 18368 12158
rect 18432 11694 18460 12718
rect 19260 12594 19288 13126
rect 19352 12918 19380 13126
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19260 12566 19380 12594
rect 18602 12336 18658 12345
rect 19352 12306 19380 12566
rect 18602 12271 18658 12280
rect 19248 12300 19300 12306
rect 18616 12170 18644 12271
rect 19248 12242 19300 12248
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18248 11614 18368 11642
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 17880 10810 17908 11086
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17972 10742 18000 10950
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 18248 9738 18276 11614
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18340 11150 18368 11494
rect 19260 11218 19288 12242
rect 19444 11898 19472 15558
rect 19628 14618 19656 18226
rect 19708 18148 19760 18154
rect 19708 18090 19760 18096
rect 19720 17814 19748 18090
rect 20180 17882 20208 22066
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20364 20602 20392 20742
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 20456 20466 20484 30110
rect 20536 30048 20588 30054
rect 20536 29990 20588 29996
rect 20548 29578 20576 29990
rect 20536 29572 20588 29578
rect 20536 29514 20588 29520
rect 20732 29306 20760 30194
rect 21732 30184 21784 30190
rect 21732 30126 21784 30132
rect 21088 30116 21140 30122
rect 21088 30058 21140 30064
rect 21100 29714 21128 30058
rect 21744 30054 21772 30126
rect 21732 30048 21784 30054
rect 21732 29990 21784 29996
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 21732 29640 21784 29646
rect 21732 29582 21784 29588
rect 20720 29300 20772 29306
rect 20720 29242 20772 29248
rect 20718 29200 20774 29209
rect 20536 29164 20588 29170
rect 20718 29135 20720 29144
rect 20536 29106 20588 29112
rect 20772 29135 20774 29144
rect 20720 29106 20772 29112
rect 20548 22420 20576 29106
rect 20812 28960 20864 28966
rect 20812 28902 20864 28908
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20732 28218 20760 28426
rect 20720 28212 20772 28218
rect 20720 28154 20772 28160
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20640 24886 20668 25094
rect 20628 24880 20680 24886
rect 20628 24822 20680 24828
rect 20824 23322 20852 28902
rect 21744 28490 21772 29582
rect 21732 28484 21784 28490
rect 21732 28426 21784 28432
rect 21744 28014 21772 28426
rect 21272 28008 21324 28014
rect 21272 27950 21324 27956
rect 21732 28008 21784 28014
rect 21732 27950 21784 27956
rect 21284 26926 21312 27950
rect 21836 27946 21864 31889
rect 22192 30388 22244 30394
rect 22192 30330 22244 30336
rect 22008 30252 22060 30258
rect 22008 30194 22060 30200
rect 22020 29170 22048 30194
rect 22100 29572 22152 29578
rect 22100 29514 22152 29520
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 22112 29034 22140 29514
rect 22204 29238 22232 30330
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22836 30252 22888 30258
rect 22836 30194 22888 30200
rect 22192 29232 22244 29238
rect 22192 29174 22244 29180
rect 22480 29186 22508 30194
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22480 29170 22600 29186
rect 22480 29164 22612 29170
rect 22480 29158 22560 29164
rect 22192 29096 22244 29102
rect 22192 29038 22244 29044
rect 22100 29028 22152 29034
rect 22100 28970 22152 28976
rect 22204 28994 22232 29038
rect 22204 28966 22324 28994
rect 22296 28558 22324 28966
rect 22480 28626 22508 29158
rect 22560 29106 22612 29112
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22296 28422 22324 28494
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 21824 27940 21876 27946
rect 21824 27882 21876 27888
rect 22008 27872 22060 27878
rect 22008 27814 22060 27820
rect 21548 27668 21600 27674
rect 21548 27610 21600 27616
rect 21456 27396 21508 27402
rect 21456 27338 21508 27344
rect 21468 27130 21496 27338
rect 21456 27124 21508 27130
rect 21456 27066 21508 27072
rect 21272 26920 21324 26926
rect 21272 26862 21324 26868
rect 20916 24670 21128 24698
rect 20916 24614 20944 24670
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 20996 24608 21048 24614
rect 20996 24550 21048 24556
rect 21008 24206 21036 24550
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 21008 23186 21036 24142
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 20904 22704 20956 22710
rect 20904 22646 20956 22652
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20628 22432 20680 22438
rect 20548 22392 20628 22420
rect 20628 22374 20680 22380
rect 20732 22098 20760 22578
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20536 21412 20588 21418
rect 20536 21354 20588 21360
rect 20548 20534 20576 21354
rect 20824 21146 20852 22034
rect 20916 21554 20944 22646
rect 21008 22642 21036 23122
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20916 20942 20944 21286
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20536 20528 20588 20534
rect 20536 20470 20588 20476
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20444 20324 20496 20330
rect 20444 20266 20496 20272
rect 20260 19712 20312 19718
rect 20258 19680 20260 19689
rect 20312 19680 20314 19689
rect 20258 19615 20314 19624
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 20272 19378 20300 19450
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20364 19174 20392 19450
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20456 18970 20484 20266
rect 20732 19446 20760 20878
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20824 20602 20852 20810
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20456 18834 20484 18906
rect 20732 18834 20760 19382
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18086 20300 18566
rect 20732 18086 20760 18634
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 19708 17808 19760 17814
rect 19708 17750 19760 17756
rect 19720 17338 19748 17750
rect 20168 17672 20220 17678
rect 20272 17660 20300 18022
rect 20220 17632 20300 17660
rect 20352 17672 20404 17678
rect 20168 17614 20220 17620
rect 20352 17614 20404 17620
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 19840 17436 20148 17456
rect 19840 17434 19846 17436
rect 19902 17434 19926 17436
rect 19982 17434 20006 17436
rect 20062 17434 20086 17436
rect 20142 17434 20148 17436
rect 19902 17382 19904 17434
rect 20084 17382 20086 17434
rect 19840 17380 19846 17382
rect 19902 17380 19926 17382
rect 19982 17380 20006 17382
rect 20062 17380 20086 17382
rect 20142 17380 20148 17382
rect 19840 17360 20148 17380
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19628 14074 19656 14554
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19720 13530 19748 16730
rect 20180 16726 20208 17614
rect 20364 17338 20392 17614
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20168 16720 20220 16726
rect 20168 16662 20220 16668
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 19840 16348 20148 16368
rect 19840 16346 19846 16348
rect 19902 16346 19926 16348
rect 19982 16346 20006 16348
rect 20062 16346 20086 16348
rect 20142 16346 20148 16348
rect 19902 16294 19904 16346
rect 20084 16294 20086 16346
rect 19840 16292 19846 16294
rect 19902 16292 19926 16294
rect 19982 16292 20006 16294
rect 20062 16292 20086 16294
rect 20142 16292 20148 16294
rect 19840 16272 20148 16292
rect 20180 15586 20208 16526
rect 20364 15910 20392 16730
rect 20548 16726 20576 17614
rect 20536 16720 20588 16726
rect 20536 16662 20588 16668
rect 20444 16516 20496 16522
rect 20444 16458 20496 16464
rect 20456 16114 20484 16458
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20548 16114 20576 16186
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20444 15972 20496 15978
rect 20444 15914 20496 15920
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20456 15722 20484 15914
rect 20364 15694 20484 15722
rect 20548 15706 20576 16050
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20536 15700 20588 15706
rect 20364 15586 20392 15694
rect 20536 15642 20588 15648
rect 20180 15558 20392 15586
rect 19840 15260 20148 15280
rect 19840 15258 19846 15260
rect 19902 15258 19926 15260
rect 19982 15258 20006 15260
rect 20062 15258 20086 15260
rect 20142 15258 20148 15260
rect 19902 15206 19904 15258
rect 20084 15206 20086 15258
rect 19840 15204 19846 15206
rect 19902 15204 19926 15206
rect 19982 15204 20006 15206
rect 20062 15204 20086 15206
rect 20142 15204 20148 15206
rect 19840 15184 20148 15204
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20180 14385 20208 14418
rect 20166 14376 20222 14385
rect 20166 14311 20222 14320
rect 19840 14172 20148 14192
rect 19840 14170 19846 14172
rect 19902 14170 19926 14172
rect 19982 14170 20006 14172
rect 20062 14170 20086 14172
rect 20142 14170 20148 14172
rect 19902 14118 19904 14170
rect 20084 14118 20086 14170
rect 19840 14116 19846 14118
rect 19902 14116 19926 14118
rect 19982 14116 20006 14118
rect 20062 14116 20086 14118
rect 20142 14116 20148 14118
rect 19840 14096 20148 14116
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19720 12986 19748 13466
rect 20260 13252 20312 13258
rect 20260 13194 20312 13200
rect 19840 13084 20148 13104
rect 19840 13082 19846 13084
rect 19902 13082 19926 13084
rect 19982 13082 20006 13084
rect 20062 13082 20086 13084
rect 20142 13082 20148 13084
rect 19902 13030 19904 13082
rect 20084 13030 20086 13082
rect 19840 13028 19846 13030
rect 19902 13028 19926 13030
rect 19982 13028 20006 13030
rect 20062 13028 20086 13030
rect 20142 13028 20148 13030
rect 19840 13008 20148 13028
rect 20272 12986 20300 13194
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19536 12442 19564 12854
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19248 11212 19300 11218
rect 19300 11172 19380 11200
rect 19248 11154 19300 11160
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18156 9710 18276 9738
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17696 7478 17724 8230
rect 17788 8022 17816 8978
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17972 8090 18000 8434
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17684 7472 17736 7478
rect 17684 7414 17736 7420
rect 17788 6866 17816 7958
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 7274 17908 7822
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17972 7410 18000 7482
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17972 6798 18000 7210
rect 18064 7206 18092 8774
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18064 7002 18092 7142
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 6322 18000 6598
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 18064 6254 18092 6938
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17604 5302 17632 5646
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 17696 5370 17724 5510
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17776 5296 17828 5302
rect 17776 5238 17828 5244
rect 17788 4622 17816 5238
rect 18064 5166 18092 5510
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17972 4214 18000 4422
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17604 3738 17632 4082
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 18064 3670 18092 5102
rect 18156 4010 18184 9710
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18248 9178 18276 9522
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 18248 7886 18276 8502
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18248 6662 18276 7346
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18064 2922 18092 3470
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 18340 2854 18368 11086
rect 19352 10674 19380 11172
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19720 10266 19748 12922
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 20088 12306 20116 12718
rect 20364 12434 20392 15558
rect 20640 15502 20668 15846
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20180 12406 20392 12434
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 19840 11996 20148 12016
rect 19840 11994 19846 11996
rect 19902 11994 19926 11996
rect 19982 11994 20006 11996
rect 20062 11994 20086 11996
rect 20142 11994 20148 11996
rect 19902 11942 19904 11994
rect 20084 11942 20086 11994
rect 19840 11940 19846 11942
rect 19902 11940 19926 11942
rect 19982 11940 20006 11942
rect 20062 11940 20086 11942
rect 20142 11940 20148 11942
rect 19840 11920 20148 11940
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19904 11354 19932 11630
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19904 11150 19932 11290
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19840 10908 20148 10928
rect 19840 10906 19846 10908
rect 19902 10906 19926 10908
rect 19982 10906 20006 10908
rect 20062 10906 20086 10908
rect 20142 10906 20148 10908
rect 19902 10854 19904 10906
rect 20084 10854 20086 10906
rect 19840 10852 19846 10854
rect 19902 10852 19926 10854
rect 19982 10852 20006 10854
rect 20062 10852 20086 10854
rect 20142 10852 20148 10854
rect 19840 10832 20148 10852
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 18972 9648 19024 9654
rect 18972 9590 19024 9596
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18892 8838 18920 9318
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18524 7818 18552 8366
rect 18616 8362 18644 8774
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18524 7410 18552 7754
rect 18708 7750 18736 8774
rect 18892 8294 18920 8774
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18708 7206 18736 7686
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18616 6322 18644 6938
rect 18708 6390 18736 7142
rect 18800 6798 18828 7346
rect 18892 6798 18920 8230
rect 18984 7478 19012 9590
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 19076 7886 19104 9386
rect 19168 8634 19196 9658
rect 19720 9654 19748 10202
rect 19840 9820 20148 9840
rect 19840 9818 19846 9820
rect 19902 9818 19926 9820
rect 19982 9818 20006 9820
rect 20062 9818 20086 9820
rect 20142 9818 20148 9820
rect 19902 9766 19904 9818
rect 20084 9766 20086 9818
rect 19840 9764 19846 9766
rect 19902 9764 19926 9766
rect 19982 9764 20006 9766
rect 20062 9764 20086 9766
rect 20142 9764 20148 9766
rect 19840 9744 20148 9764
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19352 8634 19380 8910
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19168 8514 19196 8570
rect 19168 8498 19472 8514
rect 19720 8498 19748 9318
rect 19840 8732 20148 8752
rect 19840 8730 19846 8732
rect 19902 8730 19926 8732
rect 19982 8730 20006 8732
rect 20062 8730 20086 8732
rect 20142 8730 20148 8732
rect 19902 8678 19904 8730
rect 20084 8678 20086 8730
rect 19840 8676 19846 8678
rect 19902 8676 19926 8678
rect 19982 8676 20006 8678
rect 20062 8676 20086 8678
rect 20142 8676 20148 8678
rect 19840 8656 20148 8676
rect 19168 8492 19484 8498
rect 19168 8486 19432 8492
rect 19432 8434 19484 8440
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19338 8392 19394 8401
rect 19338 8327 19340 8336
rect 19392 8327 19394 8336
rect 19708 8356 19760 8362
rect 19340 8298 19392 8304
rect 19708 8298 19760 8304
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 18984 7002 19012 7414
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18420 5704 18472 5710
rect 18616 5692 18644 6258
rect 18708 6100 18736 6326
rect 19352 6304 19380 8298
rect 19720 7410 19748 8298
rect 19840 7644 20148 7664
rect 19840 7642 19846 7644
rect 19902 7642 19926 7644
rect 19982 7642 20006 7644
rect 20062 7642 20086 7644
rect 20142 7642 20148 7644
rect 19902 7590 19904 7642
rect 20084 7590 20086 7642
rect 19840 7588 19846 7590
rect 19902 7588 19926 7590
rect 19982 7588 20006 7590
rect 20062 7588 20086 7590
rect 20142 7588 20148 7590
rect 19840 7568 20148 7588
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19720 6934 19748 7346
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19708 6928 19760 6934
rect 19708 6870 19760 6876
rect 19812 6866 19840 7278
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 20088 6730 20116 6870
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 19840 6556 20148 6576
rect 19840 6554 19846 6556
rect 19902 6554 19926 6556
rect 19982 6554 20006 6556
rect 20062 6554 20086 6556
rect 20142 6554 20148 6556
rect 19902 6502 19904 6554
rect 20084 6502 20086 6554
rect 19840 6500 19846 6502
rect 19902 6500 19926 6502
rect 19982 6500 20006 6502
rect 20062 6500 20086 6502
rect 20142 6500 20148 6502
rect 19840 6480 20148 6500
rect 20076 6384 20128 6390
rect 20076 6326 20128 6332
rect 19260 6276 19380 6304
rect 19892 6316 19944 6322
rect 18788 6112 18840 6118
rect 18708 6072 18788 6100
rect 18708 5914 18736 6072
rect 18788 6054 18840 6060
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 18696 5704 18748 5710
rect 18616 5664 18696 5692
rect 18420 5646 18472 5652
rect 18696 5646 18748 5652
rect 18432 5098 18460 5646
rect 19260 5166 19288 6276
rect 19892 6258 19944 6264
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 18420 5092 18472 5098
rect 18420 5034 18472 5040
rect 18432 4214 18460 5034
rect 19352 4758 19380 6122
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19616 5840 19668 5846
rect 19616 5782 19668 5788
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 19444 5166 19472 5714
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19536 5302 19564 5646
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 19628 4622 19656 5782
rect 19720 5370 19748 6054
rect 19904 5914 19932 6258
rect 19892 5908 19944 5914
rect 19892 5850 19944 5856
rect 20088 5846 20116 6326
rect 20076 5840 20128 5846
rect 20076 5782 20128 5788
rect 20088 5710 20116 5782
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 19840 5468 20148 5488
rect 19840 5466 19846 5468
rect 19902 5466 19926 5468
rect 19982 5466 20006 5468
rect 20062 5466 20086 5468
rect 20142 5466 20148 5468
rect 19902 5414 19904 5466
rect 20084 5414 20086 5466
rect 19840 5412 19846 5414
rect 19902 5412 19926 5414
rect 19982 5412 20006 5414
rect 20062 5412 20086 5414
rect 20142 5412 20148 5414
rect 19840 5392 20148 5412
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19720 4690 19748 5170
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19076 4214 19104 4422
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18512 4208 18564 4214
rect 18512 4150 18564 4156
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18432 3602 18460 3878
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18524 3534 18552 4150
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18892 3126 18920 3334
rect 18880 3120 18932 3126
rect 18880 3062 18932 3068
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 19076 2774 19104 3878
rect 19536 3466 19564 4422
rect 19720 4282 19748 4626
rect 19840 4380 20148 4400
rect 19840 4378 19846 4380
rect 19902 4378 19926 4380
rect 19982 4378 20006 4380
rect 20062 4378 20086 4380
rect 20142 4378 20148 4380
rect 19902 4326 19904 4378
rect 20084 4326 20086 4378
rect 19840 4324 19846 4326
rect 19902 4324 19926 4326
rect 19982 4324 20006 4326
rect 20062 4324 20086 4326
rect 20142 4324 20148 4326
rect 19840 4304 20148 4324
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19708 3460 19760 3466
rect 19708 3402 19760 3408
rect 19720 3058 19748 3402
rect 19840 3292 20148 3312
rect 19840 3290 19846 3292
rect 19902 3290 19926 3292
rect 19982 3290 20006 3292
rect 20062 3290 20086 3292
rect 20142 3290 20148 3292
rect 19902 3238 19904 3290
rect 20084 3238 20086 3290
rect 19840 3236 19846 3238
rect 19902 3236 19926 3238
rect 19982 3236 20006 3238
rect 20062 3236 20086 3238
rect 20142 3236 20148 3238
rect 19840 3216 20148 3236
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 17512 2746 17632 2774
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17604 800 17632 2746
rect 18892 2746 19104 2774
rect 18892 800 18920 2746
rect 19840 2204 20148 2224
rect 19840 2202 19846 2204
rect 19902 2202 19926 2204
rect 19982 2202 20006 2204
rect 20062 2202 20086 2204
rect 20142 2202 20148 2204
rect 19902 2150 19904 2202
rect 20084 2150 20086 2202
rect 19840 2148 19846 2150
rect 19902 2148 19926 2150
rect 19982 2148 20006 2150
rect 20062 2148 20086 2150
rect 20142 2148 20148 2150
rect 19840 2128 20148 2148
rect 20180 1986 20208 12406
rect 20456 12170 20484 12582
rect 20732 12434 20760 18022
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20916 14006 20944 14282
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21008 12986 21036 13194
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20732 12406 20944 12434
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20364 8974 20392 9318
rect 20640 8974 20668 9522
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20364 8673 20392 8774
rect 20350 8664 20406 8673
rect 20350 8599 20406 8608
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20272 7002 20300 7278
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 5710 20300 6598
rect 20364 6458 20392 8502
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20456 6866 20484 7346
rect 20548 6866 20576 8026
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20548 6662 20576 6802
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20824 5914 20852 6258
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20272 5030 20300 5646
rect 20628 5636 20680 5642
rect 20628 5578 20680 5584
rect 20640 5370 20668 5578
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20824 5234 20852 5850
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20732 3670 20760 4082
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20088 1958 20208 1986
rect 20088 800 20116 1958
rect 15304 734 15516 762
rect 16394 0 16450 800
rect 17590 0 17646 800
rect 18878 0 18934 800
rect 20074 0 20130 800
rect 20916 762 20944 12406
rect 21008 12102 21036 12922
rect 21100 12850 21128 24670
rect 21284 24614 21312 26862
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21560 20602 21588 27610
rect 22020 27606 22048 27814
rect 22008 27600 22060 27606
rect 22008 27542 22060 27548
rect 21640 26988 21692 26994
rect 21640 26930 21692 26936
rect 21652 26586 21680 26930
rect 21640 26580 21692 26586
rect 21640 26522 21692 26528
rect 21732 26308 21784 26314
rect 21732 26250 21784 26256
rect 21744 24818 21772 26250
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 21824 25696 21876 25702
rect 21824 25638 21876 25644
rect 21836 25226 21864 25638
rect 21824 25220 21876 25226
rect 21824 25162 21876 25168
rect 22020 24954 22048 25842
rect 22204 25702 22232 28018
rect 22296 27878 22324 28358
rect 22480 28218 22508 28562
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22468 28212 22520 28218
rect 22468 28154 22520 28160
rect 22468 27940 22520 27946
rect 22468 27882 22520 27888
rect 22284 27872 22336 27878
rect 22284 27814 22336 27820
rect 22192 25696 22244 25702
rect 22192 25638 22244 25644
rect 22480 25498 22508 27882
rect 22572 27606 22600 28426
rect 22560 27600 22612 27606
rect 22560 27542 22612 27548
rect 22560 27396 22612 27402
rect 22560 27338 22612 27344
rect 22468 25492 22520 25498
rect 22468 25434 22520 25440
rect 22008 24948 22060 24954
rect 22008 24890 22060 24896
rect 21732 24812 21784 24818
rect 21732 24754 21784 24760
rect 21744 22778 21772 24754
rect 22468 24336 22520 24342
rect 22468 24278 22520 24284
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 21824 23520 21876 23526
rect 21824 23462 21876 23468
rect 21836 23050 21864 23462
rect 21824 23044 21876 23050
rect 21824 22986 21876 22992
rect 22020 22778 22048 23666
rect 22204 23338 22232 24142
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22112 23322 22232 23338
rect 22100 23316 22232 23322
rect 22152 23310 22232 23316
rect 22100 23258 22152 23264
rect 22388 22930 22416 23802
rect 22480 23050 22508 24278
rect 22572 23866 22600 27338
rect 22664 26790 22692 29990
rect 22848 29306 22876 30194
rect 23112 30048 23164 30054
rect 23112 29990 23164 29996
rect 23124 29578 23152 29990
rect 23112 29572 23164 29578
rect 23112 29514 23164 29520
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 22940 29238 22968 29446
rect 22928 29232 22980 29238
rect 22742 29200 22798 29209
rect 22928 29174 22980 29180
rect 22742 29135 22744 29144
rect 22796 29135 22798 29144
rect 22744 29106 22796 29112
rect 23216 28778 23244 31889
rect 24400 29164 24452 29170
rect 24400 29106 24452 29112
rect 23848 29028 23900 29034
rect 23848 28970 23900 28976
rect 23032 28750 23244 28778
rect 22928 28484 22980 28490
rect 22848 28444 22928 28472
rect 22744 27464 22796 27470
rect 22744 27406 22796 27412
rect 22652 26784 22704 26790
rect 22652 26726 22704 26732
rect 22756 26382 22784 27406
rect 22848 27402 22876 28444
rect 22928 28426 22980 28432
rect 22928 27600 22980 27606
rect 22928 27542 22980 27548
rect 22836 27396 22888 27402
rect 22836 27338 22888 27344
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22652 25696 22704 25702
rect 22652 25638 22704 25644
rect 22664 25226 22692 25638
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22836 25288 22888 25294
rect 22836 25230 22888 25236
rect 22652 25220 22704 25226
rect 22652 25162 22704 25168
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22664 24138 22692 24346
rect 22756 24274 22784 25230
rect 22744 24268 22796 24274
rect 22744 24210 22796 24216
rect 22848 24206 22876 25230
rect 22940 25106 22968 27542
rect 23032 27470 23060 28750
rect 23204 28552 23256 28558
rect 23204 28494 23256 28500
rect 23388 28552 23440 28558
rect 23388 28494 23440 28500
rect 23216 28422 23244 28494
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 23400 28218 23428 28494
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 23572 28416 23624 28422
rect 23572 28358 23624 28364
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 23584 28150 23612 28358
rect 23676 28218 23704 28426
rect 23664 28212 23716 28218
rect 23664 28154 23716 28160
rect 23572 28144 23624 28150
rect 23572 28086 23624 28092
rect 23664 28008 23716 28014
rect 23664 27950 23716 27956
rect 23388 27872 23440 27878
rect 23440 27832 23520 27860
rect 23388 27814 23440 27820
rect 23296 27600 23348 27606
rect 23296 27542 23348 27548
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 23032 27130 23060 27406
rect 23020 27124 23072 27130
rect 23020 27066 23072 27072
rect 23308 27062 23336 27542
rect 23492 27470 23520 27832
rect 23676 27674 23704 27950
rect 23664 27668 23716 27674
rect 23716 27628 23796 27656
rect 23664 27610 23716 27616
rect 23664 27532 23716 27538
rect 23664 27474 23716 27480
rect 23480 27464 23532 27470
rect 23480 27406 23532 27412
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23492 27282 23520 27406
rect 23400 27254 23520 27282
rect 23296 27056 23348 27062
rect 23296 26998 23348 27004
rect 23020 26784 23072 26790
rect 23020 26726 23072 26732
rect 23032 26296 23060 26726
rect 23204 26376 23256 26382
rect 23204 26318 23256 26324
rect 23112 26308 23164 26314
rect 23032 26268 23112 26296
rect 23112 26250 23164 26256
rect 23020 25492 23072 25498
rect 23020 25434 23072 25440
rect 23032 25226 23060 25434
rect 23020 25220 23072 25226
rect 23020 25162 23072 25168
rect 22940 25078 23060 25106
rect 22928 24268 22980 24274
rect 22928 24210 22980 24216
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 22652 24132 22704 24138
rect 22652 24074 22704 24080
rect 22560 23860 22612 23866
rect 22560 23802 22612 23808
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22756 23322 22784 23666
rect 22744 23316 22796 23322
rect 22744 23258 22796 23264
rect 22468 23044 22520 23050
rect 22468 22986 22520 22992
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 22388 22902 22508 22930
rect 21732 22772 21784 22778
rect 21732 22714 21784 22720
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22020 21554 22048 22578
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 22020 21146 22048 21490
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 22112 20890 22140 21830
rect 22204 21690 22232 22578
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22296 21962 22324 22374
rect 22480 22234 22508 22902
rect 22572 22642 22600 22986
rect 22652 22772 22704 22778
rect 22652 22714 22704 22720
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22376 22228 22428 22234
rect 22376 22170 22428 22176
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22282 21584 22338 21593
rect 22282 21519 22284 21528
rect 22336 21519 22338 21528
rect 22284 21490 22336 21496
rect 22388 21418 22416 22170
rect 22480 21418 22508 22170
rect 22376 21412 22428 21418
rect 22376 21354 22428 21360
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 22480 21146 22508 21354
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 22192 20936 22244 20942
rect 22112 20884 22192 20890
rect 22112 20878 22244 20884
rect 22112 20862 22232 20878
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21560 19786 21588 20538
rect 22112 20534 22140 20862
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22204 19854 22232 20742
rect 22376 20528 22428 20534
rect 22376 20470 22428 20476
rect 22388 20058 22416 20470
rect 22376 20052 22428 20058
rect 22376 19994 22428 20000
rect 22572 19990 22600 22578
rect 22664 22098 22692 22714
rect 22756 22642 22784 23258
rect 22848 22778 22876 24142
rect 22940 23526 22968 24210
rect 23032 24070 23060 25078
rect 23020 24064 23072 24070
rect 23020 24006 23072 24012
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22940 22658 22968 23462
rect 23032 22982 23060 24006
rect 23020 22976 23072 22982
rect 23020 22918 23072 22924
rect 22744 22636 22796 22642
rect 22744 22578 22796 22584
rect 22848 22630 22968 22658
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 22664 21593 22692 22034
rect 22848 22030 22876 22630
rect 23124 22522 23152 26250
rect 23216 24206 23244 26318
rect 23400 26194 23428 27254
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 23492 26382 23520 27066
rect 23584 26586 23612 27406
rect 23572 26580 23624 26586
rect 23572 26522 23624 26528
rect 23676 26382 23704 27474
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 23664 26376 23716 26382
rect 23664 26318 23716 26324
rect 23400 26166 23520 26194
rect 23294 25936 23350 25945
rect 23294 25871 23296 25880
rect 23348 25871 23350 25880
rect 23296 25842 23348 25848
rect 23308 25129 23336 25842
rect 23386 25256 23442 25265
rect 23386 25191 23388 25200
rect 23440 25191 23442 25200
rect 23388 25162 23440 25168
rect 23294 25120 23350 25129
rect 23294 25055 23350 25064
rect 23308 24954 23336 25055
rect 23296 24948 23348 24954
rect 23296 24890 23348 24896
rect 23400 24410 23428 25162
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23216 23202 23244 24142
rect 23400 24070 23428 24346
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23216 23174 23336 23202
rect 23308 23118 23336 23174
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23204 22976 23256 22982
rect 23204 22918 23256 22924
rect 22940 22494 23152 22522
rect 22836 22024 22888 22030
rect 22756 21972 22836 21978
rect 22756 21966 22888 21972
rect 22756 21950 22876 21966
rect 22650 21584 22706 21593
rect 22756 21554 22784 21950
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 22848 21622 22876 21830
rect 22836 21616 22888 21622
rect 22836 21558 22888 21564
rect 22650 21519 22706 21528
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22664 21010 22692 21422
rect 22848 21350 22876 21558
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22560 19984 22612 19990
rect 22560 19926 22612 19932
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 22560 19848 22612 19854
rect 22560 19790 22612 19796
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 22572 18970 22600 19790
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 21178 18320 21234 18329
rect 21178 18255 21234 18264
rect 21192 17338 21220 18255
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 22388 16574 22416 18634
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22664 18290 22692 18566
rect 22652 18284 22704 18290
rect 22652 18226 22704 18232
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22480 16658 22508 17682
rect 22664 17678 22692 18226
rect 22756 18086 22784 18702
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22848 17898 22876 21286
rect 22940 18970 22968 22494
rect 23216 22250 23244 22918
rect 23308 22506 23336 23054
rect 23296 22500 23348 22506
rect 23296 22442 23348 22448
rect 23032 22222 23244 22250
rect 23032 19718 23060 22222
rect 23112 22092 23164 22098
rect 23112 22034 23164 22040
rect 23124 21962 23152 22034
rect 23112 21956 23164 21962
rect 23112 21898 23164 21904
rect 23124 21418 23152 21898
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 23400 21078 23428 23802
rect 23492 21894 23520 26166
rect 23676 24206 23704 26318
rect 23768 25362 23796 27628
rect 23756 25356 23808 25362
rect 23756 25298 23808 25304
rect 23756 25220 23808 25226
rect 23756 25162 23808 25168
rect 23768 25129 23796 25162
rect 23754 25120 23810 25129
rect 23754 25055 23810 25064
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23584 23066 23612 24006
rect 23676 23254 23704 24142
rect 23756 24064 23808 24070
rect 23756 24006 23808 24012
rect 23768 23662 23796 24006
rect 23756 23656 23808 23662
rect 23756 23598 23808 23604
rect 23664 23248 23716 23254
rect 23664 23190 23716 23196
rect 23768 23186 23796 23598
rect 23860 23322 23888 28970
rect 23940 28960 23992 28966
rect 23940 28902 23992 28908
rect 23952 26450 23980 28902
rect 24412 28558 24440 29106
rect 24400 28552 24452 28558
rect 24400 28494 24452 28500
rect 24032 28416 24084 28422
rect 24032 28358 24084 28364
rect 24044 27538 24072 28358
rect 24032 27532 24084 27538
rect 24032 27474 24084 27480
rect 24412 27402 24440 28494
rect 24400 27396 24452 27402
rect 24400 27338 24452 27344
rect 24032 27328 24084 27334
rect 24032 27270 24084 27276
rect 24044 27062 24072 27270
rect 24504 27130 24532 31889
rect 24563 29948 24871 29968
rect 24563 29946 24569 29948
rect 24625 29946 24649 29948
rect 24705 29946 24729 29948
rect 24785 29946 24809 29948
rect 24865 29946 24871 29948
rect 24625 29894 24627 29946
rect 24807 29894 24809 29946
rect 24563 29892 24569 29894
rect 24625 29892 24649 29894
rect 24705 29892 24729 29894
rect 24785 29892 24809 29894
rect 24865 29892 24871 29894
rect 24563 29872 24871 29892
rect 25884 28966 25912 31889
rect 26146 31648 26202 31657
rect 26146 31583 26202 31592
rect 26160 29850 26188 31583
rect 26240 30320 26292 30326
rect 26240 30262 26292 30268
rect 26148 29844 26200 29850
rect 26148 29786 26200 29792
rect 26252 29753 26280 30262
rect 26238 29744 26294 29753
rect 26238 29679 26294 29688
rect 25872 28960 25924 28966
rect 25872 28902 25924 28908
rect 24563 28860 24871 28880
rect 24563 28858 24569 28860
rect 24625 28858 24649 28860
rect 24705 28858 24729 28860
rect 24785 28858 24809 28860
rect 24865 28858 24871 28860
rect 24625 28806 24627 28858
rect 24807 28806 24809 28858
rect 24563 28804 24569 28806
rect 24625 28804 24649 28806
rect 24705 28804 24729 28806
rect 24785 28804 24809 28806
rect 24865 28804 24871 28806
rect 24563 28784 24871 28804
rect 25228 28756 25280 28762
rect 25228 28698 25280 28704
rect 24676 28416 24728 28422
rect 24676 28358 24728 28364
rect 24688 28082 24716 28358
rect 25240 28082 25268 28698
rect 26792 28144 26844 28150
rect 26792 28086 26844 28092
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25412 28076 25464 28082
rect 25412 28018 25464 28024
rect 24563 27772 24871 27792
rect 24563 27770 24569 27772
rect 24625 27770 24649 27772
rect 24705 27770 24729 27772
rect 24785 27770 24809 27772
rect 24865 27770 24871 27772
rect 24625 27718 24627 27770
rect 24807 27718 24809 27770
rect 24563 27716 24569 27718
rect 24625 27716 24649 27718
rect 24705 27716 24729 27718
rect 24785 27716 24809 27718
rect 24865 27716 24871 27718
rect 24563 27696 24871 27716
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 24492 27124 24544 27130
rect 24492 27066 24544 27072
rect 24032 27056 24084 27062
rect 24032 26998 24084 27004
rect 24964 26926 24992 27406
rect 24952 26920 25004 26926
rect 24952 26862 25004 26868
rect 24964 26790 24992 26862
rect 24952 26784 25004 26790
rect 24952 26726 25004 26732
rect 24563 26684 24871 26704
rect 24563 26682 24569 26684
rect 24625 26682 24649 26684
rect 24705 26682 24729 26684
rect 24785 26682 24809 26684
rect 24865 26682 24871 26684
rect 24625 26630 24627 26682
rect 24807 26630 24809 26682
rect 24563 26628 24569 26630
rect 24625 26628 24649 26630
rect 24705 26628 24729 26630
rect 24785 26628 24809 26630
rect 24865 26628 24871 26630
rect 24563 26608 24871 26628
rect 23940 26444 23992 26450
rect 23940 26386 23992 26392
rect 24964 25838 24992 26726
rect 25240 25922 25268 28018
rect 25424 27946 25452 28018
rect 25412 27940 25464 27946
rect 25412 27882 25464 27888
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25332 26586 25360 26862
rect 25320 26580 25372 26586
rect 25320 26522 25372 26528
rect 25056 25894 25268 25922
rect 24952 25832 25004 25838
rect 24952 25774 25004 25780
rect 24563 25596 24871 25616
rect 24563 25594 24569 25596
rect 24625 25594 24649 25596
rect 24705 25594 24729 25596
rect 24785 25594 24809 25596
rect 24865 25594 24871 25596
rect 24625 25542 24627 25594
rect 24807 25542 24809 25594
rect 24563 25540 24569 25542
rect 24625 25540 24649 25542
rect 24705 25540 24729 25542
rect 24785 25540 24809 25542
rect 24865 25540 24871 25542
rect 24563 25520 24871 25540
rect 24032 25424 24084 25430
rect 24032 25366 24084 25372
rect 24676 25424 24728 25430
rect 24676 25366 24728 25372
rect 24044 24750 24072 25366
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24412 24954 24440 25230
rect 24400 24948 24452 24954
rect 24400 24890 24452 24896
rect 24688 24886 24716 25366
rect 24676 24880 24728 24886
rect 24676 24822 24728 24828
rect 24964 24834 24992 25774
rect 25056 25498 25084 25894
rect 25228 25832 25280 25838
rect 25228 25774 25280 25780
rect 25240 25498 25268 25774
rect 25424 25702 25452 27882
rect 25780 27872 25832 27878
rect 26804 27849 26832 28086
rect 25780 27814 25832 27820
rect 26790 27840 26846 27849
rect 25792 27674 25820 27814
rect 26790 27775 26846 27784
rect 25780 27668 25832 27674
rect 25780 27610 25832 27616
rect 26804 27606 26832 27775
rect 26792 27600 26844 27606
rect 26792 27542 26844 27548
rect 25872 27396 25924 27402
rect 25872 27338 25924 27344
rect 25688 27328 25740 27334
rect 25688 27270 25740 27276
rect 25700 26994 25728 27270
rect 25884 27130 25912 27338
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25688 26988 25740 26994
rect 25688 26930 25740 26936
rect 27172 26058 27200 31889
rect 28552 28218 28580 31889
rect 29840 28694 29868 31889
rect 29828 28688 29880 28694
rect 29828 28630 29880 28636
rect 28540 28212 28592 28218
rect 28540 28154 28592 28160
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 27080 26030 27200 26058
rect 26252 25945 26280 25978
rect 26238 25936 26294 25945
rect 26238 25871 26294 25880
rect 27080 25838 27108 26030
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 27068 25832 27120 25838
rect 27068 25774 27120 25780
rect 25412 25696 25464 25702
rect 25412 25638 25464 25644
rect 25044 25492 25096 25498
rect 25044 25434 25096 25440
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25056 24970 25084 25434
rect 25056 24942 25176 24970
rect 24964 24806 25084 24834
rect 25148 24818 25176 24942
rect 25056 24750 25084 24806
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 24032 24744 24084 24750
rect 24032 24686 24084 24692
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 24124 24608 24176 24614
rect 24124 24550 24176 24556
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 24044 23798 24072 24006
rect 24032 23792 24084 23798
rect 24032 23734 24084 23740
rect 23848 23316 23900 23322
rect 23848 23258 23900 23264
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23584 23038 23704 23066
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23584 21622 23612 22034
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23388 21072 23440 21078
rect 23388 21014 23440 21020
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 23124 20806 23152 20946
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23112 20800 23164 20806
rect 23112 20742 23164 20748
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 22940 18766 22968 18906
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 22756 17870 22876 17898
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22652 17128 22704 17134
rect 22650 17096 22652 17105
rect 22704 17096 22706 17105
rect 22650 17031 22706 17040
rect 22664 16794 22692 17031
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22756 16574 22784 17870
rect 22940 16574 22968 18362
rect 22296 16546 22416 16574
rect 22664 16546 22784 16574
rect 22848 16546 22968 16574
rect 21178 16280 21234 16289
rect 21178 16215 21180 16224
rect 21232 16215 21234 16224
rect 21180 16186 21232 16192
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21652 14958 21680 15438
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21192 13870 21220 14894
rect 22020 14618 22048 15370
rect 22296 15366 22324 16546
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21192 13530 21220 13806
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21560 13376 21588 14350
rect 21652 14346 21680 14486
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21652 13938 21680 14282
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21836 13462 21864 14350
rect 22296 14278 22324 15302
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22388 14550 22416 15098
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22376 14544 22428 14550
rect 22376 14486 22428 14492
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 21824 13456 21876 13462
rect 21824 13398 21876 13404
rect 21640 13388 21692 13394
rect 21560 13348 21640 13376
rect 21692 13348 21772 13376
rect 21640 13330 21692 13336
rect 21744 13308 21772 13348
rect 22020 13326 22048 14010
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22112 13530 22140 13874
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 21824 13320 21876 13326
rect 21744 13280 21824 13308
rect 21824 13262 21876 13268
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21836 12646 21864 13262
rect 22020 12900 22048 13262
rect 22100 12912 22152 12918
rect 22020 12872 22100 12900
rect 22100 12854 22152 12860
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21178 12200 21234 12209
rect 21178 12135 21234 12144
rect 21192 12102 21220 12135
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 21192 11354 21220 12038
rect 21560 11898 21588 12378
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21836 11762 21864 12582
rect 22112 12442 22140 12854
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22204 12102 22232 13262
rect 22296 12986 22324 14214
rect 22388 13394 22416 14486
rect 22572 13530 22600 14962
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22204 11762 22232 12038
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22388 11626 22416 12106
rect 22376 11620 22428 11626
rect 22376 11562 22428 11568
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21180 9648 21232 9654
rect 21376 9636 21404 11494
rect 22480 10810 22508 12786
rect 22664 12434 22692 16546
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22756 13462 22784 13670
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22756 13190 22784 13398
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22572 12406 22692 12434
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22112 10266 22140 10610
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22204 10198 22232 10406
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 21232 9608 21404 9636
rect 21180 9590 21232 9596
rect 20996 9444 21048 9450
rect 20996 9386 21048 9392
rect 21008 9042 21036 9386
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 21192 8974 21220 9590
rect 21548 9104 21600 9110
rect 21548 9046 21600 9052
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 21008 7750 21036 8230
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 21100 7410 21128 8774
rect 21192 8090 21220 8910
rect 21272 8900 21324 8906
rect 21272 8842 21324 8848
rect 21284 8090 21312 8842
rect 21454 8664 21510 8673
rect 21454 8599 21510 8608
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21376 8401 21404 8502
rect 21468 8498 21496 8599
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21362 8392 21418 8401
rect 21560 8362 21588 9046
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21652 8430 21680 8910
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21362 8327 21418 8336
rect 21548 8356 21600 8362
rect 21548 8298 21600 8304
rect 21836 8090 21864 8978
rect 22112 8498 22140 9998
rect 22296 9654 22324 10610
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22376 10260 22428 10266
rect 22376 10202 22428 10208
rect 22284 9648 22336 9654
rect 22284 9590 22336 9596
rect 22296 9178 22324 9590
rect 22388 9382 22416 10202
rect 22480 10062 22508 10542
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22376 9376 22428 9382
rect 22376 9318 22428 9324
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22284 8900 22336 8906
rect 22284 8842 22336 8848
rect 22296 8498 22324 8842
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 21272 8084 21324 8090
rect 21824 8084 21876 8090
rect 21324 8044 21404 8072
rect 21272 8026 21324 8032
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21192 7546 21220 7822
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21376 7478 21404 8044
rect 21824 8026 21876 8032
rect 21836 7478 21864 8026
rect 21928 8022 21956 8434
rect 22008 8356 22060 8362
rect 22008 8298 22060 8304
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21364 7472 21416 7478
rect 21364 7414 21416 7420
rect 21824 7472 21876 7478
rect 21824 7414 21876 7420
rect 22020 7426 22048 8298
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 21100 6934 21128 7346
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21088 6928 21140 6934
rect 21088 6870 21140 6876
rect 21100 5914 21128 6870
rect 21284 6866 21312 7278
rect 21376 6866 21404 7414
rect 22020 7398 22140 7426
rect 21640 7268 21692 7274
rect 21640 7210 21692 7216
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21560 6662 21588 6734
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21560 6390 21588 6598
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21652 5914 21680 7210
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 22020 5846 22048 7398
rect 22112 7002 22140 7398
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 22284 7268 22336 7274
rect 22284 7210 22336 7216
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22204 6882 22232 7210
rect 22112 6866 22232 6882
rect 22100 6860 22232 6866
rect 22152 6854 22232 6860
rect 22100 6802 22152 6808
rect 22296 6798 22324 7210
rect 22284 6792 22336 6798
rect 22112 6740 22284 6746
rect 22112 6734 22336 6740
rect 22112 6718 22324 6734
rect 22468 6724 22520 6730
rect 20996 5840 21048 5846
rect 20996 5782 21048 5788
rect 22008 5840 22060 5846
rect 22008 5782 22060 5788
rect 21008 5574 21036 5782
rect 22020 5710 22048 5782
rect 22008 5704 22060 5710
rect 22008 5646 22060 5652
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21376 4622 21404 5102
rect 21468 5098 21496 5510
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 21456 5092 21508 5098
rect 21456 5034 21508 5040
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21928 4554 21956 5170
rect 22020 4622 22048 5510
rect 22112 5234 22140 6718
rect 22468 6666 22520 6672
rect 22480 6458 22508 6666
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 21916 4548 21968 4554
rect 21916 4490 21968 4496
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 21008 3058 21036 4422
rect 21928 4282 21956 4490
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21284 3738 21312 4082
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 21560 3738 21588 4014
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21560 3534 21588 3674
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 21836 3482 21864 3606
rect 22008 3528 22060 3534
rect 21836 3476 22008 3482
rect 21836 3470 22060 3476
rect 21272 3460 21324 3466
rect 21272 3402 21324 3408
rect 21836 3454 22048 3470
rect 21284 3194 21312 3402
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 21836 2446 21864 3454
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22020 2446 22048 3334
rect 22204 3058 22232 6054
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22284 5296 22336 5302
rect 22284 5238 22336 5244
rect 22296 4554 22324 5238
rect 22388 5234 22416 5850
rect 22376 5228 22428 5234
rect 22376 5170 22428 5176
rect 22468 4820 22520 4826
rect 22468 4762 22520 4768
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22284 4548 22336 4554
rect 22284 4490 22336 4496
rect 22388 4282 22416 4558
rect 22480 4486 22508 4762
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22468 4004 22520 4010
rect 22468 3946 22520 3952
rect 22480 3738 22508 3946
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 21192 870 21312 898
rect 21192 762 21220 870
rect 21284 800 21312 870
rect 22572 800 22600 12406
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22652 11756 22704 11762
rect 22756 11744 22784 12174
rect 22704 11716 22784 11744
rect 22652 11698 22704 11704
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22664 10130 22692 10610
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22756 9110 22784 9454
rect 22744 9104 22796 9110
rect 22744 9046 22796 9052
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 22664 6934 22692 7278
rect 22652 6928 22704 6934
rect 22652 6870 22704 6876
rect 22664 6458 22692 6870
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22664 5710 22692 6394
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22848 5250 22876 16546
rect 23032 14074 23060 19654
rect 23124 19334 23152 20742
rect 23216 19922 23244 20878
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23308 20058 23336 20334
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23216 19786 23244 19858
rect 23204 19780 23256 19786
rect 23204 19722 23256 19728
rect 23400 19446 23428 20538
rect 23388 19440 23440 19446
rect 23388 19382 23440 19388
rect 23124 19306 23336 19334
rect 23112 18692 23164 18698
rect 23112 18634 23164 18640
rect 23124 18426 23152 18634
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23216 17678 23244 18022
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23216 16250 23244 17478
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 23216 15434 23244 16186
rect 23204 15428 23256 15434
rect 23204 15370 23256 15376
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 23308 13734 23336 19306
rect 23400 18358 23428 19382
rect 23480 18896 23532 18902
rect 23480 18838 23532 18844
rect 23388 18352 23440 18358
rect 23388 18294 23440 18300
rect 23400 17746 23428 18294
rect 23492 18222 23520 18838
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23492 16794 23520 17070
rect 23480 16788 23532 16794
rect 23480 16730 23532 16736
rect 23388 16584 23440 16590
rect 23676 16538 23704 23038
rect 23768 22642 23796 23122
rect 23860 22982 23888 23258
rect 23848 22976 23900 22982
rect 23848 22918 23900 22924
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 24136 22098 24164 24550
rect 24563 24508 24871 24528
rect 24563 24506 24569 24508
rect 24625 24506 24649 24508
rect 24705 24506 24729 24508
rect 24785 24506 24809 24508
rect 24865 24506 24871 24508
rect 24625 24454 24627 24506
rect 24807 24454 24809 24506
rect 24563 24452 24569 24454
rect 24625 24452 24649 24454
rect 24705 24452 24729 24454
rect 24785 24452 24809 24454
rect 24865 24452 24871 24454
rect 24563 24432 24871 24452
rect 24400 24200 24452 24206
rect 24400 24142 24452 24148
rect 24412 23866 24440 24142
rect 25056 24138 25084 24686
rect 25044 24132 25096 24138
rect 25044 24074 25096 24080
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24400 23860 24452 23866
rect 24400 23802 24452 23808
rect 24596 23798 24624 24006
rect 24584 23792 24636 23798
rect 24584 23734 24636 23740
rect 24563 23420 24871 23440
rect 24563 23418 24569 23420
rect 24625 23418 24649 23420
rect 24705 23418 24729 23420
rect 24785 23418 24809 23420
rect 24865 23418 24871 23420
rect 24625 23366 24627 23418
rect 24807 23366 24809 23418
rect 24563 23364 24569 23366
rect 24625 23364 24649 23366
rect 24705 23364 24729 23366
rect 24785 23364 24809 23366
rect 24865 23364 24871 23366
rect 24563 23344 24871 23364
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 24216 22976 24268 22982
rect 24216 22918 24268 22924
rect 24228 22574 24256 22918
rect 24216 22568 24268 22574
rect 24216 22510 24268 22516
rect 24124 22092 24176 22098
rect 24176 22052 24256 22080
rect 24124 22034 24176 22040
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 23860 21690 23888 21966
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 23848 21684 23900 21690
rect 23848 21626 23900 21632
rect 24044 21622 24072 21830
rect 24032 21616 24084 21622
rect 24032 21558 24084 21564
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 23952 19854 23980 20878
rect 24136 20534 24164 21014
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 23940 19848 23992 19854
rect 23940 19790 23992 19796
rect 23952 18970 23980 19790
rect 24032 19712 24084 19718
rect 24032 19654 24084 19660
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23940 18964 23992 18970
rect 23940 18906 23992 18912
rect 23768 18834 23796 18906
rect 24044 18850 24072 19654
rect 23756 18828 23808 18834
rect 23756 18770 23808 18776
rect 23952 18822 24072 18850
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 23860 16794 23888 17206
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23388 16526 23440 16532
rect 23400 16250 23428 16526
rect 23492 16522 23704 16538
rect 23480 16516 23704 16522
rect 23532 16510 23704 16516
rect 23480 16458 23532 16464
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23584 16250 23612 16390
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23584 15502 23612 16186
rect 23676 16182 23704 16510
rect 23664 16176 23716 16182
rect 23664 16118 23716 16124
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23952 15162 23980 18822
rect 24228 18748 24256 22052
rect 24412 20058 24440 23258
rect 24563 22332 24871 22352
rect 24563 22330 24569 22332
rect 24625 22330 24649 22332
rect 24705 22330 24729 22332
rect 24785 22330 24809 22332
rect 24865 22330 24871 22332
rect 24625 22278 24627 22330
rect 24807 22278 24809 22330
rect 24563 22276 24569 22278
rect 24625 22276 24649 22278
rect 24705 22276 24729 22278
rect 24785 22276 24809 22278
rect 24865 22276 24871 22278
rect 24563 22256 24871 22276
rect 25228 21956 25280 21962
rect 25228 21898 25280 21904
rect 25240 21350 25268 21898
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 24563 21244 24871 21264
rect 24563 21242 24569 21244
rect 24625 21242 24649 21244
rect 24705 21242 24729 21244
rect 24785 21242 24809 21244
rect 24865 21242 24871 21244
rect 24625 21190 24627 21242
rect 24807 21190 24809 21242
rect 24563 21188 24569 21190
rect 24625 21188 24649 21190
rect 24705 21188 24729 21190
rect 24785 21188 24809 21190
rect 24865 21188 24871 21190
rect 24563 21168 24871 21188
rect 25136 20528 25188 20534
rect 25136 20470 25188 20476
rect 24563 20156 24871 20176
rect 24563 20154 24569 20156
rect 24625 20154 24649 20156
rect 24705 20154 24729 20156
rect 24785 20154 24809 20156
rect 24865 20154 24871 20156
rect 24625 20102 24627 20154
rect 24807 20102 24809 20154
rect 24563 20100 24569 20102
rect 24625 20100 24649 20102
rect 24705 20100 24729 20102
rect 24785 20100 24809 20102
rect 24865 20100 24871 20102
rect 24563 20080 24871 20100
rect 25148 20058 25176 20470
rect 24400 20052 24452 20058
rect 24400 19994 24452 20000
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 24412 19718 24440 19994
rect 25044 19984 25096 19990
rect 25044 19926 25096 19932
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24400 19712 24452 19718
rect 24400 19654 24452 19660
rect 24688 19514 24716 19790
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 25056 19446 25084 19926
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 24504 18766 24532 19314
rect 24563 19068 24871 19088
rect 24563 19066 24569 19068
rect 24625 19066 24649 19068
rect 24705 19066 24729 19068
rect 24785 19066 24809 19068
rect 24865 19066 24871 19068
rect 24625 19014 24627 19066
rect 24807 19014 24809 19066
rect 24563 19012 24569 19014
rect 24625 19012 24649 19014
rect 24705 19012 24729 19014
rect 24785 19012 24809 19014
rect 24865 19012 24871 19014
rect 24563 18992 24871 19012
rect 24044 18720 24256 18748
rect 24492 18760 24544 18766
rect 24044 15638 24072 18720
rect 24492 18702 24544 18708
rect 24400 17740 24452 17746
rect 24400 17682 24452 17688
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24228 17270 24256 17478
rect 24216 17264 24268 17270
rect 24216 17206 24268 17212
rect 24124 16448 24176 16454
rect 24124 16390 24176 16396
rect 24136 16182 24164 16390
rect 24228 16250 24256 17206
rect 24412 17134 24440 17682
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 24308 16992 24360 16998
rect 24308 16934 24360 16940
rect 24320 16590 24348 16934
rect 24308 16584 24360 16590
rect 24308 16526 24360 16532
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 24124 16176 24176 16182
rect 24124 16118 24176 16124
rect 24032 15632 24084 15638
rect 24032 15574 24084 15580
rect 24044 15162 24072 15574
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 23296 13728 23348 13734
rect 23296 13670 23348 13676
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12918 23336 13126
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 22940 10674 22968 12174
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 22940 9926 22968 10610
rect 23020 10532 23072 10538
rect 23020 10474 23072 10480
rect 23032 10146 23060 10474
rect 23124 10266 23152 10610
rect 23216 10606 23244 11698
rect 23204 10600 23256 10606
rect 23204 10542 23256 10548
rect 23308 10470 23336 12854
rect 23400 12306 23428 13806
rect 23676 13530 23704 13874
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 24044 13462 24072 15098
rect 24136 13734 24164 16118
rect 24228 15366 24256 16186
rect 24320 15502 24348 16526
rect 24412 16114 24440 17070
rect 24504 16708 24532 18702
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24964 18358 24992 18566
rect 24952 18352 25004 18358
rect 24952 18294 25004 18300
rect 24563 17980 24871 18000
rect 24563 17978 24569 17980
rect 24625 17978 24649 17980
rect 24705 17978 24729 17980
rect 24785 17978 24809 17980
rect 24865 17978 24871 17980
rect 24625 17926 24627 17978
rect 24807 17926 24809 17978
rect 24563 17924 24569 17926
rect 24625 17924 24649 17926
rect 24705 17924 24729 17926
rect 24785 17924 24809 17926
rect 24865 17924 24871 17926
rect 24563 17904 24871 17924
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 24780 17270 24808 17478
rect 24768 17264 24820 17270
rect 24766 17232 24768 17241
rect 24820 17232 24822 17241
rect 24766 17167 24822 17176
rect 24872 17066 24900 17546
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24860 17060 24912 17066
rect 24860 17002 24912 17008
rect 24563 16892 24871 16912
rect 24563 16890 24569 16892
rect 24625 16890 24649 16892
rect 24705 16890 24729 16892
rect 24785 16890 24809 16892
rect 24865 16890 24871 16892
rect 24625 16838 24627 16890
rect 24807 16838 24809 16890
rect 24563 16836 24569 16838
rect 24625 16836 24649 16838
rect 24705 16836 24729 16838
rect 24785 16836 24809 16838
rect 24865 16836 24871 16838
rect 24563 16816 24871 16836
rect 24504 16680 24624 16708
rect 24492 16516 24544 16522
rect 24492 16458 24544 16464
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24504 15706 24532 16458
rect 24596 16454 24624 16680
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 24563 15804 24871 15824
rect 24563 15802 24569 15804
rect 24625 15802 24649 15804
rect 24705 15802 24729 15804
rect 24785 15802 24809 15804
rect 24865 15802 24871 15804
rect 24625 15750 24627 15802
rect 24807 15750 24809 15802
rect 24563 15748 24569 15750
rect 24625 15748 24649 15750
rect 24705 15748 24729 15750
rect 24785 15748 24809 15750
rect 24865 15748 24871 15750
rect 24563 15728 24871 15748
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24308 15496 24360 15502
rect 24308 15438 24360 15444
rect 24216 15360 24268 15366
rect 24216 15302 24268 15308
rect 24504 15026 24532 15642
rect 24860 15496 24912 15502
rect 24964 15484 24992 17138
rect 25240 16574 25268 21286
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 25332 16794 25360 17138
rect 25320 16788 25372 16794
rect 25320 16730 25372 16736
rect 25240 16546 25360 16574
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 25240 15706 25268 15982
rect 25228 15700 25280 15706
rect 25228 15642 25280 15648
rect 25044 15632 25096 15638
rect 25044 15574 25096 15580
rect 24912 15456 24992 15484
rect 24860 15438 24912 15444
rect 25056 15094 25084 15574
rect 25136 15360 25188 15366
rect 25136 15302 25188 15308
rect 25044 15088 25096 15094
rect 25044 15030 25096 15036
rect 24492 15020 24544 15026
rect 24492 14962 24544 14968
rect 24563 14716 24871 14736
rect 24563 14714 24569 14716
rect 24625 14714 24649 14716
rect 24705 14714 24729 14716
rect 24785 14714 24809 14716
rect 24865 14714 24871 14716
rect 24625 14662 24627 14714
rect 24807 14662 24809 14714
rect 24563 14660 24569 14662
rect 24625 14660 24649 14662
rect 24705 14660 24729 14662
rect 24785 14660 24809 14662
rect 24865 14660 24871 14662
rect 24563 14640 24871 14660
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 24124 13728 24176 13734
rect 24124 13670 24176 13676
rect 24032 13456 24084 13462
rect 24032 13398 24084 13404
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 23952 12986 23980 13262
rect 24044 13190 24072 13398
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 23388 12300 23440 12306
rect 23388 12242 23440 12248
rect 23400 11762 23428 12242
rect 23584 12238 23612 12922
rect 23952 12850 23980 12922
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 23664 12708 23716 12714
rect 23664 12650 23716 12656
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 23676 12170 23704 12650
rect 23848 12232 23900 12238
rect 24044 12186 24072 13126
rect 24136 12918 24164 13670
rect 24563 13628 24871 13648
rect 24563 13626 24569 13628
rect 24625 13626 24649 13628
rect 24705 13626 24729 13628
rect 24785 13626 24809 13628
rect 24865 13626 24871 13628
rect 24625 13574 24627 13626
rect 24807 13574 24809 13626
rect 24563 13572 24569 13574
rect 24625 13572 24649 13574
rect 24705 13572 24729 13574
rect 24785 13572 24809 13574
rect 24865 13572 24871 13574
rect 24563 13552 24871 13572
rect 25056 13530 25084 13874
rect 25148 13734 25176 15302
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 24504 13410 24532 13466
rect 24504 13382 24624 13410
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24504 13190 24532 13262
rect 24596 13258 24624 13382
rect 25148 13258 25176 13670
rect 24584 13252 24636 13258
rect 24584 13194 24636 13200
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 25136 13252 25188 13258
rect 25136 13194 25188 13200
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24124 12912 24176 12918
rect 24124 12854 24176 12860
rect 24504 12850 24532 13126
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 24504 12730 24532 12786
rect 24412 12702 24532 12730
rect 24688 12714 24716 13194
rect 24676 12708 24728 12714
rect 24412 12238 24440 12702
rect 24676 12650 24728 12656
rect 24492 12640 24544 12646
rect 24492 12582 24544 12588
rect 23900 12180 24072 12186
rect 23848 12174 24072 12180
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 23664 12164 23716 12170
rect 23860 12158 24072 12174
rect 23664 12106 23716 12112
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23296 10464 23348 10470
rect 23296 10406 23348 10412
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23204 10192 23256 10198
rect 23032 10118 23152 10146
rect 23204 10134 23256 10140
rect 23124 9994 23152 10118
rect 23216 10062 23244 10134
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 23112 9988 23164 9994
rect 23112 9930 23164 9936
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22940 9178 22968 9862
rect 23216 9586 23244 9998
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23020 9444 23072 9450
rect 23020 9386 23072 9392
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 23032 8974 23060 9386
rect 23308 8974 23336 9590
rect 23400 9382 23428 9998
rect 23492 9874 23520 10542
rect 23572 9920 23624 9926
rect 23492 9868 23572 9874
rect 23492 9862 23624 9868
rect 23492 9846 23612 9862
rect 23492 9722 23520 9846
rect 23480 9716 23532 9722
rect 23480 9658 23532 9664
rect 23676 9489 23704 12106
rect 24044 12102 24072 12158
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24504 11898 24532 12582
rect 24563 12540 24871 12560
rect 24563 12538 24569 12540
rect 24625 12538 24649 12540
rect 24705 12538 24729 12540
rect 24785 12538 24809 12540
rect 24865 12538 24871 12540
rect 24625 12486 24627 12538
rect 24807 12486 24809 12538
rect 24563 12484 24569 12486
rect 24625 12484 24649 12486
rect 24705 12484 24729 12486
rect 24785 12484 24809 12486
rect 24865 12484 24871 12486
rect 24563 12464 24871 12484
rect 25332 12434 25360 16546
rect 25424 15366 25452 25638
rect 25780 25424 25832 25430
rect 25780 25366 25832 25372
rect 25792 25294 25820 25366
rect 27080 25362 27108 25774
rect 27172 25498 27200 25842
rect 27160 25492 27212 25498
rect 27160 25434 27212 25440
rect 27068 25356 27120 25362
rect 27068 25298 27120 25304
rect 25780 25288 25832 25294
rect 25780 25230 25832 25236
rect 25872 25288 25924 25294
rect 25872 25230 25924 25236
rect 25596 25220 25648 25226
rect 25596 25162 25648 25168
rect 25608 22234 25636 25162
rect 25688 25152 25740 25158
rect 25688 25094 25740 25100
rect 25700 24818 25728 25094
rect 25884 24954 25912 25230
rect 25872 24948 25924 24954
rect 25872 24890 25924 24896
rect 25884 24818 25912 24890
rect 26700 24880 26752 24886
rect 26700 24822 26752 24828
rect 25688 24812 25740 24818
rect 25688 24754 25740 24760
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 26712 24614 26740 24822
rect 25780 24608 25832 24614
rect 25780 24550 25832 24556
rect 26516 24608 26568 24614
rect 26516 24550 26568 24556
rect 26700 24608 26752 24614
rect 26700 24550 26752 24556
rect 25792 24274 25820 24550
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 25780 24268 25832 24274
rect 25780 24210 25832 24216
rect 26252 24041 26280 24346
rect 26528 24138 26556 24550
rect 26516 24132 26568 24138
rect 26516 24074 26568 24080
rect 26712 24070 26740 24550
rect 26700 24064 26752 24070
rect 26238 24032 26294 24041
rect 26700 24006 26752 24012
rect 27620 24064 27672 24070
rect 27620 24006 27672 24012
rect 26238 23967 26294 23976
rect 26252 23866 26280 23967
rect 26240 23860 26292 23866
rect 26240 23802 26292 23808
rect 26332 23520 26384 23526
rect 26332 23462 26384 23468
rect 26240 23044 26292 23050
rect 26240 22986 26292 22992
rect 26252 22438 26280 22986
rect 26240 22432 26292 22438
rect 26240 22374 26292 22380
rect 25596 22228 25648 22234
rect 25596 22170 25648 22176
rect 25608 21026 25636 22170
rect 25608 20998 25728 21026
rect 25596 20868 25648 20874
rect 25596 20810 25648 20816
rect 25608 20602 25636 20810
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25504 17604 25556 17610
rect 25504 17546 25556 17552
rect 25516 17338 25544 17546
rect 25700 17338 25728 20998
rect 26056 19440 26108 19446
rect 26056 19382 26108 19388
rect 26068 18970 26096 19382
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 25504 17332 25556 17338
rect 25504 17274 25556 17280
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25700 17134 25728 17274
rect 25688 17128 25740 17134
rect 25688 17070 25740 17076
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 25596 15088 25648 15094
rect 25596 15030 25648 15036
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25424 14414 25452 14758
rect 25608 14618 25636 15030
rect 25596 14612 25648 14618
rect 25596 14554 25648 14560
rect 25412 14408 25464 14414
rect 25412 14350 25464 14356
rect 25700 12850 25728 17070
rect 26252 16574 26280 22374
rect 26344 22137 26372 23462
rect 26330 22128 26386 22137
rect 26330 22063 26386 22072
rect 27526 20224 27582 20233
rect 27526 20159 27582 20168
rect 27540 19786 27568 20159
rect 26516 19780 26568 19786
rect 26516 19722 26568 19728
rect 27528 19780 27580 19786
rect 27528 19722 27580 19728
rect 26528 19514 26556 19722
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 27632 16574 27660 24006
rect 26252 16546 27108 16574
rect 27632 16546 28304 16574
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26160 16250 26188 16390
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26528 14822 26556 15506
rect 26804 15502 26832 15846
rect 26792 15496 26844 15502
rect 26792 15438 26844 15444
rect 26516 14816 26568 14822
rect 26516 14758 26568 14764
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25240 12406 25360 12434
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23952 10674 23980 11494
rect 24563 11452 24871 11472
rect 24563 11450 24569 11452
rect 24625 11450 24649 11452
rect 24705 11450 24729 11452
rect 24785 11450 24809 11452
rect 24865 11450 24871 11452
rect 24625 11398 24627 11450
rect 24807 11398 24809 11450
rect 24563 11396 24569 11398
rect 24625 11396 24649 11398
rect 24705 11396 24729 11398
rect 24785 11396 24809 11398
rect 24865 11396 24871 11398
rect 24563 11376 24871 11396
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 23768 9994 23796 10406
rect 23848 10192 23900 10198
rect 23848 10134 23900 10140
rect 23756 9988 23808 9994
rect 23756 9930 23808 9936
rect 23662 9480 23718 9489
rect 23662 9415 23718 9424
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23768 8906 23796 9930
rect 23860 8974 23888 10134
rect 23952 10062 23980 10610
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 24504 9450 24532 10542
rect 24563 10364 24871 10384
rect 24563 10362 24569 10364
rect 24625 10362 24649 10364
rect 24705 10362 24729 10364
rect 24785 10362 24809 10364
rect 24865 10362 24871 10364
rect 24625 10310 24627 10362
rect 24807 10310 24809 10362
rect 24563 10308 24569 10310
rect 24625 10308 24649 10310
rect 24705 10308 24729 10310
rect 24785 10308 24809 10310
rect 24865 10308 24871 10310
rect 24563 10288 24871 10308
rect 24964 10266 24992 10610
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24952 10260 25004 10266
rect 24952 10202 25004 10208
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24780 9586 24808 9862
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 24492 9444 24544 9450
rect 24492 9386 24544 9392
rect 24563 9276 24871 9296
rect 24563 9274 24569 9276
rect 24625 9274 24649 9276
rect 24705 9274 24729 9276
rect 24785 9274 24809 9276
rect 24865 9274 24871 9276
rect 24625 9222 24627 9274
rect 24807 9222 24809 9274
rect 24563 9220 24569 9222
rect 24625 9220 24649 9222
rect 24705 9220 24729 9222
rect 24785 9220 24809 9222
rect 24865 9220 24871 9222
rect 24563 9200 24871 9220
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23756 8900 23808 8906
rect 23756 8842 23808 8848
rect 23112 8832 23164 8838
rect 23112 8774 23164 8780
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 23032 7954 23060 8570
rect 23124 8362 23152 8774
rect 24044 8634 24072 8910
rect 24964 8906 24992 10066
rect 25056 9586 25084 10406
rect 25136 9988 25188 9994
rect 25136 9930 25188 9936
rect 25044 9580 25096 9586
rect 25044 9522 25096 9528
rect 25148 9518 25176 9930
rect 25136 9512 25188 9518
rect 25136 9454 25188 9460
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 24136 8498 24164 8774
rect 24124 8492 24176 8498
rect 24124 8434 24176 8440
rect 24492 8492 24544 8498
rect 24492 8434 24544 8440
rect 24504 8401 24532 8434
rect 24490 8392 24546 8401
rect 23112 8356 23164 8362
rect 24490 8327 24546 8336
rect 23112 8298 23164 8304
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23124 7834 23152 8298
rect 23204 8288 23256 8294
rect 23204 8230 23256 8236
rect 23032 7806 23152 7834
rect 23032 7410 23060 7806
rect 23216 7410 23244 8230
rect 24504 7954 24532 8327
rect 24563 8188 24871 8208
rect 24563 8186 24569 8188
rect 24625 8186 24649 8188
rect 24705 8186 24729 8188
rect 24785 8186 24809 8188
rect 24865 8186 24871 8188
rect 24625 8134 24627 8186
rect 24807 8134 24809 8186
rect 24563 8132 24569 8134
rect 24625 8132 24649 8134
rect 24705 8132 24729 8134
rect 24785 8132 24809 8134
rect 24865 8132 24871 8134
rect 24563 8112 24871 8132
rect 24492 7948 24544 7954
rect 24412 7908 24492 7936
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23400 7410 23428 7686
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23940 7404 23992 7410
rect 23940 7346 23992 7352
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 22940 6458 22968 6802
rect 22928 6452 22980 6458
rect 22928 6394 22980 6400
rect 23032 6186 23060 7346
rect 23480 7336 23532 7342
rect 23480 7278 23532 7284
rect 23388 7268 23440 7274
rect 23388 7210 23440 7216
rect 23400 6934 23428 7210
rect 23388 6928 23440 6934
rect 23388 6870 23440 6876
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23216 6322 23244 6734
rect 23400 6338 23428 6870
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23308 6310 23428 6338
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 22756 5222 22876 5250
rect 22756 3942 22784 5222
rect 22836 5160 22888 5166
rect 22836 5102 22888 5108
rect 22848 4826 22876 5102
rect 23032 5098 23060 6122
rect 23020 5092 23072 5098
rect 23020 5034 23072 5040
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 22940 4826 22968 4966
rect 22836 4820 22888 4826
rect 22836 4762 22888 4768
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 23216 3738 23244 6258
rect 23308 5914 23336 6310
rect 23388 6248 23440 6254
rect 23388 6190 23440 6196
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 23400 5846 23428 6190
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23400 4486 23428 5170
rect 23492 4622 23520 7278
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23768 5234 23796 5510
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23584 4690 23612 4966
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23388 4480 23440 4486
rect 23388 4422 23440 4428
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23492 4282 23520 4422
rect 23584 4282 23612 4626
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 23952 4146 23980 7346
rect 24124 6180 24176 6186
rect 24124 6122 24176 6128
rect 24136 5914 24164 6122
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24320 5778 24348 7346
rect 24412 6118 24440 7908
rect 24492 7890 24544 7896
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24688 7478 24716 7822
rect 24964 7818 24992 8842
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24780 7546 24808 7686
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 24563 7100 24871 7120
rect 24563 7098 24569 7100
rect 24625 7098 24649 7100
rect 24705 7098 24729 7100
rect 24785 7098 24809 7100
rect 24865 7098 24871 7100
rect 24625 7046 24627 7098
rect 24807 7046 24809 7098
rect 24563 7044 24569 7046
rect 24625 7044 24649 7046
rect 24705 7044 24729 7046
rect 24785 7044 24809 7046
rect 24865 7044 24871 7046
rect 24563 7024 24871 7044
rect 24860 6928 24912 6934
rect 24780 6876 24860 6882
rect 24780 6870 24912 6876
rect 24780 6854 24900 6870
rect 24780 6458 24808 6854
rect 24964 6730 24992 7754
rect 25044 6792 25096 6798
rect 25044 6734 25096 6740
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24872 6322 24900 6598
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 24492 6248 24544 6254
rect 24492 6190 24544 6196
rect 24400 6112 24452 6118
rect 24400 6054 24452 6060
rect 24412 5914 24440 6054
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24308 5772 24360 5778
rect 24308 5714 24360 5720
rect 24124 5704 24176 5710
rect 24124 5646 24176 5652
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 24136 5302 24164 5646
rect 24412 5370 24440 5646
rect 24400 5364 24452 5370
rect 24400 5306 24452 5312
rect 24124 5296 24176 5302
rect 24504 5250 24532 6190
rect 24563 6012 24871 6032
rect 24563 6010 24569 6012
rect 24625 6010 24649 6012
rect 24705 6010 24729 6012
rect 24785 6010 24809 6012
rect 24865 6010 24871 6012
rect 24625 5958 24627 6010
rect 24807 5958 24809 6010
rect 24563 5956 24569 5958
rect 24625 5956 24649 5958
rect 24705 5956 24729 5958
rect 24785 5956 24809 5958
rect 24865 5956 24871 5958
rect 24563 5936 24871 5956
rect 24768 5840 24820 5846
rect 24768 5782 24820 5788
rect 24124 5238 24176 5244
rect 24136 4622 24164 5238
rect 24412 5222 24532 5250
rect 24780 5234 24808 5782
rect 24768 5228 24820 5234
rect 24412 4690 24440 5222
rect 24768 5170 24820 5176
rect 24492 5092 24544 5098
rect 24492 5034 24544 5040
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 24124 4616 24176 4622
rect 24124 4558 24176 4564
rect 24504 4554 24532 5034
rect 24563 4924 24871 4944
rect 24563 4922 24569 4924
rect 24625 4922 24649 4924
rect 24705 4922 24729 4924
rect 24785 4922 24809 4924
rect 24865 4922 24871 4924
rect 24625 4870 24627 4922
rect 24807 4870 24809 4922
rect 24563 4868 24569 4870
rect 24625 4868 24649 4870
rect 24705 4868 24729 4870
rect 24785 4868 24809 4870
rect 24865 4868 24871 4870
rect 24563 4848 24871 4868
rect 24492 4548 24544 4554
rect 24492 4490 24544 4496
rect 24124 4480 24176 4486
rect 24124 4422 24176 4428
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 23584 3210 23612 3470
rect 23756 3460 23808 3466
rect 23756 3402 23808 3408
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23492 3194 23612 3210
rect 23492 3188 23624 3194
rect 23492 3182 23572 3188
rect 23492 2582 23520 3182
rect 23572 3130 23624 3136
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 23584 2378 23612 2994
rect 23572 2372 23624 2378
rect 23572 2314 23624 2320
rect 23676 2310 23704 3334
rect 23768 2446 23796 3402
rect 23860 2922 23888 3470
rect 23952 3194 23980 4082
rect 23940 3188 23992 3194
rect 23940 3130 23992 3136
rect 23938 3088 23994 3097
rect 24136 3058 24164 4422
rect 24964 3942 24992 6666
rect 25056 5234 25084 6734
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25148 6458 25176 6598
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 25056 4826 25084 5170
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25136 4480 25188 4486
rect 25136 4422 25188 4428
rect 25148 4214 25176 4422
rect 25136 4208 25188 4214
rect 25136 4150 25188 4156
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24563 3836 24871 3856
rect 24563 3834 24569 3836
rect 24625 3834 24649 3836
rect 24705 3834 24729 3836
rect 24785 3834 24809 3836
rect 24865 3834 24871 3836
rect 24625 3782 24627 3834
rect 24807 3782 24809 3834
rect 24563 3780 24569 3782
rect 24625 3780 24649 3782
rect 24705 3780 24729 3782
rect 24785 3780 24809 3782
rect 24865 3780 24871 3782
rect 24563 3760 24871 3780
rect 24964 3126 24992 3878
rect 24952 3120 25004 3126
rect 24952 3062 25004 3068
rect 23938 3023 23994 3032
rect 24124 3052 24176 3058
rect 23848 2916 23900 2922
rect 23848 2858 23900 2864
rect 23860 2514 23888 2858
rect 23848 2508 23900 2514
rect 23848 2450 23900 2456
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23664 2304 23716 2310
rect 23664 2246 23716 2252
rect 23952 1442 23980 3023
rect 24124 2994 24176 3000
rect 25240 2938 25268 12406
rect 25424 11558 25452 12786
rect 26528 12481 26556 14758
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26514 12472 26570 12481
rect 26514 12407 26570 12416
rect 25412 11552 25464 11558
rect 25412 11494 25464 11500
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25504 10668 25556 10674
rect 25504 10610 25556 10616
rect 25516 9926 25544 10610
rect 25504 9920 25556 9926
rect 25504 9862 25556 9868
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 25516 9722 25544 9862
rect 25504 9716 25556 9722
rect 25504 9658 25556 9664
rect 25608 9586 25636 9862
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 25516 9178 25544 9454
rect 25504 9172 25556 9178
rect 25504 9114 25556 9120
rect 25884 8090 25912 11494
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 26252 10577 26280 11290
rect 26238 10568 26294 10577
rect 26238 10503 26294 10512
rect 26712 8673 26740 14418
rect 26804 14385 26832 15438
rect 26790 14376 26846 14385
rect 26790 14311 26846 14320
rect 26698 8664 26754 8673
rect 26698 8599 26754 8608
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25780 7404 25832 7410
rect 25780 7346 25832 7352
rect 25792 7002 25820 7346
rect 25964 7200 26016 7206
rect 25964 7142 26016 7148
rect 25780 6996 25832 7002
rect 25780 6938 25832 6944
rect 25320 6792 25372 6798
rect 25320 6734 25372 6740
rect 25332 6458 25360 6734
rect 25504 6724 25556 6730
rect 25504 6666 25556 6672
rect 25688 6724 25740 6730
rect 25688 6666 25740 6672
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25516 6322 25544 6666
rect 25504 6316 25556 6322
rect 25504 6258 25556 6264
rect 25700 5778 25728 6666
rect 25976 6458 26004 7142
rect 26238 6760 26294 6769
rect 26238 6695 26294 6704
rect 25964 6452 26016 6458
rect 25964 6394 26016 6400
rect 26252 6390 26280 6695
rect 26240 6384 26292 6390
rect 26240 6326 26292 6332
rect 25964 6248 26016 6254
rect 25964 6190 26016 6196
rect 25688 5772 25740 5778
rect 25688 5714 25740 5720
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 25608 5234 25636 5646
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25608 4826 25636 5170
rect 25976 4826 26004 6190
rect 26424 5636 26476 5642
rect 26424 5578 26476 5584
rect 26436 5234 26464 5578
rect 26424 5228 26476 5234
rect 26424 5170 26476 5176
rect 26884 5024 26936 5030
rect 26884 4966 26936 4972
rect 26238 4856 26294 4865
rect 25596 4820 25648 4826
rect 25596 4762 25648 4768
rect 25964 4820 26016 4826
rect 26238 4791 26294 4800
rect 25964 4762 26016 4768
rect 26252 4758 26280 4791
rect 26240 4752 26292 4758
rect 26240 4694 26292 4700
rect 26896 4690 26924 4966
rect 25872 4684 25924 4690
rect 25872 4626 25924 4632
rect 26884 4684 26936 4690
rect 26884 4626 26936 4632
rect 25884 3602 25912 4626
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26252 4282 26280 4422
rect 26240 4276 26292 4282
rect 26240 4218 26292 4224
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 24964 2910 25268 2938
rect 24563 2748 24871 2768
rect 24563 2746 24569 2748
rect 24625 2746 24649 2748
rect 24705 2746 24729 2748
rect 24785 2746 24809 2748
rect 24865 2746 24871 2748
rect 24625 2694 24627 2746
rect 24807 2694 24809 2746
rect 24563 2692 24569 2694
rect 24625 2692 24649 2694
rect 24705 2692 24729 2694
rect 24785 2692 24809 2694
rect 24865 2692 24871 2694
rect 24563 2672 24871 2692
rect 23768 1414 23980 1442
rect 23768 800 23796 1414
rect 24964 800 24992 2910
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 25240 2582 25268 2790
rect 25792 2650 25820 2994
rect 25884 2990 25912 3538
rect 26528 3534 26556 4082
rect 26792 3732 26844 3738
rect 26792 3674 26844 3680
rect 26516 3528 26568 3534
rect 25962 3496 26018 3505
rect 26516 3470 26568 3476
rect 25962 3431 26018 3440
rect 25872 2984 25924 2990
rect 25872 2926 25924 2932
rect 25780 2644 25832 2650
rect 25780 2586 25832 2592
rect 25228 2576 25280 2582
rect 25228 2518 25280 2524
rect 25976 1442 26004 3431
rect 26056 3052 26108 3058
rect 26056 2994 26108 3000
rect 26068 2582 26096 2994
rect 26148 2984 26200 2990
rect 26148 2926 26200 2932
rect 26330 2952 26386 2961
rect 26056 2576 26108 2582
rect 26056 2518 26108 2524
rect 26160 2378 26188 2926
rect 26330 2887 26332 2896
rect 26384 2887 26386 2896
rect 26332 2858 26384 2864
rect 26528 2650 26556 3470
rect 26804 3058 26832 3674
rect 26792 3052 26844 3058
rect 26792 2994 26844 3000
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 26148 2372 26200 2378
rect 26148 2314 26200 2320
rect 25976 1414 26188 1442
rect 26160 800 26188 1414
rect 26240 1352 26292 1358
rect 26240 1294 26292 1300
rect 26252 1057 26280 1294
rect 26238 1048 26294 1057
rect 26238 983 26294 992
rect 20916 734 21220 762
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 23754 0 23810 800
rect 24950 0 25006 800
rect 26146 0 26202 800
rect 27080 762 27108 16546
rect 27712 6656 27764 6662
rect 27712 6598 27764 6604
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27264 4622 27292 5306
rect 27724 5234 27752 6598
rect 27436 5228 27488 5234
rect 27436 5170 27488 5176
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 27344 5092 27396 5098
rect 27344 5034 27396 5040
rect 27356 4758 27384 5034
rect 27344 4752 27396 4758
rect 27344 4694 27396 4700
rect 27252 4616 27304 4622
rect 27252 4558 27304 4564
rect 27264 4282 27292 4558
rect 27252 4276 27304 4282
rect 27252 4218 27304 4224
rect 27356 3738 27384 4694
rect 27448 4690 27476 5170
rect 27528 5160 27580 5166
rect 27528 5102 27580 5108
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 27540 4622 27568 5102
rect 27528 4616 27580 4622
rect 27528 4558 27580 4564
rect 27540 4214 27568 4558
rect 27528 4208 27580 4214
rect 27528 4150 27580 4156
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 27356 870 27476 898
rect 27356 762 27384 870
rect 27448 800 27476 870
rect 27080 734 27384 762
rect 27434 0 27490 800
rect 28276 762 28304 16546
rect 29828 4140 29880 4146
rect 29828 4082 29880 4088
rect 28552 870 28672 898
rect 28552 762 28580 870
rect 28644 800 28672 870
rect 29840 800 29868 4082
rect 28276 734 28580 762
rect 28630 0 28686 800
rect 29826 0 29882 800
<< via2 >>
rect 3974 32000 4030 32056
rect 4066 30640 4122 30696
rect 5678 29946 5734 29948
rect 5758 29946 5814 29948
rect 5838 29946 5894 29948
rect 5918 29946 5974 29948
rect 5678 29894 5724 29946
rect 5724 29894 5734 29946
rect 5758 29894 5788 29946
rect 5788 29894 5800 29946
rect 5800 29894 5814 29946
rect 5838 29894 5852 29946
rect 5852 29894 5864 29946
rect 5864 29894 5894 29946
rect 5918 29894 5928 29946
rect 5928 29894 5974 29946
rect 5678 29892 5734 29894
rect 5758 29892 5814 29894
rect 5838 29892 5894 29894
rect 5918 29892 5974 29894
rect 4066 29280 4122 29336
rect 4066 27920 4122 27976
rect 5678 28858 5734 28860
rect 5758 28858 5814 28860
rect 5838 28858 5894 28860
rect 5918 28858 5974 28860
rect 5678 28806 5724 28858
rect 5724 28806 5734 28858
rect 5758 28806 5788 28858
rect 5788 28806 5800 28858
rect 5800 28806 5814 28858
rect 5838 28806 5852 28858
rect 5852 28806 5864 28858
rect 5864 28806 5894 28858
rect 5918 28806 5928 28858
rect 5928 28806 5974 28858
rect 5678 28804 5734 28806
rect 5758 28804 5814 28806
rect 5838 28804 5894 28806
rect 5918 28804 5974 28806
rect 4066 26560 4122 26616
rect 4066 23840 4122 23896
rect 5678 27770 5734 27772
rect 5758 27770 5814 27772
rect 5838 27770 5894 27772
rect 5918 27770 5974 27772
rect 5678 27718 5724 27770
rect 5724 27718 5734 27770
rect 5758 27718 5788 27770
rect 5788 27718 5800 27770
rect 5800 27718 5814 27770
rect 5838 27718 5852 27770
rect 5852 27718 5864 27770
rect 5864 27718 5894 27770
rect 5918 27718 5928 27770
rect 5928 27718 5974 27770
rect 5678 27716 5734 27718
rect 5758 27716 5814 27718
rect 5838 27716 5894 27718
rect 5918 27716 5974 27718
rect 5678 26682 5734 26684
rect 5758 26682 5814 26684
rect 5838 26682 5894 26684
rect 5918 26682 5974 26684
rect 5678 26630 5724 26682
rect 5724 26630 5734 26682
rect 5758 26630 5788 26682
rect 5788 26630 5800 26682
rect 5800 26630 5814 26682
rect 5838 26630 5852 26682
rect 5852 26630 5864 26682
rect 5864 26630 5894 26682
rect 5918 26630 5928 26682
rect 5928 26630 5974 26682
rect 5678 26628 5734 26630
rect 5758 26628 5814 26630
rect 5838 26628 5894 26630
rect 5918 26628 5974 26630
rect 4066 21120 4122 21176
rect 3146 19760 3202 19816
rect 3698 18400 3754 18456
rect 3514 17040 3570 17096
rect 3698 17040 3754 17096
rect 5678 25594 5734 25596
rect 5758 25594 5814 25596
rect 5838 25594 5894 25596
rect 5918 25594 5974 25596
rect 5678 25542 5724 25594
rect 5724 25542 5734 25594
rect 5758 25542 5788 25594
rect 5788 25542 5800 25594
rect 5800 25542 5814 25594
rect 5838 25542 5852 25594
rect 5852 25542 5864 25594
rect 5864 25542 5894 25594
rect 5918 25542 5928 25594
rect 5928 25542 5974 25594
rect 5678 25540 5734 25542
rect 5758 25540 5814 25542
rect 5838 25540 5894 25542
rect 5918 25540 5974 25542
rect 5678 24506 5734 24508
rect 5758 24506 5814 24508
rect 5838 24506 5894 24508
rect 5918 24506 5974 24508
rect 5678 24454 5724 24506
rect 5724 24454 5734 24506
rect 5758 24454 5788 24506
rect 5788 24454 5800 24506
rect 5800 24454 5814 24506
rect 5838 24454 5852 24506
rect 5852 24454 5864 24506
rect 5864 24454 5894 24506
rect 5918 24454 5928 24506
rect 5928 24454 5974 24506
rect 5678 24452 5734 24454
rect 5758 24452 5814 24454
rect 5838 24452 5894 24454
rect 5918 24452 5974 24454
rect 5678 23418 5734 23420
rect 5758 23418 5814 23420
rect 5838 23418 5894 23420
rect 5918 23418 5974 23420
rect 5678 23366 5724 23418
rect 5724 23366 5734 23418
rect 5758 23366 5788 23418
rect 5788 23366 5800 23418
rect 5800 23366 5814 23418
rect 5838 23366 5852 23418
rect 5852 23366 5864 23418
rect 5864 23366 5894 23418
rect 5918 23366 5928 23418
rect 5928 23366 5974 23418
rect 5678 23364 5734 23366
rect 5758 23364 5814 23366
rect 5838 23364 5894 23366
rect 5918 23364 5974 23366
rect 5678 22330 5734 22332
rect 5758 22330 5814 22332
rect 5838 22330 5894 22332
rect 5918 22330 5974 22332
rect 5678 22278 5724 22330
rect 5724 22278 5734 22330
rect 5758 22278 5788 22330
rect 5788 22278 5800 22330
rect 5800 22278 5814 22330
rect 5838 22278 5852 22330
rect 5852 22278 5864 22330
rect 5864 22278 5894 22330
rect 5918 22278 5928 22330
rect 5928 22278 5974 22330
rect 5678 22276 5734 22278
rect 5758 22276 5814 22278
rect 5838 22276 5894 22278
rect 5918 22276 5974 22278
rect 5678 21242 5734 21244
rect 5758 21242 5814 21244
rect 5838 21242 5894 21244
rect 5918 21242 5974 21244
rect 5678 21190 5724 21242
rect 5724 21190 5734 21242
rect 5758 21190 5788 21242
rect 5788 21190 5800 21242
rect 5800 21190 5814 21242
rect 5838 21190 5852 21242
rect 5852 21190 5864 21242
rect 5864 21190 5894 21242
rect 5918 21190 5928 21242
rect 5928 21190 5974 21242
rect 5678 21188 5734 21190
rect 5758 21188 5814 21190
rect 5838 21188 5894 21190
rect 5918 21188 5974 21190
rect 5678 20154 5734 20156
rect 5758 20154 5814 20156
rect 5838 20154 5894 20156
rect 5918 20154 5974 20156
rect 5678 20102 5724 20154
rect 5724 20102 5734 20154
rect 5758 20102 5788 20154
rect 5788 20102 5800 20154
rect 5800 20102 5814 20154
rect 5838 20102 5852 20154
rect 5852 20102 5864 20154
rect 5864 20102 5894 20154
rect 5918 20102 5928 20154
rect 5928 20102 5974 20154
rect 5678 20100 5734 20102
rect 5758 20100 5814 20102
rect 5838 20100 5894 20102
rect 5918 20100 5974 20102
rect 4066 14320 4122 14376
rect 4066 12980 4122 13016
rect 4066 12960 4068 12980
rect 4068 12960 4120 12980
rect 4120 12960 4122 12980
rect 3974 11600 4030 11656
rect 5678 19066 5734 19068
rect 5758 19066 5814 19068
rect 5838 19066 5894 19068
rect 5918 19066 5974 19068
rect 5678 19014 5724 19066
rect 5724 19014 5734 19066
rect 5758 19014 5788 19066
rect 5788 19014 5800 19066
rect 5800 19014 5814 19066
rect 5838 19014 5852 19066
rect 5852 19014 5864 19066
rect 5864 19014 5894 19066
rect 5918 19014 5928 19066
rect 5928 19014 5974 19066
rect 5678 19012 5734 19014
rect 5758 19012 5814 19014
rect 5838 19012 5894 19014
rect 5918 19012 5974 19014
rect 5678 17978 5734 17980
rect 5758 17978 5814 17980
rect 5838 17978 5894 17980
rect 5918 17978 5974 17980
rect 5678 17926 5724 17978
rect 5724 17926 5734 17978
rect 5758 17926 5788 17978
rect 5788 17926 5800 17978
rect 5800 17926 5814 17978
rect 5838 17926 5852 17978
rect 5852 17926 5864 17978
rect 5864 17926 5894 17978
rect 5918 17926 5928 17978
rect 5928 17926 5974 17978
rect 5678 17924 5734 17926
rect 5758 17924 5814 17926
rect 5838 17924 5894 17926
rect 5918 17924 5974 17926
rect 5678 16890 5734 16892
rect 5758 16890 5814 16892
rect 5838 16890 5894 16892
rect 5918 16890 5974 16892
rect 5678 16838 5724 16890
rect 5724 16838 5734 16890
rect 5758 16838 5788 16890
rect 5788 16838 5800 16890
rect 5800 16838 5814 16890
rect 5838 16838 5852 16890
rect 5852 16838 5864 16890
rect 5864 16838 5894 16890
rect 5918 16838 5928 16890
rect 5928 16838 5974 16890
rect 5678 16836 5734 16838
rect 5758 16836 5814 16838
rect 5838 16836 5894 16838
rect 5918 16836 5974 16838
rect 5354 15680 5410 15736
rect 5678 15802 5734 15804
rect 5758 15802 5814 15804
rect 5838 15802 5894 15804
rect 5918 15802 5974 15804
rect 5678 15750 5724 15802
rect 5724 15750 5734 15802
rect 5758 15750 5788 15802
rect 5788 15750 5800 15802
rect 5800 15750 5814 15802
rect 5838 15750 5852 15802
rect 5852 15750 5864 15802
rect 5864 15750 5894 15802
rect 5918 15750 5928 15802
rect 5928 15750 5974 15802
rect 5678 15748 5734 15750
rect 5758 15748 5814 15750
rect 5838 15748 5894 15750
rect 5918 15748 5974 15750
rect 5678 14714 5734 14716
rect 5758 14714 5814 14716
rect 5838 14714 5894 14716
rect 5918 14714 5974 14716
rect 5678 14662 5724 14714
rect 5724 14662 5734 14714
rect 5758 14662 5788 14714
rect 5788 14662 5800 14714
rect 5800 14662 5814 14714
rect 5838 14662 5852 14714
rect 5852 14662 5864 14714
rect 5864 14662 5894 14714
rect 5918 14662 5928 14714
rect 5928 14662 5974 14714
rect 5678 14660 5734 14662
rect 5758 14660 5814 14662
rect 5838 14660 5894 14662
rect 5918 14660 5974 14662
rect 5678 13626 5734 13628
rect 5758 13626 5814 13628
rect 5838 13626 5894 13628
rect 5918 13626 5974 13628
rect 5678 13574 5724 13626
rect 5724 13574 5734 13626
rect 5758 13574 5788 13626
rect 5788 13574 5800 13626
rect 5800 13574 5814 13626
rect 5838 13574 5852 13626
rect 5852 13574 5864 13626
rect 5864 13574 5894 13626
rect 5918 13574 5928 13626
rect 5928 13574 5974 13626
rect 5678 13572 5734 13574
rect 5758 13572 5814 13574
rect 5838 13572 5894 13574
rect 5918 13572 5974 13574
rect 7102 17312 7158 17368
rect 5678 12538 5734 12540
rect 5758 12538 5814 12540
rect 5838 12538 5894 12540
rect 5918 12538 5974 12540
rect 5678 12486 5724 12538
rect 5724 12486 5734 12538
rect 5758 12486 5788 12538
rect 5788 12486 5800 12538
rect 5800 12486 5814 12538
rect 5838 12486 5852 12538
rect 5852 12486 5864 12538
rect 5864 12486 5894 12538
rect 5918 12486 5928 12538
rect 5928 12486 5974 12538
rect 5678 12484 5734 12486
rect 5758 12484 5814 12486
rect 5838 12484 5894 12486
rect 5918 12484 5974 12486
rect 4066 10260 4122 10296
rect 4066 10240 4068 10260
rect 4068 10240 4120 10260
rect 4120 10240 4122 10260
rect 4066 8900 4122 8936
rect 4066 8880 4068 8900
rect 4068 8880 4120 8900
rect 4120 8880 4122 8900
rect 3882 7520 3938 7576
rect 4066 6160 4122 6216
rect 5678 11450 5734 11452
rect 5758 11450 5814 11452
rect 5838 11450 5894 11452
rect 5918 11450 5974 11452
rect 5678 11398 5724 11450
rect 5724 11398 5734 11450
rect 5758 11398 5788 11450
rect 5788 11398 5800 11450
rect 5800 11398 5814 11450
rect 5838 11398 5852 11450
rect 5852 11398 5864 11450
rect 5864 11398 5894 11450
rect 5918 11398 5928 11450
rect 5928 11398 5974 11450
rect 5678 11396 5734 11398
rect 5758 11396 5814 11398
rect 5838 11396 5894 11398
rect 5918 11396 5974 11398
rect 5678 10362 5734 10364
rect 5758 10362 5814 10364
rect 5838 10362 5894 10364
rect 5918 10362 5974 10364
rect 5678 10310 5724 10362
rect 5724 10310 5734 10362
rect 5758 10310 5788 10362
rect 5788 10310 5800 10362
rect 5800 10310 5814 10362
rect 5838 10310 5852 10362
rect 5852 10310 5864 10362
rect 5864 10310 5894 10362
rect 5918 10310 5928 10362
rect 5928 10310 5974 10362
rect 5678 10308 5734 10310
rect 5758 10308 5814 10310
rect 5838 10308 5894 10310
rect 5918 10308 5974 10310
rect 9862 22888 9918 22944
rect 9770 22092 9826 22128
rect 9770 22072 9772 22092
rect 9772 22072 9824 22092
rect 9824 22072 9826 22092
rect 10401 30490 10457 30492
rect 10481 30490 10537 30492
rect 10561 30490 10617 30492
rect 10641 30490 10697 30492
rect 10401 30438 10447 30490
rect 10447 30438 10457 30490
rect 10481 30438 10511 30490
rect 10511 30438 10523 30490
rect 10523 30438 10537 30490
rect 10561 30438 10575 30490
rect 10575 30438 10587 30490
rect 10587 30438 10617 30490
rect 10641 30438 10651 30490
rect 10651 30438 10697 30490
rect 10401 30436 10457 30438
rect 10481 30436 10537 30438
rect 10561 30436 10617 30438
rect 10641 30436 10697 30438
rect 10401 29402 10457 29404
rect 10481 29402 10537 29404
rect 10561 29402 10617 29404
rect 10641 29402 10697 29404
rect 10401 29350 10447 29402
rect 10447 29350 10457 29402
rect 10481 29350 10511 29402
rect 10511 29350 10523 29402
rect 10523 29350 10537 29402
rect 10561 29350 10575 29402
rect 10575 29350 10587 29402
rect 10587 29350 10617 29402
rect 10641 29350 10651 29402
rect 10651 29350 10697 29402
rect 10401 29348 10457 29350
rect 10481 29348 10537 29350
rect 10561 29348 10617 29350
rect 10641 29348 10697 29350
rect 10046 26288 10102 26344
rect 10401 28314 10457 28316
rect 10481 28314 10537 28316
rect 10561 28314 10617 28316
rect 10641 28314 10697 28316
rect 10401 28262 10447 28314
rect 10447 28262 10457 28314
rect 10481 28262 10511 28314
rect 10511 28262 10523 28314
rect 10523 28262 10537 28314
rect 10561 28262 10575 28314
rect 10575 28262 10587 28314
rect 10587 28262 10617 28314
rect 10641 28262 10651 28314
rect 10651 28262 10697 28314
rect 10401 28260 10457 28262
rect 10481 28260 10537 28262
rect 10561 28260 10617 28262
rect 10641 28260 10697 28262
rect 10401 27226 10457 27228
rect 10481 27226 10537 27228
rect 10561 27226 10617 27228
rect 10641 27226 10697 27228
rect 10401 27174 10447 27226
rect 10447 27174 10457 27226
rect 10481 27174 10511 27226
rect 10511 27174 10523 27226
rect 10523 27174 10537 27226
rect 10561 27174 10575 27226
rect 10575 27174 10587 27226
rect 10587 27174 10617 27226
rect 10641 27174 10651 27226
rect 10651 27174 10697 27226
rect 10401 27172 10457 27174
rect 10481 27172 10537 27174
rect 10561 27172 10617 27174
rect 10641 27172 10697 27174
rect 10401 26138 10457 26140
rect 10481 26138 10537 26140
rect 10561 26138 10617 26140
rect 10641 26138 10697 26140
rect 10401 26086 10447 26138
rect 10447 26086 10457 26138
rect 10481 26086 10511 26138
rect 10511 26086 10523 26138
rect 10523 26086 10537 26138
rect 10561 26086 10575 26138
rect 10575 26086 10587 26138
rect 10587 26086 10617 26138
rect 10641 26086 10651 26138
rect 10651 26086 10697 26138
rect 10401 26084 10457 26086
rect 10481 26084 10537 26086
rect 10561 26084 10617 26086
rect 10641 26084 10697 26086
rect 10401 25050 10457 25052
rect 10481 25050 10537 25052
rect 10561 25050 10617 25052
rect 10641 25050 10697 25052
rect 10401 24998 10447 25050
rect 10447 24998 10457 25050
rect 10481 24998 10511 25050
rect 10511 24998 10523 25050
rect 10523 24998 10537 25050
rect 10561 24998 10575 25050
rect 10575 24998 10587 25050
rect 10587 24998 10617 25050
rect 10641 24998 10651 25050
rect 10651 24998 10697 25050
rect 10401 24996 10457 24998
rect 10481 24996 10537 24998
rect 10561 24996 10617 24998
rect 10641 24996 10697 24998
rect 10401 23962 10457 23964
rect 10481 23962 10537 23964
rect 10561 23962 10617 23964
rect 10641 23962 10697 23964
rect 10401 23910 10447 23962
rect 10447 23910 10457 23962
rect 10481 23910 10511 23962
rect 10511 23910 10523 23962
rect 10523 23910 10537 23962
rect 10561 23910 10575 23962
rect 10575 23910 10587 23962
rect 10587 23910 10617 23962
rect 10641 23910 10651 23962
rect 10651 23910 10697 23962
rect 10401 23908 10457 23910
rect 10481 23908 10537 23910
rect 10561 23908 10617 23910
rect 10641 23908 10697 23910
rect 7654 17176 7710 17232
rect 5678 9274 5734 9276
rect 5758 9274 5814 9276
rect 5838 9274 5894 9276
rect 5918 9274 5974 9276
rect 5678 9222 5724 9274
rect 5724 9222 5734 9274
rect 5758 9222 5788 9274
rect 5788 9222 5800 9274
rect 5800 9222 5814 9274
rect 5838 9222 5852 9274
rect 5852 9222 5864 9274
rect 5864 9222 5894 9274
rect 5918 9222 5928 9274
rect 5928 9222 5974 9274
rect 5678 9220 5734 9222
rect 5758 9220 5814 9222
rect 5838 9220 5894 9222
rect 5918 9220 5974 9222
rect 5678 8186 5734 8188
rect 5758 8186 5814 8188
rect 5838 8186 5894 8188
rect 5918 8186 5974 8188
rect 5678 8134 5724 8186
rect 5724 8134 5734 8186
rect 5758 8134 5788 8186
rect 5788 8134 5800 8186
rect 5800 8134 5814 8186
rect 5838 8134 5852 8186
rect 5852 8134 5864 8186
rect 5864 8134 5894 8186
rect 5918 8134 5928 8186
rect 5928 8134 5974 8186
rect 5678 8132 5734 8134
rect 5758 8132 5814 8134
rect 5838 8132 5894 8134
rect 5918 8132 5974 8134
rect 5678 7098 5734 7100
rect 5758 7098 5814 7100
rect 5838 7098 5894 7100
rect 5918 7098 5974 7100
rect 5678 7046 5724 7098
rect 5724 7046 5734 7098
rect 5758 7046 5788 7098
rect 5788 7046 5800 7098
rect 5800 7046 5814 7098
rect 5838 7046 5852 7098
rect 5852 7046 5864 7098
rect 5864 7046 5894 7098
rect 5918 7046 5928 7098
rect 5928 7046 5974 7098
rect 5678 7044 5734 7046
rect 5758 7044 5814 7046
rect 5838 7044 5894 7046
rect 5918 7044 5974 7046
rect 5678 6010 5734 6012
rect 5758 6010 5814 6012
rect 5838 6010 5894 6012
rect 5918 6010 5974 6012
rect 5678 5958 5724 6010
rect 5724 5958 5734 6010
rect 5758 5958 5788 6010
rect 5788 5958 5800 6010
rect 5800 5958 5814 6010
rect 5838 5958 5852 6010
rect 5852 5958 5864 6010
rect 5864 5958 5894 6010
rect 5918 5958 5928 6010
rect 5928 5958 5974 6010
rect 5678 5956 5734 5958
rect 5758 5956 5814 5958
rect 5838 5956 5894 5958
rect 5918 5956 5974 5958
rect 3974 4800 4030 4856
rect 5678 4922 5734 4924
rect 5758 4922 5814 4924
rect 5838 4922 5894 4924
rect 5918 4922 5974 4924
rect 5678 4870 5724 4922
rect 5724 4870 5734 4922
rect 5758 4870 5788 4922
rect 5788 4870 5800 4922
rect 5800 4870 5814 4922
rect 5838 4870 5852 4922
rect 5852 4870 5864 4922
rect 5864 4870 5894 4922
rect 5918 4870 5928 4922
rect 5928 4870 5974 4922
rect 5678 4868 5734 4870
rect 5758 4868 5814 4870
rect 5838 4868 5894 4870
rect 5918 4868 5974 4870
rect 5678 3834 5734 3836
rect 5758 3834 5814 3836
rect 5838 3834 5894 3836
rect 5918 3834 5974 3836
rect 5678 3782 5724 3834
rect 5724 3782 5734 3834
rect 5758 3782 5788 3834
rect 5788 3782 5800 3834
rect 5800 3782 5814 3834
rect 5838 3782 5852 3834
rect 5852 3782 5864 3834
rect 5864 3782 5894 3834
rect 5918 3782 5928 3834
rect 5928 3782 5974 3834
rect 5678 3780 5734 3782
rect 5758 3780 5814 3782
rect 5838 3780 5894 3782
rect 5918 3780 5974 3782
rect 1398 3440 1454 3496
rect 3054 2080 3110 2136
rect 5678 2746 5734 2748
rect 5758 2746 5814 2748
rect 5838 2746 5894 2748
rect 5918 2746 5974 2748
rect 5678 2694 5724 2746
rect 5724 2694 5734 2746
rect 5758 2694 5788 2746
rect 5788 2694 5800 2746
rect 5800 2694 5814 2746
rect 5838 2694 5852 2746
rect 5852 2694 5864 2746
rect 5864 2694 5894 2746
rect 5918 2694 5928 2746
rect 5928 2694 5974 2746
rect 5678 2692 5734 2694
rect 5758 2692 5814 2694
rect 5838 2692 5894 2694
rect 5918 2692 5974 2694
rect 10401 22874 10457 22876
rect 10481 22874 10537 22876
rect 10561 22874 10617 22876
rect 10641 22874 10697 22876
rect 10401 22822 10447 22874
rect 10447 22822 10457 22874
rect 10481 22822 10511 22874
rect 10511 22822 10523 22874
rect 10523 22822 10537 22874
rect 10561 22822 10575 22874
rect 10575 22822 10587 22874
rect 10587 22822 10617 22874
rect 10641 22822 10651 22874
rect 10651 22822 10697 22874
rect 10401 22820 10457 22822
rect 10481 22820 10537 22822
rect 10561 22820 10617 22822
rect 10641 22820 10697 22822
rect 10414 22652 10416 22672
rect 10416 22652 10468 22672
rect 10468 22652 10470 22672
rect 10414 22616 10470 22652
rect 10401 21786 10457 21788
rect 10481 21786 10537 21788
rect 10561 21786 10617 21788
rect 10641 21786 10697 21788
rect 10401 21734 10447 21786
rect 10447 21734 10457 21786
rect 10481 21734 10511 21786
rect 10511 21734 10523 21786
rect 10523 21734 10537 21786
rect 10561 21734 10575 21786
rect 10575 21734 10587 21786
rect 10587 21734 10617 21786
rect 10641 21734 10651 21786
rect 10651 21734 10697 21786
rect 10401 21732 10457 21734
rect 10481 21732 10537 21734
rect 10561 21732 10617 21734
rect 10641 21732 10697 21734
rect 10401 20698 10457 20700
rect 10481 20698 10537 20700
rect 10561 20698 10617 20700
rect 10641 20698 10697 20700
rect 10401 20646 10447 20698
rect 10447 20646 10457 20698
rect 10481 20646 10511 20698
rect 10511 20646 10523 20698
rect 10523 20646 10537 20698
rect 10561 20646 10575 20698
rect 10575 20646 10587 20698
rect 10587 20646 10617 20698
rect 10641 20646 10651 20698
rect 10651 20646 10697 20698
rect 10401 20644 10457 20646
rect 10481 20644 10537 20646
rect 10561 20644 10617 20646
rect 10641 20644 10697 20646
rect 11702 25780 11704 25800
rect 11704 25780 11756 25800
rect 11756 25780 11758 25800
rect 11702 25744 11758 25780
rect 11518 22108 11520 22128
rect 11520 22108 11572 22128
rect 11572 22108 11574 22128
rect 11518 22072 11574 22108
rect 10401 19610 10457 19612
rect 10481 19610 10537 19612
rect 10561 19610 10617 19612
rect 10641 19610 10697 19612
rect 10401 19558 10447 19610
rect 10447 19558 10457 19610
rect 10481 19558 10511 19610
rect 10511 19558 10523 19610
rect 10523 19558 10537 19610
rect 10561 19558 10575 19610
rect 10575 19558 10587 19610
rect 10587 19558 10617 19610
rect 10641 19558 10651 19610
rect 10651 19558 10697 19610
rect 10401 19556 10457 19558
rect 10481 19556 10537 19558
rect 10561 19556 10617 19558
rect 10641 19556 10697 19558
rect 10966 19352 11022 19408
rect 10401 18522 10457 18524
rect 10481 18522 10537 18524
rect 10561 18522 10617 18524
rect 10641 18522 10697 18524
rect 10401 18470 10447 18522
rect 10447 18470 10457 18522
rect 10481 18470 10511 18522
rect 10511 18470 10523 18522
rect 10523 18470 10537 18522
rect 10561 18470 10575 18522
rect 10575 18470 10587 18522
rect 10587 18470 10617 18522
rect 10641 18470 10651 18522
rect 10651 18470 10697 18522
rect 10401 18468 10457 18470
rect 10481 18468 10537 18470
rect 10561 18468 10617 18470
rect 10641 18468 10697 18470
rect 10874 17620 10876 17640
rect 10876 17620 10928 17640
rect 10928 17620 10930 17640
rect 10401 17434 10457 17436
rect 10481 17434 10537 17436
rect 10561 17434 10617 17436
rect 10641 17434 10697 17436
rect 10401 17382 10447 17434
rect 10447 17382 10457 17434
rect 10481 17382 10511 17434
rect 10511 17382 10523 17434
rect 10523 17382 10537 17434
rect 10561 17382 10575 17434
rect 10575 17382 10587 17434
rect 10587 17382 10617 17434
rect 10641 17382 10651 17434
rect 10651 17382 10697 17434
rect 10401 17380 10457 17382
rect 10481 17380 10537 17382
rect 10561 17380 10617 17382
rect 10641 17380 10697 17382
rect 10874 17584 10930 17620
rect 12622 27124 12678 27160
rect 12622 27104 12624 27124
rect 12624 27104 12676 27124
rect 12676 27104 12678 27124
rect 12530 25644 12532 25664
rect 12532 25644 12584 25664
rect 12584 25644 12586 25664
rect 12530 25608 12586 25644
rect 13174 25764 13230 25800
rect 13174 25744 13176 25764
rect 13176 25744 13228 25764
rect 13228 25744 13230 25764
rect 15124 29946 15180 29948
rect 15204 29946 15260 29948
rect 15284 29946 15340 29948
rect 15364 29946 15420 29948
rect 15124 29894 15170 29946
rect 15170 29894 15180 29946
rect 15204 29894 15234 29946
rect 15234 29894 15246 29946
rect 15246 29894 15260 29946
rect 15284 29894 15298 29946
rect 15298 29894 15310 29946
rect 15310 29894 15340 29946
rect 15364 29894 15374 29946
rect 15374 29894 15420 29946
rect 15124 29892 15180 29894
rect 15204 29892 15260 29894
rect 15284 29892 15340 29894
rect 15364 29892 15420 29894
rect 15124 28858 15180 28860
rect 15204 28858 15260 28860
rect 15284 28858 15340 28860
rect 15364 28858 15420 28860
rect 15124 28806 15170 28858
rect 15170 28806 15180 28858
rect 15204 28806 15234 28858
rect 15234 28806 15246 28858
rect 15246 28806 15260 28858
rect 15284 28806 15298 28858
rect 15298 28806 15310 28858
rect 15310 28806 15340 28858
rect 15364 28806 15374 28858
rect 15374 28806 15420 28858
rect 15124 28804 15180 28806
rect 15204 28804 15260 28806
rect 15284 28804 15340 28806
rect 15364 28804 15420 28806
rect 15124 27770 15180 27772
rect 15204 27770 15260 27772
rect 15284 27770 15340 27772
rect 15364 27770 15420 27772
rect 15124 27718 15170 27770
rect 15170 27718 15180 27770
rect 15204 27718 15234 27770
rect 15234 27718 15246 27770
rect 15246 27718 15260 27770
rect 15284 27718 15298 27770
rect 15298 27718 15310 27770
rect 15310 27718 15340 27770
rect 15364 27718 15374 27770
rect 15374 27718 15420 27770
rect 15124 27716 15180 27718
rect 15204 27716 15260 27718
rect 15284 27716 15340 27718
rect 15364 27716 15420 27718
rect 15198 27104 15254 27160
rect 11794 20984 11850 21040
rect 10401 16346 10457 16348
rect 10481 16346 10537 16348
rect 10561 16346 10617 16348
rect 10641 16346 10697 16348
rect 10401 16294 10447 16346
rect 10447 16294 10457 16346
rect 10481 16294 10511 16346
rect 10511 16294 10523 16346
rect 10523 16294 10537 16346
rect 10561 16294 10575 16346
rect 10575 16294 10587 16346
rect 10587 16294 10617 16346
rect 10641 16294 10651 16346
rect 10651 16294 10697 16346
rect 10401 16292 10457 16294
rect 10481 16292 10537 16294
rect 10561 16292 10617 16294
rect 10641 16292 10697 16294
rect 10401 15258 10457 15260
rect 10481 15258 10537 15260
rect 10561 15258 10617 15260
rect 10641 15258 10697 15260
rect 10401 15206 10447 15258
rect 10447 15206 10457 15258
rect 10481 15206 10511 15258
rect 10511 15206 10523 15258
rect 10523 15206 10537 15258
rect 10561 15206 10575 15258
rect 10575 15206 10587 15258
rect 10587 15206 10617 15258
rect 10641 15206 10651 15258
rect 10651 15206 10697 15258
rect 10401 15204 10457 15206
rect 10481 15204 10537 15206
rect 10561 15204 10617 15206
rect 10641 15204 10697 15206
rect 10401 14170 10457 14172
rect 10481 14170 10537 14172
rect 10561 14170 10617 14172
rect 10641 14170 10697 14172
rect 10401 14118 10447 14170
rect 10447 14118 10457 14170
rect 10481 14118 10511 14170
rect 10511 14118 10523 14170
rect 10523 14118 10537 14170
rect 10561 14118 10575 14170
rect 10575 14118 10587 14170
rect 10587 14118 10617 14170
rect 10641 14118 10651 14170
rect 10651 14118 10697 14170
rect 10401 14116 10457 14118
rect 10481 14116 10537 14118
rect 10561 14116 10617 14118
rect 10641 14116 10697 14118
rect 10401 13082 10457 13084
rect 10481 13082 10537 13084
rect 10561 13082 10617 13084
rect 10641 13082 10697 13084
rect 10401 13030 10447 13082
rect 10447 13030 10457 13082
rect 10481 13030 10511 13082
rect 10511 13030 10523 13082
rect 10523 13030 10537 13082
rect 10561 13030 10575 13082
rect 10575 13030 10587 13082
rect 10587 13030 10617 13082
rect 10641 13030 10651 13082
rect 10651 13030 10697 13082
rect 10401 13028 10457 13030
rect 10481 13028 10537 13030
rect 10561 13028 10617 13030
rect 10641 13028 10697 13030
rect 10401 11994 10457 11996
rect 10481 11994 10537 11996
rect 10561 11994 10617 11996
rect 10641 11994 10697 11996
rect 10401 11942 10447 11994
rect 10447 11942 10457 11994
rect 10481 11942 10511 11994
rect 10511 11942 10523 11994
rect 10523 11942 10537 11994
rect 10561 11942 10575 11994
rect 10575 11942 10587 11994
rect 10587 11942 10617 11994
rect 10641 11942 10651 11994
rect 10651 11942 10697 11994
rect 10401 11940 10457 11942
rect 10481 11940 10537 11942
rect 10561 11940 10617 11942
rect 10641 11940 10697 11942
rect 10401 10906 10457 10908
rect 10481 10906 10537 10908
rect 10561 10906 10617 10908
rect 10641 10906 10697 10908
rect 10401 10854 10447 10906
rect 10447 10854 10457 10906
rect 10481 10854 10511 10906
rect 10511 10854 10523 10906
rect 10523 10854 10537 10906
rect 10561 10854 10575 10906
rect 10575 10854 10587 10906
rect 10587 10854 10617 10906
rect 10641 10854 10651 10906
rect 10651 10854 10697 10906
rect 10401 10852 10457 10854
rect 10481 10852 10537 10854
rect 10561 10852 10617 10854
rect 10641 10852 10697 10854
rect 10401 9818 10457 9820
rect 10481 9818 10537 9820
rect 10561 9818 10617 9820
rect 10641 9818 10697 9820
rect 10401 9766 10447 9818
rect 10447 9766 10457 9818
rect 10481 9766 10511 9818
rect 10511 9766 10523 9818
rect 10523 9766 10537 9818
rect 10561 9766 10575 9818
rect 10575 9766 10587 9818
rect 10587 9766 10617 9818
rect 10641 9766 10651 9818
rect 10651 9766 10697 9818
rect 10401 9764 10457 9766
rect 10481 9764 10537 9766
rect 10561 9764 10617 9766
rect 10641 9764 10697 9766
rect 12162 20304 12218 20360
rect 11978 17620 11980 17640
rect 11980 17620 12032 17640
rect 12032 17620 12034 17640
rect 11978 17584 12034 17620
rect 12254 17856 12310 17912
rect 12162 17176 12218 17232
rect 12806 17720 12862 17776
rect 15124 26682 15180 26684
rect 15204 26682 15260 26684
rect 15284 26682 15340 26684
rect 15364 26682 15420 26684
rect 15124 26630 15170 26682
rect 15170 26630 15180 26682
rect 15204 26630 15234 26682
rect 15234 26630 15246 26682
rect 15246 26630 15260 26682
rect 15284 26630 15298 26682
rect 15298 26630 15310 26682
rect 15310 26630 15340 26682
rect 15364 26630 15374 26682
rect 15374 26630 15420 26682
rect 15124 26628 15180 26630
rect 15204 26628 15260 26630
rect 15284 26628 15340 26630
rect 15364 26628 15420 26630
rect 15566 26288 15622 26344
rect 15124 25594 15180 25596
rect 15204 25594 15260 25596
rect 15284 25594 15340 25596
rect 15364 25594 15420 25596
rect 15124 25542 15170 25594
rect 15170 25542 15180 25594
rect 15204 25542 15234 25594
rect 15234 25542 15246 25594
rect 15246 25542 15260 25594
rect 15284 25542 15298 25594
rect 15298 25542 15310 25594
rect 15310 25542 15340 25594
rect 15364 25542 15374 25594
rect 15374 25542 15420 25594
rect 15124 25540 15180 25542
rect 15204 25540 15260 25542
rect 15284 25540 15340 25542
rect 15364 25540 15420 25542
rect 15566 25236 15568 25256
rect 15568 25236 15620 25256
rect 15620 25236 15622 25256
rect 15566 25200 15622 25236
rect 13818 19352 13874 19408
rect 13266 17720 13322 17776
rect 13082 17312 13138 17368
rect 10401 8730 10457 8732
rect 10481 8730 10537 8732
rect 10561 8730 10617 8732
rect 10641 8730 10697 8732
rect 10401 8678 10447 8730
rect 10447 8678 10457 8730
rect 10481 8678 10511 8730
rect 10511 8678 10523 8730
rect 10523 8678 10537 8730
rect 10561 8678 10575 8730
rect 10575 8678 10587 8730
rect 10587 8678 10617 8730
rect 10641 8678 10651 8730
rect 10651 8678 10697 8730
rect 10401 8676 10457 8678
rect 10481 8676 10537 8678
rect 10561 8676 10617 8678
rect 10641 8676 10697 8678
rect 3330 720 3386 776
rect 10401 7642 10457 7644
rect 10481 7642 10537 7644
rect 10561 7642 10617 7644
rect 10641 7642 10697 7644
rect 10401 7590 10447 7642
rect 10447 7590 10457 7642
rect 10481 7590 10511 7642
rect 10511 7590 10523 7642
rect 10523 7590 10537 7642
rect 10561 7590 10575 7642
rect 10575 7590 10587 7642
rect 10587 7590 10617 7642
rect 10641 7590 10651 7642
rect 10651 7590 10697 7642
rect 10401 7588 10457 7590
rect 10481 7588 10537 7590
rect 10561 7588 10617 7590
rect 10641 7588 10697 7590
rect 10401 6554 10457 6556
rect 10481 6554 10537 6556
rect 10561 6554 10617 6556
rect 10641 6554 10697 6556
rect 10401 6502 10447 6554
rect 10447 6502 10457 6554
rect 10481 6502 10511 6554
rect 10511 6502 10523 6554
rect 10523 6502 10537 6554
rect 10561 6502 10575 6554
rect 10575 6502 10587 6554
rect 10587 6502 10617 6554
rect 10641 6502 10651 6554
rect 10651 6502 10697 6554
rect 10401 6500 10457 6502
rect 10481 6500 10537 6502
rect 10561 6500 10617 6502
rect 10641 6500 10697 6502
rect 10401 5466 10457 5468
rect 10481 5466 10537 5468
rect 10561 5466 10617 5468
rect 10641 5466 10697 5468
rect 10401 5414 10447 5466
rect 10447 5414 10457 5466
rect 10481 5414 10511 5466
rect 10511 5414 10523 5466
rect 10523 5414 10537 5466
rect 10561 5414 10575 5466
rect 10575 5414 10587 5466
rect 10587 5414 10617 5466
rect 10641 5414 10651 5466
rect 10651 5414 10697 5466
rect 10401 5412 10457 5414
rect 10481 5412 10537 5414
rect 10561 5412 10617 5414
rect 10641 5412 10697 5414
rect 10401 4378 10457 4380
rect 10481 4378 10537 4380
rect 10561 4378 10617 4380
rect 10641 4378 10697 4380
rect 10401 4326 10447 4378
rect 10447 4326 10457 4378
rect 10481 4326 10511 4378
rect 10511 4326 10523 4378
rect 10523 4326 10537 4378
rect 10561 4326 10575 4378
rect 10575 4326 10587 4378
rect 10587 4326 10617 4378
rect 10641 4326 10651 4378
rect 10651 4326 10697 4378
rect 10401 4324 10457 4326
rect 10481 4324 10537 4326
rect 10561 4324 10617 4326
rect 10641 4324 10697 4326
rect 10401 3290 10457 3292
rect 10481 3290 10537 3292
rect 10561 3290 10617 3292
rect 10641 3290 10697 3292
rect 10401 3238 10447 3290
rect 10447 3238 10457 3290
rect 10481 3238 10511 3290
rect 10511 3238 10523 3290
rect 10523 3238 10537 3290
rect 10561 3238 10575 3290
rect 10575 3238 10587 3290
rect 10587 3238 10617 3290
rect 10641 3238 10651 3290
rect 10651 3238 10697 3290
rect 10401 3236 10457 3238
rect 10481 3236 10537 3238
rect 10561 3236 10617 3238
rect 10641 3236 10697 3238
rect 12714 14048 12770 14104
rect 13726 14048 13782 14104
rect 12990 12164 13046 12200
rect 12990 12144 12992 12164
rect 12992 12144 13044 12164
rect 13044 12144 13046 12164
rect 12162 9424 12218 9480
rect 11978 9288 12034 9344
rect 12346 9288 12402 9344
rect 12898 9460 12900 9480
rect 12900 9460 12952 9480
rect 12952 9460 12954 9480
rect 12898 9424 12954 9460
rect 14094 20304 14150 20360
rect 14186 17856 14242 17912
rect 15124 24506 15180 24508
rect 15204 24506 15260 24508
rect 15284 24506 15340 24508
rect 15364 24506 15420 24508
rect 15124 24454 15170 24506
rect 15170 24454 15180 24506
rect 15204 24454 15234 24506
rect 15234 24454 15246 24506
rect 15246 24454 15260 24506
rect 15284 24454 15298 24506
rect 15298 24454 15310 24506
rect 15310 24454 15340 24506
rect 15364 24454 15374 24506
rect 15374 24454 15420 24506
rect 15124 24452 15180 24454
rect 15204 24452 15260 24454
rect 15284 24452 15340 24454
rect 15364 24452 15420 24454
rect 15842 25200 15898 25256
rect 15124 23418 15180 23420
rect 15204 23418 15260 23420
rect 15284 23418 15340 23420
rect 15364 23418 15420 23420
rect 15124 23366 15170 23418
rect 15170 23366 15180 23418
rect 15204 23366 15234 23418
rect 15234 23366 15246 23418
rect 15246 23366 15260 23418
rect 15284 23366 15298 23418
rect 15298 23366 15310 23418
rect 15310 23366 15340 23418
rect 15364 23366 15374 23418
rect 15374 23366 15420 23418
rect 15124 23364 15180 23366
rect 15204 23364 15260 23366
rect 15284 23364 15340 23366
rect 15364 23364 15420 23366
rect 15124 22330 15180 22332
rect 15204 22330 15260 22332
rect 15284 22330 15340 22332
rect 15364 22330 15420 22332
rect 15124 22278 15170 22330
rect 15170 22278 15180 22330
rect 15204 22278 15234 22330
rect 15234 22278 15246 22330
rect 15246 22278 15260 22330
rect 15284 22278 15298 22330
rect 15298 22278 15310 22330
rect 15310 22278 15340 22330
rect 15364 22278 15374 22330
rect 15374 22278 15420 22330
rect 15124 22276 15180 22278
rect 15204 22276 15260 22278
rect 15284 22276 15340 22278
rect 15364 22276 15420 22278
rect 10401 2202 10457 2204
rect 10481 2202 10537 2204
rect 10561 2202 10617 2204
rect 10641 2202 10697 2204
rect 10401 2150 10447 2202
rect 10447 2150 10457 2202
rect 10481 2150 10511 2202
rect 10511 2150 10523 2202
rect 10523 2150 10537 2202
rect 10561 2150 10575 2202
rect 10575 2150 10587 2202
rect 10587 2150 10617 2202
rect 10641 2150 10651 2202
rect 10651 2150 10697 2202
rect 10401 2148 10457 2150
rect 10481 2148 10537 2150
rect 10561 2148 10617 2150
rect 10641 2148 10697 2150
rect 14922 17312 14978 17368
rect 15124 21242 15180 21244
rect 15204 21242 15260 21244
rect 15284 21242 15340 21244
rect 15364 21242 15420 21244
rect 15124 21190 15170 21242
rect 15170 21190 15180 21242
rect 15204 21190 15234 21242
rect 15234 21190 15246 21242
rect 15246 21190 15260 21242
rect 15284 21190 15298 21242
rect 15298 21190 15310 21242
rect 15310 21190 15340 21242
rect 15364 21190 15374 21242
rect 15374 21190 15420 21242
rect 15124 21188 15180 21190
rect 15204 21188 15260 21190
rect 15284 21188 15340 21190
rect 15364 21188 15420 21190
rect 15124 20154 15180 20156
rect 15204 20154 15260 20156
rect 15284 20154 15340 20156
rect 15364 20154 15420 20156
rect 15124 20102 15170 20154
rect 15170 20102 15180 20154
rect 15204 20102 15234 20154
rect 15234 20102 15246 20154
rect 15246 20102 15260 20154
rect 15284 20102 15298 20154
rect 15298 20102 15310 20154
rect 15310 20102 15340 20154
rect 15364 20102 15374 20154
rect 15374 20102 15420 20154
rect 15124 20100 15180 20102
rect 15204 20100 15260 20102
rect 15284 20100 15340 20102
rect 15364 20100 15420 20102
rect 15658 20984 15714 21040
rect 15124 19066 15180 19068
rect 15204 19066 15260 19068
rect 15284 19066 15340 19068
rect 15364 19066 15420 19068
rect 15124 19014 15170 19066
rect 15170 19014 15180 19066
rect 15204 19014 15234 19066
rect 15234 19014 15246 19066
rect 15246 19014 15260 19066
rect 15284 19014 15298 19066
rect 15298 19014 15310 19066
rect 15310 19014 15340 19066
rect 15364 19014 15374 19066
rect 15374 19014 15420 19066
rect 15124 19012 15180 19014
rect 15204 19012 15260 19014
rect 15284 19012 15340 19014
rect 15364 19012 15420 19014
rect 15124 17978 15180 17980
rect 15204 17978 15260 17980
rect 15284 17978 15340 17980
rect 15364 17978 15420 17980
rect 15124 17926 15170 17978
rect 15170 17926 15180 17978
rect 15204 17926 15234 17978
rect 15234 17926 15246 17978
rect 15246 17926 15260 17978
rect 15284 17926 15298 17978
rect 15298 17926 15310 17978
rect 15310 17926 15340 17978
rect 15364 17926 15374 17978
rect 15374 17926 15420 17978
rect 15124 17924 15180 17926
rect 15204 17924 15260 17926
rect 15284 17924 15340 17926
rect 15364 17924 15420 17926
rect 17406 26988 17462 27024
rect 17406 26968 17408 26988
rect 17408 26968 17460 26988
rect 17460 26968 17462 26988
rect 15124 16890 15180 16892
rect 15204 16890 15260 16892
rect 15284 16890 15340 16892
rect 15364 16890 15420 16892
rect 15124 16838 15170 16890
rect 15170 16838 15180 16890
rect 15204 16838 15234 16890
rect 15234 16838 15246 16890
rect 15246 16838 15260 16890
rect 15284 16838 15298 16890
rect 15298 16838 15310 16890
rect 15310 16838 15340 16890
rect 15364 16838 15374 16890
rect 15374 16838 15420 16890
rect 15124 16836 15180 16838
rect 15204 16836 15260 16838
rect 15284 16836 15340 16838
rect 15364 16836 15420 16838
rect 14278 7948 14334 7984
rect 14278 7928 14280 7948
rect 14280 7928 14332 7948
rect 14332 7928 14334 7948
rect 15124 15802 15180 15804
rect 15204 15802 15260 15804
rect 15284 15802 15340 15804
rect 15364 15802 15420 15804
rect 15124 15750 15170 15802
rect 15170 15750 15180 15802
rect 15204 15750 15234 15802
rect 15234 15750 15246 15802
rect 15246 15750 15260 15802
rect 15284 15750 15298 15802
rect 15298 15750 15310 15802
rect 15310 15750 15340 15802
rect 15364 15750 15374 15802
rect 15374 15750 15420 15802
rect 15124 15748 15180 15750
rect 15204 15748 15260 15750
rect 15284 15748 15340 15750
rect 15364 15748 15420 15750
rect 16210 17312 16266 17368
rect 15124 14714 15180 14716
rect 15204 14714 15260 14716
rect 15284 14714 15340 14716
rect 15364 14714 15420 14716
rect 15124 14662 15170 14714
rect 15170 14662 15180 14714
rect 15204 14662 15234 14714
rect 15234 14662 15246 14714
rect 15246 14662 15260 14714
rect 15284 14662 15298 14714
rect 15298 14662 15310 14714
rect 15310 14662 15340 14714
rect 15364 14662 15374 14714
rect 15374 14662 15420 14714
rect 15124 14660 15180 14662
rect 15204 14660 15260 14662
rect 15284 14660 15340 14662
rect 15364 14660 15420 14662
rect 15124 13626 15180 13628
rect 15204 13626 15260 13628
rect 15284 13626 15340 13628
rect 15364 13626 15420 13628
rect 15124 13574 15170 13626
rect 15170 13574 15180 13626
rect 15204 13574 15234 13626
rect 15234 13574 15246 13626
rect 15246 13574 15260 13626
rect 15284 13574 15298 13626
rect 15298 13574 15310 13626
rect 15310 13574 15340 13626
rect 15364 13574 15374 13626
rect 15374 13574 15420 13626
rect 15124 13572 15180 13574
rect 15204 13572 15260 13574
rect 15284 13572 15340 13574
rect 15364 13572 15420 13574
rect 15124 12538 15180 12540
rect 15204 12538 15260 12540
rect 15284 12538 15340 12540
rect 15364 12538 15420 12540
rect 15124 12486 15170 12538
rect 15170 12486 15180 12538
rect 15204 12486 15234 12538
rect 15234 12486 15246 12538
rect 15246 12486 15260 12538
rect 15284 12486 15298 12538
rect 15298 12486 15310 12538
rect 15310 12486 15340 12538
rect 15364 12486 15374 12538
rect 15374 12486 15420 12538
rect 15124 12484 15180 12486
rect 15204 12484 15260 12486
rect 15284 12484 15340 12486
rect 15364 12484 15420 12486
rect 15658 12316 15660 12336
rect 15660 12316 15712 12336
rect 15712 12316 15714 12336
rect 15658 12280 15714 12316
rect 15124 11450 15180 11452
rect 15204 11450 15260 11452
rect 15284 11450 15340 11452
rect 15364 11450 15420 11452
rect 15124 11398 15170 11450
rect 15170 11398 15180 11450
rect 15204 11398 15234 11450
rect 15234 11398 15246 11450
rect 15246 11398 15260 11450
rect 15284 11398 15298 11450
rect 15298 11398 15310 11450
rect 15310 11398 15340 11450
rect 15364 11398 15374 11450
rect 15374 11398 15420 11450
rect 15124 11396 15180 11398
rect 15204 11396 15260 11398
rect 15284 11396 15340 11398
rect 15364 11396 15420 11398
rect 15124 10362 15180 10364
rect 15204 10362 15260 10364
rect 15284 10362 15340 10364
rect 15364 10362 15420 10364
rect 15124 10310 15170 10362
rect 15170 10310 15180 10362
rect 15204 10310 15234 10362
rect 15234 10310 15246 10362
rect 15246 10310 15260 10362
rect 15284 10310 15298 10362
rect 15298 10310 15310 10362
rect 15310 10310 15340 10362
rect 15364 10310 15374 10362
rect 15374 10310 15420 10362
rect 15124 10308 15180 10310
rect 15204 10308 15260 10310
rect 15284 10308 15340 10310
rect 15364 10308 15420 10310
rect 17866 27396 17922 27432
rect 17866 27376 17868 27396
rect 17868 27376 17920 27396
rect 17920 27376 17922 27396
rect 18786 27004 18788 27024
rect 18788 27004 18840 27024
rect 18840 27004 18842 27024
rect 18786 26968 18842 27004
rect 19846 30490 19902 30492
rect 19926 30490 19982 30492
rect 20006 30490 20062 30492
rect 20086 30490 20142 30492
rect 19846 30438 19892 30490
rect 19892 30438 19902 30490
rect 19926 30438 19956 30490
rect 19956 30438 19968 30490
rect 19968 30438 19982 30490
rect 20006 30438 20020 30490
rect 20020 30438 20032 30490
rect 20032 30438 20062 30490
rect 20086 30438 20096 30490
rect 20096 30438 20142 30490
rect 19846 30436 19902 30438
rect 19926 30436 19982 30438
rect 20006 30436 20062 30438
rect 20086 30436 20142 30438
rect 19846 29402 19902 29404
rect 19926 29402 19982 29404
rect 20006 29402 20062 29404
rect 20086 29402 20142 29404
rect 19846 29350 19892 29402
rect 19892 29350 19902 29402
rect 19926 29350 19956 29402
rect 19956 29350 19968 29402
rect 19968 29350 19982 29402
rect 20006 29350 20020 29402
rect 20020 29350 20032 29402
rect 20032 29350 20062 29402
rect 20086 29350 20096 29402
rect 20096 29350 20142 29402
rect 19846 29348 19902 29350
rect 19926 29348 19982 29350
rect 20006 29348 20062 29350
rect 20086 29348 20142 29350
rect 19846 28314 19902 28316
rect 19926 28314 19982 28316
rect 20006 28314 20062 28316
rect 20086 28314 20142 28316
rect 19846 28262 19892 28314
rect 19892 28262 19902 28314
rect 19926 28262 19956 28314
rect 19956 28262 19968 28314
rect 19968 28262 19982 28314
rect 20006 28262 20020 28314
rect 20020 28262 20032 28314
rect 20032 28262 20062 28314
rect 20086 28262 20096 28314
rect 20096 28262 20142 28314
rect 19846 28260 19902 28262
rect 19926 28260 19982 28262
rect 20006 28260 20062 28262
rect 20086 28260 20142 28262
rect 19706 27376 19762 27432
rect 19846 27226 19902 27228
rect 19926 27226 19982 27228
rect 20006 27226 20062 27228
rect 20086 27226 20142 27228
rect 19846 27174 19892 27226
rect 19892 27174 19902 27226
rect 19926 27174 19956 27226
rect 19956 27174 19968 27226
rect 19968 27174 19982 27226
rect 20006 27174 20020 27226
rect 20020 27174 20032 27226
rect 20032 27174 20062 27226
rect 20086 27174 20096 27226
rect 20096 27174 20142 27226
rect 19846 27172 19902 27174
rect 19926 27172 19982 27174
rect 20006 27172 20062 27174
rect 20086 27172 20142 27174
rect 17682 17856 17738 17912
rect 18694 23044 18750 23080
rect 18694 23024 18696 23044
rect 18696 23024 18748 23044
rect 18748 23024 18750 23044
rect 15124 9274 15180 9276
rect 15204 9274 15260 9276
rect 15284 9274 15340 9276
rect 15364 9274 15420 9276
rect 15124 9222 15170 9274
rect 15170 9222 15180 9274
rect 15204 9222 15234 9274
rect 15234 9222 15246 9274
rect 15246 9222 15260 9274
rect 15284 9222 15298 9274
rect 15298 9222 15310 9274
rect 15310 9222 15340 9274
rect 15364 9222 15374 9274
rect 15374 9222 15420 9274
rect 15124 9220 15180 9222
rect 15204 9220 15260 9222
rect 15284 9220 15340 9222
rect 15364 9220 15420 9222
rect 15124 8186 15180 8188
rect 15204 8186 15260 8188
rect 15284 8186 15340 8188
rect 15364 8186 15420 8188
rect 15124 8134 15170 8186
rect 15170 8134 15180 8186
rect 15204 8134 15234 8186
rect 15234 8134 15246 8186
rect 15246 8134 15260 8186
rect 15284 8134 15298 8186
rect 15298 8134 15310 8186
rect 15310 8134 15340 8186
rect 15364 8134 15374 8186
rect 15374 8134 15420 8186
rect 15124 8132 15180 8134
rect 15204 8132 15260 8134
rect 15284 8132 15340 8134
rect 15364 8132 15420 8134
rect 15124 7098 15180 7100
rect 15204 7098 15260 7100
rect 15284 7098 15340 7100
rect 15364 7098 15420 7100
rect 15124 7046 15170 7098
rect 15170 7046 15180 7098
rect 15204 7046 15234 7098
rect 15234 7046 15246 7098
rect 15246 7046 15260 7098
rect 15284 7046 15298 7098
rect 15298 7046 15310 7098
rect 15310 7046 15340 7098
rect 15364 7046 15374 7098
rect 15374 7046 15420 7098
rect 15124 7044 15180 7046
rect 15204 7044 15260 7046
rect 15284 7044 15340 7046
rect 15364 7044 15420 7046
rect 15124 6010 15180 6012
rect 15204 6010 15260 6012
rect 15284 6010 15340 6012
rect 15364 6010 15420 6012
rect 15124 5958 15170 6010
rect 15170 5958 15180 6010
rect 15204 5958 15234 6010
rect 15234 5958 15246 6010
rect 15246 5958 15260 6010
rect 15284 5958 15298 6010
rect 15298 5958 15310 6010
rect 15310 5958 15340 6010
rect 15364 5958 15374 6010
rect 15374 5958 15420 6010
rect 15124 5956 15180 5958
rect 15204 5956 15260 5958
rect 15284 5956 15340 5958
rect 15364 5956 15420 5958
rect 15124 4922 15180 4924
rect 15204 4922 15260 4924
rect 15284 4922 15340 4924
rect 15364 4922 15420 4924
rect 15124 4870 15170 4922
rect 15170 4870 15180 4922
rect 15204 4870 15234 4922
rect 15234 4870 15246 4922
rect 15246 4870 15260 4922
rect 15284 4870 15298 4922
rect 15298 4870 15310 4922
rect 15310 4870 15340 4922
rect 15364 4870 15374 4922
rect 15374 4870 15420 4922
rect 15124 4868 15180 4870
rect 15204 4868 15260 4870
rect 15284 4868 15340 4870
rect 15364 4868 15420 4870
rect 15124 3834 15180 3836
rect 15204 3834 15260 3836
rect 15284 3834 15340 3836
rect 15364 3834 15420 3836
rect 15124 3782 15170 3834
rect 15170 3782 15180 3834
rect 15204 3782 15234 3834
rect 15234 3782 15246 3834
rect 15246 3782 15260 3834
rect 15284 3782 15298 3834
rect 15298 3782 15310 3834
rect 15310 3782 15340 3834
rect 15364 3782 15374 3834
rect 15374 3782 15420 3834
rect 15124 3780 15180 3782
rect 15204 3780 15260 3782
rect 15284 3780 15340 3782
rect 15364 3780 15420 3782
rect 17222 7948 17278 7984
rect 17222 7928 17224 7948
rect 17224 7928 17276 7948
rect 17276 7928 17278 7948
rect 15124 2746 15180 2748
rect 15204 2746 15260 2748
rect 15284 2746 15340 2748
rect 15364 2746 15420 2748
rect 15124 2694 15170 2746
rect 15170 2694 15180 2746
rect 15204 2694 15234 2746
rect 15234 2694 15246 2746
rect 15246 2694 15260 2746
rect 15284 2694 15298 2746
rect 15298 2694 15310 2746
rect 15310 2694 15340 2746
rect 15364 2694 15374 2746
rect 15374 2694 15420 2746
rect 15124 2692 15180 2694
rect 15204 2692 15260 2694
rect 15284 2692 15340 2694
rect 15364 2692 15420 2694
rect 19846 26138 19902 26140
rect 19926 26138 19982 26140
rect 20006 26138 20062 26140
rect 20086 26138 20142 26140
rect 19846 26086 19892 26138
rect 19892 26086 19902 26138
rect 19926 26086 19956 26138
rect 19956 26086 19968 26138
rect 19968 26086 19982 26138
rect 20006 26086 20020 26138
rect 20020 26086 20032 26138
rect 20032 26086 20062 26138
rect 20086 26086 20096 26138
rect 20096 26086 20142 26138
rect 19846 26084 19902 26086
rect 19926 26084 19982 26086
rect 20006 26084 20062 26086
rect 20086 26084 20142 26086
rect 19706 25100 19708 25120
rect 19708 25100 19760 25120
rect 19760 25100 19762 25120
rect 19338 21972 19340 21992
rect 19340 21972 19392 21992
rect 19392 21972 19394 21992
rect 19338 21936 19394 21972
rect 19706 25064 19762 25100
rect 19846 25050 19902 25052
rect 19926 25050 19982 25052
rect 20006 25050 20062 25052
rect 20086 25050 20142 25052
rect 19846 24998 19892 25050
rect 19892 24998 19902 25050
rect 19926 24998 19956 25050
rect 19956 24998 19968 25050
rect 19968 24998 19982 25050
rect 20006 24998 20020 25050
rect 20020 24998 20032 25050
rect 20032 24998 20062 25050
rect 20086 24998 20096 25050
rect 20096 24998 20142 25050
rect 19846 24996 19902 24998
rect 19926 24996 19982 24998
rect 20006 24996 20062 24998
rect 20086 24996 20142 24998
rect 19846 23962 19902 23964
rect 19926 23962 19982 23964
rect 20006 23962 20062 23964
rect 20086 23962 20142 23964
rect 19846 23910 19892 23962
rect 19892 23910 19902 23962
rect 19926 23910 19956 23962
rect 19956 23910 19968 23962
rect 19968 23910 19982 23962
rect 20006 23910 20020 23962
rect 20020 23910 20032 23962
rect 20032 23910 20062 23962
rect 20086 23910 20096 23962
rect 20096 23910 20142 23962
rect 19846 23908 19902 23910
rect 19926 23908 19982 23910
rect 20006 23908 20062 23910
rect 20086 23908 20142 23910
rect 19846 22874 19902 22876
rect 19926 22874 19982 22876
rect 20006 22874 20062 22876
rect 20086 22874 20142 22876
rect 19846 22822 19892 22874
rect 19892 22822 19902 22874
rect 19926 22822 19956 22874
rect 19956 22822 19968 22874
rect 19968 22822 19982 22874
rect 20006 22822 20020 22874
rect 20020 22822 20032 22874
rect 20032 22822 20062 22874
rect 20086 22822 20096 22874
rect 20096 22822 20142 22874
rect 19846 22820 19902 22822
rect 19926 22820 19982 22822
rect 20006 22820 20062 22822
rect 20086 22820 20142 22822
rect 19846 21786 19902 21788
rect 19926 21786 19982 21788
rect 20006 21786 20062 21788
rect 20086 21786 20142 21788
rect 19846 21734 19892 21786
rect 19892 21734 19902 21786
rect 19926 21734 19956 21786
rect 19956 21734 19968 21786
rect 19968 21734 19982 21786
rect 20006 21734 20020 21786
rect 20020 21734 20032 21786
rect 20032 21734 20062 21786
rect 20086 21734 20096 21786
rect 20096 21734 20142 21786
rect 19846 21732 19902 21734
rect 19926 21732 19982 21734
rect 20006 21732 20062 21734
rect 20086 21732 20142 21734
rect 19846 20698 19902 20700
rect 19926 20698 19982 20700
rect 20006 20698 20062 20700
rect 20086 20698 20142 20700
rect 19846 20646 19892 20698
rect 19892 20646 19902 20698
rect 19926 20646 19956 20698
rect 19956 20646 19968 20698
rect 19968 20646 19982 20698
rect 20006 20646 20020 20698
rect 20020 20646 20032 20698
rect 20032 20646 20062 20698
rect 20086 20646 20096 20698
rect 20096 20646 20142 20698
rect 19846 20644 19902 20646
rect 19926 20644 19982 20646
rect 20006 20644 20062 20646
rect 20086 20644 20142 20646
rect 19846 19610 19902 19612
rect 19926 19610 19982 19612
rect 20006 19610 20062 19612
rect 20086 19610 20142 19612
rect 19846 19558 19892 19610
rect 19892 19558 19902 19610
rect 19926 19558 19956 19610
rect 19956 19558 19968 19610
rect 19968 19558 19982 19610
rect 20006 19558 20020 19610
rect 20020 19558 20032 19610
rect 20032 19558 20062 19610
rect 20086 19558 20096 19610
rect 20096 19558 20142 19610
rect 19846 19556 19902 19558
rect 19926 19556 19982 19558
rect 20006 19556 20062 19558
rect 20086 19556 20142 19558
rect 19846 18522 19902 18524
rect 19926 18522 19982 18524
rect 20006 18522 20062 18524
rect 20086 18522 20142 18524
rect 19846 18470 19892 18522
rect 19892 18470 19902 18522
rect 19926 18470 19956 18522
rect 19956 18470 19968 18522
rect 19968 18470 19982 18522
rect 20006 18470 20020 18522
rect 20020 18470 20032 18522
rect 20032 18470 20062 18522
rect 20086 18470 20096 18522
rect 20096 18470 20142 18522
rect 19846 18468 19902 18470
rect 19926 18468 19982 18470
rect 20006 18468 20062 18470
rect 20086 18468 20142 18470
rect 19338 14356 19340 14376
rect 19340 14356 19392 14376
rect 19392 14356 19394 14376
rect 19338 14320 19394 14356
rect 18602 12280 18658 12336
rect 20718 29164 20774 29200
rect 20718 29144 20720 29164
rect 20720 29144 20772 29164
rect 20772 29144 20774 29164
rect 20258 19660 20260 19680
rect 20260 19660 20312 19680
rect 20312 19660 20314 19680
rect 20258 19624 20314 19660
rect 19846 17434 19902 17436
rect 19926 17434 19982 17436
rect 20006 17434 20062 17436
rect 20086 17434 20142 17436
rect 19846 17382 19892 17434
rect 19892 17382 19902 17434
rect 19926 17382 19956 17434
rect 19956 17382 19968 17434
rect 19968 17382 19982 17434
rect 20006 17382 20020 17434
rect 20020 17382 20032 17434
rect 20032 17382 20062 17434
rect 20086 17382 20096 17434
rect 20096 17382 20142 17434
rect 19846 17380 19902 17382
rect 19926 17380 19982 17382
rect 20006 17380 20062 17382
rect 20086 17380 20142 17382
rect 19846 16346 19902 16348
rect 19926 16346 19982 16348
rect 20006 16346 20062 16348
rect 20086 16346 20142 16348
rect 19846 16294 19892 16346
rect 19892 16294 19902 16346
rect 19926 16294 19956 16346
rect 19956 16294 19968 16346
rect 19968 16294 19982 16346
rect 20006 16294 20020 16346
rect 20020 16294 20032 16346
rect 20032 16294 20062 16346
rect 20086 16294 20096 16346
rect 20096 16294 20142 16346
rect 19846 16292 19902 16294
rect 19926 16292 19982 16294
rect 20006 16292 20062 16294
rect 20086 16292 20142 16294
rect 19846 15258 19902 15260
rect 19926 15258 19982 15260
rect 20006 15258 20062 15260
rect 20086 15258 20142 15260
rect 19846 15206 19892 15258
rect 19892 15206 19902 15258
rect 19926 15206 19956 15258
rect 19956 15206 19968 15258
rect 19968 15206 19982 15258
rect 20006 15206 20020 15258
rect 20020 15206 20032 15258
rect 20032 15206 20062 15258
rect 20086 15206 20096 15258
rect 20096 15206 20142 15258
rect 19846 15204 19902 15206
rect 19926 15204 19982 15206
rect 20006 15204 20062 15206
rect 20086 15204 20142 15206
rect 20166 14320 20222 14376
rect 19846 14170 19902 14172
rect 19926 14170 19982 14172
rect 20006 14170 20062 14172
rect 20086 14170 20142 14172
rect 19846 14118 19892 14170
rect 19892 14118 19902 14170
rect 19926 14118 19956 14170
rect 19956 14118 19968 14170
rect 19968 14118 19982 14170
rect 20006 14118 20020 14170
rect 20020 14118 20032 14170
rect 20032 14118 20062 14170
rect 20086 14118 20096 14170
rect 20096 14118 20142 14170
rect 19846 14116 19902 14118
rect 19926 14116 19982 14118
rect 20006 14116 20062 14118
rect 20086 14116 20142 14118
rect 19846 13082 19902 13084
rect 19926 13082 19982 13084
rect 20006 13082 20062 13084
rect 20086 13082 20142 13084
rect 19846 13030 19892 13082
rect 19892 13030 19902 13082
rect 19926 13030 19956 13082
rect 19956 13030 19968 13082
rect 19968 13030 19982 13082
rect 20006 13030 20020 13082
rect 20020 13030 20032 13082
rect 20032 13030 20062 13082
rect 20086 13030 20096 13082
rect 20096 13030 20142 13082
rect 19846 13028 19902 13030
rect 19926 13028 19982 13030
rect 20006 13028 20062 13030
rect 20086 13028 20142 13030
rect 19846 11994 19902 11996
rect 19926 11994 19982 11996
rect 20006 11994 20062 11996
rect 20086 11994 20142 11996
rect 19846 11942 19892 11994
rect 19892 11942 19902 11994
rect 19926 11942 19956 11994
rect 19956 11942 19968 11994
rect 19968 11942 19982 11994
rect 20006 11942 20020 11994
rect 20020 11942 20032 11994
rect 20032 11942 20062 11994
rect 20086 11942 20096 11994
rect 20096 11942 20142 11994
rect 19846 11940 19902 11942
rect 19926 11940 19982 11942
rect 20006 11940 20062 11942
rect 20086 11940 20142 11942
rect 19846 10906 19902 10908
rect 19926 10906 19982 10908
rect 20006 10906 20062 10908
rect 20086 10906 20142 10908
rect 19846 10854 19892 10906
rect 19892 10854 19902 10906
rect 19926 10854 19956 10906
rect 19956 10854 19968 10906
rect 19968 10854 19982 10906
rect 20006 10854 20020 10906
rect 20020 10854 20032 10906
rect 20032 10854 20062 10906
rect 20086 10854 20096 10906
rect 20096 10854 20142 10906
rect 19846 10852 19902 10854
rect 19926 10852 19982 10854
rect 20006 10852 20062 10854
rect 20086 10852 20142 10854
rect 19846 9818 19902 9820
rect 19926 9818 19982 9820
rect 20006 9818 20062 9820
rect 20086 9818 20142 9820
rect 19846 9766 19892 9818
rect 19892 9766 19902 9818
rect 19926 9766 19956 9818
rect 19956 9766 19968 9818
rect 19968 9766 19982 9818
rect 20006 9766 20020 9818
rect 20020 9766 20032 9818
rect 20032 9766 20062 9818
rect 20086 9766 20096 9818
rect 20096 9766 20142 9818
rect 19846 9764 19902 9766
rect 19926 9764 19982 9766
rect 20006 9764 20062 9766
rect 20086 9764 20142 9766
rect 19846 8730 19902 8732
rect 19926 8730 19982 8732
rect 20006 8730 20062 8732
rect 20086 8730 20142 8732
rect 19846 8678 19892 8730
rect 19892 8678 19902 8730
rect 19926 8678 19956 8730
rect 19956 8678 19968 8730
rect 19968 8678 19982 8730
rect 20006 8678 20020 8730
rect 20020 8678 20032 8730
rect 20032 8678 20062 8730
rect 20086 8678 20096 8730
rect 20096 8678 20142 8730
rect 19846 8676 19902 8678
rect 19926 8676 19982 8678
rect 20006 8676 20062 8678
rect 20086 8676 20142 8678
rect 19338 8356 19394 8392
rect 19338 8336 19340 8356
rect 19340 8336 19392 8356
rect 19392 8336 19394 8356
rect 19846 7642 19902 7644
rect 19926 7642 19982 7644
rect 20006 7642 20062 7644
rect 20086 7642 20142 7644
rect 19846 7590 19892 7642
rect 19892 7590 19902 7642
rect 19926 7590 19956 7642
rect 19956 7590 19968 7642
rect 19968 7590 19982 7642
rect 20006 7590 20020 7642
rect 20020 7590 20032 7642
rect 20032 7590 20062 7642
rect 20086 7590 20096 7642
rect 20096 7590 20142 7642
rect 19846 7588 19902 7590
rect 19926 7588 19982 7590
rect 20006 7588 20062 7590
rect 20086 7588 20142 7590
rect 19846 6554 19902 6556
rect 19926 6554 19982 6556
rect 20006 6554 20062 6556
rect 20086 6554 20142 6556
rect 19846 6502 19892 6554
rect 19892 6502 19902 6554
rect 19926 6502 19956 6554
rect 19956 6502 19968 6554
rect 19968 6502 19982 6554
rect 20006 6502 20020 6554
rect 20020 6502 20032 6554
rect 20032 6502 20062 6554
rect 20086 6502 20096 6554
rect 20096 6502 20142 6554
rect 19846 6500 19902 6502
rect 19926 6500 19982 6502
rect 20006 6500 20062 6502
rect 20086 6500 20142 6502
rect 19846 5466 19902 5468
rect 19926 5466 19982 5468
rect 20006 5466 20062 5468
rect 20086 5466 20142 5468
rect 19846 5414 19892 5466
rect 19892 5414 19902 5466
rect 19926 5414 19956 5466
rect 19956 5414 19968 5466
rect 19968 5414 19982 5466
rect 20006 5414 20020 5466
rect 20020 5414 20032 5466
rect 20032 5414 20062 5466
rect 20086 5414 20096 5466
rect 20096 5414 20142 5466
rect 19846 5412 19902 5414
rect 19926 5412 19982 5414
rect 20006 5412 20062 5414
rect 20086 5412 20142 5414
rect 19846 4378 19902 4380
rect 19926 4378 19982 4380
rect 20006 4378 20062 4380
rect 20086 4378 20142 4380
rect 19846 4326 19892 4378
rect 19892 4326 19902 4378
rect 19926 4326 19956 4378
rect 19956 4326 19968 4378
rect 19968 4326 19982 4378
rect 20006 4326 20020 4378
rect 20020 4326 20032 4378
rect 20032 4326 20062 4378
rect 20086 4326 20096 4378
rect 20096 4326 20142 4378
rect 19846 4324 19902 4326
rect 19926 4324 19982 4326
rect 20006 4324 20062 4326
rect 20086 4324 20142 4326
rect 19846 3290 19902 3292
rect 19926 3290 19982 3292
rect 20006 3290 20062 3292
rect 20086 3290 20142 3292
rect 19846 3238 19892 3290
rect 19892 3238 19902 3290
rect 19926 3238 19956 3290
rect 19956 3238 19968 3290
rect 19968 3238 19982 3290
rect 20006 3238 20020 3290
rect 20020 3238 20032 3290
rect 20032 3238 20062 3290
rect 20086 3238 20096 3290
rect 20096 3238 20142 3290
rect 19846 3236 19902 3238
rect 19926 3236 19982 3238
rect 20006 3236 20062 3238
rect 20086 3236 20142 3238
rect 19846 2202 19902 2204
rect 19926 2202 19982 2204
rect 20006 2202 20062 2204
rect 20086 2202 20142 2204
rect 19846 2150 19892 2202
rect 19892 2150 19902 2202
rect 19926 2150 19956 2202
rect 19956 2150 19968 2202
rect 19968 2150 19982 2202
rect 20006 2150 20020 2202
rect 20020 2150 20032 2202
rect 20032 2150 20062 2202
rect 20086 2150 20096 2202
rect 20096 2150 20142 2202
rect 19846 2148 19902 2150
rect 19926 2148 19982 2150
rect 20006 2148 20062 2150
rect 20086 2148 20142 2150
rect 20350 8608 20406 8664
rect 22742 29164 22798 29200
rect 22742 29144 22744 29164
rect 22744 29144 22796 29164
rect 22796 29144 22798 29164
rect 22282 21548 22338 21584
rect 22282 21528 22284 21548
rect 22284 21528 22336 21548
rect 22336 21528 22338 21548
rect 23294 25900 23350 25936
rect 23294 25880 23296 25900
rect 23296 25880 23348 25900
rect 23348 25880 23350 25900
rect 23386 25220 23442 25256
rect 23386 25200 23388 25220
rect 23388 25200 23440 25220
rect 23440 25200 23442 25220
rect 23294 25064 23350 25120
rect 22650 21528 22706 21584
rect 21178 18264 21234 18320
rect 23754 25064 23810 25120
rect 24569 29946 24625 29948
rect 24649 29946 24705 29948
rect 24729 29946 24785 29948
rect 24809 29946 24865 29948
rect 24569 29894 24615 29946
rect 24615 29894 24625 29946
rect 24649 29894 24679 29946
rect 24679 29894 24691 29946
rect 24691 29894 24705 29946
rect 24729 29894 24743 29946
rect 24743 29894 24755 29946
rect 24755 29894 24785 29946
rect 24809 29894 24819 29946
rect 24819 29894 24865 29946
rect 24569 29892 24625 29894
rect 24649 29892 24705 29894
rect 24729 29892 24785 29894
rect 24809 29892 24865 29894
rect 26146 31592 26202 31648
rect 26238 29688 26294 29744
rect 24569 28858 24625 28860
rect 24649 28858 24705 28860
rect 24729 28858 24785 28860
rect 24809 28858 24865 28860
rect 24569 28806 24615 28858
rect 24615 28806 24625 28858
rect 24649 28806 24679 28858
rect 24679 28806 24691 28858
rect 24691 28806 24705 28858
rect 24729 28806 24743 28858
rect 24743 28806 24755 28858
rect 24755 28806 24785 28858
rect 24809 28806 24819 28858
rect 24819 28806 24865 28858
rect 24569 28804 24625 28806
rect 24649 28804 24705 28806
rect 24729 28804 24785 28806
rect 24809 28804 24865 28806
rect 24569 27770 24625 27772
rect 24649 27770 24705 27772
rect 24729 27770 24785 27772
rect 24809 27770 24865 27772
rect 24569 27718 24615 27770
rect 24615 27718 24625 27770
rect 24649 27718 24679 27770
rect 24679 27718 24691 27770
rect 24691 27718 24705 27770
rect 24729 27718 24743 27770
rect 24743 27718 24755 27770
rect 24755 27718 24785 27770
rect 24809 27718 24819 27770
rect 24819 27718 24865 27770
rect 24569 27716 24625 27718
rect 24649 27716 24705 27718
rect 24729 27716 24785 27718
rect 24809 27716 24865 27718
rect 24569 26682 24625 26684
rect 24649 26682 24705 26684
rect 24729 26682 24785 26684
rect 24809 26682 24865 26684
rect 24569 26630 24615 26682
rect 24615 26630 24625 26682
rect 24649 26630 24679 26682
rect 24679 26630 24691 26682
rect 24691 26630 24705 26682
rect 24729 26630 24743 26682
rect 24743 26630 24755 26682
rect 24755 26630 24785 26682
rect 24809 26630 24819 26682
rect 24819 26630 24865 26682
rect 24569 26628 24625 26630
rect 24649 26628 24705 26630
rect 24729 26628 24785 26630
rect 24809 26628 24865 26630
rect 24569 25594 24625 25596
rect 24649 25594 24705 25596
rect 24729 25594 24785 25596
rect 24809 25594 24865 25596
rect 24569 25542 24615 25594
rect 24615 25542 24625 25594
rect 24649 25542 24679 25594
rect 24679 25542 24691 25594
rect 24691 25542 24705 25594
rect 24729 25542 24743 25594
rect 24743 25542 24755 25594
rect 24755 25542 24785 25594
rect 24809 25542 24819 25594
rect 24819 25542 24865 25594
rect 24569 25540 24625 25542
rect 24649 25540 24705 25542
rect 24729 25540 24785 25542
rect 24809 25540 24865 25542
rect 26790 27784 26846 27840
rect 26238 25880 26294 25936
rect 22650 17076 22652 17096
rect 22652 17076 22704 17096
rect 22704 17076 22706 17096
rect 22650 17040 22706 17076
rect 21178 16244 21234 16280
rect 21178 16224 21180 16244
rect 21180 16224 21232 16244
rect 21232 16224 21234 16244
rect 21178 12144 21234 12200
rect 21454 8608 21510 8664
rect 21362 8336 21418 8392
rect 24569 24506 24625 24508
rect 24649 24506 24705 24508
rect 24729 24506 24785 24508
rect 24809 24506 24865 24508
rect 24569 24454 24615 24506
rect 24615 24454 24625 24506
rect 24649 24454 24679 24506
rect 24679 24454 24691 24506
rect 24691 24454 24705 24506
rect 24729 24454 24743 24506
rect 24743 24454 24755 24506
rect 24755 24454 24785 24506
rect 24809 24454 24819 24506
rect 24819 24454 24865 24506
rect 24569 24452 24625 24454
rect 24649 24452 24705 24454
rect 24729 24452 24785 24454
rect 24809 24452 24865 24454
rect 24569 23418 24625 23420
rect 24649 23418 24705 23420
rect 24729 23418 24785 23420
rect 24809 23418 24865 23420
rect 24569 23366 24615 23418
rect 24615 23366 24625 23418
rect 24649 23366 24679 23418
rect 24679 23366 24691 23418
rect 24691 23366 24705 23418
rect 24729 23366 24743 23418
rect 24743 23366 24755 23418
rect 24755 23366 24785 23418
rect 24809 23366 24819 23418
rect 24819 23366 24865 23418
rect 24569 23364 24625 23366
rect 24649 23364 24705 23366
rect 24729 23364 24785 23366
rect 24809 23364 24865 23366
rect 24569 22330 24625 22332
rect 24649 22330 24705 22332
rect 24729 22330 24785 22332
rect 24809 22330 24865 22332
rect 24569 22278 24615 22330
rect 24615 22278 24625 22330
rect 24649 22278 24679 22330
rect 24679 22278 24691 22330
rect 24691 22278 24705 22330
rect 24729 22278 24743 22330
rect 24743 22278 24755 22330
rect 24755 22278 24785 22330
rect 24809 22278 24819 22330
rect 24819 22278 24865 22330
rect 24569 22276 24625 22278
rect 24649 22276 24705 22278
rect 24729 22276 24785 22278
rect 24809 22276 24865 22278
rect 24569 21242 24625 21244
rect 24649 21242 24705 21244
rect 24729 21242 24785 21244
rect 24809 21242 24865 21244
rect 24569 21190 24615 21242
rect 24615 21190 24625 21242
rect 24649 21190 24679 21242
rect 24679 21190 24691 21242
rect 24691 21190 24705 21242
rect 24729 21190 24743 21242
rect 24743 21190 24755 21242
rect 24755 21190 24785 21242
rect 24809 21190 24819 21242
rect 24819 21190 24865 21242
rect 24569 21188 24625 21190
rect 24649 21188 24705 21190
rect 24729 21188 24785 21190
rect 24809 21188 24865 21190
rect 24569 20154 24625 20156
rect 24649 20154 24705 20156
rect 24729 20154 24785 20156
rect 24809 20154 24865 20156
rect 24569 20102 24615 20154
rect 24615 20102 24625 20154
rect 24649 20102 24679 20154
rect 24679 20102 24691 20154
rect 24691 20102 24705 20154
rect 24729 20102 24743 20154
rect 24743 20102 24755 20154
rect 24755 20102 24785 20154
rect 24809 20102 24819 20154
rect 24819 20102 24865 20154
rect 24569 20100 24625 20102
rect 24649 20100 24705 20102
rect 24729 20100 24785 20102
rect 24809 20100 24865 20102
rect 24569 19066 24625 19068
rect 24649 19066 24705 19068
rect 24729 19066 24785 19068
rect 24809 19066 24865 19068
rect 24569 19014 24615 19066
rect 24615 19014 24625 19066
rect 24649 19014 24679 19066
rect 24679 19014 24691 19066
rect 24691 19014 24705 19066
rect 24729 19014 24743 19066
rect 24743 19014 24755 19066
rect 24755 19014 24785 19066
rect 24809 19014 24819 19066
rect 24819 19014 24865 19066
rect 24569 19012 24625 19014
rect 24649 19012 24705 19014
rect 24729 19012 24785 19014
rect 24809 19012 24865 19014
rect 24569 17978 24625 17980
rect 24649 17978 24705 17980
rect 24729 17978 24785 17980
rect 24809 17978 24865 17980
rect 24569 17926 24615 17978
rect 24615 17926 24625 17978
rect 24649 17926 24679 17978
rect 24679 17926 24691 17978
rect 24691 17926 24705 17978
rect 24729 17926 24743 17978
rect 24743 17926 24755 17978
rect 24755 17926 24785 17978
rect 24809 17926 24819 17978
rect 24819 17926 24865 17978
rect 24569 17924 24625 17926
rect 24649 17924 24705 17926
rect 24729 17924 24785 17926
rect 24809 17924 24865 17926
rect 24766 17212 24768 17232
rect 24768 17212 24820 17232
rect 24820 17212 24822 17232
rect 24766 17176 24822 17212
rect 24569 16890 24625 16892
rect 24649 16890 24705 16892
rect 24729 16890 24785 16892
rect 24809 16890 24865 16892
rect 24569 16838 24615 16890
rect 24615 16838 24625 16890
rect 24649 16838 24679 16890
rect 24679 16838 24691 16890
rect 24691 16838 24705 16890
rect 24729 16838 24743 16890
rect 24743 16838 24755 16890
rect 24755 16838 24785 16890
rect 24809 16838 24819 16890
rect 24819 16838 24865 16890
rect 24569 16836 24625 16838
rect 24649 16836 24705 16838
rect 24729 16836 24785 16838
rect 24809 16836 24865 16838
rect 24569 15802 24625 15804
rect 24649 15802 24705 15804
rect 24729 15802 24785 15804
rect 24809 15802 24865 15804
rect 24569 15750 24615 15802
rect 24615 15750 24625 15802
rect 24649 15750 24679 15802
rect 24679 15750 24691 15802
rect 24691 15750 24705 15802
rect 24729 15750 24743 15802
rect 24743 15750 24755 15802
rect 24755 15750 24785 15802
rect 24809 15750 24819 15802
rect 24819 15750 24865 15802
rect 24569 15748 24625 15750
rect 24649 15748 24705 15750
rect 24729 15748 24785 15750
rect 24809 15748 24865 15750
rect 24569 14714 24625 14716
rect 24649 14714 24705 14716
rect 24729 14714 24785 14716
rect 24809 14714 24865 14716
rect 24569 14662 24615 14714
rect 24615 14662 24625 14714
rect 24649 14662 24679 14714
rect 24679 14662 24691 14714
rect 24691 14662 24705 14714
rect 24729 14662 24743 14714
rect 24743 14662 24755 14714
rect 24755 14662 24785 14714
rect 24809 14662 24819 14714
rect 24819 14662 24865 14714
rect 24569 14660 24625 14662
rect 24649 14660 24705 14662
rect 24729 14660 24785 14662
rect 24809 14660 24865 14662
rect 24569 13626 24625 13628
rect 24649 13626 24705 13628
rect 24729 13626 24785 13628
rect 24809 13626 24865 13628
rect 24569 13574 24615 13626
rect 24615 13574 24625 13626
rect 24649 13574 24679 13626
rect 24679 13574 24691 13626
rect 24691 13574 24705 13626
rect 24729 13574 24743 13626
rect 24743 13574 24755 13626
rect 24755 13574 24785 13626
rect 24809 13574 24819 13626
rect 24819 13574 24865 13626
rect 24569 13572 24625 13574
rect 24649 13572 24705 13574
rect 24729 13572 24785 13574
rect 24809 13572 24865 13574
rect 24569 12538 24625 12540
rect 24649 12538 24705 12540
rect 24729 12538 24785 12540
rect 24809 12538 24865 12540
rect 24569 12486 24615 12538
rect 24615 12486 24625 12538
rect 24649 12486 24679 12538
rect 24679 12486 24691 12538
rect 24691 12486 24705 12538
rect 24729 12486 24743 12538
rect 24743 12486 24755 12538
rect 24755 12486 24785 12538
rect 24809 12486 24819 12538
rect 24819 12486 24865 12538
rect 24569 12484 24625 12486
rect 24649 12484 24705 12486
rect 24729 12484 24785 12486
rect 24809 12484 24865 12486
rect 26238 23976 26294 24032
rect 26330 22072 26386 22128
rect 27526 20168 27582 20224
rect 24569 11450 24625 11452
rect 24649 11450 24705 11452
rect 24729 11450 24785 11452
rect 24809 11450 24865 11452
rect 24569 11398 24615 11450
rect 24615 11398 24625 11450
rect 24649 11398 24679 11450
rect 24679 11398 24691 11450
rect 24691 11398 24705 11450
rect 24729 11398 24743 11450
rect 24743 11398 24755 11450
rect 24755 11398 24785 11450
rect 24809 11398 24819 11450
rect 24819 11398 24865 11450
rect 24569 11396 24625 11398
rect 24649 11396 24705 11398
rect 24729 11396 24785 11398
rect 24809 11396 24865 11398
rect 23662 9424 23718 9480
rect 24569 10362 24625 10364
rect 24649 10362 24705 10364
rect 24729 10362 24785 10364
rect 24809 10362 24865 10364
rect 24569 10310 24615 10362
rect 24615 10310 24625 10362
rect 24649 10310 24679 10362
rect 24679 10310 24691 10362
rect 24691 10310 24705 10362
rect 24729 10310 24743 10362
rect 24743 10310 24755 10362
rect 24755 10310 24785 10362
rect 24809 10310 24819 10362
rect 24819 10310 24865 10362
rect 24569 10308 24625 10310
rect 24649 10308 24705 10310
rect 24729 10308 24785 10310
rect 24809 10308 24865 10310
rect 24569 9274 24625 9276
rect 24649 9274 24705 9276
rect 24729 9274 24785 9276
rect 24809 9274 24865 9276
rect 24569 9222 24615 9274
rect 24615 9222 24625 9274
rect 24649 9222 24679 9274
rect 24679 9222 24691 9274
rect 24691 9222 24705 9274
rect 24729 9222 24743 9274
rect 24743 9222 24755 9274
rect 24755 9222 24785 9274
rect 24809 9222 24819 9274
rect 24819 9222 24865 9274
rect 24569 9220 24625 9222
rect 24649 9220 24705 9222
rect 24729 9220 24785 9222
rect 24809 9220 24865 9222
rect 24490 8336 24546 8392
rect 24569 8186 24625 8188
rect 24649 8186 24705 8188
rect 24729 8186 24785 8188
rect 24809 8186 24865 8188
rect 24569 8134 24615 8186
rect 24615 8134 24625 8186
rect 24649 8134 24679 8186
rect 24679 8134 24691 8186
rect 24691 8134 24705 8186
rect 24729 8134 24743 8186
rect 24743 8134 24755 8186
rect 24755 8134 24785 8186
rect 24809 8134 24819 8186
rect 24819 8134 24865 8186
rect 24569 8132 24625 8134
rect 24649 8132 24705 8134
rect 24729 8132 24785 8134
rect 24809 8132 24865 8134
rect 24569 7098 24625 7100
rect 24649 7098 24705 7100
rect 24729 7098 24785 7100
rect 24809 7098 24865 7100
rect 24569 7046 24615 7098
rect 24615 7046 24625 7098
rect 24649 7046 24679 7098
rect 24679 7046 24691 7098
rect 24691 7046 24705 7098
rect 24729 7046 24743 7098
rect 24743 7046 24755 7098
rect 24755 7046 24785 7098
rect 24809 7046 24819 7098
rect 24819 7046 24865 7098
rect 24569 7044 24625 7046
rect 24649 7044 24705 7046
rect 24729 7044 24785 7046
rect 24809 7044 24865 7046
rect 24569 6010 24625 6012
rect 24649 6010 24705 6012
rect 24729 6010 24785 6012
rect 24809 6010 24865 6012
rect 24569 5958 24615 6010
rect 24615 5958 24625 6010
rect 24649 5958 24679 6010
rect 24679 5958 24691 6010
rect 24691 5958 24705 6010
rect 24729 5958 24743 6010
rect 24743 5958 24755 6010
rect 24755 5958 24785 6010
rect 24809 5958 24819 6010
rect 24819 5958 24865 6010
rect 24569 5956 24625 5958
rect 24649 5956 24705 5958
rect 24729 5956 24785 5958
rect 24809 5956 24865 5958
rect 24569 4922 24625 4924
rect 24649 4922 24705 4924
rect 24729 4922 24785 4924
rect 24809 4922 24865 4924
rect 24569 4870 24615 4922
rect 24615 4870 24625 4922
rect 24649 4870 24679 4922
rect 24679 4870 24691 4922
rect 24691 4870 24705 4922
rect 24729 4870 24743 4922
rect 24743 4870 24755 4922
rect 24755 4870 24785 4922
rect 24809 4870 24819 4922
rect 24819 4870 24865 4922
rect 24569 4868 24625 4870
rect 24649 4868 24705 4870
rect 24729 4868 24785 4870
rect 24809 4868 24865 4870
rect 23938 3032 23994 3088
rect 24569 3834 24625 3836
rect 24649 3834 24705 3836
rect 24729 3834 24785 3836
rect 24809 3834 24865 3836
rect 24569 3782 24615 3834
rect 24615 3782 24625 3834
rect 24649 3782 24679 3834
rect 24679 3782 24691 3834
rect 24691 3782 24705 3834
rect 24729 3782 24743 3834
rect 24743 3782 24755 3834
rect 24755 3782 24785 3834
rect 24809 3782 24819 3834
rect 24819 3782 24865 3834
rect 24569 3780 24625 3782
rect 24649 3780 24705 3782
rect 24729 3780 24785 3782
rect 24809 3780 24865 3782
rect 26514 12416 26570 12472
rect 26238 10512 26294 10568
rect 26790 14320 26846 14376
rect 26698 8608 26754 8664
rect 26238 6704 26294 6760
rect 26238 4800 26294 4856
rect 24569 2746 24625 2748
rect 24649 2746 24705 2748
rect 24729 2746 24785 2748
rect 24809 2746 24865 2748
rect 24569 2694 24615 2746
rect 24615 2694 24625 2746
rect 24649 2694 24679 2746
rect 24679 2694 24691 2746
rect 24691 2694 24705 2746
rect 24729 2694 24743 2746
rect 24743 2694 24755 2746
rect 24755 2694 24785 2746
rect 24809 2694 24819 2746
rect 24819 2694 24865 2746
rect 24569 2692 24625 2694
rect 24649 2692 24705 2694
rect 24729 2692 24785 2694
rect 24809 2692 24865 2694
rect 25962 3440 26018 3496
rect 26330 2916 26386 2952
rect 26330 2896 26332 2916
rect 26332 2896 26384 2916
rect 26384 2896 26386 2916
rect 26238 992 26294 1048
<< metal3 >>
rect 0 32058 800 32088
rect 3969 32058 4035 32061
rect 0 32056 4035 32058
rect 0 32000 3974 32056
rect 4030 32000 4035 32056
rect 0 31998 4035 32000
rect 0 31968 800 31998
rect 3969 31995 4035 31998
rect 26141 31650 26207 31653
rect 29745 31650 30545 31680
rect 26141 31648 30545 31650
rect 26141 31592 26146 31648
rect 26202 31592 30545 31648
rect 26141 31590 30545 31592
rect 26141 31587 26207 31590
rect 29745 31560 30545 31590
rect 0 30698 800 30728
rect 4061 30698 4127 30701
rect 0 30696 4127 30698
rect 0 30640 4066 30696
rect 4122 30640 4127 30696
rect 0 30638 4127 30640
rect 0 30608 800 30638
rect 4061 30635 4127 30638
rect 10389 30496 10709 30497
rect 10389 30432 10397 30496
rect 10461 30432 10477 30496
rect 10541 30432 10557 30496
rect 10621 30432 10637 30496
rect 10701 30432 10709 30496
rect 10389 30431 10709 30432
rect 19834 30496 20154 30497
rect 19834 30432 19842 30496
rect 19906 30432 19922 30496
rect 19986 30432 20002 30496
rect 20066 30432 20082 30496
rect 20146 30432 20154 30496
rect 19834 30431 20154 30432
rect 5666 29952 5986 29953
rect 5666 29888 5674 29952
rect 5738 29888 5754 29952
rect 5818 29888 5834 29952
rect 5898 29888 5914 29952
rect 5978 29888 5986 29952
rect 5666 29887 5986 29888
rect 15112 29952 15432 29953
rect 15112 29888 15120 29952
rect 15184 29888 15200 29952
rect 15264 29888 15280 29952
rect 15344 29888 15360 29952
rect 15424 29888 15432 29952
rect 15112 29887 15432 29888
rect 24557 29952 24877 29953
rect 24557 29888 24565 29952
rect 24629 29888 24645 29952
rect 24709 29888 24725 29952
rect 24789 29888 24805 29952
rect 24869 29888 24877 29952
rect 24557 29887 24877 29888
rect 26233 29746 26299 29749
rect 29745 29746 30545 29776
rect 26233 29744 30545 29746
rect 26233 29688 26238 29744
rect 26294 29688 30545 29744
rect 26233 29686 30545 29688
rect 26233 29683 26299 29686
rect 29745 29656 30545 29686
rect 10389 29408 10709 29409
rect 0 29338 800 29368
rect 10389 29344 10397 29408
rect 10461 29344 10477 29408
rect 10541 29344 10557 29408
rect 10621 29344 10637 29408
rect 10701 29344 10709 29408
rect 10389 29343 10709 29344
rect 19834 29408 20154 29409
rect 19834 29344 19842 29408
rect 19906 29344 19922 29408
rect 19986 29344 20002 29408
rect 20066 29344 20082 29408
rect 20146 29344 20154 29408
rect 19834 29343 20154 29344
rect 4061 29338 4127 29341
rect 0 29336 4127 29338
rect 0 29280 4066 29336
rect 4122 29280 4127 29336
rect 0 29278 4127 29280
rect 0 29248 800 29278
rect 4061 29275 4127 29278
rect 20713 29202 20779 29205
rect 22737 29202 22803 29205
rect 20713 29200 22803 29202
rect 20713 29144 20718 29200
rect 20774 29144 22742 29200
rect 22798 29144 22803 29200
rect 20713 29142 22803 29144
rect 20713 29139 20779 29142
rect 22737 29139 22803 29142
rect 5666 28864 5986 28865
rect 5666 28800 5674 28864
rect 5738 28800 5754 28864
rect 5818 28800 5834 28864
rect 5898 28800 5914 28864
rect 5978 28800 5986 28864
rect 5666 28799 5986 28800
rect 15112 28864 15432 28865
rect 15112 28800 15120 28864
rect 15184 28800 15200 28864
rect 15264 28800 15280 28864
rect 15344 28800 15360 28864
rect 15424 28800 15432 28864
rect 15112 28799 15432 28800
rect 24557 28864 24877 28865
rect 24557 28800 24565 28864
rect 24629 28800 24645 28864
rect 24709 28800 24725 28864
rect 24789 28800 24805 28864
rect 24869 28800 24877 28864
rect 24557 28799 24877 28800
rect 10389 28320 10709 28321
rect 10389 28256 10397 28320
rect 10461 28256 10477 28320
rect 10541 28256 10557 28320
rect 10621 28256 10637 28320
rect 10701 28256 10709 28320
rect 10389 28255 10709 28256
rect 19834 28320 20154 28321
rect 19834 28256 19842 28320
rect 19906 28256 19922 28320
rect 19986 28256 20002 28320
rect 20066 28256 20082 28320
rect 20146 28256 20154 28320
rect 19834 28255 20154 28256
rect 0 27978 800 28008
rect 4061 27978 4127 27981
rect 0 27976 4127 27978
rect 0 27920 4066 27976
rect 4122 27920 4127 27976
rect 0 27918 4127 27920
rect 0 27888 800 27918
rect 4061 27915 4127 27918
rect 26785 27842 26851 27845
rect 29745 27842 30545 27872
rect 26785 27840 30545 27842
rect 26785 27784 26790 27840
rect 26846 27784 30545 27840
rect 26785 27782 30545 27784
rect 26785 27779 26851 27782
rect 5666 27776 5986 27777
rect 5666 27712 5674 27776
rect 5738 27712 5754 27776
rect 5818 27712 5834 27776
rect 5898 27712 5914 27776
rect 5978 27712 5986 27776
rect 5666 27711 5986 27712
rect 15112 27776 15432 27777
rect 15112 27712 15120 27776
rect 15184 27712 15200 27776
rect 15264 27712 15280 27776
rect 15344 27712 15360 27776
rect 15424 27712 15432 27776
rect 15112 27711 15432 27712
rect 24557 27776 24877 27777
rect 24557 27712 24565 27776
rect 24629 27712 24645 27776
rect 24709 27712 24725 27776
rect 24789 27712 24805 27776
rect 24869 27712 24877 27776
rect 29745 27752 30545 27782
rect 24557 27711 24877 27712
rect 17861 27434 17927 27437
rect 19701 27434 19767 27437
rect 17861 27432 19767 27434
rect 17861 27376 17866 27432
rect 17922 27376 19706 27432
rect 19762 27376 19767 27432
rect 17861 27374 19767 27376
rect 17861 27371 17927 27374
rect 19701 27371 19767 27374
rect 10389 27232 10709 27233
rect 10389 27168 10397 27232
rect 10461 27168 10477 27232
rect 10541 27168 10557 27232
rect 10621 27168 10637 27232
rect 10701 27168 10709 27232
rect 10389 27167 10709 27168
rect 19834 27232 20154 27233
rect 19834 27168 19842 27232
rect 19906 27168 19922 27232
rect 19986 27168 20002 27232
rect 20066 27168 20082 27232
rect 20146 27168 20154 27232
rect 19834 27167 20154 27168
rect 12617 27162 12683 27165
rect 15193 27162 15259 27165
rect 12617 27160 15259 27162
rect 12617 27104 12622 27160
rect 12678 27104 15198 27160
rect 15254 27104 15259 27160
rect 12617 27102 15259 27104
rect 12617 27099 12683 27102
rect 15193 27099 15259 27102
rect 17401 27026 17467 27029
rect 18781 27026 18847 27029
rect 17401 27024 18847 27026
rect 17401 26968 17406 27024
rect 17462 26968 18786 27024
rect 18842 26968 18847 27024
rect 17401 26966 18847 26968
rect 17401 26963 17467 26966
rect 18781 26963 18847 26966
rect 5666 26688 5986 26689
rect 0 26618 800 26648
rect 5666 26624 5674 26688
rect 5738 26624 5754 26688
rect 5818 26624 5834 26688
rect 5898 26624 5914 26688
rect 5978 26624 5986 26688
rect 5666 26623 5986 26624
rect 15112 26688 15432 26689
rect 15112 26624 15120 26688
rect 15184 26624 15200 26688
rect 15264 26624 15280 26688
rect 15344 26624 15360 26688
rect 15424 26624 15432 26688
rect 15112 26623 15432 26624
rect 24557 26688 24877 26689
rect 24557 26624 24565 26688
rect 24629 26624 24645 26688
rect 24709 26624 24725 26688
rect 24789 26624 24805 26688
rect 24869 26624 24877 26688
rect 24557 26623 24877 26624
rect 4061 26618 4127 26621
rect 0 26616 4127 26618
rect 0 26560 4066 26616
rect 4122 26560 4127 26616
rect 0 26558 4127 26560
rect 0 26528 800 26558
rect 4061 26555 4127 26558
rect 10041 26346 10107 26349
rect 15561 26346 15627 26349
rect 10041 26344 15627 26346
rect 10041 26288 10046 26344
rect 10102 26288 15566 26344
rect 15622 26288 15627 26344
rect 10041 26286 15627 26288
rect 10041 26283 10107 26286
rect 15561 26283 15627 26286
rect 10389 26144 10709 26145
rect 10389 26080 10397 26144
rect 10461 26080 10477 26144
rect 10541 26080 10557 26144
rect 10621 26080 10637 26144
rect 10701 26080 10709 26144
rect 10389 26079 10709 26080
rect 19834 26144 20154 26145
rect 19834 26080 19842 26144
rect 19906 26080 19922 26144
rect 19986 26080 20002 26144
rect 20066 26080 20082 26144
rect 20146 26080 20154 26144
rect 19834 26079 20154 26080
rect 23289 25938 23355 25941
rect 2730 25936 23355 25938
rect 2730 25880 23294 25936
rect 23350 25880 23355 25936
rect 2730 25878 23355 25880
rect 0 25258 800 25288
rect 2730 25258 2790 25878
rect 23289 25875 23355 25878
rect 26233 25938 26299 25941
rect 29745 25938 30545 25968
rect 26233 25936 30545 25938
rect 26233 25880 26238 25936
rect 26294 25880 30545 25936
rect 26233 25878 30545 25880
rect 26233 25875 26299 25878
rect 29745 25848 30545 25878
rect 11697 25802 11763 25805
rect 13169 25802 13235 25805
rect 11697 25800 13235 25802
rect 11697 25744 11702 25800
rect 11758 25744 13174 25800
rect 13230 25744 13235 25800
rect 11697 25742 13235 25744
rect 11697 25739 11763 25742
rect 13169 25739 13235 25742
rect 12525 25668 12591 25669
rect 12525 25666 12572 25668
rect 12480 25664 12572 25666
rect 12480 25608 12530 25664
rect 12480 25606 12572 25608
rect 12525 25604 12572 25606
rect 12636 25604 12642 25668
rect 12525 25603 12591 25604
rect 5666 25600 5986 25601
rect 5666 25536 5674 25600
rect 5738 25536 5754 25600
rect 5818 25536 5834 25600
rect 5898 25536 5914 25600
rect 5978 25536 5986 25600
rect 5666 25535 5986 25536
rect 15112 25600 15432 25601
rect 15112 25536 15120 25600
rect 15184 25536 15200 25600
rect 15264 25536 15280 25600
rect 15344 25536 15360 25600
rect 15424 25536 15432 25600
rect 15112 25535 15432 25536
rect 24557 25600 24877 25601
rect 24557 25536 24565 25600
rect 24629 25536 24645 25600
rect 24709 25536 24725 25600
rect 24789 25536 24805 25600
rect 24869 25536 24877 25600
rect 24557 25535 24877 25536
rect 0 25198 2790 25258
rect 15561 25258 15627 25261
rect 15837 25258 15903 25261
rect 23381 25258 23447 25261
rect 15561 25256 23447 25258
rect 15561 25200 15566 25256
rect 15622 25200 15842 25256
rect 15898 25200 23386 25256
rect 23442 25200 23447 25256
rect 15561 25198 23447 25200
rect 0 25168 800 25198
rect 15561 25195 15627 25198
rect 15837 25195 15903 25198
rect 23381 25195 23447 25198
rect 19374 25060 19380 25124
rect 19444 25122 19450 25124
rect 19701 25122 19767 25125
rect 19444 25120 19767 25122
rect 19444 25064 19706 25120
rect 19762 25064 19767 25120
rect 19444 25062 19767 25064
rect 19444 25060 19450 25062
rect 19701 25059 19767 25062
rect 23289 25122 23355 25125
rect 23749 25122 23815 25125
rect 23289 25120 23815 25122
rect 23289 25064 23294 25120
rect 23350 25064 23754 25120
rect 23810 25064 23815 25120
rect 23289 25062 23815 25064
rect 23289 25059 23355 25062
rect 23749 25059 23815 25062
rect 10389 25056 10709 25057
rect 10389 24992 10397 25056
rect 10461 24992 10477 25056
rect 10541 24992 10557 25056
rect 10621 24992 10637 25056
rect 10701 24992 10709 25056
rect 10389 24991 10709 24992
rect 19834 25056 20154 25057
rect 19834 24992 19842 25056
rect 19906 24992 19922 25056
rect 19986 24992 20002 25056
rect 20066 24992 20082 25056
rect 20146 24992 20154 25056
rect 19834 24991 20154 24992
rect 5666 24512 5986 24513
rect 5666 24448 5674 24512
rect 5738 24448 5754 24512
rect 5818 24448 5834 24512
rect 5898 24448 5914 24512
rect 5978 24448 5986 24512
rect 5666 24447 5986 24448
rect 15112 24512 15432 24513
rect 15112 24448 15120 24512
rect 15184 24448 15200 24512
rect 15264 24448 15280 24512
rect 15344 24448 15360 24512
rect 15424 24448 15432 24512
rect 15112 24447 15432 24448
rect 24557 24512 24877 24513
rect 24557 24448 24565 24512
rect 24629 24448 24645 24512
rect 24709 24448 24725 24512
rect 24789 24448 24805 24512
rect 24869 24448 24877 24512
rect 24557 24447 24877 24448
rect 26233 24034 26299 24037
rect 29745 24034 30545 24064
rect 26233 24032 30545 24034
rect 26233 23976 26238 24032
rect 26294 23976 30545 24032
rect 26233 23974 30545 23976
rect 26233 23971 26299 23974
rect 10389 23968 10709 23969
rect 0 23898 800 23928
rect 10389 23904 10397 23968
rect 10461 23904 10477 23968
rect 10541 23904 10557 23968
rect 10621 23904 10637 23968
rect 10701 23904 10709 23968
rect 10389 23903 10709 23904
rect 19834 23968 20154 23969
rect 19834 23904 19842 23968
rect 19906 23904 19922 23968
rect 19986 23904 20002 23968
rect 20066 23904 20082 23968
rect 20146 23904 20154 23968
rect 29745 23944 30545 23974
rect 19834 23903 20154 23904
rect 4061 23898 4127 23901
rect 0 23896 4127 23898
rect 0 23840 4066 23896
rect 4122 23840 4127 23896
rect 0 23838 4127 23840
rect 0 23808 800 23838
rect 4061 23835 4127 23838
rect 5666 23424 5986 23425
rect 5666 23360 5674 23424
rect 5738 23360 5754 23424
rect 5818 23360 5834 23424
rect 5898 23360 5914 23424
rect 5978 23360 5986 23424
rect 5666 23359 5986 23360
rect 15112 23424 15432 23425
rect 15112 23360 15120 23424
rect 15184 23360 15200 23424
rect 15264 23360 15280 23424
rect 15344 23360 15360 23424
rect 15424 23360 15432 23424
rect 15112 23359 15432 23360
rect 24557 23424 24877 23425
rect 24557 23360 24565 23424
rect 24629 23360 24645 23424
rect 24709 23360 24725 23424
rect 24789 23360 24805 23424
rect 24869 23360 24877 23424
rect 24557 23359 24877 23360
rect 18689 23082 18755 23085
rect 2730 23080 18755 23082
rect 2730 23024 18694 23080
rect 18750 23024 18755 23080
rect 2730 23022 18755 23024
rect 0 22538 800 22568
rect 2730 22538 2790 23022
rect 18689 23019 18755 23022
rect 9857 22946 9923 22949
rect 9857 22944 10058 22946
rect 9857 22888 9862 22944
rect 9918 22888 10058 22944
rect 9857 22886 10058 22888
rect 9857 22883 9923 22886
rect 9998 22674 10058 22886
rect 10389 22880 10709 22881
rect 10389 22816 10397 22880
rect 10461 22816 10477 22880
rect 10541 22816 10557 22880
rect 10621 22816 10637 22880
rect 10701 22816 10709 22880
rect 10389 22815 10709 22816
rect 19834 22880 20154 22881
rect 19834 22816 19842 22880
rect 19906 22816 19922 22880
rect 19986 22816 20002 22880
rect 20066 22816 20082 22880
rect 20146 22816 20154 22880
rect 19834 22815 20154 22816
rect 10409 22674 10475 22677
rect 9998 22672 10475 22674
rect 9998 22616 10414 22672
rect 10470 22616 10475 22672
rect 9998 22614 10475 22616
rect 10409 22611 10475 22614
rect 0 22478 2790 22538
rect 0 22448 800 22478
rect 5666 22336 5986 22337
rect 5666 22272 5674 22336
rect 5738 22272 5754 22336
rect 5818 22272 5834 22336
rect 5898 22272 5914 22336
rect 5978 22272 5986 22336
rect 5666 22271 5986 22272
rect 15112 22336 15432 22337
rect 15112 22272 15120 22336
rect 15184 22272 15200 22336
rect 15264 22272 15280 22336
rect 15344 22272 15360 22336
rect 15424 22272 15432 22336
rect 15112 22271 15432 22272
rect 24557 22336 24877 22337
rect 24557 22272 24565 22336
rect 24629 22272 24645 22336
rect 24709 22272 24725 22336
rect 24789 22272 24805 22336
rect 24869 22272 24877 22336
rect 24557 22271 24877 22272
rect 9765 22130 9831 22133
rect 11513 22130 11579 22133
rect 9765 22128 11579 22130
rect 9765 22072 9770 22128
rect 9826 22072 11518 22128
rect 11574 22072 11579 22128
rect 9765 22070 11579 22072
rect 9765 22067 9831 22070
rect 11513 22067 11579 22070
rect 26325 22130 26391 22133
rect 29745 22130 30545 22160
rect 26325 22128 30545 22130
rect 26325 22072 26330 22128
rect 26386 22072 30545 22128
rect 26325 22070 30545 22072
rect 26325 22067 26391 22070
rect 29745 22040 30545 22070
rect 19333 21994 19399 21997
rect 19558 21994 19564 21996
rect 19333 21992 19564 21994
rect 19333 21936 19338 21992
rect 19394 21936 19564 21992
rect 19333 21934 19564 21936
rect 19333 21931 19399 21934
rect 19558 21932 19564 21934
rect 19628 21932 19634 21996
rect 10389 21792 10709 21793
rect 10389 21728 10397 21792
rect 10461 21728 10477 21792
rect 10541 21728 10557 21792
rect 10621 21728 10637 21792
rect 10701 21728 10709 21792
rect 10389 21727 10709 21728
rect 19834 21792 20154 21793
rect 19834 21728 19842 21792
rect 19906 21728 19922 21792
rect 19986 21728 20002 21792
rect 20066 21728 20082 21792
rect 20146 21728 20154 21792
rect 19834 21727 20154 21728
rect 22277 21586 22343 21589
rect 22645 21586 22711 21589
rect 22277 21584 22711 21586
rect 22277 21528 22282 21584
rect 22338 21528 22650 21584
rect 22706 21528 22711 21584
rect 22277 21526 22711 21528
rect 22277 21523 22343 21526
rect 22645 21523 22711 21526
rect 5666 21248 5986 21249
rect 0 21178 800 21208
rect 5666 21184 5674 21248
rect 5738 21184 5754 21248
rect 5818 21184 5834 21248
rect 5898 21184 5914 21248
rect 5978 21184 5986 21248
rect 5666 21183 5986 21184
rect 15112 21248 15432 21249
rect 15112 21184 15120 21248
rect 15184 21184 15200 21248
rect 15264 21184 15280 21248
rect 15344 21184 15360 21248
rect 15424 21184 15432 21248
rect 15112 21183 15432 21184
rect 24557 21248 24877 21249
rect 24557 21184 24565 21248
rect 24629 21184 24645 21248
rect 24709 21184 24725 21248
rect 24789 21184 24805 21248
rect 24869 21184 24877 21248
rect 24557 21183 24877 21184
rect 4061 21178 4127 21181
rect 0 21176 4127 21178
rect 0 21120 4066 21176
rect 4122 21120 4127 21176
rect 0 21118 4127 21120
rect 0 21088 800 21118
rect 4061 21115 4127 21118
rect 11789 21042 11855 21045
rect 15653 21042 15719 21045
rect 11789 21040 15719 21042
rect 11789 20984 11794 21040
rect 11850 20984 15658 21040
rect 15714 20984 15719 21040
rect 11789 20982 15719 20984
rect 11789 20979 11855 20982
rect 15653 20979 15719 20982
rect 10389 20704 10709 20705
rect 10389 20640 10397 20704
rect 10461 20640 10477 20704
rect 10541 20640 10557 20704
rect 10621 20640 10637 20704
rect 10701 20640 10709 20704
rect 10389 20639 10709 20640
rect 19834 20704 20154 20705
rect 19834 20640 19842 20704
rect 19906 20640 19922 20704
rect 19986 20640 20002 20704
rect 20066 20640 20082 20704
rect 20146 20640 20154 20704
rect 19834 20639 20154 20640
rect 12157 20362 12223 20365
rect 14089 20362 14155 20365
rect 12157 20360 14155 20362
rect 12157 20304 12162 20360
rect 12218 20304 14094 20360
rect 14150 20304 14155 20360
rect 12157 20302 14155 20304
rect 12157 20299 12223 20302
rect 14089 20299 14155 20302
rect 27521 20226 27587 20229
rect 29745 20226 30545 20256
rect 27521 20224 30545 20226
rect 27521 20168 27526 20224
rect 27582 20168 30545 20224
rect 27521 20166 30545 20168
rect 27521 20163 27587 20166
rect 5666 20160 5986 20161
rect 5666 20096 5674 20160
rect 5738 20096 5754 20160
rect 5818 20096 5834 20160
rect 5898 20096 5914 20160
rect 5978 20096 5986 20160
rect 5666 20095 5986 20096
rect 15112 20160 15432 20161
rect 15112 20096 15120 20160
rect 15184 20096 15200 20160
rect 15264 20096 15280 20160
rect 15344 20096 15360 20160
rect 15424 20096 15432 20160
rect 15112 20095 15432 20096
rect 24557 20160 24877 20161
rect 24557 20096 24565 20160
rect 24629 20096 24645 20160
rect 24709 20096 24725 20160
rect 24789 20096 24805 20160
rect 24869 20096 24877 20160
rect 29745 20136 30545 20166
rect 24557 20095 24877 20096
rect 0 19818 800 19848
rect 3141 19818 3207 19821
rect 0 19816 3207 19818
rect 0 19760 3146 19816
rect 3202 19760 3207 19816
rect 0 19758 3207 19760
rect 0 19728 800 19758
rect 3141 19755 3207 19758
rect 20253 19684 20319 19685
rect 20253 19680 20300 19684
rect 20364 19682 20370 19684
rect 20253 19624 20258 19680
rect 20253 19620 20300 19624
rect 20364 19622 20410 19682
rect 20364 19620 20370 19622
rect 20253 19619 20319 19620
rect 10389 19616 10709 19617
rect 10389 19552 10397 19616
rect 10461 19552 10477 19616
rect 10541 19552 10557 19616
rect 10621 19552 10637 19616
rect 10701 19552 10709 19616
rect 10389 19551 10709 19552
rect 19834 19616 20154 19617
rect 19834 19552 19842 19616
rect 19906 19552 19922 19616
rect 19986 19552 20002 19616
rect 20066 19552 20082 19616
rect 20146 19552 20154 19616
rect 19834 19551 20154 19552
rect 10961 19410 11027 19413
rect 13813 19410 13879 19413
rect 10961 19408 13879 19410
rect 10961 19352 10966 19408
rect 11022 19352 13818 19408
rect 13874 19352 13879 19408
rect 10961 19350 13879 19352
rect 10961 19347 11027 19350
rect 13813 19347 13879 19350
rect 5666 19072 5986 19073
rect 5666 19008 5674 19072
rect 5738 19008 5754 19072
rect 5818 19008 5834 19072
rect 5898 19008 5914 19072
rect 5978 19008 5986 19072
rect 5666 19007 5986 19008
rect 15112 19072 15432 19073
rect 15112 19008 15120 19072
rect 15184 19008 15200 19072
rect 15264 19008 15280 19072
rect 15344 19008 15360 19072
rect 15424 19008 15432 19072
rect 15112 19007 15432 19008
rect 24557 19072 24877 19073
rect 24557 19008 24565 19072
rect 24629 19008 24645 19072
rect 24709 19008 24725 19072
rect 24789 19008 24805 19072
rect 24869 19008 24877 19072
rect 24557 19007 24877 19008
rect 10389 18528 10709 18529
rect 0 18458 800 18488
rect 10389 18464 10397 18528
rect 10461 18464 10477 18528
rect 10541 18464 10557 18528
rect 10621 18464 10637 18528
rect 10701 18464 10709 18528
rect 10389 18463 10709 18464
rect 19834 18528 20154 18529
rect 19834 18464 19842 18528
rect 19906 18464 19922 18528
rect 19986 18464 20002 18528
rect 20066 18464 20082 18528
rect 20146 18464 20154 18528
rect 19834 18463 20154 18464
rect 3693 18458 3759 18461
rect 0 18456 3759 18458
rect 0 18400 3698 18456
rect 3754 18400 3759 18456
rect 0 18398 3759 18400
rect 0 18368 800 18398
rect 3693 18395 3759 18398
rect 21173 18322 21239 18325
rect 29745 18322 30545 18352
rect 21173 18320 30545 18322
rect 21173 18264 21178 18320
rect 21234 18264 30545 18320
rect 21173 18262 30545 18264
rect 21173 18259 21239 18262
rect 29745 18232 30545 18262
rect 5666 17984 5986 17985
rect 5666 17920 5674 17984
rect 5738 17920 5754 17984
rect 5818 17920 5834 17984
rect 5898 17920 5914 17984
rect 5978 17920 5986 17984
rect 5666 17919 5986 17920
rect 15112 17984 15432 17985
rect 15112 17920 15120 17984
rect 15184 17920 15200 17984
rect 15264 17920 15280 17984
rect 15344 17920 15360 17984
rect 15424 17920 15432 17984
rect 15112 17919 15432 17920
rect 24557 17984 24877 17985
rect 24557 17920 24565 17984
rect 24629 17920 24645 17984
rect 24709 17920 24725 17984
rect 24789 17920 24805 17984
rect 24869 17920 24877 17984
rect 24557 17919 24877 17920
rect 12249 17914 12315 17917
rect 14181 17914 14247 17917
rect 12249 17912 14247 17914
rect 12249 17856 12254 17912
rect 12310 17856 14186 17912
rect 14242 17856 14247 17912
rect 12249 17854 14247 17856
rect 12249 17851 12315 17854
rect 14181 17851 14247 17854
rect 17677 17914 17743 17917
rect 19374 17914 19380 17916
rect 17677 17912 19380 17914
rect 17677 17856 17682 17912
rect 17738 17856 19380 17912
rect 17677 17854 19380 17856
rect 17677 17851 17743 17854
rect 19374 17852 19380 17854
rect 19444 17852 19450 17916
rect 12801 17778 12867 17781
rect 13261 17778 13327 17781
rect 12801 17776 13327 17778
rect 12801 17720 12806 17776
rect 12862 17720 13266 17776
rect 13322 17720 13327 17776
rect 12801 17718 13327 17720
rect 12801 17715 12867 17718
rect 13261 17715 13327 17718
rect 10869 17642 10935 17645
rect 11973 17642 12039 17645
rect 10869 17640 12039 17642
rect 10869 17584 10874 17640
rect 10930 17584 11978 17640
rect 12034 17584 12039 17640
rect 10869 17582 12039 17584
rect 10869 17579 10935 17582
rect 11973 17579 12039 17582
rect 10389 17440 10709 17441
rect 10389 17376 10397 17440
rect 10461 17376 10477 17440
rect 10541 17376 10557 17440
rect 10621 17376 10637 17440
rect 10701 17376 10709 17440
rect 10389 17375 10709 17376
rect 19834 17440 20154 17441
rect 19834 17376 19842 17440
rect 19906 17376 19922 17440
rect 19986 17376 20002 17440
rect 20066 17376 20082 17440
rect 20146 17376 20154 17440
rect 19834 17375 20154 17376
rect 7097 17370 7163 17373
rect 13077 17370 13143 17373
rect 14917 17370 14983 17373
rect 16205 17370 16271 17373
rect 7097 17368 7298 17370
rect 7097 17312 7102 17368
rect 7158 17312 7298 17368
rect 7097 17310 7298 17312
rect 7097 17307 7163 17310
rect 7238 17234 7298 17310
rect 13077 17368 16271 17370
rect 13077 17312 13082 17368
rect 13138 17312 14922 17368
rect 14978 17312 16210 17368
rect 16266 17312 16271 17368
rect 13077 17310 16271 17312
rect 13077 17307 13143 17310
rect 14917 17307 14983 17310
rect 16205 17307 16271 17310
rect 7649 17234 7715 17237
rect 7238 17232 7715 17234
rect 7238 17176 7654 17232
rect 7710 17176 7715 17232
rect 7238 17174 7715 17176
rect 7649 17171 7715 17174
rect 12157 17234 12223 17237
rect 24761 17234 24827 17237
rect 12157 17232 24827 17234
rect 12157 17176 12162 17232
rect 12218 17176 24766 17232
rect 24822 17176 24827 17232
rect 12157 17174 24827 17176
rect 12157 17171 12223 17174
rect 24761 17171 24827 17174
rect 0 17098 800 17128
rect 3509 17098 3575 17101
rect 0 17096 3575 17098
rect 0 17040 3514 17096
rect 3570 17040 3575 17096
rect 0 17038 3575 17040
rect 0 17008 800 17038
rect 3509 17035 3575 17038
rect 3693 17098 3759 17101
rect 22645 17098 22711 17101
rect 3693 17096 22711 17098
rect 3693 17040 3698 17096
rect 3754 17040 22650 17096
rect 22706 17040 22711 17096
rect 3693 17038 22711 17040
rect 3693 17035 3759 17038
rect 22645 17035 22711 17038
rect 5666 16896 5986 16897
rect 5666 16832 5674 16896
rect 5738 16832 5754 16896
rect 5818 16832 5834 16896
rect 5898 16832 5914 16896
rect 5978 16832 5986 16896
rect 5666 16831 5986 16832
rect 15112 16896 15432 16897
rect 15112 16832 15120 16896
rect 15184 16832 15200 16896
rect 15264 16832 15280 16896
rect 15344 16832 15360 16896
rect 15424 16832 15432 16896
rect 15112 16831 15432 16832
rect 24557 16896 24877 16897
rect 24557 16832 24565 16896
rect 24629 16832 24645 16896
rect 24709 16832 24725 16896
rect 24789 16832 24805 16896
rect 24869 16832 24877 16896
rect 24557 16831 24877 16832
rect 10389 16352 10709 16353
rect 10389 16288 10397 16352
rect 10461 16288 10477 16352
rect 10541 16288 10557 16352
rect 10621 16288 10637 16352
rect 10701 16288 10709 16352
rect 10389 16287 10709 16288
rect 19834 16352 20154 16353
rect 19834 16288 19842 16352
rect 19906 16288 19922 16352
rect 19986 16288 20002 16352
rect 20066 16288 20082 16352
rect 20146 16288 20154 16352
rect 19834 16287 20154 16288
rect 21173 16282 21239 16285
rect 29745 16282 30545 16312
rect 21173 16280 30545 16282
rect 21173 16224 21178 16280
rect 21234 16224 30545 16280
rect 21173 16222 30545 16224
rect 21173 16219 21239 16222
rect 29745 16192 30545 16222
rect 5666 15808 5986 15809
rect 0 15738 800 15768
rect 5666 15744 5674 15808
rect 5738 15744 5754 15808
rect 5818 15744 5834 15808
rect 5898 15744 5914 15808
rect 5978 15744 5986 15808
rect 5666 15743 5986 15744
rect 15112 15808 15432 15809
rect 15112 15744 15120 15808
rect 15184 15744 15200 15808
rect 15264 15744 15280 15808
rect 15344 15744 15360 15808
rect 15424 15744 15432 15808
rect 15112 15743 15432 15744
rect 24557 15808 24877 15809
rect 24557 15744 24565 15808
rect 24629 15744 24645 15808
rect 24709 15744 24725 15808
rect 24789 15744 24805 15808
rect 24869 15744 24877 15808
rect 24557 15743 24877 15744
rect 5349 15738 5415 15741
rect 0 15736 5415 15738
rect 0 15680 5354 15736
rect 5410 15680 5415 15736
rect 0 15678 5415 15680
rect 0 15648 800 15678
rect 5349 15675 5415 15678
rect 10389 15264 10709 15265
rect 10389 15200 10397 15264
rect 10461 15200 10477 15264
rect 10541 15200 10557 15264
rect 10621 15200 10637 15264
rect 10701 15200 10709 15264
rect 10389 15199 10709 15200
rect 19834 15264 20154 15265
rect 19834 15200 19842 15264
rect 19906 15200 19922 15264
rect 19986 15200 20002 15264
rect 20066 15200 20082 15264
rect 20146 15200 20154 15264
rect 19834 15199 20154 15200
rect 5666 14720 5986 14721
rect 5666 14656 5674 14720
rect 5738 14656 5754 14720
rect 5818 14656 5834 14720
rect 5898 14656 5914 14720
rect 5978 14656 5986 14720
rect 5666 14655 5986 14656
rect 15112 14720 15432 14721
rect 15112 14656 15120 14720
rect 15184 14656 15200 14720
rect 15264 14656 15280 14720
rect 15344 14656 15360 14720
rect 15424 14656 15432 14720
rect 15112 14655 15432 14656
rect 24557 14720 24877 14721
rect 24557 14656 24565 14720
rect 24629 14656 24645 14720
rect 24709 14656 24725 14720
rect 24789 14656 24805 14720
rect 24869 14656 24877 14720
rect 24557 14655 24877 14656
rect 0 14378 800 14408
rect 4061 14378 4127 14381
rect 0 14376 4127 14378
rect 0 14320 4066 14376
rect 4122 14320 4127 14376
rect 0 14318 4127 14320
rect 0 14288 800 14318
rect 4061 14315 4127 14318
rect 19333 14378 19399 14381
rect 20161 14378 20227 14381
rect 19333 14376 20227 14378
rect 19333 14320 19338 14376
rect 19394 14320 20166 14376
rect 20222 14320 20227 14376
rect 19333 14318 20227 14320
rect 19333 14315 19399 14318
rect 20161 14315 20227 14318
rect 26785 14378 26851 14381
rect 29745 14378 30545 14408
rect 26785 14376 30545 14378
rect 26785 14320 26790 14376
rect 26846 14320 30545 14376
rect 26785 14318 30545 14320
rect 26785 14315 26851 14318
rect 29745 14288 30545 14318
rect 10389 14176 10709 14177
rect 10389 14112 10397 14176
rect 10461 14112 10477 14176
rect 10541 14112 10557 14176
rect 10621 14112 10637 14176
rect 10701 14112 10709 14176
rect 10389 14111 10709 14112
rect 19834 14176 20154 14177
rect 19834 14112 19842 14176
rect 19906 14112 19922 14176
rect 19986 14112 20002 14176
rect 20066 14112 20082 14176
rect 20146 14112 20154 14176
rect 19834 14111 20154 14112
rect 12566 14044 12572 14108
rect 12636 14106 12642 14108
rect 12709 14106 12775 14109
rect 13721 14106 13787 14109
rect 12636 14104 13787 14106
rect 12636 14048 12714 14104
rect 12770 14048 13726 14104
rect 13782 14048 13787 14104
rect 12636 14046 13787 14048
rect 12636 14044 12642 14046
rect 12709 14043 12775 14046
rect 13721 14043 13787 14046
rect 5666 13632 5986 13633
rect 5666 13568 5674 13632
rect 5738 13568 5754 13632
rect 5818 13568 5834 13632
rect 5898 13568 5914 13632
rect 5978 13568 5986 13632
rect 5666 13567 5986 13568
rect 15112 13632 15432 13633
rect 15112 13568 15120 13632
rect 15184 13568 15200 13632
rect 15264 13568 15280 13632
rect 15344 13568 15360 13632
rect 15424 13568 15432 13632
rect 15112 13567 15432 13568
rect 24557 13632 24877 13633
rect 24557 13568 24565 13632
rect 24629 13568 24645 13632
rect 24709 13568 24725 13632
rect 24789 13568 24805 13632
rect 24869 13568 24877 13632
rect 24557 13567 24877 13568
rect 10389 13088 10709 13089
rect 0 13018 800 13048
rect 10389 13024 10397 13088
rect 10461 13024 10477 13088
rect 10541 13024 10557 13088
rect 10621 13024 10637 13088
rect 10701 13024 10709 13088
rect 10389 13023 10709 13024
rect 19834 13088 20154 13089
rect 19834 13024 19842 13088
rect 19906 13024 19922 13088
rect 19986 13024 20002 13088
rect 20066 13024 20082 13088
rect 20146 13024 20154 13088
rect 19834 13023 20154 13024
rect 4061 13018 4127 13021
rect 0 13016 4127 13018
rect 0 12960 4066 13016
rect 4122 12960 4127 13016
rect 0 12958 4127 12960
rect 0 12928 800 12958
rect 4061 12955 4127 12958
rect 5666 12544 5986 12545
rect 5666 12480 5674 12544
rect 5738 12480 5754 12544
rect 5818 12480 5834 12544
rect 5898 12480 5914 12544
rect 5978 12480 5986 12544
rect 5666 12479 5986 12480
rect 15112 12544 15432 12545
rect 15112 12480 15120 12544
rect 15184 12480 15200 12544
rect 15264 12480 15280 12544
rect 15344 12480 15360 12544
rect 15424 12480 15432 12544
rect 15112 12479 15432 12480
rect 24557 12544 24877 12545
rect 24557 12480 24565 12544
rect 24629 12480 24645 12544
rect 24709 12480 24725 12544
rect 24789 12480 24805 12544
rect 24869 12480 24877 12544
rect 24557 12479 24877 12480
rect 26509 12474 26575 12477
rect 29745 12474 30545 12504
rect 26509 12472 30545 12474
rect 26509 12416 26514 12472
rect 26570 12416 30545 12472
rect 26509 12414 30545 12416
rect 26509 12411 26575 12414
rect 29745 12384 30545 12414
rect 15653 12338 15719 12341
rect 18597 12338 18663 12341
rect 15653 12336 18663 12338
rect 15653 12280 15658 12336
rect 15714 12280 18602 12336
rect 18658 12280 18663 12336
rect 15653 12278 18663 12280
rect 15653 12275 15719 12278
rect 18597 12275 18663 12278
rect 12985 12202 13051 12205
rect 21173 12202 21239 12205
rect 12985 12200 21239 12202
rect 12985 12144 12990 12200
rect 13046 12144 21178 12200
rect 21234 12144 21239 12200
rect 12985 12142 21239 12144
rect 12985 12139 13051 12142
rect 21173 12139 21239 12142
rect 10389 12000 10709 12001
rect 10389 11936 10397 12000
rect 10461 11936 10477 12000
rect 10541 11936 10557 12000
rect 10621 11936 10637 12000
rect 10701 11936 10709 12000
rect 10389 11935 10709 11936
rect 19834 12000 20154 12001
rect 19834 11936 19842 12000
rect 19906 11936 19922 12000
rect 19986 11936 20002 12000
rect 20066 11936 20082 12000
rect 20146 11936 20154 12000
rect 19834 11935 20154 11936
rect 0 11658 800 11688
rect 3969 11658 4035 11661
rect 0 11656 4035 11658
rect 0 11600 3974 11656
rect 4030 11600 4035 11656
rect 0 11598 4035 11600
rect 0 11568 800 11598
rect 3969 11595 4035 11598
rect 5666 11456 5986 11457
rect 5666 11392 5674 11456
rect 5738 11392 5754 11456
rect 5818 11392 5834 11456
rect 5898 11392 5914 11456
rect 5978 11392 5986 11456
rect 5666 11391 5986 11392
rect 15112 11456 15432 11457
rect 15112 11392 15120 11456
rect 15184 11392 15200 11456
rect 15264 11392 15280 11456
rect 15344 11392 15360 11456
rect 15424 11392 15432 11456
rect 15112 11391 15432 11392
rect 24557 11456 24877 11457
rect 24557 11392 24565 11456
rect 24629 11392 24645 11456
rect 24709 11392 24725 11456
rect 24789 11392 24805 11456
rect 24869 11392 24877 11456
rect 24557 11391 24877 11392
rect 10389 10912 10709 10913
rect 10389 10848 10397 10912
rect 10461 10848 10477 10912
rect 10541 10848 10557 10912
rect 10621 10848 10637 10912
rect 10701 10848 10709 10912
rect 10389 10847 10709 10848
rect 19834 10912 20154 10913
rect 19834 10848 19842 10912
rect 19906 10848 19922 10912
rect 19986 10848 20002 10912
rect 20066 10848 20082 10912
rect 20146 10848 20154 10912
rect 19834 10847 20154 10848
rect 26233 10570 26299 10573
rect 29745 10570 30545 10600
rect 26233 10568 30545 10570
rect 26233 10512 26238 10568
rect 26294 10512 30545 10568
rect 26233 10510 30545 10512
rect 26233 10507 26299 10510
rect 29745 10480 30545 10510
rect 5666 10368 5986 10369
rect 0 10298 800 10328
rect 5666 10304 5674 10368
rect 5738 10304 5754 10368
rect 5818 10304 5834 10368
rect 5898 10304 5914 10368
rect 5978 10304 5986 10368
rect 5666 10303 5986 10304
rect 15112 10368 15432 10369
rect 15112 10304 15120 10368
rect 15184 10304 15200 10368
rect 15264 10304 15280 10368
rect 15344 10304 15360 10368
rect 15424 10304 15432 10368
rect 15112 10303 15432 10304
rect 24557 10368 24877 10369
rect 24557 10304 24565 10368
rect 24629 10304 24645 10368
rect 24709 10304 24725 10368
rect 24789 10304 24805 10368
rect 24869 10304 24877 10368
rect 24557 10303 24877 10304
rect 4061 10298 4127 10301
rect 0 10296 4127 10298
rect 0 10240 4066 10296
rect 4122 10240 4127 10296
rect 0 10238 4127 10240
rect 0 10208 800 10238
rect 4061 10235 4127 10238
rect 10389 9824 10709 9825
rect 10389 9760 10397 9824
rect 10461 9760 10477 9824
rect 10541 9760 10557 9824
rect 10621 9760 10637 9824
rect 10701 9760 10709 9824
rect 10389 9759 10709 9760
rect 19834 9824 20154 9825
rect 19834 9760 19842 9824
rect 19906 9760 19922 9824
rect 19986 9760 20002 9824
rect 20066 9760 20082 9824
rect 20146 9760 20154 9824
rect 19834 9759 20154 9760
rect 12157 9482 12223 9485
rect 12893 9482 12959 9485
rect 23657 9482 23723 9485
rect 12157 9480 23723 9482
rect 12157 9424 12162 9480
rect 12218 9424 12898 9480
rect 12954 9424 23662 9480
rect 23718 9424 23723 9480
rect 12157 9422 23723 9424
rect 12157 9419 12223 9422
rect 12893 9419 12959 9422
rect 23657 9419 23723 9422
rect 11973 9346 12039 9349
rect 12341 9346 12407 9349
rect 11973 9344 12407 9346
rect 11973 9288 11978 9344
rect 12034 9288 12346 9344
rect 12402 9288 12407 9344
rect 11973 9286 12407 9288
rect 11973 9283 12039 9286
rect 12341 9283 12407 9286
rect 5666 9280 5986 9281
rect 5666 9216 5674 9280
rect 5738 9216 5754 9280
rect 5818 9216 5834 9280
rect 5898 9216 5914 9280
rect 5978 9216 5986 9280
rect 5666 9215 5986 9216
rect 15112 9280 15432 9281
rect 15112 9216 15120 9280
rect 15184 9216 15200 9280
rect 15264 9216 15280 9280
rect 15344 9216 15360 9280
rect 15424 9216 15432 9280
rect 15112 9215 15432 9216
rect 24557 9280 24877 9281
rect 24557 9216 24565 9280
rect 24629 9216 24645 9280
rect 24709 9216 24725 9280
rect 24789 9216 24805 9280
rect 24869 9216 24877 9280
rect 24557 9215 24877 9216
rect 0 8938 800 8968
rect 4061 8938 4127 8941
rect 0 8936 4127 8938
rect 0 8880 4066 8936
rect 4122 8880 4127 8936
rect 0 8878 4127 8880
rect 0 8848 800 8878
rect 4061 8875 4127 8878
rect 10389 8736 10709 8737
rect 10389 8672 10397 8736
rect 10461 8672 10477 8736
rect 10541 8672 10557 8736
rect 10621 8672 10637 8736
rect 10701 8672 10709 8736
rect 10389 8671 10709 8672
rect 19834 8736 20154 8737
rect 19834 8672 19842 8736
rect 19906 8672 19922 8736
rect 19986 8672 20002 8736
rect 20066 8672 20082 8736
rect 20146 8672 20154 8736
rect 19834 8671 20154 8672
rect 20345 8666 20411 8669
rect 21449 8666 21515 8669
rect 20345 8664 21515 8666
rect 20345 8608 20350 8664
rect 20406 8608 21454 8664
rect 21510 8608 21515 8664
rect 20345 8606 21515 8608
rect 20345 8603 20411 8606
rect 21449 8603 21515 8606
rect 26693 8666 26759 8669
rect 29745 8666 30545 8696
rect 26693 8664 30545 8666
rect 26693 8608 26698 8664
rect 26754 8608 30545 8664
rect 26693 8606 30545 8608
rect 26693 8603 26759 8606
rect 29745 8576 30545 8606
rect 19333 8394 19399 8397
rect 21357 8394 21423 8397
rect 24485 8394 24551 8397
rect 19333 8392 24551 8394
rect 19333 8336 19338 8392
rect 19394 8336 21362 8392
rect 21418 8336 24490 8392
rect 24546 8336 24551 8392
rect 19333 8334 24551 8336
rect 19333 8331 19399 8334
rect 21357 8331 21423 8334
rect 24485 8331 24551 8334
rect 5666 8192 5986 8193
rect 5666 8128 5674 8192
rect 5738 8128 5754 8192
rect 5818 8128 5834 8192
rect 5898 8128 5914 8192
rect 5978 8128 5986 8192
rect 5666 8127 5986 8128
rect 15112 8192 15432 8193
rect 15112 8128 15120 8192
rect 15184 8128 15200 8192
rect 15264 8128 15280 8192
rect 15344 8128 15360 8192
rect 15424 8128 15432 8192
rect 15112 8127 15432 8128
rect 24557 8192 24877 8193
rect 24557 8128 24565 8192
rect 24629 8128 24645 8192
rect 24709 8128 24725 8192
rect 24789 8128 24805 8192
rect 24869 8128 24877 8192
rect 24557 8127 24877 8128
rect 14273 7986 14339 7989
rect 17217 7986 17283 7989
rect 14273 7984 17283 7986
rect 14273 7928 14278 7984
rect 14334 7928 17222 7984
rect 17278 7928 17283 7984
rect 14273 7926 17283 7928
rect 14273 7923 14339 7926
rect 17217 7923 17283 7926
rect 10389 7648 10709 7649
rect 0 7578 800 7608
rect 10389 7584 10397 7648
rect 10461 7584 10477 7648
rect 10541 7584 10557 7648
rect 10621 7584 10637 7648
rect 10701 7584 10709 7648
rect 10389 7583 10709 7584
rect 19834 7648 20154 7649
rect 19834 7584 19842 7648
rect 19906 7584 19922 7648
rect 19986 7584 20002 7648
rect 20066 7584 20082 7648
rect 20146 7584 20154 7648
rect 19834 7583 20154 7584
rect 3877 7578 3943 7581
rect 0 7576 3943 7578
rect 0 7520 3882 7576
rect 3938 7520 3943 7576
rect 0 7518 3943 7520
rect 0 7488 800 7518
rect 3877 7515 3943 7518
rect 5666 7104 5986 7105
rect 5666 7040 5674 7104
rect 5738 7040 5754 7104
rect 5818 7040 5834 7104
rect 5898 7040 5914 7104
rect 5978 7040 5986 7104
rect 5666 7039 5986 7040
rect 15112 7104 15432 7105
rect 15112 7040 15120 7104
rect 15184 7040 15200 7104
rect 15264 7040 15280 7104
rect 15344 7040 15360 7104
rect 15424 7040 15432 7104
rect 15112 7039 15432 7040
rect 24557 7104 24877 7105
rect 24557 7040 24565 7104
rect 24629 7040 24645 7104
rect 24709 7040 24725 7104
rect 24789 7040 24805 7104
rect 24869 7040 24877 7104
rect 24557 7039 24877 7040
rect 26233 6762 26299 6765
rect 29745 6762 30545 6792
rect 26233 6760 30545 6762
rect 26233 6704 26238 6760
rect 26294 6704 30545 6760
rect 26233 6702 30545 6704
rect 26233 6699 26299 6702
rect 29745 6672 30545 6702
rect 10389 6560 10709 6561
rect 10389 6496 10397 6560
rect 10461 6496 10477 6560
rect 10541 6496 10557 6560
rect 10621 6496 10637 6560
rect 10701 6496 10709 6560
rect 10389 6495 10709 6496
rect 19834 6560 20154 6561
rect 19834 6496 19842 6560
rect 19906 6496 19922 6560
rect 19986 6496 20002 6560
rect 20066 6496 20082 6560
rect 20146 6496 20154 6560
rect 19834 6495 20154 6496
rect 0 6218 800 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 800 6158
rect 4061 6155 4127 6158
rect 5666 6016 5986 6017
rect 5666 5952 5674 6016
rect 5738 5952 5754 6016
rect 5818 5952 5834 6016
rect 5898 5952 5914 6016
rect 5978 5952 5986 6016
rect 5666 5951 5986 5952
rect 15112 6016 15432 6017
rect 15112 5952 15120 6016
rect 15184 5952 15200 6016
rect 15264 5952 15280 6016
rect 15344 5952 15360 6016
rect 15424 5952 15432 6016
rect 15112 5951 15432 5952
rect 24557 6016 24877 6017
rect 24557 5952 24565 6016
rect 24629 5952 24645 6016
rect 24709 5952 24725 6016
rect 24789 5952 24805 6016
rect 24869 5952 24877 6016
rect 24557 5951 24877 5952
rect 10389 5472 10709 5473
rect 10389 5408 10397 5472
rect 10461 5408 10477 5472
rect 10541 5408 10557 5472
rect 10621 5408 10637 5472
rect 10701 5408 10709 5472
rect 10389 5407 10709 5408
rect 19834 5472 20154 5473
rect 19834 5408 19842 5472
rect 19906 5408 19922 5472
rect 19986 5408 20002 5472
rect 20066 5408 20082 5472
rect 20146 5408 20154 5472
rect 19834 5407 20154 5408
rect 5666 4928 5986 4929
rect 0 4858 800 4888
rect 5666 4864 5674 4928
rect 5738 4864 5754 4928
rect 5818 4864 5834 4928
rect 5898 4864 5914 4928
rect 5978 4864 5986 4928
rect 5666 4863 5986 4864
rect 15112 4928 15432 4929
rect 15112 4864 15120 4928
rect 15184 4864 15200 4928
rect 15264 4864 15280 4928
rect 15344 4864 15360 4928
rect 15424 4864 15432 4928
rect 15112 4863 15432 4864
rect 24557 4928 24877 4929
rect 24557 4864 24565 4928
rect 24629 4864 24645 4928
rect 24709 4864 24725 4928
rect 24789 4864 24805 4928
rect 24869 4864 24877 4928
rect 24557 4863 24877 4864
rect 3969 4858 4035 4861
rect 0 4856 4035 4858
rect 0 4800 3974 4856
rect 4030 4800 4035 4856
rect 0 4798 4035 4800
rect 0 4768 800 4798
rect 3969 4795 4035 4798
rect 26233 4858 26299 4861
rect 29745 4858 30545 4888
rect 26233 4856 30545 4858
rect 26233 4800 26238 4856
rect 26294 4800 30545 4856
rect 26233 4798 30545 4800
rect 26233 4795 26299 4798
rect 29745 4768 30545 4798
rect 10389 4384 10709 4385
rect 10389 4320 10397 4384
rect 10461 4320 10477 4384
rect 10541 4320 10557 4384
rect 10621 4320 10637 4384
rect 10701 4320 10709 4384
rect 10389 4319 10709 4320
rect 19834 4384 20154 4385
rect 19834 4320 19842 4384
rect 19906 4320 19922 4384
rect 19986 4320 20002 4384
rect 20066 4320 20082 4384
rect 20146 4320 20154 4384
rect 19834 4319 20154 4320
rect 5666 3840 5986 3841
rect 5666 3776 5674 3840
rect 5738 3776 5754 3840
rect 5818 3776 5834 3840
rect 5898 3776 5914 3840
rect 5978 3776 5986 3840
rect 5666 3775 5986 3776
rect 15112 3840 15432 3841
rect 15112 3776 15120 3840
rect 15184 3776 15200 3840
rect 15264 3776 15280 3840
rect 15344 3776 15360 3840
rect 15424 3776 15432 3840
rect 15112 3775 15432 3776
rect 24557 3840 24877 3841
rect 24557 3776 24565 3840
rect 24629 3776 24645 3840
rect 24709 3776 24725 3840
rect 24789 3776 24805 3840
rect 24869 3776 24877 3840
rect 24557 3775 24877 3776
rect 0 3498 800 3528
rect 1393 3498 1459 3501
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3408 800 3438
rect 1393 3435 1459 3438
rect 19558 3436 19564 3500
rect 19628 3498 19634 3500
rect 25957 3498 26023 3501
rect 19628 3496 26023 3498
rect 19628 3440 25962 3496
rect 26018 3440 26023 3496
rect 19628 3438 26023 3440
rect 19628 3436 19634 3438
rect 25957 3435 26023 3438
rect 10389 3296 10709 3297
rect 10389 3232 10397 3296
rect 10461 3232 10477 3296
rect 10541 3232 10557 3296
rect 10621 3232 10637 3296
rect 10701 3232 10709 3296
rect 10389 3231 10709 3232
rect 19834 3296 20154 3297
rect 19834 3232 19842 3296
rect 19906 3232 19922 3296
rect 19986 3232 20002 3296
rect 20066 3232 20082 3296
rect 20146 3232 20154 3296
rect 19834 3231 20154 3232
rect 20294 3028 20300 3092
rect 20364 3090 20370 3092
rect 23933 3090 23999 3093
rect 20364 3088 23999 3090
rect 20364 3032 23938 3088
rect 23994 3032 23999 3088
rect 20364 3030 23999 3032
rect 20364 3028 20370 3030
rect 23933 3027 23999 3030
rect 26325 2954 26391 2957
rect 29745 2954 30545 2984
rect 26325 2952 30545 2954
rect 26325 2896 26330 2952
rect 26386 2896 30545 2952
rect 26325 2894 30545 2896
rect 26325 2891 26391 2894
rect 29745 2864 30545 2894
rect 5666 2752 5986 2753
rect 5666 2688 5674 2752
rect 5738 2688 5754 2752
rect 5818 2688 5834 2752
rect 5898 2688 5914 2752
rect 5978 2688 5986 2752
rect 5666 2687 5986 2688
rect 15112 2752 15432 2753
rect 15112 2688 15120 2752
rect 15184 2688 15200 2752
rect 15264 2688 15280 2752
rect 15344 2688 15360 2752
rect 15424 2688 15432 2752
rect 15112 2687 15432 2688
rect 24557 2752 24877 2753
rect 24557 2688 24565 2752
rect 24629 2688 24645 2752
rect 24709 2688 24725 2752
rect 24789 2688 24805 2752
rect 24869 2688 24877 2752
rect 24557 2687 24877 2688
rect 10389 2208 10709 2209
rect 0 2138 800 2168
rect 10389 2144 10397 2208
rect 10461 2144 10477 2208
rect 10541 2144 10557 2208
rect 10621 2144 10637 2208
rect 10701 2144 10709 2208
rect 10389 2143 10709 2144
rect 19834 2208 20154 2209
rect 19834 2144 19842 2208
rect 19906 2144 19922 2208
rect 19986 2144 20002 2208
rect 20066 2144 20082 2208
rect 20146 2144 20154 2208
rect 19834 2143 20154 2144
rect 3049 2138 3115 2141
rect 0 2136 3115 2138
rect 0 2080 3054 2136
rect 3110 2080 3115 2136
rect 0 2078 3115 2080
rect 0 2048 800 2078
rect 3049 2075 3115 2078
rect 26233 1050 26299 1053
rect 29745 1050 30545 1080
rect 26233 1048 30545 1050
rect 26233 992 26238 1048
rect 26294 992 30545 1048
rect 26233 990 30545 992
rect 26233 987 26299 990
rect 29745 960 30545 990
rect 0 778 800 808
rect 3325 778 3391 781
rect 0 776 3391 778
rect 0 720 3330 776
rect 3386 720 3391 776
rect 0 718 3391 720
rect 0 688 800 718
rect 3325 715 3391 718
<< via3 >>
rect 10397 30492 10461 30496
rect 10397 30436 10401 30492
rect 10401 30436 10457 30492
rect 10457 30436 10461 30492
rect 10397 30432 10461 30436
rect 10477 30492 10541 30496
rect 10477 30436 10481 30492
rect 10481 30436 10537 30492
rect 10537 30436 10541 30492
rect 10477 30432 10541 30436
rect 10557 30492 10621 30496
rect 10557 30436 10561 30492
rect 10561 30436 10617 30492
rect 10617 30436 10621 30492
rect 10557 30432 10621 30436
rect 10637 30492 10701 30496
rect 10637 30436 10641 30492
rect 10641 30436 10697 30492
rect 10697 30436 10701 30492
rect 10637 30432 10701 30436
rect 19842 30492 19906 30496
rect 19842 30436 19846 30492
rect 19846 30436 19902 30492
rect 19902 30436 19906 30492
rect 19842 30432 19906 30436
rect 19922 30492 19986 30496
rect 19922 30436 19926 30492
rect 19926 30436 19982 30492
rect 19982 30436 19986 30492
rect 19922 30432 19986 30436
rect 20002 30492 20066 30496
rect 20002 30436 20006 30492
rect 20006 30436 20062 30492
rect 20062 30436 20066 30492
rect 20002 30432 20066 30436
rect 20082 30492 20146 30496
rect 20082 30436 20086 30492
rect 20086 30436 20142 30492
rect 20142 30436 20146 30492
rect 20082 30432 20146 30436
rect 5674 29948 5738 29952
rect 5674 29892 5678 29948
rect 5678 29892 5734 29948
rect 5734 29892 5738 29948
rect 5674 29888 5738 29892
rect 5754 29948 5818 29952
rect 5754 29892 5758 29948
rect 5758 29892 5814 29948
rect 5814 29892 5818 29948
rect 5754 29888 5818 29892
rect 5834 29948 5898 29952
rect 5834 29892 5838 29948
rect 5838 29892 5894 29948
rect 5894 29892 5898 29948
rect 5834 29888 5898 29892
rect 5914 29948 5978 29952
rect 5914 29892 5918 29948
rect 5918 29892 5974 29948
rect 5974 29892 5978 29948
rect 5914 29888 5978 29892
rect 15120 29948 15184 29952
rect 15120 29892 15124 29948
rect 15124 29892 15180 29948
rect 15180 29892 15184 29948
rect 15120 29888 15184 29892
rect 15200 29948 15264 29952
rect 15200 29892 15204 29948
rect 15204 29892 15260 29948
rect 15260 29892 15264 29948
rect 15200 29888 15264 29892
rect 15280 29948 15344 29952
rect 15280 29892 15284 29948
rect 15284 29892 15340 29948
rect 15340 29892 15344 29948
rect 15280 29888 15344 29892
rect 15360 29948 15424 29952
rect 15360 29892 15364 29948
rect 15364 29892 15420 29948
rect 15420 29892 15424 29948
rect 15360 29888 15424 29892
rect 24565 29948 24629 29952
rect 24565 29892 24569 29948
rect 24569 29892 24625 29948
rect 24625 29892 24629 29948
rect 24565 29888 24629 29892
rect 24645 29948 24709 29952
rect 24645 29892 24649 29948
rect 24649 29892 24705 29948
rect 24705 29892 24709 29948
rect 24645 29888 24709 29892
rect 24725 29948 24789 29952
rect 24725 29892 24729 29948
rect 24729 29892 24785 29948
rect 24785 29892 24789 29948
rect 24725 29888 24789 29892
rect 24805 29948 24869 29952
rect 24805 29892 24809 29948
rect 24809 29892 24865 29948
rect 24865 29892 24869 29948
rect 24805 29888 24869 29892
rect 10397 29404 10461 29408
rect 10397 29348 10401 29404
rect 10401 29348 10457 29404
rect 10457 29348 10461 29404
rect 10397 29344 10461 29348
rect 10477 29404 10541 29408
rect 10477 29348 10481 29404
rect 10481 29348 10537 29404
rect 10537 29348 10541 29404
rect 10477 29344 10541 29348
rect 10557 29404 10621 29408
rect 10557 29348 10561 29404
rect 10561 29348 10617 29404
rect 10617 29348 10621 29404
rect 10557 29344 10621 29348
rect 10637 29404 10701 29408
rect 10637 29348 10641 29404
rect 10641 29348 10697 29404
rect 10697 29348 10701 29404
rect 10637 29344 10701 29348
rect 19842 29404 19906 29408
rect 19842 29348 19846 29404
rect 19846 29348 19902 29404
rect 19902 29348 19906 29404
rect 19842 29344 19906 29348
rect 19922 29404 19986 29408
rect 19922 29348 19926 29404
rect 19926 29348 19982 29404
rect 19982 29348 19986 29404
rect 19922 29344 19986 29348
rect 20002 29404 20066 29408
rect 20002 29348 20006 29404
rect 20006 29348 20062 29404
rect 20062 29348 20066 29404
rect 20002 29344 20066 29348
rect 20082 29404 20146 29408
rect 20082 29348 20086 29404
rect 20086 29348 20142 29404
rect 20142 29348 20146 29404
rect 20082 29344 20146 29348
rect 5674 28860 5738 28864
rect 5674 28804 5678 28860
rect 5678 28804 5734 28860
rect 5734 28804 5738 28860
rect 5674 28800 5738 28804
rect 5754 28860 5818 28864
rect 5754 28804 5758 28860
rect 5758 28804 5814 28860
rect 5814 28804 5818 28860
rect 5754 28800 5818 28804
rect 5834 28860 5898 28864
rect 5834 28804 5838 28860
rect 5838 28804 5894 28860
rect 5894 28804 5898 28860
rect 5834 28800 5898 28804
rect 5914 28860 5978 28864
rect 5914 28804 5918 28860
rect 5918 28804 5974 28860
rect 5974 28804 5978 28860
rect 5914 28800 5978 28804
rect 15120 28860 15184 28864
rect 15120 28804 15124 28860
rect 15124 28804 15180 28860
rect 15180 28804 15184 28860
rect 15120 28800 15184 28804
rect 15200 28860 15264 28864
rect 15200 28804 15204 28860
rect 15204 28804 15260 28860
rect 15260 28804 15264 28860
rect 15200 28800 15264 28804
rect 15280 28860 15344 28864
rect 15280 28804 15284 28860
rect 15284 28804 15340 28860
rect 15340 28804 15344 28860
rect 15280 28800 15344 28804
rect 15360 28860 15424 28864
rect 15360 28804 15364 28860
rect 15364 28804 15420 28860
rect 15420 28804 15424 28860
rect 15360 28800 15424 28804
rect 24565 28860 24629 28864
rect 24565 28804 24569 28860
rect 24569 28804 24625 28860
rect 24625 28804 24629 28860
rect 24565 28800 24629 28804
rect 24645 28860 24709 28864
rect 24645 28804 24649 28860
rect 24649 28804 24705 28860
rect 24705 28804 24709 28860
rect 24645 28800 24709 28804
rect 24725 28860 24789 28864
rect 24725 28804 24729 28860
rect 24729 28804 24785 28860
rect 24785 28804 24789 28860
rect 24725 28800 24789 28804
rect 24805 28860 24869 28864
rect 24805 28804 24809 28860
rect 24809 28804 24865 28860
rect 24865 28804 24869 28860
rect 24805 28800 24869 28804
rect 10397 28316 10461 28320
rect 10397 28260 10401 28316
rect 10401 28260 10457 28316
rect 10457 28260 10461 28316
rect 10397 28256 10461 28260
rect 10477 28316 10541 28320
rect 10477 28260 10481 28316
rect 10481 28260 10537 28316
rect 10537 28260 10541 28316
rect 10477 28256 10541 28260
rect 10557 28316 10621 28320
rect 10557 28260 10561 28316
rect 10561 28260 10617 28316
rect 10617 28260 10621 28316
rect 10557 28256 10621 28260
rect 10637 28316 10701 28320
rect 10637 28260 10641 28316
rect 10641 28260 10697 28316
rect 10697 28260 10701 28316
rect 10637 28256 10701 28260
rect 19842 28316 19906 28320
rect 19842 28260 19846 28316
rect 19846 28260 19902 28316
rect 19902 28260 19906 28316
rect 19842 28256 19906 28260
rect 19922 28316 19986 28320
rect 19922 28260 19926 28316
rect 19926 28260 19982 28316
rect 19982 28260 19986 28316
rect 19922 28256 19986 28260
rect 20002 28316 20066 28320
rect 20002 28260 20006 28316
rect 20006 28260 20062 28316
rect 20062 28260 20066 28316
rect 20002 28256 20066 28260
rect 20082 28316 20146 28320
rect 20082 28260 20086 28316
rect 20086 28260 20142 28316
rect 20142 28260 20146 28316
rect 20082 28256 20146 28260
rect 5674 27772 5738 27776
rect 5674 27716 5678 27772
rect 5678 27716 5734 27772
rect 5734 27716 5738 27772
rect 5674 27712 5738 27716
rect 5754 27772 5818 27776
rect 5754 27716 5758 27772
rect 5758 27716 5814 27772
rect 5814 27716 5818 27772
rect 5754 27712 5818 27716
rect 5834 27772 5898 27776
rect 5834 27716 5838 27772
rect 5838 27716 5894 27772
rect 5894 27716 5898 27772
rect 5834 27712 5898 27716
rect 5914 27772 5978 27776
rect 5914 27716 5918 27772
rect 5918 27716 5974 27772
rect 5974 27716 5978 27772
rect 5914 27712 5978 27716
rect 15120 27772 15184 27776
rect 15120 27716 15124 27772
rect 15124 27716 15180 27772
rect 15180 27716 15184 27772
rect 15120 27712 15184 27716
rect 15200 27772 15264 27776
rect 15200 27716 15204 27772
rect 15204 27716 15260 27772
rect 15260 27716 15264 27772
rect 15200 27712 15264 27716
rect 15280 27772 15344 27776
rect 15280 27716 15284 27772
rect 15284 27716 15340 27772
rect 15340 27716 15344 27772
rect 15280 27712 15344 27716
rect 15360 27772 15424 27776
rect 15360 27716 15364 27772
rect 15364 27716 15420 27772
rect 15420 27716 15424 27772
rect 15360 27712 15424 27716
rect 24565 27772 24629 27776
rect 24565 27716 24569 27772
rect 24569 27716 24625 27772
rect 24625 27716 24629 27772
rect 24565 27712 24629 27716
rect 24645 27772 24709 27776
rect 24645 27716 24649 27772
rect 24649 27716 24705 27772
rect 24705 27716 24709 27772
rect 24645 27712 24709 27716
rect 24725 27772 24789 27776
rect 24725 27716 24729 27772
rect 24729 27716 24785 27772
rect 24785 27716 24789 27772
rect 24725 27712 24789 27716
rect 24805 27772 24869 27776
rect 24805 27716 24809 27772
rect 24809 27716 24865 27772
rect 24865 27716 24869 27772
rect 24805 27712 24869 27716
rect 10397 27228 10461 27232
rect 10397 27172 10401 27228
rect 10401 27172 10457 27228
rect 10457 27172 10461 27228
rect 10397 27168 10461 27172
rect 10477 27228 10541 27232
rect 10477 27172 10481 27228
rect 10481 27172 10537 27228
rect 10537 27172 10541 27228
rect 10477 27168 10541 27172
rect 10557 27228 10621 27232
rect 10557 27172 10561 27228
rect 10561 27172 10617 27228
rect 10617 27172 10621 27228
rect 10557 27168 10621 27172
rect 10637 27228 10701 27232
rect 10637 27172 10641 27228
rect 10641 27172 10697 27228
rect 10697 27172 10701 27228
rect 10637 27168 10701 27172
rect 19842 27228 19906 27232
rect 19842 27172 19846 27228
rect 19846 27172 19902 27228
rect 19902 27172 19906 27228
rect 19842 27168 19906 27172
rect 19922 27228 19986 27232
rect 19922 27172 19926 27228
rect 19926 27172 19982 27228
rect 19982 27172 19986 27228
rect 19922 27168 19986 27172
rect 20002 27228 20066 27232
rect 20002 27172 20006 27228
rect 20006 27172 20062 27228
rect 20062 27172 20066 27228
rect 20002 27168 20066 27172
rect 20082 27228 20146 27232
rect 20082 27172 20086 27228
rect 20086 27172 20142 27228
rect 20142 27172 20146 27228
rect 20082 27168 20146 27172
rect 5674 26684 5738 26688
rect 5674 26628 5678 26684
rect 5678 26628 5734 26684
rect 5734 26628 5738 26684
rect 5674 26624 5738 26628
rect 5754 26684 5818 26688
rect 5754 26628 5758 26684
rect 5758 26628 5814 26684
rect 5814 26628 5818 26684
rect 5754 26624 5818 26628
rect 5834 26684 5898 26688
rect 5834 26628 5838 26684
rect 5838 26628 5894 26684
rect 5894 26628 5898 26684
rect 5834 26624 5898 26628
rect 5914 26684 5978 26688
rect 5914 26628 5918 26684
rect 5918 26628 5974 26684
rect 5974 26628 5978 26684
rect 5914 26624 5978 26628
rect 15120 26684 15184 26688
rect 15120 26628 15124 26684
rect 15124 26628 15180 26684
rect 15180 26628 15184 26684
rect 15120 26624 15184 26628
rect 15200 26684 15264 26688
rect 15200 26628 15204 26684
rect 15204 26628 15260 26684
rect 15260 26628 15264 26684
rect 15200 26624 15264 26628
rect 15280 26684 15344 26688
rect 15280 26628 15284 26684
rect 15284 26628 15340 26684
rect 15340 26628 15344 26684
rect 15280 26624 15344 26628
rect 15360 26684 15424 26688
rect 15360 26628 15364 26684
rect 15364 26628 15420 26684
rect 15420 26628 15424 26684
rect 15360 26624 15424 26628
rect 24565 26684 24629 26688
rect 24565 26628 24569 26684
rect 24569 26628 24625 26684
rect 24625 26628 24629 26684
rect 24565 26624 24629 26628
rect 24645 26684 24709 26688
rect 24645 26628 24649 26684
rect 24649 26628 24705 26684
rect 24705 26628 24709 26684
rect 24645 26624 24709 26628
rect 24725 26684 24789 26688
rect 24725 26628 24729 26684
rect 24729 26628 24785 26684
rect 24785 26628 24789 26684
rect 24725 26624 24789 26628
rect 24805 26684 24869 26688
rect 24805 26628 24809 26684
rect 24809 26628 24865 26684
rect 24865 26628 24869 26684
rect 24805 26624 24869 26628
rect 10397 26140 10461 26144
rect 10397 26084 10401 26140
rect 10401 26084 10457 26140
rect 10457 26084 10461 26140
rect 10397 26080 10461 26084
rect 10477 26140 10541 26144
rect 10477 26084 10481 26140
rect 10481 26084 10537 26140
rect 10537 26084 10541 26140
rect 10477 26080 10541 26084
rect 10557 26140 10621 26144
rect 10557 26084 10561 26140
rect 10561 26084 10617 26140
rect 10617 26084 10621 26140
rect 10557 26080 10621 26084
rect 10637 26140 10701 26144
rect 10637 26084 10641 26140
rect 10641 26084 10697 26140
rect 10697 26084 10701 26140
rect 10637 26080 10701 26084
rect 19842 26140 19906 26144
rect 19842 26084 19846 26140
rect 19846 26084 19902 26140
rect 19902 26084 19906 26140
rect 19842 26080 19906 26084
rect 19922 26140 19986 26144
rect 19922 26084 19926 26140
rect 19926 26084 19982 26140
rect 19982 26084 19986 26140
rect 19922 26080 19986 26084
rect 20002 26140 20066 26144
rect 20002 26084 20006 26140
rect 20006 26084 20062 26140
rect 20062 26084 20066 26140
rect 20002 26080 20066 26084
rect 20082 26140 20146 26144
rect 20082 26084 20086 26140
rect 20086 26084 20142 26140
rect 20142 26084 20146 26140
rect 20082 26080 20146 26084
rect 12572 25664 12636 25668
rect 12572 25608 12586 25664
rect 12586 25608 12636 25664
rect 12572 25604 12636 25608
rect 5674 25596 5738 25600
rect 5674 25540 5678 25596
rect 5678 25540 5734 25596
rect 5734 25540 5738 25596
rect 5674 25536 5738 25540
rect 5754 25596 5818 25600
rect 5754 25540 5758 25596
rect 5758 25540 5814 25596
rect 5814 25540 5818 25596
rect 5754 25536 5818 25540
rect 5834 25596 5898 25600
rect 5834 25540 5838 25596
rect 5838 25540 5894 25596
rect 5894 25540 5898 25596
rect 5834 25536 5898 25540
rect 5914 25596 5978 25600
rect 5914 25540 5918 25596
rect 5918 25540 5974 25596
rect 5974 25540 5978 25596
rect 5914 25536 5978 25540
rect 15120 25596 15184 25600
rect 15120 25540 15124 25596
rect 15124 25540 15180 25596
rect 15180 25540 15184 25596
rect 15120 25536 15184 25540
rect 15200 25596 15264 25600
rect 15200 25540 15204 25596
rect 15204 25540 15260 25596
rect 15260 25540 15264 25596
rect 15200 25536 15264 25540
rect 15280 25596 15344 25600
rect 15280 25540 15284 25596
rect 15284 25540 15340 25596
rect 15340 25540 15344 25596
rect 15280 25536 15344 25540
rect 15360 25596 15424 25600
rect 15360 25540 15364 25596
rect 15364 25540 15420 25596
rect 15420 25540 15424 25596
rect 15360 25536 15424 25540
rect 24565 25596 24629 25600
rect 24565 25540 24569 25596
rect 24569 25540 24625 25596
rect 24625 25540 24629 25596
rect 24565 25536 24629 25540
rect 24645 25596 24709 25600
rect 24645 25540 24649 25596
rect 24649 25540 24705 25596
rect 24705 25540 24709 25596
rect 24645 25536 24709 25540
rect 24725 25596 24789 25600
rect 24725 25540 24729 25596
rect 24729 25540 24785 25596
rect 24785 25540 24789 25596
rect 24725 25536 24789 25540
rect 24805 25596 24869 25600
rect 24805 25540 24809 25596
rect 24809 25540 24865 25596
rect 24865 25540 24869 25596
rect 24805 25536 24869 25540
rect 19380 25060 19444 25124
rect 10397 25052 10461 25056
rect 10397 24996 10401 25052
rect 10401 24996 10457 25052
rect 10457 24996 10461 25052
rect 10397 24992 10461 24996
rect 10477 25052 10541 25056
rect 10477 24996 10481 25052
rect 10481 24996 10537 25052
rect 10537 24996 10541 25052
rect 10477 24992 10541 24996
rect 10557 25052 10621 25056
rect 10557 24996 10561 25052
rect 10561 24996 10617 25052
rect 10617 24996 10621 25052
rect 10557 24992 10621 24996
rect 10637 25052 10701 25056
rect 10637 24996 10641 25052
rect 10641 24996 10697 25052
rect 10697 24996 10701 25052
rect 10637 24992 10701 24996
rect 19842 25052 19906 25056
rect 19842 24996 19846 25052
rect 19846 24996 19902 25052
rect 19902 24996 19906 25052
rect 19842 24992 19906 24996
rect 19922 25052 19986 25056
rect 19922 24996 19926 25052
rect 19926 24996 19982 25052
rect 19982 24996 19986 25052
rect 19922 24992 19986 24996
rect 20002 25052 20066 25056
rect 20002 24996 20006 25052
rect 20006 24996 20062 25052
rect 20062 24996 20066 25052
rect 20002 24992 20066 24996
rect 20082 25052 20146 25056
rect 20082 24996 20086 25052
rect 20086 24996 20142 25052
rect 20142 24996 20146 25052
rect 20082 24992 20146 24996
rect 5674 24508 5738 24512
rect 5674 24452 5678 24508
rect 5678 24452 5734 24508
rect 5734 24452 5738 24508
rect 5674 24448 5738 24452
rect 5754 24508 5818 24512
rect 5754 24452 5758 24508
rect 5758 24452 5814 24508
rect 5814 24452 5818 24508
rect 5754 24448 5818 24452
rect 5834 24508 5898 24512
rect 5834 24452 5838 24508
rect 5838 24452 5894 24508
rect 5894 24452 5898 24508
rect 5834 24448 5898 24452
rect 5914 24508 5978 24512
rect 5914 24452 5918 24508
rect 5918 24452 5974 24508
rect 5974 24452 5978 24508
rect 5914 24448 5978 24452
rect 15120 24508 15184 24512
rect 15120 24452 15124 24508
rect 15124 24452 15180 24508
rect 15180 24452 15184 24508
rect 15120 24448 15184 24452
rect 15200 24508 15264 24512
rect 15200 24452 15204 24508
rect 15204 24452 15260 24508
rect 15260 24452 15264 24508
rect 15200 24448 15264 24452
rect 15280 24508 15344 24512
rect 15280 24452 15284 24508
rect 15284 24452 15340 24508
rect 15340 24452 15344 24508
rect 15280 24448 15344 24452
rect 15360 24508 15424 24512
rect 15360 24452 15364 24508
rect 15364 24452 15420 24508
rect 15420 24452 15424 24508
rect 15360 24448 15424 24452
rect 24565 24508 24629 24512
rect 24565 24452 24569 24508
rect 24569 24452 24625 24508
rect 24625 24452 24629 24508
rect 24565 24448 24629 24452
rect 24645 24508 24709 24512
rect 24645 24452 24649 24508
rect 24649 24452 24705 24508
rect 24705 24452 24709 24508
rect 24645 24448 24709 24452
rect 24725 24508 24789 24512
rect 24725 24452 24729 24508
rect 24729 24452 24785 24508
rect 24785 24452 24789 24508
rect 24725 24448 24789 24452
rect 24805 24508 24869 24512
rect 24805 24452 24809 24508
rect 24809 24452 24865 24508
rect 24865 24452 24869 24508
rect 24805 24448 24869 24452
rect 10397 23964 10461 23968
rect 10397 23908 10401 23964
rect 10401 23908 10457 23964
rect 10457 23908 10461 23964
rect 10397 23904 10461 23908
rect 10477 23964 10541 23968
rect 10477 23908 10481 23964
rect 10481 23908 10537 23964
rect 10537 23908 10541 23964
rect 10477 23904 10541 23908
rect 10557 23964 10621 23968
rect 10557 23908 10561 23964
rect 10561 23908 10617 23964
rect 10617 23908 10621 23964
rect 10557 23904 10621 23908
rect 10637 23964 10701 23968
rect 10637 23908 10641 23964
rect 10641 23908 10697 23964
rect 10697 23908 10701 23964
rect 10637 23904 10701 23908
rect 19842 23964 19906 23968
rect 19842 23908 19846 23964
rect 19846 23908 19902 23964
rect 19902 23908 19906 23964
rect 19842 23904 19906 23908
rect 19922 23964 19986 23968
rect 19922 23908 19926 23964
rect 19926 23908 19982 23964
rect 19982 23908 19986 23964
rect 19922 23904 19986 23908
rect 20002 23964 20066 23968
rect 20002 23908 20006 23964
rect 20006 23908 20062 23964
rect 20062 23908 20066 23964
rect 20002 23904 20066 23908
rect 20082 23964 20146 23968
rect 20082 23908 20086 23964
rect 20086 23908 20142 23964
rect 20142 23908 20146 23964
rect 20082 23904 20146 23908
rect 5674 23420 5738 23424
rect 5674 23364 5678 23420
rect 5678 23364 5734 23420
rect 5734 23364 5738 23420
rect 5674 23360 5738 23364
rect 5754 23420 5818 23424
rect 5754 23364 5758 23420
rect 5758 23364 5814 23420
rect 5814 23364 5818 23420
rect 5754 23360 5818 23364
rect 5834 23420 5898 23424
rect 5834 23364 5838 23420
rect 5838 23364 5894 23420
rect 5894 23364 5898 23420
rect 5834 23360 5898 23364
rect 5914 23420 5978 23424
rect 5914 23364 5918 23420
rect 5918 23364 5974 23420
rect 5974 23364 5978 23420
rect 5914 23360 5978 23364
rect 15120 23420 15184 23424
rect 15120 23364 15124 23420
rect 15124 23364 15180 23420
rect 15180 23364 15184 23420
rect 15120 23360 15184 23364
rect 15200 23420 15264 23424
rect 15200 23364 15204 23420
rect 15204 23364 15260 23420
rect 15260 23364 15264 23420
rect 15200 23360 15264 23364
rect 15280 23420 15344 23424
rect 15280 23364 15284 23420
rect 15284 23364 15340 23420
rect 15340 23364 15344 23420
rect 15280 23360 15344 23364
rect 15360 23420 15424 23424
rect 15360 23364 15364 23420
rect 15364 23364 15420 23420
rect 15420 23364 15424 23420
rect 15360 23360 15424 23364
rect 24565 23420 24629 23424
rect 24565 23364 24569 23420
rect 24569 23364 24625 23420
rect 24625 23364 24629 23420
rect 24565 23360 24629 23364
rect 24645 23420 24709 23424
rect 24645 23364 24649 23420
rect 24649 23364 24705 23420
rect 24705 23364 24709 23420
rect 24645 23360 24709 23364
rect 24725 23420 24789 23424
rect 24725 23364 24729 23420
rect 24729 23364 24785 23420
rect 24785 23364 24789 23420
rect 24725 23360 24789 23364
rect 24805 23420 24869 23424
rect 24805 23364 24809 23420
rect 24809 23364 24865 23420
rect 24865 23364 24869 23420
rect 24805 23360 24869 23364
rect 10397 22876 10461 22880
rect 10397 22820 10401 22876
rect 10401 22820 10457 22876
rect 10457 22820 10461 22876
rect 10397 22816 10461 22820
rect 10477 22876 10541 22880
rect 10477 22820 10481 22876
rect 10481 22820 10537 22876
rect 10537 22820 10541 22876
rect 10477 22816 10541 22820
rect 10557 22876 10621 22880
rect 10557 22820 10561 22876
rect 10561 22820 10617 22876
rect 10617 22820 10621 22876
rect 10557 22816 10621 22820
rect 10637 22876 10701 22880
rect 10637 22820 10641 22876
rect 10641 22820 10697 22876
rect 10697 22820 10701 22876
rect 10637 22816 10701 22820
rect 19842 22876 19906 22880
rect 19842 22820 19846 22876
rect 19846 22820 19902 22876
rect 19902 22820 19906 22876
rect 19842 22816 19906 22820
rect 19922 22876 19986 22880
rect 19922 22820 19926 22876
rect 19926 22820 19982 22876
rect 19982 22820 19986 22876
rect 19922 22816 19986 22820
rect 20002 22876 20066 22880
rect 20002 22820 20006 22876
rect 20006 22820 20062 22876
rect 20062 22820 20066 22876
rect 20002 22816 20066 22820
rect 20082 22876 20146 22880
rect 20082 22820 20086 22876
rect 20086 22820 20142 22876
rect 20142 22820 20146 22876
rect 20082 22816 20146 22820
rect 5674 22332 5738 22336
rect 5674 22276 5678 22332
rect 5678 22276 5734 22332
rect 5734 22276 5738 22332
rect 5674 22272 5738 22276
rect 5754 22332 5818 22336
rect 5754 22276 5758 22332
rect 5758 22276 5814 22332
rect 5814 22276 5818 22332
rect 5754 22272 5818 22276
rect 5834 22332 5898 22336
rect 5834 22276 5838 22332
rect 5838 22276 5894 22332
rect 5894 22276 5898 22332
rect 5834 22272 5898 22276
rect 5914 22332 5978 22336
rect 5914 22276 5918 22332
rect 5918 22276 5974 22332
rect 5974 22276 5978 22332
rect 5914 22272 5978 22276
rect 15120 22332 15184 22336
rect 15120 22276 15124 22332
rect 15124 22276 15180 22332
rect 15180 22276 15184 22332
rect 15120 22272 15184 22276
rect 15200 22332 15264 22336
rect 15200 22276 15204 22332
rect 15204 22276 15260 22332
rect 15260 22276 15264 22332
rect 15200 22272 15264 22276
rect 15280 22332 15344 22336
rect 15280 22276 15284 22332
rect 15284 22276 15340 22332
rect 15340 22276 15344 22332
rect 15280 22272 15344 22276
rect 15360 22332 15424 22336
rect 15360 22276 15364 22332
rect 15364 22276 15420 22332
rect 15420 22276 15424 22332
rect 15360 22272 15424 22276
rect 24565 22332 24629 22336
rect 24565 22276 24569 22332
rect 24569 22276 24625 22332
rect 24625 22276 24629 22332
rect 24565 22272 24629 22276
rect 24645 22332 24709 22336
rect 24645 22276 24649 22332
rect 24649 22276 24705 22332
rect 24705 22276 24709 22332
rect 24645 22272 24709 22276
rect 24725 22332 24789 22336
rect 24725 22276 24729 22332
rect 24729 22276 24785 22332
rect 24785 22276 24789 22332
rect 24725 22272 24789 22276
rect 24805 22332 24869 22336
rect 24805 22276 24809 22332
rect 24809 22276 24865 22332
rect 24865 22276 24869 22332
rect 24805 22272 24869 22276
rect 19564 21932 19628 21996
rect 10397 21788 10461 21792
rect 10397 21732 10401 21788
rect 10401 21732 10457 21788
rect 10457 21732 10461 21788
rect 10397 21728 10461 21732
rect 10477 21788 10541 21792
rect 10477 21732 10481 21788
rect 10481 21732 10537 21788
rect 10537 21732 10541 21788
rect 10477 21728 10541 21732
rect 10557 21788 10621 21792
rect 10557 21732 10561 21788
rect 10561 21732 10617 21788
rect 10617 21732 10621 21788
rect 10557 21728 10621 21732
rect 10637 21788 10701 21792
rect 10637 21732 10641 21788
rect 10641 21732 10697 21788
rect 10697 21732 10701 21788
rect 10637 21728 10701 21732
rect 19842 21788 19906 21792
rect 19842 21732 19846 21788
rect 19846 21732 19902 21788
rect 19902 21732 19906 21788
rect 19842 21728 19906 21732
rect 19922 21788 19986 21792
rect 19922 21732 19926 21788
rect 19926 21732 19982 21788
rect 19982 21732 19986 21788
rect 19922 21728 19986 21732
rect 20002 21788 20066 21792
rect 20002 21732 20006 21788
rect 20006 21732 20062 21788
rect 20062 21732 20066 21788
rect 20002 21728 20066 21732
rect 20082 21788 20146 21792
rect 20082 21732 20086 21788
rect 20086 21732 20142 21788
rect 20142 21732 20146 21788
rect 20082 21728 20146 21732
rect 5674 21244 5738 21248
rect 5674 21188 5678 21244
rect 5678 21188 5734 21244
rect 5734 21188 5738 21244
rect 5674 21184 5738 21188
rect 5754 21244 5818 21248
rect 5754 21188 5758 21244
rect 5758 21188 5814 21244
rect 5814 21188 5818 21244
rect 5754 21184 5818 21188
rect 5834 21244 5898 21248
rect 5834 21188 5838 21244
rect 5838 21188 5894 21244
rect 5894 21188 5898 21244
rect 5834 21184 5898 21188
rect 5914 21244 5978 21248
rect 5914 21188 5918 21244
rect 5918 21188 5974 21244
rect 5974 21188 5978 21244
rect 5914 21184 5978 21188
rect 15120 21244 15184 21248
rect 15120 21188 15124 21244
rect 15124 21188 15180 21244
rect 15180 21188 15184 21244
rect 15120 21184 15184 21188
rect 15200 21244 15264 21248
rect 15200 21188 15204 21244
rect 15204 21188 15260 21244
rect 15260 21188 15264 21244
rect 15200 21184 15264 21188
rect 15280 21244 15344 21248
rect 15280 21188 15284 21244
rect 15284 21188 15340 21244
rect 15340 21188 15344 21244
rect 15280 21184 15344 21188
rect 15360 21244 15424 21248
rect 15360 21188 15364 21244
rect 15364 21188 15420 21244
rect 15420 21188 15424 21244
rect 15360 21184 15424 21188
rect 24565 21244 24629 21248
rect 24565 21188 24569 21244
rect 24569 21188 24625 21244
rect 24625 21188 24629 21244
rect 24565 21184 24629 21188
rect 24645 21244 24709 21248
rect 24645 21188 24649 21244
rect 24649 21188 24705 21244
rect 24705 21188 24709 21244
rect 24645 21184 24709 21188
rect 24725 21244 24789 21248
rect 24725 21188 24729 21244
rect 24729 21188 24785 21244
rect 24785 21188 24789 21244
rect 24725 21184 24789 21188
rect 24805 21244 24869 21248
rect 24805 21188 24809 21244
rect 24809 21188 24865 21244
rect 24865 21188 24869 21244
rect 24805 21184 24869 21188
rect 10397 20700 10461 20704
rect 10397 20644 10401 20700
rect 10401 20644 10457 20700
rect 10457 20644 10461 20700
rect 10397 20640 10461 20644
rect 10477 20700 10541 20704
rect 10477 20644 10481 20700
rect 10481 20644 10537 20700
rect 10537 20644 10541 20700
rect 10477 20640 10541 20644
rect 10557 20700 10621 20704
rect 10557 20644 10561 20700
rect 10561 20644 10617 20700
rect 10617 20644 10621 20700
rect 10557 20640 10621 20644
rect 10637 20700 10701 20704
rect 10637 20644 10641 20700
rect 10641 20644 10697 20700
rect 10697 20644 10701 20700
rect 10637 20640 10701 20644
rect 19842 20700 19906 20704
rect 19842 20644 19846 20700
rect 19846 20644 19902 20700
rect 19902 20644 19906 20700
rect 19842 20640 19906 20644
rect 19922 20700 19986 20704
rect 19922 20644 19926 20700
rect 19926 20644 19982 20700
rect 19982 20644 19986 20700
rect 19922 20640 19986 20644
rect 20002 20700 20066 20704
rect 20002 20644 20006 20700
rect 20006 20644 20062 20700
rect 20062 20644 20066 20700
rect 20002 20640 20066 20644
rect 20082 20700 20146 20704
rect 20082 20644 20086 20700
rect 20086 20644 20142 20700
rect 20142 20644 20146 20700
rect 20082 20640 20146 20644
rect 5674 20156 5738 20160
rect 5674 20100 5678 20156
rect 5678 20100 5734 20156
rect 5734 20100 5738 20156
rect 5674 20096 5738 20100
rect 5754 20156 5818 20160
rect 5754 20100 5758 20156
rect 5758 20100 5814 20156
rect 5814 20100 5818 20156
rect 5754 20096 5818 20100
rect 5834 20156 5898 20160
rect 5834 20100 5838 20156
rect 5838 20100 5894 20156
rect 5894 20100 5898 20156
rect 5834 20096 5898 20100
rect 5914 20156 5978 20160
rect 5914 20100 5918 20156
rect 5918 20100 5974 20156
rect 5974 20100 5978 20156
rect 5914 20096 5978 20100
rect 15120 20156 15184 20160
rect 15120 20100 15124 20156
rect 15124 20100 15180 20156
rect 15180 20100 15184 20156
rect 15120 20096 15184 20100
rect 15200 20156 15264 20160
rect 15200 20100 15204 20156
rect 15204 20100 15260 20156
rect 15260 20100 15264 20156
rect 15200 20096 15264 20100
rect 15280 20156 15344 20160
rect 15280 20100 15284 20156
rect 15284 20100 15340 20156
rect 15340 20100 15344 20156
rect 15280 20096 15344 20100
rect 15360 20156 15424 20160
rect 15360 20100 15364 20156
rect 15364 20100 15420 20156
rect 15420 20100 15424 20156
rect 15360 20096 15424 20100
rect 24565 20156 24629 20160
rect 24565 20100 24569 20156
rect 24569 20100 24625 20156
rect 24625 20100 24629 20156
rect 24565 20096 24629 20100
rect 24645 20156 24709 20160
rect 24645 20100 24649 20156
rect 24649 20100 24705 20156
rect 24705 20100 24709 20156
rect 24645 20096 24709 20100
rect 24725 20156 24789 20160
rect 24725 20100 24729 20156
rect 24729 20100 24785 20156
rect 24785 20100 24789 20156
rect 24725 20096 24789 20100
rect 24805 20156 24869 20160
rect 24805 20100 24809 20156
rect 24809 20100 24865 20156
rect 24865 20100 24869 20156
rect 24805 20096 24869 20100
rect 20300 19680 20364 19684
rect 20300 19624 20314 19680
rect 20314 19624 20364 19680
rect 20300 19620 20364 19624
rect 10397 19612 10461 19616
rect 10397 19556 10401 19612
rect 10401 19556 10457 19612
rect 10457 19556 10461 19612
rect 10397 19552 10461 19556
rect 10477 19612 10541 19616
rect 10477 19556 10481 19612
rect 10481 19556 10537 19612
rect 10537 19556 10541 19612
rect 10477 19552 10541 19556
rect 10557 19612 10621 19616
rect 10557 19556 10561 19612
rect 10561 19556 10617 19612
rect 10617 19556 10621 19612
rect 10557 19552 10621 19556
rect 10637 19612 10701 19616
rect 10637 19556 10641 19612
rect 10641 19556 10697 19612
rect 10697 19556 10701 19612
rect 10637 19552 10701 19556
rect 19842 19612 19906 19616
rect 19842 19556 19846 19612
rect 19846 19556 19902 19612
rect 19902 19556 19906 19612
rect 19842 19552 19906 19556
rect 19922 19612 19986 19616
rect 19922 19556 19926 19612
rect 19926 19556 19982 19612
rect 19982 19556 19986 19612
rect 19922 19552 19986 19556
rect 20002 19612 20066 19616
rect 20002 19556 20006 19612
rect 20006 19556 20062 19612
rect 20062 19556 20066 19612
rect 20002 19552 20066 19556
rect 20082 19612 20146 19616
rect 20082 19556 20086 19612
rect 20086 19556 20142 19612
rect 20142 19556 20146 19612
rect 20082 19552 20146 19556
rect 5674 19068 5738 19072
rect 5674 19012 5678 19068
rect 5678 19012 5734 19068
rect 5734 19012 5738 19068
rect 5674 19008 5738 19012
rect 5754 19068 5818 19072
rect 5754 19012 5758 19068
rect 5758 19012 5814 19068
rect 5814 19012 5818 19068
rect 5754 19008 5818 19012
rect 5834 19068 5898 19072
rect 5834 19012 5838 19068
rect 5838 19012 5894 19068
rect 5894 19012 5898 19068
rect 5834 19008 5898 19012
rect 5914 19068 5978 19072
rect 5914 19012 5918 19068
rect 5918 19012 5974 19068
rect 5974 19012 5978 19068
rect 5914 19008 5978 19012
rect 15120 19068 15184 19072
rect 15120 19012 15124 19068
rect 15124 19012 15180 19068
rect 15180 19012 15184 19068
rect 15120 19008 15184 19012
rect 15200 19068 15264 19072
rect 15200 19012 15204 19068
rect 15204 19012 15260 19068
rect 15260 19012 15264 19068
rect 15200 19008 15264 19012
rect 15280 19068 15344 19072
rect 15280 19012 15284 19068
rect 15284 19012 15340 19068
rect 15340 19012 15344 19068
rect 15280 19008 15344 19012
rect 15360 19068 15424 19072
rect 15360 19012 15364 19068
rect 15364 19012 15420 19068
rect 15420 19012 15424 19068
rect 15360 19008 15424 19012
rect 24565 19068 24629 19072
rect 24565 19012 24569 19068
rect 24569 19012 24625 19068
rect 24625 19012 24629 19068
rect 24565 19008 24629 19012
rect 24645 19068 24709 19072
rect 24645 19012 24649 19068
rect 24649 19012 24705 19068
rect 24705 19012 24709 19068
rect 24645 19008 24709 19012
rect 24725 19068 24789 19072
rect 24725 19012 24729 19068
rect 24729 19012 24785 19068
rect 24785 19012 24789 19068
rect 24725 19008 24789 19012
rect 24805 19068 24869 19072
rect 24805 19012 24809 19068
rect 24809 19012 24865 19068
rect 24865 19012 24869 19068
rect 24805 19008 24869 19012
rect 10397 18524 10461 18528
rect 10397 18468 10401 18524
rect 10401 18468 10457 18524
rect 10457 18468 10461 18524
rect 10397 18464 10461 18468
rect 10477 18524 10541 18528
rect 10477 18468 10481 18524
rect 10481 18468 10537 18524
rect 10537 18468 10541 18524
rect 10477 18464 10541 18468
rect 10557 18524 10621 18528
rect 10557 18468 10561 18524
rect 10561 18468 10617 18524
rect 10617 18468 10621 18524
rect 10557 18464 10621 18468
rect 10637 18524 10701 18528
rect 10637 18468 10641 18524
rect 10641 18468 10697 18524
rect 10697 18468 10701 18524
rect 10637 18464 10701 18468
rect 19842 18524 19906 18528
rect 19842 18468 19846 18524
rect 19846 18468 19902 18524
rect 19902 18468 19906 18524
rect 19842 18464 19906 18468
rect 19922 18524 19986 18528
rect 19922 18468 19926 18524
rect 19926 18468 19982 18524
rect 19982 18468 19986 18524
rect 19922 18464 19986 18468
rect 20002 18524 20066 18528
rect 20002 18468 20006 18524
rect 20006 18468 20062 18524
rect 20062 18468 20066 18524
rect 20002 18464 20066 18468
rect 20082 18524 20146 18528
rect 20082 18468 20086 18524
rect 20086 18468 20142 18524
rect 20142 18468 20146 18524
rect 20082 18464 20146 18468
rect 5674 17980 5738 17984
rect 5674 17924 5678 17980
rect 5678 17924 5734 17980
rect 5734 17924 5738 17980
rect 5674 17920 5738 17924
rect 5754 17980 5818 17984
rect 5754 17924 5758 17980
rect 5758 17924 5814 17980
rect 5814 17924 5818 17980
rect 5754 17920 5818 17924
rect 5834 17980 5898 17984
rect 5834 17924 5838 17980
rect 5838 17924 5894 17980
rect 5894 17924 5898 17980
rect 5834 17920 5898 17924
rect 5914 17980 5978 17984
rect 5914 17924 5918 17980
rect 5918 17924 5974 17980
rect 5974 17924 5978 17980
rect 5914 17920 5978 17924
rect 15120 17980 15184 17984
rect 15120 17924 15124 17980
rect 15124 17924 15180 17980
rect 15180 17924 15184 17980
rect 15120 17920 15184 17924
rect 15200 17980 15264 17984
rect 15200 17924 15204 17980
rect 15204 17924 15260 17980
rect 15260 17924 15264 17980
rect 15200 17920 15264 17924
rect 15280 17980 15344 17984
rect 15280 17924 15284 17980
rect 15284 17924 15340 17980
rect 15340 17924 15344 17980
rect 15280 17920 15344 17924
rect 15360 17980 15424 17984
rect 15360 17924 15364 17980
rect 15364 17924 15420 17980
rect 15420 17924 15424 17980
rect 15360 17920 15424 17924
rect 24565 17980 24629 17984
rect 24565 17924 24569 17980
rect 24569 17924 24625 17980
rect 24625 17924 24629 17980
rect 24565 17920 24629 17924
rect 24645 17980 24709 17984
rect 24645 17924 24649 17980
rect 24649 17924 24705 17980
rect 24705 17924 24709 17980
rect 24645 17920 24709 17924
rect 24725 17980 24789 17984
rect 24725 17924 24729 17980
rect 24729 17924 24785 17980
rect 24785 17924 24789 17980
rect 24725 17920 24789 17924
rect 24805 17980 24869 17984
rect 24805 17924 24809 17980
rect 24809 17924 24865 17980
rect 24865 17924 24869 17980
rect 24805 17920 24869 17924
rect 19380 17852 19444 17916
rect 10397 17436 10461 17440
rect 10397 17380 10401 17436
rect 10401 17380 10457 17436
rect 10457 17380 10461 17436
rect 10397 17376 10461 17380
rect 10477 17436 10541 17440
rect 10477 17380 10481 17436
rect 10481 17380 10537 17436
rect 10537 17380 10541 17436
rect 10477 17376 10541 17380
rect 10557 17436 10621 17440
rect 10557 17380 10561 17436
rect 10561 17380 10617 17436
rect 10617 17380 10621 17436
rect 10557 17376 10621 17380
rect 10637 17436 10701 17440
rect 10637 17380 10641 17436
rect 10641 17380 10697 17436
rect 10697 17380 10701 17436
rect 10637 17376 10701 17380
rect 19842 17436 19906 17440
rect 19842 17380 19846 17436
rect 19846 17380 19902 17436
rect 19902 17380 19906 17436
rect 19842 17376 19906 17380
rect 19922 17436 19986 17440
rect 19922 17380 19926 17436
rect 19926 17380 19982 17436
rect 19982 17380 19986 17436
rect 19922 17376 19986 17380
rect 20002 17436 20066 17440
rect 20002 17380 20006 17436
rect 20006 17380 20062 17436
rect 20062 17380 20066 17436
rect 20002 17376 20066 17380
rect 20082 17436 20146 17440
rect 20082 17380 20086 17436
rect 20086 17380 20142 17436
rect 20142 17380 20146 17436
rect 20082 17376 20146 17380
rect 5674 16892 5738 16896
rect 5674 16836 5678 16892
rect 5678 16836 5734 16892
rect 5734 16836 5738 16892
rect 5674 16832 5738 16836
rect 5754 16892 5818 16896
rect 5754 16836 5758 16892
rect 5758 16836 5814 16892
rect 5814 16836 5818 16892
rect 5754 16832 5818 16836
rect 5834 16892 5898 16896
rect 5834 16836 5838 16892
rect 5838 16836 5894 16892
rect 5894 16836 5898 16892
rect 5834 16832 5898 16836
rect 5914 16892 5978 16896
rect 5914 16836 5918 16892
rect 5918 16836 5974 16892
rect 5974 16836 5978 16892
rect 5914 16832 5978 16836
rect 15120 16892 15184 16896
rect 15120 16836 15124 16892
rect 15124 16836 15180 16892
rect 15180 16836 15184 16892
rect 15120 16832 15184 16836
rect 15200 16892 15264 16896
rect 15200 16836 15204 16892
rect 15204 16836 15260 16892
rect 15260 16836 15264 16892
rect 15200 16832 15264 16836
rect 15280 16892 15344 16896
rect 15280 16836 15284 16892
rect 15284 16836 15340 16892
rect 15340 16836 15344 16892
rect 15280 16832 15344 16836
rect 15360 16892 15424 16896
rect 15360 16836 15364 16892
rect 15364 16836 15420 16892
rect 15420 16836 15424 16892
rect 15360 16832 15424 16836
rect 24565 16892 24629 16896
rect 24565 16836 24569 16892
rect 24569 16836 24625 16892
rect 24625 16836 24629 16892
rect 24565 16832 24629 16836
rect 24645 16892 24709 16896
rect 24645 16836 24649 16892
rect 24649 16836 24705 16892
rect 24705 16836 24709 16892
rect 24645 16832 24709 16836
rect 24725 16892 24789 16896
rect 24725 16836 24729 16892
rect 24729 16836 24785 16892
rect 24785 16836 24789 16892
rect 24725 16832 24789 16836
rect 24805 16892 24869 16896
rect 24805 16836 24809 16892
rect 24809 16836 24865 16892
rect 24865 16836 24869 16892
rect 24805 16832 24869 16836
rect 10397 16348 10461 16352
rect 10397 16292 10401 16348
rect 10401 16292 10457 16348
rect 10457 16292 10461 16348
rect 10397 16288 10461 16292
rect 10477 16348 10541 16352
rect 10477 16292 10481 16348
rect 10481 16292 10537 16348
rect 10537 16292 10541 16348
rect 10477 16288 10541 16292
rect 10557 16348 10621 16352
rect 10557 16292 10561 16348
rect 10561 16292 10617 16348
rect 10617 16292 10621 16348
rect 10557 16288 10621 16292
rect 10637 16348 10701 16352
rect 10637 16292 10641 16348
rect 10641 16292 10697 16348
rect 10697 16292 10701 16348
rect 10637 16288 10701 16292
rect 19842 16348 19906 16352
rect 19842 16292 19846 16348
rect 19846 16292 19902 16348
rect 19902 16292 19906 16348
rect 19842 16288 19906 16292
rect 19922 16348 19986 16352
rect 19922 16292 19926 16348
rect 19926 16292 19982 16348
rect 19982 16292 19986 16348
rect 19922 16288 19986 16292
rect 20002 16348 20066 16352
rect 20002 16292 20006 16348
rect 20006 16292 20062 16348
rect 20062 16292 20066 16348
rect 20002 16288 20066 16292
rect 20082 16348 20146 16352
rect 20082 16292 20086 16348
rect 20086 16292 20142 16348
rect 20142 16292 20146 16348
rect 20082 16288 20146 16292
rect 5674 15804 5738 15808
rect 5674 15748 5678 15804
rect 5678 15748 5734 15804
rect 5734 15748 5738 15804
rect 5674 15744 5738 15748
rect 5754 15804 5818 15808
rect 5754 15748 5758 15804
rect 5758 15748 5814 15804
rect 5814 15748 5818 15804
rect 5754 15744 5818 15748
rect 5834 15804 5898 15808
rect 5834 15748 5838 15804
rect 5838 15748 5894 15804
rect 5894 15748 5898 15804
rect 5834 15744 5898 15748
rect 5914 15804 5978 15808
rect 5914 15748 5918 15804
rect 5918 15748 5974 15804
rect 5974 15748 5978 15804
rect 5914 15744 5978 15748
rect 15120 15804 15184 15808
rect 15120 15748 15124 15804
rect 15124 15748 15180 15804
rect 15180 15748 15184 15804
rect 15120 15744 15184 15748
rect 15200 15804 15264 15808
rect 15200 15748 15204 15804
rect 15204 15748 15260 15804
rect 15260 15748 15264 15804
rect 15200 15744 15264 15748
rect 15280 15804 15344 15808
rect 15280 15748 15284 15804
rect 15284 15748 15340 15804
rect 15340 15748 15344 15804
rect 15280 15744 15344 15748
rect 15360 15804 15424 15808
rect 15360 15748 15364 15804
rect 15364 15748 15420 15804
rect 15420 15748 15424 15804
rect 15360 15744 15424 15748
rect 24565 15804 24629 15808
rect 24565 15748 24569 15804
rect 24569 15748 24625 15804
rect 24625 15748 24629 15804
rect 24565 15744 24629 15748
rect 24645 15804 24709 15808
rect 24645 15748 24649 15804
rect 24649 15748 24705 15804
rect 24705 15748 24709 15804
rect 24645 15744 24709 15748
rect 24725 15804 24789 15808
rect 24725 15748 24729 15804
rect 24729 15748 24785 15804
rect 24785 15748 24789 15804
rect 24725 15744 24789 15748
rect 24805 15804 24869 15808
rect 24805 15748 24809 15804
rect 24809 15748 24865 15804
rect 24865 15748 24869 15804
rect 24805 15744 24869 15748
rect 10397 15260 10461 15264
rect 10397 15204 10401 15260
rect 10401 15204 10457 15260
rect 10457 15204 10461 15260
rect 10397 15200 10461 15204
rect 10477 15260 10541 15264
rect 10477 15204 10481 15260
rect 10481 15204 10537 15260
rect 10537 15204 10541 15260
rect 10477 15200 10541 15204
rect 10557 15260 10621 15264
rect 10557 15204 10561 15260
rect 10561 15204 10617 15260
rect 10617 15204 10621 15260
rect 10557 15200 10621 15204
rect 10637 15260 10701 15264
rect 10637 15204 10641 15260
rect 10641 15204 10697 15260
rect 10697 15204 10701 15260
rect 10637 15200 10701 15204
rect 19842 15260 19906 15264
rect 19842 15204 19846 15260
rect 19846 15204 19902 15260
rect 19902 15204 19906 15260
rect 19842 15200 19906 15204
rect 19922 15260 19986 15264
rect 19922 15204 19926 15260
rect 19926 15204 19982 15260
rect 19982 15204 19986 15260
rect 19922 15200 19986 15204
rect 20002 15260 20066 15264
rect 20002 15204 20006 15260
rect 20006 15204 20062 15260
rect 20062 15204 20066 15260
rect 20002 15200 20066 15204
rect 20082 15260 20146 15264
rect 20082 15204 20086 15260
rect 20086 15204 20142 15260
rect 20142 15204 20146 15260
rect 20082 15200 20146 15204
rect 5674 14716 5738 14720
rect 5674 14660 5678 14716
rect 5678 14660 5734 14716
rect 5734 14660 5738 14716
rect 5674 14656 5738 14660
rect 5754 14716 5818 14720
rect 5754 14660 5758 14716
rect 5758 14660 5814 14716
rect 5814 14660 5818 14716
rect 5754 14656 5818 14660
rect 5834 14716 5898 14720
rect 5834 14660 5838 14716
rect 5838 14660 5894 14716
rect 5894 14660 5898 14716
rect 5834 14656 5898 14660
rect 5914 14716 5978 14720
rect 5914 14660 5918 14716
rect 5918 14660 5974 14716
rect 5974 14660 5978 14716
rect 5914 14656 5978 14660
rect 15120 14716 15184 14720
rect 15120 14660 15124 14716
rect 15124 14660 15180 14716
rect 15180 14660 15184 14716
rect 15120 14656 15184 14660
rect 15200 14716 15264 14720
rect 15200 14660 15204 14716
rect 15204 14660 15260 14716
rect 15260 14660 15264 14716
rect 15200 14656 15264 14660
rect 15280 14716 15344 14720
rect 15280 14660 15284 14716
rect 15284 14660 15340 14716
rect 15340 14660 15344 14716
rect 15280 14656 15344 14660
rect 15360 14716 15424 14720
rect 15360 14660 15364 14716
rect 15364 14660 15420 14716
rect 15420 14660 15424 14716
rect 15360 14656 15424 14660
rect 24565 14716 24629 14720
rect 24565 14660 24569 14716
rect 24569 14660 24625 14716
rect 24625 14660 24629 14716
rect 24565 14656 24629 14660
rect 24645 14716 24709 14720
rect 24645 14660 24649 14716
rect 24649 14660 24705 14716
rect 24705 14660 24709 14716
rect 24645 14656 24709 14660
rect 24725 14716 24789 14720
rect 24725 14660 24729 14716
rect 24729 14660 24785 14716
rect 24785 14660 24789 14716
rect 24725 14656 24789 14660
rect 24805 14716 24869 14720
rect 24805 14660 24809 14716
rect 24809 14660 24865 14716
rect 24865 14660 24869 14716
rect 24805 14656 24869 14660
rect 10397 14172 10461 14176
rect 10397 14116 10401 14172
rect 10401 14116 10457 14172
rect 10457 14116 10461 14172
rect 10397 14112 10461 14116
rect 10477 14172 10541 14176
rect 10477 14116 10481 14172
rect 10481 14116 10537 14172
rect 10537 14116 10541 14172
rect 10477 14112 10541 14116
rect 10557 14172 10621 14176
rect 10557 14116 10561 14172
rect 10561 14116 10617 14172
rect 10617 14116 10621 14172
rect 10557 14112 10621 14116
rect 10637 14172 10701 14176
rect 10637 14116 10641 14172
rect 10641 14116 10697 14172
rect 10697 14116 10701 14172
rect 10637 14112 10701 14116
rect 19842 14172 19906 14176
rect 19842 14116 19846 14172
rect 19846 14116 19902 14172
rect 19902 14116 19906 14172
rect 19842 14112 19906 14116
rect 19922 14172 19986 14176
rect 19922 14116 19926 14172
rect 19926 14116 19982 14172
rect 19982 14116 19986 14172
rect 19922 14112 19986 14116
rect 20002 14172 20066 14176
rect 20002 14116 20006 14172
rect 20006 14116 20062 14172
rect 20062 14116 20066 14172
rect 20002 14112 20066 14116
rect 20082 14172 20146 14176
rect 20082 14116 20086 14172
rect 20086 14116 20142 14172
rect 20142 14116 20146 14172
rect 20082 14112 20146 14116
rect 12572 14044 12636 14108
rect 5674 13628 5738 13632
rect 5674 13572 5678 13628
rect 5678 13572 5734 13628
rect 5734 13572 5738 13628
rect 5674 13568 5738 13572
rect 5754 13628 5818 13632
rect 5754 13572 5758 13628
rect 5758 13572 5814 13628
rect 5814 13572 5818 13628
rect 5754 13568 5818 13572
rect 5834 13628 5898 13632
rect 5834 13572 5838 13628
rect 5838 13572 5894 13628
rect 5894 13572 5898 13628
rect 5834 13568 5898 13572
rect 5914 13628 5978 13632
rect 5914 13572 5918 13628
rect 5918 13572 5974 13628
rect 5974 13572 5978 13628
rect 5914 13568 5978 13572
rect 15120 13628 15184 13632
rect 15120 13572 15124 13628
rect 15124 13572 15180 13628
rect 15180 13572 15184 13628
rect 15120 13568 15184 13572
rect 15200 13628 15264 13632
rect 15200 13572 15204 13628
rect 15204 13572 15260 13628
rect 15260 13572 15264 13628
rect 15200 13568 15264 13572
rect 15280 13628 15344 13632
rect 15280 13572 15284 13628
rect 15284 13572 15340 13628
rect 15340 13572 15344 13628
rect 15280 13568 15344 13572
rect 15360 13628 15424 13632
rect 15360 13572 15364 13628
rect 15364 13572 15420 13628
rect 15420 13572 15424 13628
rect 15360 13568 15424 13572
rect 24565 13628 24629 13632
rect 24565 13572 24569 13628
rect 24569 13572 24625 13628
rect 24625 13572 24629 13628
rect 24565 13568 24629 13572
rect 24645 13628 24709 13632
rect 24645 13572 24649 13628
rect 24649 13572 24705 13628
rect 24705 13572 24709 13628
rect 24645 13568 24709 13572
rect 24725 13628 24789 13632
rect 24725 13572 24729 13628
rect 24729 13572 24785 13628
rect 24785 13572 24789 13628
rect 24725 13568 24789 13572
rect 24805 13628 24869 13632
rect 24805 13572 24809 13628
rect 24809 13572 24865 13628
rect 24865 13572 24869 13628
rect 24805 13568 24869 13572
rect 10397 13084 10461 13088
rect 10397 13028 10401 13084
rect 10401 13028 10457 13084
rect 10457 13028 10461 13084
rect 10397 13024 10461 13028
rect 10477 13084 10541 13088
rect 10477 13028 10481 13084
rect 10481 13028 10537 13084
rect 10537 13028 10541 13084
rect 10477 13024 10541 13028
rect 10557 13084 10621 13088
rect 10557 13028 10561 13084
rect 10561 13028 10617 13084
rect 10617 13028 10621 13084
rect 10557 13024 10621 13028
rect 10637 13084 10701 13088
rect 10637 13028 10641 13084
rect 10641 13028 10697 13084
rect 10697 13028 10701 13084
rect 10637 13024 10701 13028
rect 19842 13084 19906 13088
rect 19842 13028 19846 13084
rect 19846 13028 19902 13084
rect 19902 13028 19906 13084
rect 19842 13024 19906 13028
rect 19922 13084 19986 13088
rect 19922 13028 19926 13084
rect 19926 13028 19982 13084
rect 19982 13028 19986 13084
rect 19922 13024 19986 13028
rect 20002 13084 20066 13088
rect 20002 13028 20006 13084
rect 20006 13028 20062 13084
rect 20062 13028 20066 13084
rect 20002 13024 20066 13028
rect 20082 13084 20146 13088
rect 20082 13028 20086 13084
rect 20086 13028 20142 13084
rect 20142 13028 20146 13084
rect 20082 13024 20146 13028
rect 5674 12540 5738 12544
rect 5674 12484 5678 12540
rect 5678 12484 5734 12540
rect 5734 12484 5738 12540
rect 5674 12480 5738 12484
rect 5754 12540 5818 12544
rect 5754 12484 5758 12540
rect 5758 12484 5814 12540
rect 5814 12484 5818 12540
rect 5754 12480 5818 12484
rect 5834 12540 5898 12544
rect 5834 12484 5838 12540
rect 5838 12484 5894 12540
rect 5894 12484 5898 12540
rect 5834 12480 5898 12484
rect 5914 12540 5978 12544
rect 5914 12484 5918 12540
rect 5918 12484 5974 12540
rect 5974 12484 5978 12540
rect 5914 12480 5978 12484
rect 15120 12540 15184 12544
rect 15120 12484 15124 12540
rect 15124 12484 15180 12540
rect 15180 12484 15184 12540
rect 15120 12480 15184 12484
rect 15200 12540 15264 12544
rect 15200 12484 15204 12540
rect 15204 12484 15260 12540
rect 15260 12484 15264 12540
rect 15200 12480 15264 12484
rect 15280 12540 15344 12544
rect 15280 12484 15284 12540
rect 15284 12484 15340 12540
rect 15340 12484 15344 12540
rect 15280 12480 15344 12484
rect 15360 12540 15424 12544
rect 15360 12484 15364 12540
rect 15364 12484 15420 12540
rect 15420 12484 15424 12540
rect 15360 12480 15424 12484
rect 24565 12540 24629 12544
rect 24565 12484 24569 12540
rect 24569 12484 24625 12540
rect 24625 12484 24629 12540
rect 24565 12480 24629 12484
rect 24645 12540 24709 12544
rect 24645 12484 24649 12540
rect 24649 12484 24705 12540
rect 24705 12484 24709 12540
rect 24645 12480 24709 12484
rect 24725 12540 24789 12544
rect 24725 12484 24729 12540
rect 24729 12484 24785 12540
rect 24785 12484 24789 12540
rect 24725 12480 24789 12484
rect 24805 12540 24869 12544
rect 24805 12484 24809 12540
rect 24809 12484 24865 12540
rect 24865 12484 24869 12540
rect 24805 12480 24869 12484
rect 10397 11996 10461 12000
rect 10397 11940 10401 11996
rect 10401 11940 10457 11996
rect 10457 11940 10461 11996
rect 10397 11936 10461 11940
rect 10477 11996 10541 12000
rect 10477 11940 10481 11996
rect 10481 11940 10537 11996
rect 10537 11940 10541 11996
rect 10477 11936 10541 11940
rect 10557 11996 10621 12000
rect 10557 11940 10561 11996
rect 10561 11940 10617 11996
rect 10617 11940 10621 11996
rect 10557 11936 10621 11940
rect 10637 11996 10701 12000
rect 10637 11940 10641 11996
rect 10641 11940 10697 11996
rect 10697 11940 10701 11996
rect 10637 11936 10701 11940
rect 19842 11996 19906 12000
rect 19842 11940 19846 11996
rect 19846 11940 19902 11996
rect 19902 11940 19906 11996
rect 19842 11936 19906 11940
rect 19922 11996 19986 12000
rect 19922 11940 19926 11996
rect 19926 11940 19982 11996
rect 19982 11940 19986 11996
rect 19922 11936 19986 11940
rect 20002 11996 20066 12000
rect 20002 11940 20006 11996
rect 20006 11940 20062 11996
rect 20062 11940 20066 11996
rect 20002 11936 20066 11940
rect 20082 11996 20146 12000
rect 20082 11940 20086 11996
rect 20086 11940 20142 11996
rect 20142 11940 20146 11996
rect 20082 11936 20146 11940
rect 5674 11452 5738 11456
rect 5674 11396 5678 11452
rect 5678 11396 5734 11452
rect 5734 11396 5738 11452
rect 5674 11392 5738 11396
rect 5754 11452 5818 11456
rect 5754 11396 5758 11452
rect 5758 11396 5814 11452
rect 5814 11396 5818 11452
rect 5754 11392 5818 11396
rect 5834 11452 5898 11456
rect 5834 11396 5838 11452
rect 5838 11396 5894 11452
rect 5894 11396 5898 11452
rect 5834 11392 5898 11396
rect 5914 11452 5978 11456
rect 5914 11396 5918 11452
rect 5918 11396 5974 11452
rect 5974 11396 5978 11452
rect 5914 11392 5978 11396
rect 15120 11452 15184 11456
rect 15120 11396 15124 11452
rect 15124 11396 15180 11452
rect 15180 11396 15184 11452
rect 15120 11392 15184 11396
rect 15200 11452 15264 11456
rect 15200 11396 15204 11452
rect 15204 11396 15260 11452
rect 15260 11396 15264 11452
rect 15200 11392 15264 11396
rect 15280 11452 15344 11456
rect 15280 11396 15284 11452
rect 15284 11396 15340 11452
rect 15340 11396 15344 11452
rect 15280 11392 15344 11396
rect 15360 11452 15424 11456
rect 15360 11396 15364 11452
rect 15364 11396 15420 11452
rect 15420 11396 15424 11452
rect 15360 11392 15424 11396
rect 24565 11452 24629 11456
rect 24565 11396 24569 11452
rect 24569 11396 24625 11452
rect 24625 11396 24629 11452
rect 24565 11392 24629 11396
rect 24645 11452 24709 11456
rect 24645 11396 24649 11452
rect 24649 11396 24705 11452
rect 24705 11396 24709 11452
rect 24645 11392 24709 11396
rect 24725 11452 24789 11456
rect 24725 11396 24729 11452
rect 24729 11396 24785 11452
rect 24785 11396 24789 11452
rect 24725 11392 24789 11396
rect 24805 11452 24869 11456
rect 24805 11396 24809 11452
rect 24809 11396 24865 11452
rect 24865 11396 24869 11452
rect 24805 11392 24869 11396
rect 10397 10908 10461 10912
rect 10397 10852 10401 10908
rect 10401 10852 10457 10908
rect 10457 10852 10461 10908
rect 10397 10848 10461 10852
rect 10477 10908 10541 10912
rect 10477 10852 10481 10908
rect 10481 10852 10537 10908
rect 10537 10852 10541 10908
rect 10477 10848 10541 10852
rect 10557 10908 10621 10912
rect 10557 10852 10561 10908
rect 10561 10852 10617 10908
rect 10617 10852 10621 10908
rect 10557 10848 10621 10852
rect 10637 10908 10701 10912
rect 10637 10852 10641 10908
rect 10641 10852 10697 10908
rect 10697 10852 10701 10908
rect 10637 10848 10701 10852
rect 19842 10908 19906 10912
rect 19842 10852 19846 10908
rect 19846 10852 19902 10908
rect 19902 10852 19906 10908
rect 19842 10848 19906 10852
rect 19922 10908 19986 10912
rect 19922 10852 19926 10908
rect 19926 10852 19982 10908
rect 19982 10852 19986 10908
rect 19922 10848 19986 10852
rect 20002 10908 20066 10912
rect 20002 10852 20006 10908
rect 20006 10852 20062 10908
rect 20062 10852 20066 10908
rect 20002 10848 20066 10852
rect 20082 10908 20146 10912
rect 20082 10852 20086 10908
rect 20086 10852 20142 10908
rect 20142 10852 20146 10908
rect 20082 10848 20146 10852
rect 5674 10364 5738 10368
rect 5674 10308 5678 10364
rect 5678 10308 5734 10364
rect 5734 10308 5738 10364
rect 5674 10304 5738 10308
rect 5754 10364 5818 10368
rect 5754 10308 5758 10364
rect 5758 10308 5814 10364
rect 5814 10308 5818 10364
rect 5754 10304 5818 10308
rect 5834 10364 5898 10368
rect 5834 10308 5838 10364
rect 5838 10308 5894 10364
rect 5894 10308 5898 10364
rect 5834 10304 5898 10308
rect 5914 10364 5978 10368
rect 5914 10308 5918 10364
rect 5918 10308 5974 10364
rect 5974 10308 5978 10364
rect 5914 10304 5978 10308
rect 15120 10364 15184 10368
rect 15120 10308 15124 10364
rect 15124 10308 15180 10364
rect 15180 10308 15184 10364
rect 15120 10304 15184 10308
rect 15200 10364 15264 10368
rect 15200 10308 15204 10364
rect 15204 10308 15260 10364
rect 15260 10308 15264 10364
rect 15200 10304 15264 10308
rect 15280 10364 15344 10368
rect 15280 10308 15284 10364
rect 15284 10308 15340 10364
rect 15340 10308 15344 10364
rect 15280 10304 15344 10308
rect 15360 10364 15424 10368
rect 15360 10308 15364 10364
rect 15364 10308 15420 10364
rect 15420 10308 15424 10364
rect 15360 10304 15424 10308
rect 24565 10364 24629 10368
rect 24565 10308 24569 10364
rect 24569 10308 24625 10364
rect 24625 10308 24629 10364
rect 24565 10304 24629 10308
rect 24645 10364 24709 10368
rect 24645 10308 24649 10364
rect 24649 10308 24705 10364
rect 24705 10308 24709 10364
rect 24645 10304 24709 10308
rect 24725 10364 24789 10368
rect 24725 10308 24729 10364
rect 24729 10308 24785 10364
rect 24785 10308 24789 10364
rect 24725 10304 24789 10308
rect 24805 10364 24869 10368
rect 24805 10308 24809 10364
rect 24809 10308 24865 10364
rect 24865 10308 24869 10364
rect 24805 10304 24869 10308
rect 10397 9820 10461 9824
rect 10397 9764 10401 9820
rect 10401 9764 10457 9820
rect 10457 9764 10461 9820
rect 10397 9760 10461 9764
rect 10477 9820 10541 9824
rect 10477 9764 10481 9820
rect 10481 9764 10537 9820
rect 10537 9764 10541 9820
rect 10477 9760 10541 9764
rect 10557 9820 10621 9824
rect 10557 9764 10561 9820
rect 10561 9764 10617 9820
rect 10617 9764 10621 9820
rect 10557 9760 10621 9764
rect 10637 9820 10701 9824
rect 10637 9764 10641 9820
rect 10641 9764 10697 9820
rect 10697 9764 10701 9820
rect 10637 9760 10701 9764
rect 19842 9820 19906 9824
rect 19842 9764 19846 9820
rect 19846 9764 19902 9820
rect 19902 9764 19906 9820
rect 19842 9760 19906 9764
rect 19922 9820 19986 9824
rect 19922 9764 19926 9820
rect 19926 9764 19982 9820
rect 19982 9764 19986 9820
rect 19922 9760 19986 9764
rect 20002 9820 20066 9824
rect 20002 9764 20006 9820
rect 20006 9764 20062 9820
rect 20062 9764 20066 9820
rect 20002 9760 20066 9764
rect 20082 9820 20146 9824
rect 20082 9764 20086 9820
rect 20086 9764 20142 9820
rect 20142 9764 20146 9820
rect 20082 9760 20146 9764
rect 5674 9276 5738 9280
rect 5674 9220 5678 9276
rect 5678 9220 5734 9276
rect 5734 9220 5738 9276
rect 5674 9216 5738 9220
rect 5754 9276 5818 9280
rect 5754 9220 5758 9276
rect 5758 9220 5814 9276
rect 5814 9220 5818 9276
rect 5754 9216 5818 9220
rect 5834 9276 5898 9280
rect 5834 9220 5838 9276
rect 5838 9220 5894 9276
rect 5894 9220 5898 9276
rect 5834 9216 5898 9220
rect 5914 9276 5978 9280
rect 5914 9220 5918 9276
rect 5918 9220 5974 9276
rect 5974 9220 5978 9276
rect 5914 9216 5978 9220
rect 15120 9276 15184 9280
rect 15120 9220 15124 9276
rect 15124 9220 15180 9276
rect 15180 9220 15184 9276
rect 15120 9216 15184 9220
rect 15200 9276 15264 9280
rect 15200 9220 15204 9276
rect 15204 9220 15260 9276
rect 15260 9220 15264 9276
rect 15200 9216 15264 9220
rect 15280 9276 15344 9280
rect 15280 9220 15284 9276
rect 15284 9220 15340 9276
rect 15340 9220 15344 9276
rect 15280 9216 15344 9220
rect 15360 9276 15424 9280
rect 15360 9220 15364 9276
rect 15364 9220 15420 9276
rect 15420 9220 15424 9276
rect 15360 9216 15424 9220
rect 24565 9276 24629 9280
rect 24565 9220 24569 9276
rect 24569 9220 24625 9276
rect 24625 9220 24629 9276
rect 24565 9216 24629 9220
rect 24645 9276 24709 9280
rect 24645 9220 24649 9276
rect 24649 9220 24705 9276
rect 24705 9220 24709 9276
rect 24645 9216 24709 9220
rect 24725 9276 24789 9280
rect 24725 9220 24729 9276
rect 24729 9220 24785 9276
rect 24785 9220 24789 9276
rect 24725 9216 24789 9220
rect 24805 9276 24869 9280
rect 24805 9220 24809 9276
rect 24809 9220 24865 9276
rect 24865 9220 24869 9276
rect 24805 9216 24869 9220
rect 10397 8732 10461 8736
rect 10397 8676 10401 8732
rect 10401 8676 10457 8732
rect 10457 8676 10461 8732
rect 10397 8672 10461 8676
rect 10477 8732 10541 8736
rect 10477 8676 10481 8732
rect 10481 8676 10537 8732
rect 10537 8676 10541 8732
rect 10477 8672 10541 8676
rect 10557 8732 10621 8736
rect 10557 8676 10561 8732
rect 10561 8676 10617 8732
rect 10617 8676 10621 8732
rect 10557 8672 10621 8676
rect 10637 8732 10701 8736
rect 10637 8676 10641 8732
rect 10641 8676 10697 8732
rect 10697 8676 10701 8732
rect 10637 8672 10701 8676
rect 19842 8732 19906 8736
rect 19842 8676 19846 8732
rect 19846 8676 19902 8732
rect 19902 8676 19906 8732
rect 19842 8672 19906 8676
rect 19922 8732 19986 8736
rect 19922 8676 19926 8732
rect 19926 8676 19982 8732
rect 19982 8676 19986 8732
rect 19922 8672 19986 8676
rect 20002 8732 20066 8736
rect 20002 8676 20006 8732
rect 20006 8676 20062 8732
rect 20062 8676 20066 8732
rect 20002 8672 20066 8676
rect 20082 8732 20146 8736
rect 20082 8676 20086 8732
rect 20086 8676 20142 8732
rect 20142 8676 20146 8732
rect 20082 8672 20146 8676
rect 5674 8188 5738 8192
rect 5674 8132 5678 8188
rect 5678 8132 5734 8188
rect 5734 8132 5738 8188
rect 5674 8128 5738 8132
rect 5754 8188 5818 8192
rect 5754 8132 5758 8188
rect 5758 8132 5814 8188
rect 5814 8132 5818 8188
rect 5754 8128 5818 8132
rect 5834 8188 5898 8192
rect 5834 8132 5838 8188
rect 5838 8132 5894 8188
rect 5894 8132 5898 8188
rect 5834 8128 5898 8132
rect 5914 8188 5978 8192
rect 5914 8132 5918 8188
rect 5918 8132 5974 8188
rect 5974 8132 5978 8188
rect 5914 8128 5978 8132
rect 15120 8188 15184 8192
rect 15120 8132 15124 8188
rect 15124 8132 15180 8188
rect 15180 8132 15184 8188
rect 15120 8128 15184 8132
rect 15200 8188 15264 8192
rect 15200 8132 15204 8188
rect 15204 8132 15260 8188
rect 15260 8132 15264 8188
rect 15200 8128 15264 8132
rect 15280 8188 15344 8192
rect 15280 8132 15284 8188
rect 15284 8132 15340 8188
rect 15340 8132 15344 8188
rect 15280 8128 15344 8132
rect 15360 8188 15424 8192
rect 15360 8132 15364 8188
rect 15364 8132 15420 8188
rect 15420 8132 15424 8188
rect 15360 8128 15424 8132
rect 24565 8188 24629 8192
rect 24565 8132 24569 8188
rect 24569 8132 24625 8188
rect 24625 8132 24629 8188
rect 24565 8128 24629 8132
rect 24645 8188 24709 8192
rect 24645 8132 24649 8188
rect 24649 8132 24705 8188
rect 24705 8132 24709 8188
rect 24645 8128 24709 8132
rect 24725 8188 24789 8192
rect 24725 8132 24729 8188
rect 24729 8132 24785 8188
rect 24785 8132 24789 8188
rect 24725 8128 24789 8132
rect 24805 8188 24869 8192
rect 24805 8132 24809 8188
rect 24809 8132 24865 8188
rect 24865 8132 24869 8188
rect 24805 8128 24869 8132
rect 10397 7644 10461 7648
rect 10397 7588 10401 7644
rect 10401 7588 10457 7644
rect 10457 7588 10461 7644
rect 10397 7584 10461 7588
rect 10477 7644 10541 7648
rect 10477 7588 10481 7644
rect 10481 7588 10537 7644
rect 10537 7588 10541 7644
rect 10477 7584 10541 7588
rect 10557 7644 10621 7648
rect 10557 7588 10561 7644
rect 10561 7588 10617 7644
rect 10617 7588 10621 7644
rect 10557 7584 10621 7588
rect 10637 7644 10701 7648
rect 10637 7588 10641 7644
rect 10641 7588 10697 7644
rect 10697 7588 10701 7644
rect 10637 7584 10701 7588
rect 19842 7644 19906 7648
rect 19842 7588 19846 7644
rect 19846 7588 19902 7644
rect 19902 7588 19906 7644
rect 19842 7584 19906 7588
rect 19922 7644 19986 7648
rect 19922 7588 19926 7644
rect 19926 7588 19982 7644
rect 19982 7588 19986 7644
rect 19922 7584 19986 7588
rect 20002 7644 20066 7648
rect 20002 7588 20006 7644
rect 20006 7588 20062 7644
rect 20062 7588 20066 7644
rect 20002 7584 20066 7588
rect 20082 7644 20146 7648
rect 20082 7588 20086 7644
rect 20086 7588 20142 7644
rect 20142 7588 20146 7644
rect 20082 7584 20146 7588
rect 5674 7100 5738 7104
rect 5674 7044 5678 7100
rect 5678 7044 5734 7100
rect 5734 7044 5738 7100
rect 5674 7040 5738 7044
rect 5754 7100 5818 7104
rect 5754 7044 5758 7100
rect 5758 7044 5814 7100
rect 5814 7044 5818 7100
rect 5754 7040 5818 7044
rect 5834 7100 5898 7104
rect 5834 7044 5838 7100
rect 5838 7044 5894 7100
rect 5894 7044 5898 7100
rect 5834 7040 5898 7044
rect 5914 7100 5978 7104
rect 5914 7044 5918 7100
rect 5918 7044 5974 7100
rect 5974 7044 5978 7100
rect 5914 7040 5978 7044
rect 15120 7100 15184 7104
rect 15120 7044 15124 7100
rect 15124 7044 15180 7100
rect 15180 7044 15184 7100
rect 15120 7040 15184 7044
rect 15200 7100 15264 7104
rect 15200 7044 15204 7100
rect 15204 7044 15260 7100
rect 15260 7044 15264 7100
rect 15200 7040 15264 7044
rect 15280 7100 15344 7104
rect 15280 7044 15284 7100
rect 15284 7044 15340 7100
rect 15340 7044 15344 7100
rect 15280 7040 15344 7044
rect 15360 7100 15424 7104
rect 15360 7044 15364 7100
rect 15364 7044 15420 7100
rect 15420 7044 15424 7100
rect 15360 7040 15424 7044
rect 24565 7100 24629 7104
rect 24565 7044 24569 7100
rect 24569 7044 24625 7100
rect 24625 7044 24629 7100
rect 24565 7040 24629 7044
rect 24645 7100 24709 7104
rect 24645 7044 24649 7100
rect 24649 7044 24705 7100
rect 24705 7044 24709 7100
rect 24645 7040 24709 7044
rect 24725 7100 24789 7104
rect 24725 7044 24729 7100
rect 24729 7044 24785 7100
rect 24785 7044 24789 7100
rect 24725 7040 24789 7044
rect 24805 7100 24869 7104
rect 24805 7044 24809 7100
rect 24809 7044 24865 7100
rect 24865 7044 24869 7100
rect 24805 7040 24869 7044
rect 10397 6556 10461 6560
rect 10397 6500 10401 6556
rect 10401 6500 10457 6556
rect 10457 6500 10461 6556
rect 10397 6496 10461 6500
rect 10477 6556 10541 6560
rect 10477 6500 10481 6556
rect 10481 6500 10537 6556
rect 10537 6500 10541 6556
rect 10477 6496 10541 6500
rect 10557 6556 10621 6560
rect 10557 6500 10561 6556
rect 10561 6500 10617 6556
rect 10617 6500 10621 6556
rect 10557 6496 10621 6500
rect 10637 6556 10701 6560
rect 10637 6500 10641 6556
rect 10641 6500 10697 6556
rect 10697 6500 10701 6556
rect 10637 6496 10701 6500
rect 19842 6556 19906 6560
rect 19842 6500 19846 6556
rect 19846 6500 19902 6556
rect 19902 6500 19906 6556
rect 19842 6496 19906 6500
rect 19922 6556 19986 6560
rect 19922 6500 19926 6556
rect 19926 6500 19982 6556
rect 19982 6500 19986 6556
rect 19922 6496 19986 6500
rect 20002 6556 20066 6560
rect 20002 6500 20006 6556
rect 20006 6500 20062 6556
rect 20062 6500 20066 6556
rect 20002 6496 20066 6500
rect 20082 6556 20146 6560
rect 20082 6500 20086 6556
rect 20086 6500 20142 6556
rect 20142 6500 20146 6556
rect 20082 6496 20146 6500
rect 5674 6012 5738 6016
rect 5674 5956 5678 6012
rect 5678 5956 5734 6012
rect 5734 5956 5738 6012
rect 5674 5952 5738 5956
rect 5754 6012 5818 6016
rect 5754 5956 5758 6012
rect 5758 5956 5814 6012
rect 5814 5956 5818 6012
rect 5754 5952 5818 5956
rect 5834 6012 5898 6016
rect 5834 5956 5838 6012
rect 5838 5956 5894 6012
rect 5894 5956 5898 6012
rect 5834 5952 5898 5956
rect 5914 6012 5978 6016
rect 5914 5956 5918 6012
rect 5918 5956 5974 6012
rect 5974 5956 5978 6012
rect 5914 5952 5978 5956
rect 15120 6012 15184 6016
rect 15120 5956 15124 6012
rect 15124 5956 15180 6012
rect 15180 5956 15184 6012
rect 15120 5952 15184 5956
rect 15200 6012 15264 6016
rect 15200 5956 15204 6012
rect 15204 5956 15260 6012
rect 15260 5956 15264 6012
rect 15200 5952 15264 5956
rect 15280 6012 15344 6016
rect 15280 5956 15284 6012
rect 15284 5956 15340 6012
rect 15340 5956 15344 6012
rect 15280 5952 15344 5956
rect 15360 6012 15424 6016
rect 15360 5956 15364 6012
rect 15364 5956 15420 6012
rect 15420 5956 15424 6012
rect 15360 5952 15424 5956
rect 24565 6012 24629 6016
rect 24565 5956 24569 6012
rect 24569 5956 24625 6012
rect 24625 5956 24629 6012
rect 24565 5952 24629 5956
rect 24645 6012 24709 6016
rect 24645 5956 24649 6012
rect 24649 5956 24705 6012
rect 24705 5956 24709 6012
rect 24645 5952 24709 5956
rect 24725 6012 24789 6016
rect 24725 5956 24729 6012
rect 24729 5956 24785 6012
rect 24785 5956 24789 6012
rect 24725 5952 24789 5956
rect 24805 6012 24869 6016
rect 24805 5956 24809 6012
rect 24809 5956 24865 6012
rect 24865 5956 24869 6012
rect 24805 5952 24869 5956
rect 10397 5468 10461 5472
rect 10397 5412 10401 5468
rect 10401 5412 10457 5468
rect 10457 5412 10461 5468
rect 10397 5408 10461 5412
rect 10477 5468 10541 5472
rect 10477 5412 10481 5468
rect 10481 5412 10537 5468
rect 10537 5412 10541 5468
rect 10477 5408 10541 5412
rect 10557 5468 10621 5472
rect 10557 5412 10561 5468
rect 10561 5412 10617 5468
rect 10617 5412 10621 5468
rect 10557 5408 10621 5412
rect 10637 5468 10701 5472
rect 10637 5412 10641 5468
rect 10641 5412 10697 5468
rect 10697 5412 10701 5468
rect 10637 5408 10701 5412
rect 19842 5468 19906 5472
rect 19842 5412 19846 5468
rect 19846 5412 19902 5468
rect 19902 5412 19906 5468
rect 19842 5408 19906 5412
rect 19922 5468 19986 5472
rect 19922 5412 19926 5468
rect 19926 5412 19982 5468
rect 19982 5412 19986 5468
rect 19922 5408 19986 5412
rect 20002 5468 20066 5472
rect 20002 5412 20006 5468
rect 20006 5412 20062 5468
rect 20062 5412 20066 5468
rect 20002 5408 20066 5412
rect 20082 5468 20146 5472
rect 20082 5412 20086 5468
rect 20086 5412 20142 5468
rect 20142 5412 20146 5468
rect 20082 5408 20146 5412
rect 5674 4924 5738 4928
rect 5674 4868 5678 4924
rect 5678 4868 5734 4924
rect 5734 4868 5738 4924
rect 5674 4864 5738 4868
rect 5754 4924 5818 4928
rect 5754 4868 5758 4924
rect 5758 4868 5814 4924
rect 5814 4868 5818 4924
rect 5754 4864 5818 4868
rect 5834 4924 5898 4928
rect 5834 4868 5838 4924
rect 5838 4868 5894 4924
rect 5894 4868 5898 4924
rect 5834 4864 5898 4868
rect 5914 4924 5978 4928
rect 5914 4868 5918 4924
rect 5918 4868 5974 4924
rect 5974 4868 5978 4924
rect 5914 4864 5978 4868
rect 15120 4924 15184 4928
rect 15120 4868 15124 4924
rect 15124 4868 15180 4924
rect 15180 4868 15184 4924
rect 15120 4864 15184 4868
rect 15200 4924 15264 4928
rect 15200 4868 15204 4924
rect 15204 4868 15260 4924
rect 15260 4868 15264 4924
rect 15200 4864 15264 4868
rect 15280 4924 15344 4928
rect 15280 4868 15284 4924
rect 15284 4868 15340 4924
rect 15340 4868 15344 4924
rect 15280 4864 15344 4868
rect 15360 4924 15424 4928
rect 15360 4868 15364 4924
rect 15364 4868 15420 4924
rect 15420 4868 15424 4924
rect 15360 4864 15424 4868
rect 24565 4924 24629 4928
rect 24565 4868 24569 4924
rect 24569 4868 24625 4924
rect 24625 4868 24629 4924
rect 24565 4864 24629 4868
rect 24645 4924 24709 4928
rect 24645 4868 24649 4924
rect 24649 4868 24705 4924
rect 24705 4868 24709 4924
rect 24645 4864 24709 4868
rect 24725 4924 24789 4928
rect 24725 4868 24729 4924
rect 24729 4868 24785 4924
rect 24785 4868 24789 4924
rect 24725 4864 24789 4868
rect 24805 4924 24869 4928
rect 24805 4868 24809 4924
rect 24809 4868 24865 4924
rect 24865 4868 24869 4924
rect 24805 4864 24869 4868
rect 10397 4380 10461 4384
rect 10397 4324 10401 4380
rect 10401 4324 10457 4380
rect 10457 4324 10461 4380
rect 10397 4320 10461 4324
rect 10477 4380 10541 4384
rect 10477 4324 10481 4380
rect 10481 4324 10537 4380
rect 10537 4324 10541 4380
rect 10477 4320 10541 4324
rect 10557 4380 10621 4384
rect 10557 4324 10561 4380
rect 10561 4324 10617 4380
rect 10617 4324 10621 4380
rect 10557 4320 10621 4324
rect 10637 4380 10701 4384
rect 10637 4324 10641 4380
rect 10641 4324 10697 4380
rect 10697 4324 10701 4380
rect 10637 4320 10701 4324
rect 19842 4380 19906 4384
rect 19842 4324 19846 4380
rect 19846 4324 19902 4380
rect 19902 4324 19906 4380
rect 19842 4320 19906 4324
rect 19922 4380 19986 4384
rect 19922 4324 19926 4380
rect 19926 4324 19982 4380
rect 19982 4324 19986 4380
rect 19922 4320 19986 4324
rect 20002 4380 20066 4384
rect 20002 4324 20006 4380
rect 20006 4324 20062 4380
rect 20062 4324 20066 4380
rect 20002 4320 20066 4324
rect 20082 4380 20146 4384
rect 20082 4324 20086 4380
rect 20086 4324 20142 4380
rect 20142 4324 20146 4380
rect 20082 4320 20146 4324
rect 5674 3836 5738 3840
rect 5674 3780 5678 3836
rect 5678 3780 5734 3836
rect 5734 3780 5738 3836
rect 5674 3776 5738 3780
rect 5754 3836 5818 3840
rect 5754 3780 5758 3836
rect 5758 3780 5814 3836
rect 5814 3780 5818 3836
rect 5754 3776 5818 3780
rect 5834 3836 5898 3840
rect 5834 3780 5838 3836
rect 5838 3780 5894 3836
rect 5894 3780 5898 3836
rect 5834 3776 5898 3780
rect 5914 3836 5978 3840
rect 5914 3780 5918 3836
rect 5918 3780 5974 3836
rect 5974 3780 5978 3836
rect 5914 3776 5978 3780
rect 15120 3836 15184 3840
rect 15120 3780 15124 3836
rect 15124 3780 15180 3836
rect 15180 3780 15184 3836
rect 15120 3776 15184 3780
rect 15200 3836 15264 3840
rect 15200 3780 15204 3836
rect 15204 3780 15260 3836
rect 15260 3780 15264 3836
rect 15200 3776 15264 3780
rect 15280 3836 15344 3840
rect 15280 3780 15284 3836
rect 15284 3780 15340 3836
rect 15340 3780 15344 3836
rect 15280 3776 15344 3780
rect 15360 3836 15424 3840
rect 15360 3780 15364 3836
rect 15364 3780 15420 3836
rect 15420 3780 15424 3836
rect 15360 3776 15424 3780
rect 24565 3836 24629 3840
rect 24565 3780 24569 3836
rect 24569 3780 24625 3836
rect 24625 3780 24629 3836
rect 24565 3776 24629 3780
rect 24645 3836 24709 3840
rect 24645 3780 24649 3836
rect 24649 3780 24705 3836
rect 24705 3780 24709 3836
rect 24645 3776 24709 3780
rect 24725 3836 24789 3840
rect 24725 3780 24729 3836
rect 24729 3780 24785 3836
rect 24785 3780 24789 3836
rect 24725 3776 24789 3780
rect 24805 3836 24869 3840
rect 24805 3780 24809 3836
rect 24809 3780 24865 3836
rect 24865 3780 24869 3836
rect 24805 3776 24869 3780
rect 19564 3436 19628 3500
rect 10397 3292 10461 3296
rect 10397 3236 10401 3292
rect 10401 3236 10457 3292
rect 10457 3236 10461 3292
rect 10397 3232 10461 3236
rect 10477 3292 10541 3296
rect 10477 3236 10481 3292
rect 10481 3236 10537 3292
rect 10537 3236 10541 3292
rect 10477 3232 10541 3236
rect 10557 3292 10621 3296
rect 10557 3236 10561 3292
rect 10561 3236 10617 3292
rect 10617 3236 10621 3292
rect 10557 3232 10621 3236
rect 10637 3292 10701 3296
rect 10637 3236 10641 3292
rect 10641 3236 10697 3292
rect 10697 3236 10701 3292
rect 10637 3232 10701 3236
rect 19842 3292 19906 3296
rect 19842 3236 19846 3292
rect 19846 3236 19902 3292
rect 19902 3236 19906 3292
rect 19842 3232 19906 3236
rect 19922 3292 19986 3296
rect 19922 3236 19926 3292
rect 19926 3236 19982 3292
rect 19982 3236 19986 3292
rect 19922 3232 19986 3236
rect 20002 3292 20066 3296
rect 20002 3236 20006 3292
rect 20006 3236 20062 3292
rect 20062 3236 20066 3292
rect 20002 3232 20066 3236
rect 20082 3292 20146 3296
rect 20082 3236 20086 3292
rect 20086 3236 20142 3292
rect 20142 3236 20146 3292
rect 20082 3232 20146 3236
rect 20300 3028 20364 3092
rect 5674 2748 5738 2752
rect 5674 2692 5678 2748
rect 5678 2692 5734 2748
rect 5734 2692 5738 2748
rect 5674 2688 5738 2692
rect 5754 2748 5818 2752
rect 5754 2692 5758 2748
rect 5758 2692 5814 2748
rect 5814 2692 5818 2748
rect 5754 2688 5818 2692
rect 5834 2748 5898 2752
rect 5834 2692 5838 2748
rect 5838 2692 5894 2748
rect 5894 2692 5898 2748
rect 5834 2688 5898 2692
rect 5914 2748 5978 2752
rect 5914 2692 5918 2748
rect 5918 2692 5974 2748
rect 5974 2692 5978 2748
rect 5914 2688 5978 2692
rect 15120 2748 15184 2752
rect 15120 2692 15124 2748
rect 15124 2692 15180 2748
rect 15180 2692 15184 2748
rect 15120 2688 15184 2692
rect 15200 2748 15264 2752
rect 15200 2692 15204 2748
rect 15204 2692 15260 2748
rect 15260 2692 15264 2748
rect 15200 2688 15264 2692
rect 15280 2748 15344 2752
rect 15280 2692 15284 2748
rect 15284 2692 15340 2748
rect 15340 2692 15344 2748
rect 15280 2688 15344 2692
rect 15360 2748 15424 2752
rect 15360 2692 15364 2748
rect 15364 2692 15420 2748
rect 15420 2692 15424 2748
rect 15360 2688 15424 2692
rect 24565 2748 24629 2752
rect 24565 2692 24569 2748
rect 24569 2692 24625 2748
rect 24625 2692 24629 2748
rect 24565 2688 24629 2692
rect 24645 2748 24709 2752
rect 24645 2692 24649 2748
rect 24649 2692 24705 2748
rect 24705 2692 24709 2748
rect 24645 2688 24709 2692
rect 24725 2748 24789 2752
rect 24725 2692 24729 2748
rect 24729 2692 24785 2748
rect 24785 2692 24789 2748
rect 24725 2688 24789 2692
rect 24805 2748 24869 2752
rect 24805 2692 24809 2748
rect 24809 2692 24865 2748
rect 24865 2692 24869 2748
rect 24805 2688 24869 2692
rect 10397 2204 10461 2208
rect 10397 2148 10401 2204
rect 10401 2148 10457 2204
rect 10457 2148 10461 2204
rect 10397 2144 10461 2148
rect 10477 2204 10541 2208
rect 10477 2148 10481 2204
rect 10481 2148 10537 2204
rect 10537 2148 10541 2204
rect 10477 2144 10541 2148
rect 10557 2204 10621 2208
rect 10557 2148 10561 2204
rect 10561 2148 10617 2204
rect 10617 2148 10621 2204
rect 10557 2144 10621 2148
rect 10637 2204 10701 2208
rect 10637 2148 10641 2204
rect 10641 2148 10697 2204
rect 10697 2148 10701 2204
rect 10637 2144 10701 2148
rect 19842 2204 19906 2208
rect 19842 2148 19846 2204
rect 19846 2148 19902 2204
rect 19902 2148 19906 2204
rect 19842 2144 19906 2148
rect 19922 2204 19986 2208
rect 19922 2148 19926 2204
rect 19926 2148 19982 2204
rect 19982 2148 19986 2204
rect 19922 2144 19986 2148
rect 20002 2204 20066 2208
rect 20002 2148 20006 2204
rect 20006 2148 20062 2204
rect 20062 2148 20066 2204
rect 20002 2144 20066 2148
rect 20082 2204 20146 2208
rect 20082 2148 20086 2204
rect 20086 2148 20142 2204
rect 20142 2148 20146 2204
rect 20082 2144 20146 2148
<< metal4 >>
rect 5666 29952 5987 30512
rect 5666 29888 5674 29952
rect 5738 29888 5754 29952
rect 5818 29888 5834 29952
rect 5898 29888 5914 29952
rect 5978 29888 5987 29952
rect 5666 28864 5987 29888
rect 5666 28800 5674 28864
rect 5738 28800 5754 28864
rect 5818 28800 5834 28864
rect 5898 28800 5914 28864
rect 5978 28800 5987 28864
rect 5666 27776 5987 28800
rect 5666 27712 5674 27776
rect 5738 27712 5754 27776
rect 5818 27712 5834 27776
rect 5898 27712 5914 27776
rect 5978 27712 5987 27776
rect 5666 26688 5987 27712
rect 5666 26624 5674 26688
rect 5738 26624 5754 26688
rect 5818 26624 5834 26688
rect 5898 26624 5914 26688
rect 5978 26624 5987 26688
rect 5666 25600 5987 26624
rect 5666 25536 5674 25600
rect 5738 25536 5754 25600
rect 5818 25536 5834 25600
rect 5898 25536 5914 25600
rect 5978 25536 5987 25600
rect 5666 24512 5987 25536
rect 5666 24448 5674 24512
rect 5738 24448 5754 24512
rect 5818 24448 5834 24512
rect 5898 24448 5914 24512
rect 5978 24448 5987 24512
rect 5666 23424 5987 24448
rect 5666 23360 5674 23424
rect 5738 23360 5754 23424
rect 5818 23360 5834 23424
rect 5898 23360 5914 23424
rect 5978 23360 5987 23424
rect 5666 22336 5987 23360
rect 5666 22272 5674 22336
rect 5738 22272 5754 22336
rect 5818 22272 5834 22336
rect 5898 22272 5914 22336
rect 5978 22272 5987 22336
rect 5666 21248 5987 22272
rect 5666 21184 5674 21248
rect 5738 21184 5754 21248
rect 5818 21184 5834 21248
rect 5898 21184 5914 21248
rect 5978 21184 5987 21248
rect 5666 20160 5987 21184
rect 5666 20096 5674 20160
rect 5738 20096 5754 20160
rect 5818 20096 5834 20160
rect 5898 20096 5914 20160
rect 5978 20096 5987 20160
rect 5666 19072 5987 20096
rect 5666 19008 5674 19072
rect 5738 19008 5754 19072
rect 5818 19008 5834 19072
rect 5898 19008 5914 19072
rect 5978 19008 5987 19072
rect 5666 17984 5987 19008
rect 5666 17920 5674 17984
rect 5738 17920 5754 17984
rect 5818 17920 5834 17984
rect 5898 17920 5914 17984
rect 5978 17920 5987 17984
rect 5666 16896 5987 17920
rect 5666 16832 5674 16896
rect 5738 16832 5754 16896
rect 5818 16832 5834 16896
rect 5898 16832 5914 16896
rect 5978 16832 5987 16896
rect 5666 15808 5987 16832
rect 5666 15744 5674 15808
rect 5738 15744 5754 15808
rect 5818 15744 5834 15808
rect 5898 15744 5914 15808
rect 5978 15744 5987 15808
rect 5666 14720 5987 15744
rect 5666 14656 5674 14720
rect 5738 14656 5754 14720
rect 5818 14656 5834 14720
rect 5898 14656 5914 14720
rect 5978 14656 5987 14720
rect 5666 13632 5987 14656
rect 5666 13568 5674 13632
rect 5738 13568 5754 13632
rect 5818 13568 5834 13632
rect 5898 13568 5914 13632
rect 5978 13568 5987 13632
rect 5666 12544 5987 13568
rect 5666 12480 5674 12544
rect 5738 12480 5754 12544
rect 5818 12480 5834 12544
rect 5898 12480 5914 12544
rect 5978 12480 5987 12544
rect 5666 11456 5987 12480
rect 5666 11392 5674 11456
rect 5738 11392 5754 11456
rect 5818 11392 5834 11456
rect 5898 11392 5914 11456
rect 5978 11392 5987 11456
rect 5666 10368 5987 11392
rect 5666 10304 5674 10368
rect 5738 10304 5754 10368
rect 5818 10304 5834 10368
rect 5898 10304 5914 10368
rect 5978 10304 5987 10368
rect 5666 9280 5987 10304
rect 5666 9216 5674 9280
rect 5738 9216 5754 9280
rect 5818 9216 5834 9280
rect 5898 9216 5914 9280
rect 5978 9216 5987 9280
rect 5666 8192 5987 9216
rect 5666 8128 5674 8192
rect 5738 8128 5754 8192
rect 5818 8128 5834 8192
rect 5898 8128 5914 8192
rect 5978 8128 5987 8192
rect 5666 7104 5987 8128
rect 5666 7040 5674 7104
rect 5738 7040 5754 7104
rect 5818 7040 5834 7104
rect 5898 7040 5914 7104
rect 5978 7040 5987 7104
rect 5666 6016 5987 7040
rect 5666 5952 5674 6016
rect 5738 5952 5754 6016
rect 5818 5952 5834 6016
rect 5898 5952 5914 6016
rect 5978 5952 5987 6016
rect 5666 4928 5987 5952
rect 5666 4864 5674 4928
rect 5738 4864 5754 4928
rect 5818 4864 5834 4928
rect 5898 4864 5914 4928
rect 5978 4864 5987 4928
rect 5666 3840 5987 4864
rect 5666 3776 5674 3840
rect 5738 3776 5754 3840
rect 5818 3776 5834 3840
rect 5898 3776 5914 3840
rect 5978 3776 5987 3840
rect 5666 2752 5987 3776
rect 5666 2688 5674 2752
rect 5738 2688 5754 2752
rect 5818 2688 5834 2752
rect 5898 2688 5914 2752
rect 5978 2688 5987 2752
rect 5666 2128 5987 2688
rect 10389 30496 10709 30512
rect 10389 30432 10397 30496
rect 10461 30432 10477 30496
rect 10541 30432 10557 30496
rect 10621 30432 10637 30496
rect 10701 30432 10709 30496
rect 10389 29408 10709 30432
rect 10389 29344 10397 29408
rect 10461 29344 10477 29408
rect 10541 29344 10557 29408
rect 10621 29344 10637 29408
rect 10701 29344 10709 29408
rect 10389 28320 10709 29344
rect 10389 28256 10397 28320
rect 10461 28256 10477 28320
rect 10541 28256 10557 28320
rect 10621 28256 10637 28320
rect 10701 28256 10709 28320
rect 10389 27232 10709 28256
rect 10389 27168 10397 27232
rect 10461 27168 10477 27232
rect 10541 27168 10557 27232
rect 10621 27168 10637 27232
rect 10701 27168 10709 27232
rect 10389 26144 10709 27168
rect 10389 26080 10397 26144
rect 10461 26080 10477 26144
rect 10541 26080 10557 26144
rect 10621 26080 10637 26144
rect 10701 26080 10709 26144
rect 10389 25056 10709 26080
rect 15112 29952 15432 30512
rect 15112 29888 15120 29952
rect 15184 29888 15200 29952
rect 15264 29888 15280 29952
rect 15344 29888 15360 29952
rect 15424 29888 15432 29952
rect 15112 28864 15432 29888
rect 15112 28800 15120 28864
rect 15184 28800 15200 28864
rect 15264 28800 15280 28864
rect 15344 28800 15360 28864
rect 15424 28800 15432 28864
rect 15112 27776 15432 28800
rect 15112 27712 15120 27776
rect 15184 27712 15200 27776
rect 15264 27712 15280 27776
rect 15344 27712 15360 27776
rect 15424 27712 15432 27776
rect 15112 26688 15432 27712
rect 15112 26624 15120 26688
rect 15184 26624 15200 26688
rect 15264 26624 15280 26688
rect 15344 26624 15360 26688
rect 15424 26624 15432 26688
rect 12571 25668 12637 25669
rect 12571 25604 12572 25668
rect 12636 25604 12637 25668
rect 12571 25603 12637 25604
rect 10389 24992 10397 25056
rect 10461 24992 10477 25056
rect 10541 24992 10557 25056
rect 10621 24992 10637 25056
rect 10701 24992 10709 25056
rect 10389 23968 10709 24992
rect 10389 23904 10397 23968
rect 10461 23904 10477 23968
rect 10541 23904 10557 23968
rect 10621 23904 10637 23968
rect 10701 23904 10709 23968
rect 10389 22880 10709 23904
rect 10389 22816 10397 22880
rect 10461 22816 10477 22880
rect 10541 22816 10557 22880
rect 10621 22816 10637 22880
rect 10701 22816 10709 22880
rect 10389 21792 10709 22816
rect 10389 21728 10397 21792
rect 10461 21728 10477 21792
rect 10541 21728 10557 21792
rect 10621 21728 10637 21792
rect 10701 21728 10709 21792
rect 10389 20704 10709 21728
rect 10389 20640 10397 20704
rect 10461 20640 10477 20704
rect 10541 20640 10557 20704
rect 10621 20640 10637 20704
rect 10701 20640 10709 20704
rect 10389 19616 10709 20640
rect 10389 19552 10397 19616
rect 10461 19552 10477 19616
rect 10541 19552 10557 19616
rect 10621 19552 10637 19616
rect 10701 19552 10709 19616
rect 10389 18528 10709 19552
rect 10389 18464 10397 18528
rect 10461 18464 10477 18528
rect 10541 18464 10557 18528
rect 10621 18464 10637 18528
rect 10701 18464 10709 18528
rect 10389 17440 10709 18464
rect 10389 17376 10397 17440
rect 10461 17376 10477 17440
rect 10541 17376 10557 17440
rect 10621 17376 10637 17440
rect 10701 17376 10709 17440
rect 10389 16352 10709 17376
rect 10389 16288 10397 16352
rect 10461 16288 10477 16352
rect 10541 16288 10557 16352
rect 10621 16288 10637 16352
rect 10701 16288 10709 16352
rect 10389 15264 10709 16288
rect 10389 15200 10397 15264
rect 10461 15200 10477 15264
rect 10541 15200 10557 15264
rect 10621 15200 10637 15264
rect 10701 15200 10709 15264
rect 10389 14176 10709 15200
rect 10389 14112 10397 14176
rect 10461 14112 10477 14176
rect 10541 14112 10557 14176
rect 10621 14112 10637 14176
rect 10701 14112 10709 14176
rect 10389 13088 10709 14112
rect 12574 14109 12634 25603
rect 15112 25600 15432 26624
rect 15112 25536 15120 25600
rect 15184 25536 15200 25600
rect 15264 25536 15280 25600
rect 15344 25536 15360 25600
rect 15424 25536 15432 25600
rect 15112 24512 15432 25536
rect 19834 30496 20154 30512
rect 19834 30432 19842 30496
rect 19906 30432 19922 30496
rect 19986 30432 20002 30496
rect 20066 30432 20082 30496
rect 20146 30432 20154 30496
rect 19834 29408 20154 30432
rect 19834 29344 19842 29408
rect 19906 29344 19922 29408
rect 19986 29344 20002 29408
rect 20066 29344 20082 29408
rect 20146 29344 20154 29408
rect 19834 28320 20154 29344
rect 19834 28256 19842 28320
rect 19906 28256 19922 28320
rect 19986 28256 20002 28320
rect 20066 28256 20082 28320
rect 20146 28256 20154 28320
rect 19834 27232 20154 28256
rect 19834 27168 19842 27232
rect 19906 27168 19922 27232
rect 19986 27168 20002 27232
rect 20066 27168 20082 27232
rect 20146 27168 20154 27232
rect 19834 26144 20154 27168
rect 19834 26080 19842 26144
rect 19906 26080 19922 26144
rect 19986 26080 20002 26144
rect 20066 26080 20082 26144
rect 20146 26080 20154 26144
rect 19379 25124 19445 25125
rect 19379 25060 19380 25124
rect 19444 25060 19445 25124
rect 19379 25059 19445 25060
rect 15112 24448 15120 24512
rect 15184 24448 15200 24512
rect 15264 24448 15280 24512
rect 15344 24448 15360 24512
rect 15424 24448 15432 24512
rect 15112 23424 15432 24448
rect 15112 23360 15120 23424
rect 15184 23360 15200 23424
rect 15264 23360 15280 23424
rect 15344 23360 15360 23424
rect 15424 23360 15432 23424
rect 15112 22336 15432 23360
rect 15112 22272 15120 22336
rect 15184 22272 15200 22336
rect 15264 22272 15280 22336
rect 15344 22272 15360 22336
rect 15424 22272 15432 22336
rect 15112 21248 15432 22272
rect 15112 21184 15120 21248
rect 15184 21184 15200 21248
rect 15264 21184 15280 21248
rect 15344 21184 15360 21248
rect 15424 21184 15432 21248
rect 15112 20160 15432 21184
rect 15112 20096 15120 20160
rect 15184 20096 15200 20160
rect 15264 20096 15280 20160
rect 15344 20096 15360 20160
rect 15424 20096 15432 20160
rect 15112 19072 15432 20096
rect 15112 19008 15120 19072
rect 15184 19008 15200 19072
rect 15264 19008 15280 19072
rect 15344 19008 15360 19072
rect 15424 19008 15432 19072
rect 15112 17984 15432 19008
rect 15112 17920 15120 17984
rect 15184 17920 15200 17984
rect 15264 17920 15280 17984
rect 15344 17920 15360 17984
rect 15424 17920 15432 17984
rect 15112 16896 15432 17920
rect 19382 17917 19442 25059
rect 19834 25056 20154 26080
rect 19834 24992 19842 25056
rect 19906 24992 19922 25056
rect 19986 24992 20002 25056
rect 20066 24992 20082 25056
rect 20146 24992 20154 25056
rect 19834 23968 20154 24992
rect 19834 23904 19842 23968
rect 19906 23904 19922 23968
rect 19986 23904 20002 23968
rect 20066 23904 20082 23968
rect 20146 23904 20154 23968
rect 19834 22880 20154 23904
rect 19834 22816 19842 22880
rect 19906 22816 19922 22880
rect 19986 22816 20002 22880
rect 20066 22816 20082 22880
rect 20146 22816 20154 22880
rect 19563 21996 19629 21997
rect 19563 21932 19564 21996
rect 19628 21932 19629 21996
rect 19563 21931 19629 21932
rect 19379 17916 19445 17917
rect 19379 17852 19380 17916
rect 19444 17852 19445 17916
rect 19379 17851 19445 17852
rect 15112 16832 15120 16896
rect 15184 16832 15200 16896
rect 15264 16832 15280 16896
rect 15344 16832 15360 16896
rect 15424 16832 15432 16896
rect 15112 15808 15432 16832
rect 15112 15744 15120 15808
rect 15184 15744 15200 15808
rect 15264 15744 15280 15808
rect 15344 15744 15360 15808
rect 15424 15744 15432 15808
rect 15112 14720 15432 15744
rect 15112 14656 15120 14720
rect 15184 14656 15200 14720
rect 15264 14656 15280 14720
rect 15344 14656 15360 14720
rect 15424 14656 15432 14720
rect 12571 14108 12637 14109
rect 12571 14044 12572 14108
rect 12636 14044 12637 14108
rect 12571 14043 12637 14044
rect 10389 13024 10397 13088
rect 10461 13024 10477 13088
rect 10541 13024 10557 13088
rect 10621 13024 10637 13088
rect 10701 13024 10709 13088
rect 10389 12000 10709 13024
rect 10389 11936 10397 12000
rect 10461 11936 10477 12000
rect 10541 11936 10557 12000
rect 10621 11936 10637 12000
rect 10701 11936 10709 12000
rect 10389 10912 10709 11936
rect 10389 10848 10397 10912
rect 10461 10848 10477 10912
rect 10541 10848 10557 10912
rect 10621 10848 10637 10912
rect 10701 10848 10709 10912
rect 10389 9824 10709 10848
rect 10389 9760 10397 9824
rect 10461 9760 10477 9824
rect 10541 9760 10557 9824
rect 10621 9760 10637 9824
rect 10701 9760 10709 9824
rect 10389 8736 10709 9760
rect 10389 8672 10397 8736
rect 10461 8672 10477 8736
rect 10541 8672 10557 8736
rect 10621 8672 10637 8736
rect 10701 8672 10709 8736
rect 10389 7648 10709 8672
rect 10389 7584 10397 7648
rect 10461 7584 10477 7648
rect 10541 7584 10557 7648
rect 10621 7584 10637 7648
rect 10701 7584 10709 7648
rect 10389 6560 10709 7584
rect 10389 6496 10397 6560
rect 10461 6496 10477 6560
rect 10541 6496 10557 6560
rect 10621 6496 10637 6560
rect 10701 6496 10709 6560
rect 10389 5472 10709 6496
rect 10389 5408 10397 5472
rect 10461 5408 10477 5472
rect 10541 5408 10557 5472
rect 10621 5408 10637 5472
rect 10701 5408 10709 5472
rect 10389 4384 10709 5408
rect 10389 4320 10397 4384
rect 10461 4320 10477 4384
rect 10541 4320 10557 4384
rect 10621 4320 10637 4384
rect 10701 4320 10709 4384
rect 10389 3296 10709 4320
rect 10389 3232 10397 3296
rect 10461 3232 10477 3296
rect 10541 3232 10557 3296
rect 10621 3232 10637 3296
rect 10701 3232 10709 3296
rect 10389 2208 10709 3232
rect 10389 2144 10397 2208
rect 10461 2144 10477 2208
rect 10541 2144 10557 2208
rect 10621 2144 10637 2208
rect 10701 2144 10709 2208
rect 10389 2128 10709 2144
rect 15112 13632 15432 14656
rect 15112 13568 15120 13632
rect 15184 13568 15200 13632
rect 15264 13568 15280 13632
rect 15344 13568 15360 13632
rect 15424 13568 15432 13632
rect 15112 12544 15432 13568
rect 15112 12480 15120 12544
rect 15184 12480 15200 12544
rect 15264 12480 15280 12544
rect 15344 12480 15360 12544
rect 15424 12480 15432 12544
rect 15112 11456 15432 12480
rect 15112 11392 15120 11456
rect 15184 11392 15200 11456
rect 15264 11392 15280 11456
rect 15344 11392 15360 11456
rect 15424 11392 15432 11456
rect 15112 10368 15432 11392
rect 15112 10304 15120 10368
rect 15184 10304 15200 10368
rect 15264 10304 15280 10368
rect 15344 10304 15360 10368
rect 15424 10304 15432 10368
rect 15112 9280 15432 10304
rect 15112 9216 15120 9280
rect 15184 9216 15200 9280
rect 15264 9216 15280 9280
rect 15344 9216 15360 9280
rect 15424 9216 15432 9280
rect 15112 8192 15432 9216
rect 15112 8128 15120 8192
rect 15184 8128 15200 8192
rect 15264 8128 15280 8192
rect 15344 8128 15360 8192
rect 15424 8128 15432 8192
rect 15112 7104 15432 8128
rect 15112 7040 15120 7104
rect 15184 7040 15200 7104
rect 15264 7040 15280 7104
rect 15344 7040 15360 7104
rect 15424 7040 15432 7104
rect 15112 6016 15432 7040
rect 15112 5952 15120 6016
rect 15184 5952 15200 6016
rect 15264 5952 15280 6016
rect 15344 5952 15360 6016
rect 15424 5952 15432 6016
rect 15112 4928 15432 5952
rect 15112 4864 15120 4928
rect 15184 4864 15200 4928
rect 15264 4864 15280 4928
rect 15344 4864 15360 4928
rect 15424 4864 15432 4928
rect 15112 3840 15432 4864
rect 15112 3776 15120 3840
rect 15184 3776 15200 3840
rect 15264 3776 15280 3840
rect 15344 3776 15360 3840
rect 15424 3776 15432 3840
rect 15112 2752 15432 3776
rect 19566 3501 19626 21931
rect 19834 21792 20154 22816
rect 19834 21728 19842 21792
rect 19906 21728 19922 21792
rect 19986 21728 20002 21792
rect 20066 21728 20082 21792
rect 20146 21728 20154 21792
rect 19834 20704 20154 21728
rect 19834 20640 19842 20704
rect 19906 20640 19922 20704
rect 19986 20640 20002 20704
rect 20066 20640 20082 20704
rect 20146 20640 20154 20704
rect 19834 19616 20154 20640
rect 24557 29952 24877 30512
rect 24557 29888 24565 29952
rect 24629 29888 24645 29952
rect 24709 29888 24725 29952
rect 24789 29888 24805 29952
rect 24869 29888 24877 29952
rect 24557 28864 24877 29888
rect 24557 28800 24565 28864
rect 24629 28800 24645 28864
rect 24709 28800 24725 28864
rect 24789 28800 24805 28864
rect 24869 28800 24877 28864
rect 24557 27776 24877 28800
rect 24557 27712 24565 27776
rect 24629 27712 24645 27776
rect 24709 27712 24725 27776
rect 24789 27712 24805 27776
rect 24869 27712 24877 27776
rect 24557 26688 24877 27712
rect 24557 26624 24565 26688
rect 24629 26624 24645 26688
rect 24709 26624 24725 26688
rect 24789 26624 24805 26688
rect 24869 26624 24877 26688
rect 24557 25600 24877 26624
rect 24557 25536 24565 25600
rect 24629 25536 24645 25600
rect 24709 25536 24725 25600
rect 24789 25536 24805 25600
rect 24869 25536 24877 25600
rect 24557 24512 24877 25536
rect 24557 24448 24565 24512
rect 24629 24448 24645 24512
rect 24709 24448 24725 24512
rect 24789 24448 24805 24512
rect 24869 24448 24877 24512
rect 24557 23424 24877 24448
rect 24557 23360 24565 23424
rect 24629 23360 24645 23424
rect 24709 23360 24725 23424
rect 24789 23360 24805 23424
rect 24869 23360 24877 23424
rect 24557 22336 24877 23360
rect 24557 22272 24565 22336
rect 24629 22272 24645 22336
rect 24709 22272 24725 22336
rect 24789 22272 24805 22336
rect 24869 22272 24877 22336
rect 24557 21248 24877 22272
rect 24557 21184 24565 21248
rect 24629 21184 24645 21248
rect 24709 21184 24725 21248
rect 24789 21184 24805 21248
rect 24869 21184 24877 21248
rect 24557 20160 24877 21184
rect 24557 20096 24565 20160
rect 24629 20096 24645 20160
rect 24709 20096 24725 20160
rect 24789 20096 24805 20160
rect 24869 20096 24877 20160
rect 20299 19684 20365 19685
rect 20299 19620 20300 19684
rect 20364 19620 20365 19684
rect 20299 19619 20365 19620
rect 19834 19552 19842 19616
rect 19906 19552 19922 19616
rect 19986 19552 20002 19616
rect 20066 19552 20082 19616
rect 20146 19552 20154 19616
rect 19834 18528 20154 19552
rect 19834 18464 19842 18528
rect 19906 18464 19922 18528
rect 19986 18464 20002 18528
rect 20066 18464 20082 18528
rect 20146 18464 20154 18528
rect 19834 17440 20154 18464
rect 19834 17376 19842 17440
rect 19906 17376 19922 17440
rect 19986 17376 20002 17440
rect 20066 17376 20082 17440
rect 20146 17376 20154 17440
rect 19834 16352 20154 17376
rect 19834 16288 19842 16352
rect 19906 16288 19922 16352
rect 19986 16288 20002 16352
rect 20066 16288 20082 16352
rect 20146 16288 20154 16352
rect 19834 15264 20154 16288
rect 19834 15200 19842 15264
rect 19906 15200 19922 15264
rect 19986 15200 20002 15264
rect 20066 15200 20082 15264
rect 20146 15200 20154 15264
rect 19834 14176 20154 15200
rect 19834 14112 19842 14176
rect 19906 14112 19922 14176
rect 19986 14112 20002 14176
rect 20066 14112 20082 14176
rect 20146 14112 20154 14176
rect 19834 13088 20154 14112
rect 19834 13024 19842 13088
rect 19906 13024 19922 13088
rect 19986 13024 20002 13088
rect 20066 13024 20082 13088
rect 20146 13024 20154 13088
rect 19834 12000 20154 13024
rect 19834 11936 19842 12000
rect 19906 11936 19922 12000
rect 19986 11936 20002 12000
rect 20066 11936 20082 12000
rect 20146 11936 20154 12000
rect 19834 10912 20154 11936
rect 19834 10848 19842 10912
rect 19906 10848 19922 10912
rect 19986 10848 20002 10912
rect 20066 10848 20082 10912
rect 20146 10848 20154 10912
rect 19834 9824 20154 10848
rect 19834 9760 19842 9824
rect 19906 9760 19922 9824
rect 19986 9760 20002 9824
rect 20066 9760 20082 9824
rect 20146 9760 20154 9824
rect 19834 8736 20154 9760
rect 19834 8672 19842 8736
rect 19906 8672 19922 8736
rect 19986 8672 20002 8736
rect 20066 8672 20082 8736
rect 20146 8672 20154 8736
rect 19834 7648 20154 8672
rect 19834 7584 19842 7648
rect 19906 7584 19922 7648
rect 19986 7584 20002 7648
rect 20066 7584 20082 7648
rect 20146 7584 20154 7648
rect 19834 6560 20154 7584
rect 19834 6496 19842 6560
rect 19906 6496 19922 6560
rect 19986 6496 20002 6560
rect 20066 6496 20082 6560
rect 20146 6496 20154 6560
rect 19834 5472 20154 6496
rect 19834 5408 19842 5472
rect 19906 5408 19922 5472
rect 19986 5408 20002 5472
rect 20066 5408 20082 5472
rect 20146 5408 20154 5472
rect 19834 4384 20154 5408
rect 19834 4320 19842 4384
rect 19906 4320 19922 4384
rect 19986 4320 20002 4384
rect 20066 4320 20082 4384
rect 20146 4320 20154 4384
rect 19563 3500 19629 3501
rect 19563 3436 19564 3500
rect 19628 3436 19629 3500
rect 19563 3435 19629 3436
rect 15112 2688 15120 2752
rect 15184 2688 15200 2752
rect 15264 2688 15280 2752
rect 15344 2688 15360 2752
rect 15424 2688 15432 2752
rect 15112 2128 15432 2688
rect 19834 3296 20154 4320
rect 19834 3232 19842 3296
rect 19906 3232 19922 3296
rect 19986 3232 20002 3296
rect 20066 3232 20082 3296
rect 20146 3232 20154 3296
rect 19834 2208 20154 3232
rect 20302 3093 20362 19619
rect 24557 19072 24877 20096
rect 24557 19008 24565 19072
rect 24629 19008 24645 19072
rect 24709 19008 24725 19072
rect 24789 19008 24805 19072
rect 24869 19008 24877 19072
rect 24557 17984 24877 19008
rect 24557 17920 24565 17984
rect 24629 17920 24645 17984
rect 24709 17920 24725 17984
rect 24789 17920 24805 17984
rect 24869 17920 24877 17984
rect 24557 16896 24877 17920
rect 24557 16832 24565 16896
rect 24629 16832 24645 16896
rect 24709 16832 24725 16896
rect 24789 16832 24805 16896
rect 24869 16832 24877 16896
rect 24557 15808 24877 16832
rect 24557 15744 24565 15808
rect 24629 15744 24645 15808
rect 24709 15744 24725 15808
rect 24789 15744 24805 15808
rect 24869 15744 24877 15808
rect 24557 14720 24877 15744
rect 24557 14656 24565 14720
rect 24629 14656 24645 14720
rect 24709 14656 24725 14720
rect 24789 14656 24805 14720
rect 24869 14656 24877 14720
rect 24557 13632 24877 14656
rect 24557 13568 24565 13632
rect 24629 13568 24645 13632
rect 24709 13568 24725 13632
rect 24789 13568 24805 13632
rect 24869 13568 24877 13632
rect 24557 12544 24877 13568
rect 24557 12480 24565 12544
rect 24629 12480 24645 12544
rect 24709 12480 24725 12544
rect 24789 12480 24805 12544
rect 24869 12480 24877 12544
rect 24557 11456 24877 12480
rect 24557 11392 24565 11456
rect 24629 11392 24645 11456
rect 24709 11392 24725 11456
rect 24789 11392 24805 11456
rect 24869 11392 24877 11456
rect 24557 10368 24877 11392
rect 24557 10304 24565 10368
rect 24629 10304 24645 10368
rect 24709 10304 24725 10368
rect 24789 10304 24805 10368
rect 24869 10304 24877 10368
rect 24557 9280 24877 10304
rect 24557 9216 24565 9280
rect 24629 9216 24645 9280
rect 24709 9216 24725 9280
rect 24789 9216 24805 9280
rect 24869 9216 24877 9280
rect 24557 8192 24877 9216
rect 24557 8128 24565 8192
rect 24629 8128 24645 8192
rect 24709 8128 24725 8192
rect 24789 8128 24805 8192
rect 24869 8128 24877 8192
rect 24557 7104 24877 8128
rect 24557 7040 24565 7104
rect 24629 7040 24645 7104
rect 24709 7040 24725 7104
rect 24789 7040 24805 7104
rect 24869 7040 24877 7104
rect 24557 6016 24877 7040
rect 24557 5952 24565 6016
rect 24629 5952 24645 6016
rect 24709 5952 24725 6016
rect 24789 5952 24805 6016
rect 24869 5952 24877 6016
rect 24557 4928 24877 5952
rect 24557 4864 24565 4928
rect 24629 4864 24645 4928
rect 24709 4864 24725 4928
rect 24789 4864 24805 4928
rect 24869 4864 24877 4928
rect 24557 3840 24877 4864
rect 24557 3776 24565 3840
rect 24629 3776 24645 3840
rect 24709 3776 24725 3840
rect 24789 3776 24805 3840
rect 24869 3776 24877 3840
rect 20299 3092 20365 3093
rect 20299 3028 20300 3092
rect 20364 3028 20365 3092
rect 20299 3027 20365 3028
rect 19834 2144 19842 2208
rect 19906 2144 19922 2208
rect 19986 2144 20002 2208
rect 20066 2144 20082 2208
rect 20146 2144 20154 2208
rect 19834 2128 20154 2144
rect 24557 2752 24877 3776
rect 24557 2688 24565 2752
rect 24629 2688 24645 2752
rect 24709 2688 24725 2752
rect 24789 2688 24805 2752
rect 24869 2688 24877 2752
rect 24557 2128 24877 2688
use sky130_fd_sc_hd__decap_12  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1639504043
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 2852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1639504043
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1639504043
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1630_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 2944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1639504043
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1639504043
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1639504043
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_23
timestamp 1639504043
transform 1 0 3220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_35
timestamp 1639504043
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1639504043
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1639504043
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1639504043
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1639504043
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1639504043
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1639504043
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1639504043
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1639504043
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1639504043
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_76
timestamp 1639504043
transform 1 0 8096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_84 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1639504043
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1499_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1632_
timestamp 1639504043
transform 1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101
timestamp 1639504043
transform 1 0 10396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1639504043
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1639504043
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1639504043
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1732_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 9568 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 9292 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1733_
timestamp 1639504043
transform 1 0 11684 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1493_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 11684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1639504043
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1639504043
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1639504043
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1734_
timestamp 1639504043
transform -1 0 13708 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1494_
timestamp 1639504043
transform -1 0 12788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_127
timestamp 1639504043
transform 1 0 12788 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_121
timestamp 1639504043
transform 1 0 12236 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_129
timestamp 1639504043
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__A
timestamp 1639504043
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1639504043
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_146
timestamp 1639504043
transform 1 0 14536 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1639504043
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1487_
timestamp 1639504043
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1488_
timestamp 1639504043
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1768_
timestamp 1639504043
transform 1 0 13708 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_0_158
timestamp 1639504043
transform 1 0 15640 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1639504043
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1639504043
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_154
timestamp 1639504043
transform 1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1639504043
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1639504043
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1639504043
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 16008 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1766_
timestamp 1639504043
transform 1 0 16652 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_0_180
timestamp 1639504043
transform 1 0 17664 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1639504043
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1639504043
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 17664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1767_
timestamp 1639504043
transform -1 0 19780 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1639504043
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1639504043
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_203
timestamp 1639504043
transform 1 0 19780 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1746_
timestamp 1639504043
transform 1 0 19872 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_2  _1440_
timestamp 1639504043
transform 1 0 21804 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1639504043
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1639504043
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1639504043
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1639504043
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1639504043
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1445_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 23184 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_0_238
timestamp 1639504043
transform 1 0 23000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_230
timestamp 1639504043
transform 1 0 22264 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1748_
timestamp 1639504043
transform 1 0 21896 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1639504043
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_246
timestamp 1639504043
transform 1 0 23736 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1639504043
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1441_
timestamp 1639504043
transform -1 0 23736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1444_
timestamp 1639504043
transform 1 0 23828 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1749_
timestamp 1639504043
transform 1 0 23828 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1691_
timestamp 1639504043
transform 1 0 25392 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _1447_
timestamp 1639504043
transform 1 0 25852 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1446_
timestamp 1639504043
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_265
timestamp 1639504043
transform 1 0 25484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1449_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 26220 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1639504043
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1639504043
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1639504043
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1639504043
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1639504043
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1639504043
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1639504043
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1639504043
transform -1 0 29440 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1639504043
transform -1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1639504043
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1639504043
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1639504043
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1639504043
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1639504043
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1639504043
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1639504043
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1639504043
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 1639504043
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_61
timestamp 1639504043
transform 1 0 6716 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1555_
timestamp 1639504043
transform 1 0 6440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 1639504043
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1639504043
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1639504043
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1639504043
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__A
timestamp 1639504043
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1639504043
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1639504043
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 10488 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1497_
timestamp 1639504043
transform -1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1498_
timestamp 1639504043
transform -1 0 10120 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_110
timestamp 1639504043
transform 1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1491_
timestamp 1639504043
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1769_
timestamp 1639504043
transform 1 0 11500 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1639504043
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1639504043
transform 1 0 14352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1639504043
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1486_
timestamp 1639504043
transform 1 0 14720 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1489_
timestamp 1639504043
transform -1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_163
timestamp 1639504043
transform 1 0 16100 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 16100 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1480_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 17756 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1736_
timestamp 1639504043
transform -1 0 17020 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_184
timestamp 1639504043
transform 1 0 18032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1639504043
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1639504043
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1246_
timestamp 1639504043
transform -1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1735_
timestamp 1639504043
transform -1 0 18952 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_214
timestamp 1639504043
transform 1 0 20792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_2  _1250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 21160 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1747_
timestamp 1639504043
transform 1 0 19228 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_2_234
timestamp 1639504043
transform 1 0 22632 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _1442_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 22632 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1692_
timestamp 1639504043
transform 1 0 23184 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1639504043
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1639504043
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1443_
timestamp 1639504043
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_265
timestamp 1639504043
transform 1 0 25484 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_273
timestamp 1639504043
transform 1 0 26220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_279
timestamp 1639504043
transform 1 0 26772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1448_
timestamp 1639504043
transform 1 0 26496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_291
timestamp 1639504043
transform 1 0 27876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_303
timestamp 1639504043
transform 1 0 28980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1639504043
transform -1 0 29440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1639504043
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1639504043
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1639504043
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1639504043
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1761_
timestamp 1639504043
transform -1 0 6256 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1639504043
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1719_
timestamp 1639504043
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1719__S
timestamp 1639504043
transform -1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_74
timestamp 1639504043
transform 1 0 7912 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_82
timestamp 1639504043
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1554_
timestamp 1639504043
transform -1 0 7728 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1731_
timestamp 1639504043
transform 1 0 8924 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1639504043
transform 1 0 9752 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1495_
timestamp 1639504043
transform -1 0 11316 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__A
timestamp 1639504043
transform 1 0 12604 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1639504043
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1639504043
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp 1639504043
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1639504043
transform 1 0 12420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_127
timestamp 1639504043
transform 1 0 12788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1639504043
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1492_
timestamp 1639504043
transform -1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_138
timestamp 1639504043
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_150
timestamp 1639504043
transform 1 0 14904 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1241_
timestamp 1639504043
transform -1 0 15548 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1242_
timestamp 1639504043
transform -1 0 13800 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_3_157
timestamp 1639504043
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1639504043
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_174
timestamp 1639504043
transform 1 0 17112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1639504043
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 17112 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_3_178
timestamp 1639504043
transform 1 0 17480 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1639504043
transform 1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1481_
timestamp 1639504043
transform 1 0 17572 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1482_
timestamp 1639504043
transform -1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1484_
timestamp 1639504043
transform -1 0 18676 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1485_
timestamp 1639504043
transform -1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_197
timestamp 1639504043
transform 1 0 19228 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_218
timestamp 1639504043
transform 1 0 21160 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 1639504043
transform 1 0 20332 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1639504043
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1639504043
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_237
timestamp 1639504043
transform 1 0 22908 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1639504043
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1251_
timestamp 1639504043
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_248
timestamp 1639504043
transform 1 0 23920 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_254
timestamp 1639504043
transform 1 0 24472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1234_
timestamp 1639504043
transform -1 0 23920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1750_
timestamp 1639504043
transform 1 0 24564 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_3_272
timestamp 1639504043
transform 1 0 26128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1639504043
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _1450_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 26956 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1451_
timestamp 1639504043
transform 1 0 26404 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_3_286
timestamp 1639504043
transform 1 0 27416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_298
timestamp 1639504043
transform 1 0 28520 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_304
timestamp 1639504043
transform 1 0 29072 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1639504043
transform -1 0 29440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1634__A
timestamp 1639504043
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1639504043
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_9
timestamp 1639504043
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1639504043
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1634_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1639504043
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1639504043
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1759_
timestamp 1639504043
transform 1 0 3772 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1720__S
timestamp 1639504043
transform 1 0 6992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_46
timestamp 1639504043
transform 1 0 5336 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_52
timestamp 1639504043
transform 1 0 5888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_56
timestamp 1639504043
transform 1 0 6256 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1553_
timestamp 1639504043
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1639504043
transform 1 0 7176 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_78
timestamp 1639504043
transform 1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1639504043
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1504_
timestamp 1639504043
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1771_
timestamp 1639504043
transform 1 0 8924 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__a21bo_2  _1501_
timestamp 1639504043
transform 1 0 10488 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1639504043
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_126
timestamp 1639504043
transform 1 0 12696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1239_
timestamp 1639504043
transform 1 0 11224 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1510_
timestamp 1639504043
transform 1 0 12236 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1517_
timestamp 1639504043
transform -1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1639504043
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1639504043
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_147
timestamp 1639504043
transform 1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_151
timestamp 1639504043
transform 1 0 14996 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1639504043
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1248_
timestamp 1639504043
transform 1 0 15088 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1490_
timestamp 1639504043
transform -1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1514_
timestamp 1639504043
transform 1 0 14168 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1776_
timestamp 1639504043
transform -1 0 17296 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_4_176
timestamp 1639504043
transform 1 0 17296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_182
timestamp 1639504043
transform 1 0 17848 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1639504043
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1639504043
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1249_
timestamp 1639504043
transform -1 0 17848 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1639504043
transform 1 0 20056 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_214
timestamp 1639504043
transform 1 0 20792 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1658_
timestamp 1639504043
transform 1 0 20976 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1659_
timestamp 1639504043
transform 1 0 19228 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_225
timestamp 1639504043
transform 1 0 21804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1639504043
transform 1 0 22908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1252_
timestamp 1639504043
transform -1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1589_
timestamp 1639504043
transform 1 0 21896 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1590_
timestamp 1639504043
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1639504043
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_262
timestamp 1639504043
transform 1 0 25208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1639504043
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1661_
timestamp 1639504043
transform -1 0 24104 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1662_
timestamp 1639504043
transform -1 0 25208 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1688_
timestamp 1639504043
transform 1 0 26404 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1690_
timestamp 1639504043
transform 1 0 25576 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_291
timestamp 1639504043
transform 1 0 27876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_303
timestamp 1639504043
transform 1 0 28980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1639504043
transform -1 0 29440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1452_
timestamp 1639504043
transform -1 0 27876 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_5_15
timestamp 1639504043
transform 1 0 2484 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_19
timestamp 1639504043
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1639504043
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1639504043
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1539_
timestamp 1639504043
transform -1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1721__S
timestamp 1639504043
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 1639504043
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1544_
timestamp 1639504043
transform -1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1721_
timestamp 1639504043
transform 1 0 3864 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_44
timestamp 1639504043
transform 1 0 5152 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_50
timestamp 1639504043
transform 1 0 5704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp 1639504043
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1639504043
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1545_
timestamp 1639504043
transform 1 0 5796 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1549_
timestamp 1639504043
transform 1 0 6624 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__A
timestamp 1639504043
transform 1 0 8648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1639504043
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1503_
timestamp 1639504043
transform -1 0 9384 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1550_
timestamp 1639504043
transform -1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1720_
timestamp 1639504043
transform -1 0 8004 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_102
timestamp 1639504043
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_90
timestamp 1639504043
transform 1 0 9384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_94
timestamp 1639504043
transform 1 0 9752 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1500_
timestamp 1639504043
transform -1 0 11132 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1502_
timestamp 1639504043
transform -1 0 9752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1509_
timestamp 1639504043
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1639504043
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1506_
timestamp 1639504043
transform 1 0 11500 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 12144 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1728_
timestamp 1639504043
transform 1 0 12788 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_136
timestamp 1639504043
transform 1 0 13616 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_146
timestamp 1639504043
transform 1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__nor4_2  _1243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 15640 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_2  _1515_
timestamp 1639504043
transform 1 0 13800 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_158
timestamp 1639504043
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1639504043
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1639504043
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_2  _1244_
timestamp 1639504043
transform -1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__A1
timestamp 1639504043
transform 1 0 19044 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_190
timestamp 1639504043
transform 1 0 18584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_194
timestamp 1639504043
transform 1 0 18952 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1245_
timestamp 1639504043
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1726_
timestamp 1639504043
transform 1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__A
timestamp 1639504043
transform 1 0 20884 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_209
timestamp 1639504043
transform 1 0 20332 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1639504043
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1594_
timestamp 1639504043
transform 1 0 20056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1595_
timestamp 1639504043
transform -1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 1639504043
transform -1 0 20056 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1639504043
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1639504043
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o22ai_2  _1593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 21804 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1682_
timestamp 1639504043
transform 1 0 22724 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1237_
timestamp 1639504043
transform -1 0 24472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1253_
timestamp 1639504043
transform 1 0 23552 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_2  _1609_
timestamp 1639504043
transform 1 0 24472 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1639504043
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1639504043
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_2  _1454_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 26956 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1608_
timestamp 1639504043
transform -1 0 26496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1673_
timestamp 1639504043
transform 1 0 25392 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1639504043
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1639504043
transform -1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1453_
timestamp 1639504043
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1639504043
transform 1 0 2116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1639504043
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1639504043
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1639504043
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1639504043
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1537_
timestamp 1639504043
transform -1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1538_
timestamp 1639504043
transform -1 0 3588 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1722_
timestamp 1639504043
transform 1 0 2208 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1758_
timestamp 1639504043
transform 1 0 1472 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1639504043
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_24
timestamp 1639504043
transform 1 0 3312 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1639504043
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1722__S
timestamp 1639504043
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__and2_2  _1543_
timestamp 1639504043
transform 1 0 3956 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _1541_
timestamp 1639504043
transform -1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1540_
timestamp 1639504043
transform 1 0 4600 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_7_32
timestamp 1639504043
transform 1 0 4048 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_37
timestamp 1639504043
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1542_
timestamp 1639504043
transform -1 0 5336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_43
timestamp 1639504043
transform 1 0 5060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1639504043
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_63
timestamp 1639504043
transform 1 0 6900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1639504043
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1169_
timestamp 1639504043
transform -1 0 6072 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1546_
timestamp 1639504043
transform -1 0 6808 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1547_
timestamp 1639504043
transform 1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1551_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _1552_
timestamp 1639504043
transform -1 0 6072 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1760_
timestamp 1639504043
transform -1 0 8648 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1639504043
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1639504043
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_75
timestamp 1639504043
transform 1 0 8004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_83
timestamp 1639504043
transform 1 0 8740 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1639504043
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1513_
timestamp 1639504043
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1773_
timestamp 1639504043
transform 1 0 9108 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1639504043
transform 1 0 10120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1639504043
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1729_
timestamp 1639504043
transform 1 0 9292 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1508_
timestamp 1639504043
transform -1 0 12144 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1507_
timestamp 1639504043
transform 1 0 12144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1505_
timestamp 1639504043
transform 1 0 11224 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1639504043
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1639504043
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1518_
timestamp 1639504043
transform 1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1639504043
transform 1 0 12420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_127
timestamp 1639504043
transform 1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1774_
timestamp 1639504043
transform 1 0 12604 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_6_115
timestamp 1639504043
transform 1 0 11684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_132
timestamp 1639504043
transform 1 0 13248 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1639504043
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1639504043
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1639504043
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1516_
timestamp 1639504043
transform -1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1519_
timestamp 1639504043
transform 1 0 14628 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1775_
timestamp 1639504043
transform 1 0 14168 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_6_157
timestamp 1639504043
transform 1 0 15548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_169
timestamp 1639504043
transform 1 0 16652 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1639504043
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp 1639504043
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1639504043
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1520_
timestamp 1639504043
transform -1 0 15548 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1521_
timestamp 1639504043
transform -1 0 16192 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1681_
timestamp 1639504043
transform -1 0 18492 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1522_
timestamp 1639504043
transform -1 0 17848 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_7_177
timestamp 1639504043
transform 1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1639504043
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _1598_
timestamp 1639504043
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1478_
timestamp 1639504043
transform -1 0 18584 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1477_
timestamp 1639504043
transform 1 0 18492 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_186
timestamp 1639504043
transform 1 0 18216 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1639504043
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_195
timestamp 1639504043
transform 1 0 19044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1597_
timestamp 1639504043
transform -1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_205
timestamp 1639504043
transform 1 0 19964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_201
timestamp 1639504043
transform 1 0 19596 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1596_
timestamp 1639504043
transform 1 0 20332 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1591_
timestamp 1639504043
transform 1 0 20608 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1475_
timestamp 1639504043
transform -1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1474_
timestamp 1639504043
transform 1 0 20792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1639504043
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_211
timestamp 1639504043
transform 1 0 20516 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_2  _1599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1660_
timestamp 1639504043
transform 1 0 22080 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1584_
timestamp 1639504043
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1483_
timestamp 1639504043
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1639504043
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1639504043
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1639504043
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_226
timestamp 1639504043
transform 1 0 21896 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1695_
timestamp 1639504043
transform 1 0 22908 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1600_
timestamp 1639504043
transform 1 0 22356 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_6_236
timestamp 1639504043
transform 1 0 22816 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_230
timestamp 1639504043
transform 1 0 22264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1238_
timestamp 1639504043
transform -1 0 24196 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_246
timestamp 1639504043
transform 1 0 23736 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_244
timestamp 1639504043
transform 1 0 23552 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1663_
timestamp 1639504043
transform -1 0 25208 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1254_
timestamp 1639504043
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1639504043
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_252
timestamp 1639504043
transform 1 0 24288 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_256
timestamp 1639504043
transform 1 0 24656 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1639504043
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1236_
timestamp 1639504043
transform -1 0 25484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_262
timestamp 1639504043
transform 1 0 25208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_268
timestamp 1639504043
transform 1 0 25760 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_280
timestamp 1639504043
transform 1 0 26864 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 1639504043
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1639504043
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1639504043
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1607_
timestamp 1639504043
transform 1 0 25300 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 1639504043
transform 1 0 25484 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_292
timestamp 1639504043
transform 1 0 27968 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_304
timestamp 1639504043
transform 1 0 29072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1639504043
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1639504043
transform -1 0 29440 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1639504043
transform -1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1723__S
timestamp 1639504043
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_18
timestamp 1639504043
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1639504043
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1639504043
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1639504043
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1534_
timestamp 1639504043
transform -1 0 2576 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1639504043
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_37
timestamp 1639504043
transform 1 0 4508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1639504043
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1170_
timestamp 1639504043
transform 1 0 4692 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1536_
timestamp 1639504043
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1718__S
timestamp 1639504043
transform 1 0 6808 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_44
timestamp 1639504043
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_56
timestamp 1639504043
transform 1 0 6256 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _1556_
timestamp 1639504043
transform 1 0 5520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1762_
timestamp 1639504043
transform -1 0 8556 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__A
timestamp 1639504043
transform 1 0 9016 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1639504043
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1639504043
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1639504043
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_94
timestamp 1639504043
transform 1 0 9752 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1512_
timestamp 1639504043
transform -1 0 9752 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1772_
timestamp 1639504043
transform -1 0 12052 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_8_128
timestamp 1639504043
transform 1 0 12880 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1730_
timestamp 1639504043
transform 1 0 12052 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1639504043
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1639504043
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1727_
timestamp 1639504043
transform 1 0 14444 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1639504043
transform 1 0 15272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1655_
timestamp 1639504043
transform 1 0 17112 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1753_
timestamp 1639504043
transform -1 0 17112 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_8_183
timestamp 1639504043
transform 1 0 17940 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1639504043
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1639504043
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1639504043
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1439_
timestamp 1639504043
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1694__A1
timestamp 1639504043
transform 1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_203
timestamp 1639504043
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_217
timestamp 1639504043
transform 1 0 21068 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1581_
timestamp 1639504043
transform -1 0 19780 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1694_
timestamp 1639504043
transform 1 0 20240 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_238
timestamp 1639504043
transform 1 0 23000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _1235_
timestamp 1639504043
transform 1 0 23092 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1592_
timestamp 1639504043
transform 1 0 21344 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_2  _1602_
timestamp 1639504043
transform 1 0 21896 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp 1639504043
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1639504043
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1639504043
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o22ai_2  _1612_
timestamp 1639504043
transform 1 0 24564 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _1610_
timestamp 1639504043
transform 1 0 25484 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1751_
timestamp 1639504043
transform 1 0 25944 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_8_287
timestamp 1639504043
transform 1 0 27508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_299
timestamp 1639504043
transform 1 0 28612 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1639504043
transform -1 0 29440 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_19
timestamp 1639504043
transform 1 0 2852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1639504043
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1639504043
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1531_
timestamp 1639504043
transform 1 0 2944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1532_
timestamp 1639504043
transform -1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1723_
timestamp 1639504043
transform 1 0 1748 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1168_
timestamp 1639504043
transform 1 0 4324 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1175_
timestamp 1639504043
transform -1 0 4324 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1530_
timestamp 1639504043
transform 1 0 4876 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_9_46
timestamp 1639504043
transform 1 0 5336 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_52
timestamp 1639504043
transform 1 0 5888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1639504043
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1639504043
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1557_
timestamp 1639504043
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1558_
timestamp 1639504043
transform 1 0 6440 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1718_
timestamp 1639504043
transform -1 0 7820 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp 1639504043
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1807_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 9936 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_9_104
timestamp 1639504043
transform 1 0 10672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_96
timestamp 1639504043
transform 1 0 9936 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 10856 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1639504043
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1639504043
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1639504043
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1887_
timestamp 1639504043
transform 1 0 12236 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_9_142
timestamp 1639504043
transform 1 0 14168 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1639504043
transform 1 0 15272 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1639504043
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1639504043
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1639504043
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1639504043
transform 1 0 18492 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__or3_2  _1228_
timestamp 1639504043
transform 1 0 18676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1230_
timestamp 1639504043
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1231_
timestamp 1639504043
transform 1 0 18032 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 17480 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1222_
timestamp 1639504043
transform -1 0 19504 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_2  _1585_
timestamp 1639504043
transform 1 0 19504 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1693_
timestamp 1639504043
transform 1 0 20608 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1639504043
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_225
timestamp 1639504043
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_233
timestamp 1639504043
transform 1 0 22540 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1639504043
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _1601_
timestamp 1639504043
transform -1 0 22540 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_2  _1606_
timestamp 1639504043
transform 1 0 23092 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_9_249
timestamp 1639504043
transform 1 0 24012 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_258
timestamp 1639504043
transform 1 0 24840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1603_
timestamp 1639504043
transform 1 0 24104 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1604_
timestamp 1639504043
transform 1 0 24564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_266
timestamp 1639504043
transform 1 0 25576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_271
timestamp 1639504043
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1639504043
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1639504043
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1639504043
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1611_
timestamp 1639504043
transform 1 0 25760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1639504043
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1639504043
transform -1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1639504043
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1639504043
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1639504043
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1757_
timestamp 1639504043
transform 1 0 1472 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1639504043
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1639504043
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1639504043
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1763_
timestamp 1639504043
transform 1 0 3864 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_10_59
timestamp 1639504043
transform 1 0 6532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1560_
timestamp 1639504043
transform 1 0 5428 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1565_
timestamp 1639504043
transform 1 0 5888 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_10_67
timestamp 1639504043
transform 1 0 7268 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1639504043
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1639504043
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1639504043
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1363_
timestamp 1639504043
transform -1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1559_
timestamp 1639504043
transform -1 0 8004 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_clk_i
timestamp 1639504043
transform -1 0 7728 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_i_A
timestamp 1639504043
transform -1 0 9568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp 1639504043
transform 1 0 9200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_92
timestamp 1639504043
transform 1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_96
timestamp 1639504043
transform 1 0 9936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1805_
timestamp 1639504043
transform 1 0 10028 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_10_118
timestamp 1639504043
transform 1 0 11960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0967_
timestamp 1639504043
transform 1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 12236 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1639504043
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B1
timestamp 1639504043
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A
timestamp 1639504043
transform 1 0 14996 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_143
timestamp 1639504043
transform 1 0 14260 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_147
timestamp 1639504043
transform 1 0 14628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1639504043
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0968_
timestamp 1639504043
transform 1 0 13248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0973_
timestamp 1639504043
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0988_
timestamp 1639504043
transform -1 0 14996 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_158
timestamp 1639504043
transform 1 0 15640 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_167
timestamp 1639504043
transform 1 0 16468 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1224_
timestamp 1639504043
transform 1 0 15916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1226_
timestamp 1639504043
transform 1 0 15180 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1227_
timestamp 1639504043
transform 1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1587_
timestamp 1639504043
transform 1 0 16652 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_10_176
timestamp 1639504043
transform 1 0 17296 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_184
timestamp 1639504043
transform 1 0 18032 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1639504043
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1639504043
transform 1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1577_
timestamp 1639504043
transform -1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1639504043
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_209
timestamp 1639504043
transform 1 0 20332 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp 1639504043
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1261_
timestamp 1639504043
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_clk_i
timestamp 1639504043
transform 1 0 20516 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1639504043
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_226
timestamp 1639504043
transform 1 0 21896 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1229_
timestamp 1639504043
transform 1 0 21620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1605_
timestamp 1639504043
transform 1 0 23000 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1639504043
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_262
timestamp 1639504043
transform 1 0 25208 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1639504043
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1646_
timestamp 1639504043
transform 1 0 24380 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_274
timestamp 1639504043
transform 1 0 26312 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_286
timestamp 1639504043
transform 1 0 27416 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_298
timestamp 1639504043
transform 1 0 28520 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_304
timestamp 1639504043
transform 1 0 29072 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1639504043
transform -1 0 29440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_14
timestamp 1639504043
transform 1 0 2392 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1639504043
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1639504043
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1535_
timestamp 1639504043
transform -1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_26
timestamp 1639504043
transform 1 0 3496 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_38
timestamp 1639504043
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_42
timestamp 1639504043
transform 1 0 4968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1561_
timestamp 1639504043
transform 1 0 5060 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1716__S
timestamp 1639504043
transform 1 0 6624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1639504043
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1171_
timestamp 1639504043
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1564_
timestamp 1639504043
transform -1 0 6624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1716_
timestamp 1639504043
transform -1 0 7636 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_71
timestamp 1639504043
transform 1 0 7636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1362_
timestamp 1639504043
transform 1 0 8740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clk_i
timestamp 1639504043
transform -1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _1364_
timestamp 1639504043
transform -1 0 10120 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1368_
timestamp 1639504043
transform 1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1369_
timestamp 1639504043
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1370_
timestamp 1639504043
transform -1 0 10856 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__B1
timestamp 1639504043
transform -1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__B1
timestamp 1639504043
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_117
timestamp 1639504043
transform 1 0 11868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1639504043
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0969_
timestamp 1639504043
transform 1 0 12052 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1885_
timestamp 1639504043
transform 1 0 12788 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__and3_2  _0987_
timestamp 1639504043
transform -1 0 15272 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1639504043
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1639504043
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1223_
timestamp 1639504043
transform 1 0 15272 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1586_
timestamp 1639504043
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1664_
timestamp 1639504043
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__B1
timestamp 1639504043
transform 1 0 19044 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_178
timestamp 1639504043
transform 1 0 17480 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_2  _1588_
timestamp 1639504043
transform 1 0 17940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_clk_i
timestamp 1639504043
transform -1 0 17940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1639504043
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1639504043
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_2  _1582_
timestamp 1639504043
transform 1 0 19228 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_233
timestamp 1639504043
transform 1 0 22540 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1639504043
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1232_
timestamp 1639504043
transform 1 0 21252 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1262_
timestamp 1639504043
transform 1 0 21804 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1580_
timestamp 1639504043
transform 1 0 22264 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_245
timestamp 1639504043
transform 1 0 23644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_251
timestamp 1639504043
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1216_
timestamp 1639504043
transform -1 0 24196 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_266
timestamp 1639504043
transform 1 0 25576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1639504043
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1639504043
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1639504043
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1255_
timestamp 1639504043
transform 1 0 25300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1639504043
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1639504043
transform -1 0 29440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_15
timestamp 1639504043
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_21
timestamp 1639504043
transform 1 0 3036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1639504043
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1639504043
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1639504043
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1639504043
transform 1 0 4048 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1639504043
transform 1 0 4784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1639504043
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1167_
timestamp 1639504043
transform 1 0 3128 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1174_
timestamp 1639504043
transform -1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1562_
timestamp 1639504043
transform -1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_44
timestamp 1639504043
transform 1 0 5152 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_52
timestamp 1639504043
transform 1 0 5888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1566_
timestamp 1639504043
transform -1 0 6716 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1764_
timestamp 1639504043
transform -1 0 8280 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_12_78
timestamp 1639504043
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1639504043
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1365_
timestamp 1639504043
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_88
timestamp 1639504043
transform 1 0 9200 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_96
timestamp 1639504043
transform 1 0 9936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1886_
timestamp 1639504043
transform -1 0 12052 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A1
timestamp 1639504043
transform -1 0 12972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__B1
timestamp 1639504043
transform 1 0 12972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_119
timestamp 1639504043
transform 1 0 12052 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_131
timestamp 1639504043
transform 1 0 13156 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A
timestamp 1639504043
transform 1 0 14996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 1639504043
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1639504043
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1639504043
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0974_
timestamp 1639504043
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__A
timestamp 1639504043
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_155
timestamp 1639504043
transform 1 0 15364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1752_
timestamp 1639504043
transform -1 0 17296 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_12_176
timestamp 1639504043
transform 1 0 17296 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1639504043
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1639504043
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1654_
timestamp 1639504043
transform 1 0 17388 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1656_
timestamp 1639504043
transform 1 0 18216 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1639504043
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_2  _1583_
timestamp 1639504043
transform 1 0 19320 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1639_
timestamp 1639504043
transform 1 0 20424 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1639504043
transform 1 0 21252 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_232
timestamp 1639504043
transform 1 0 22448 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1233_
timestamp 1639504043
transform 1 0 21344 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1256_
timestamp 1639504043
transform 1 0 21804 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _1259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 23276 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1639504043
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1639504043
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o22ai_2  _1260_
timestamp 1639504043
transform 1 0 23276 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_2  _1830_
timestamp 1639504043
transform -1 0 25944 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_12_270
timestamp 1639504043
transform 1 0 25944 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_282
timestamp 1639504043
transform 1 0 27048 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_294
timestamp 1639504043
transform 1 0 28152 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_302
timestamp 1639504043
transform 1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1639504043
transform -1 0 29440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1639504043
transform 1 0 2116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_17
timestamp 1639504043
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1639504043
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1639504043
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1639504043
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1524_
timestamp 1639504043
transform 1 0 3036 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1525_
timestamp 1639504043
transform 1 0 2944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1526_
timestamp 1639504043
transform -1 0 2668 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1756_
timestamp 1639504043
transform 1 0 1380 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1725__S
timestamp 1639504043
transform 1 0 4600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1639504043
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_40
timestamp 1639504043
transform 1 0 4784 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1639504043
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1176_
timestamp 1639504043
transform 1 0 3680 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1717_
timestamp 1639504043
transform 1 0 4324 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1725_
timestamp 1639504043
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1717__S
timestamp 1639504043
transform 1 0 5612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1639504043
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1639504043
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_48
timestamp 1639504043
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1639504043
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_2  _1172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1563_
timestamp 1639504043
transform -1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1765_
timestamp 1639504043
transform 1 0 5796 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1639504043
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1639504043
transform 1 0 7360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1639504043
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1639504043
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1366_
timestamp 1639504043
transform -1 0 9200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1567_
timestamp 1639504043
transform -1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1806_
timestamp 1639504043
transform -1 0 9752 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__B1
timestamp 1639504043
transform -1 0 10672 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_100
timestamp 1639504043
transform 1 0 10304 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_88
timestamp 1639504043
transform 1 0 9200 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _0972_
timestamp 1639504043
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1367_
timestamp 1639504043
transform -1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0971_
timestamp 1639504043
transform -1 0 12052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1639504043
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0965_
timestamp 1639504043
transform 1 0 12052 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1639504043
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_118
timestamp 1639504043
transform 1 0 11960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_114
timestamp 1639504043
transform 1 0 11592 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__B1
timestamp 1639504043
transform 1 0 11408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1639504043
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__B1
timestamp 1639504043
transform -1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1888_
timestamp 1639504043
transform -1 0 13984 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _0962_
timestamp 1639504043
transform -1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1639504043
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_137
timestamp 1639504043
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_133
timestamp 1639504043
transform 1 0 13340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__B1
timestamp 1639504043
transform -1 0 14076 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__a41o_2  _1007_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1002_
timestamp 1639504043
transform -1 0 14904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0870_
timestamp 1639504043
transform 1 0 14904 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1639504043
transform -1 0 15180 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_141
timestamp 1639504043
transform 1 0 14076 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1639504043
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 1639504043
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1639504043
transform 1 0 15456 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_168
timestamp 1639504043
transform 1 0 16560 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1639504043
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1639504043
transform -1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1220_
timestamp 1639504043
transform 1 0 15180 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1221_
timestamp 1639504043
transform 1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1687__A1
timestamp 1639504043
transform 1 0 19044 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_177
timestamp 1639504043
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1639504043
transform 1 0 17664 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1639504043
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1639504043
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1754_
timestamp 1639504043
transform 1 0 17480 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_i_A
timestamp 1639504043
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1639504043
transform 1 0 19596 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_199
timestamp 1639504043
transform 1 0 19412 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_211
timestamp 1639504043
transform 1 0 20516 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1638_
timestamp 1639504043
transform 1 0 20516 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1687_
timestamp 1639504043
transform 1 0 19688 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clk_i
timestamp 1639504043
transform -1 0 19596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1579_
timestamp 1639504043
transform -1 0 21620 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1263_
timestamp 1639504043
transform 1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1639504043
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_223
timestamp 1639504043
transform 1 0 21620 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_227
timestamp 1639504043
transform 1 0 21988 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1639504043
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A
timestamp 1639504043
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__or4_2  _1578_
timestamp 1639504043
transform -1 0 23460 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1268_
timestamp 1639504043
transform -1 0 23460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1639504043
transform 1 0 22172 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_232
timestamp 1639504043
transform 1 0 22448 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_235
timestamp 1639504043
transform 1 0 22724 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1257_
timestamp 1639504043
transform 1 0 23460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1219_
timestamp 1639504043
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1218_
timestamp 1639504043
transform 1 0 23460 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_14_248
timestamp 1639504043
transform 1 0 23920 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_246
timestamp 1639504043
transform 1 0 23736 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_2  _1265_
timestamp 1639504043
transform -1 0 25392 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _1258_
timestamp 1639504043
transform -1 0 25024 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1639504043
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_253
timestamp 1639504043
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1829_
timestamp 1639504043
transform 1 0 25024 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_13_267
timestamp 1639504043
transform 1 0 25668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1639504043
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1639504043
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1639504043
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1639504043
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1217_
timestamp 1639504043
transform -1 0 25668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1639504043
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1639504043
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_301
timestamp 1639504043
transform 1 0 28796 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1639504043
transform -1 0 29440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1639504043
transform -1 0 29440 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1639504043
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1527_
timestamp 1639504043
transform -1 0 2760 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1529_
timestamp 1639504043
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1724_
timestamp 1639504043
transform 1 0 1656 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1755_
timestamp 1639504043
transform -1 0 4324 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_15_35
timestamp 1639504043
transform 1 0 4324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_42
timestamp 1639504043
transform 1 0 4968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1177_
timestamp 1639504043
transform -1 0 4968 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1715__S
timestamp 1639504043
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_60
timestamp 1639504043
transform 1 0 6624 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1639504043
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1173_
timestamp 1639504043
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1715_
timestamp 1639504043
transform -1 0 6072 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_68
timestamp 1639504043
transform 1 0 7360 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1808_
timestamp 1639504043
transform 1 0 7544 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__B1
timestamp 1639504043
transform 1 0 10488 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_104
timestamp 1639504043
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1359_
timestamp 1639504043
transform -1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1360_
timestamp 1639504043
transform -1 0 10212 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1639504043
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1639504043
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_129
timestamp 1639504043
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1639504043
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1639504043
transform -1 0 12420 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0963_
timestamp 1639504043
transform -1 0 12696 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0964_
timestamp 1639504043
transform -1 0 12972 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_133
timestamp 1639504043
transform 1 0 13340 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1639504043
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1639504043
transform 1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0961_
timestamp 1639504043
transform -1 0 13708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1842_
timestamp 1639504043
transform 1 0 14996 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__B1
timestamp 1639504043
transform 1 0 17112 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1639504043
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 1639504043
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1639504043
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_176
timestamp 1639504043
transform 1 0 17296 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_194
timestamp 1639504043
transform 1 0 18952 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1851_
timestamp 1639504043
transform 1 0 17388 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_15_206
timestamp 1639504043
transform 1 0 20056 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1827_
timestamp 1639504043
transform 1 0 20148 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1639504043
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o22ai_2  _1269_
timestamp 1639504043
transform 1 0 22816 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1270_
timestamp 1639504043
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1271_
timestamp 1639504043
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_249
timestamp 1639504043
transform 1 0 24012 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_255
timestamp 1639504043
transform 1 0 24564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1264_
timestamp 1639504043
transform -1 0 25392 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1266_
timestamp 1639504043
transform -1 0 24012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_264
timestamp 1639504043
transform 1 0 25392 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1639504043
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1639504043
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1639504043
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1639504043
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1639504043
transform -1 0 29440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1724__S
timestamp 1639504043
transform 1 0 2484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_17
timestamp 1639504043
transform 1 0 2668 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1639504043
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1639504043
transform 1 0 1932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1639504043
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1528_
timestamp 1639504043
transform -1 0 2484 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1639504043
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_34
timestamp 1639504043
transform 1 0 4232 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1639504043
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1523_
timestamp 1639504043
transform 1 0 3772 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1533_
timestamp 1639504043
transform -1 0 5244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_45
timestamp 1639504043
transform 1 0 5244 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_52
timestamp 1639504043
transform 1 0 5888 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_60
timestamp 1639504043
transform 1 0 6624 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1193_
timestamp 1639504043
transform 1 0 6716 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1568_
timestamp 1639504043
transform 1 0 5428 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_16_70
timestamp 1639504043
transform 1 0 7544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1639504043
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1639504043
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1356_
timestamp 1639504043
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1548_
timestamp 1639504043
transform 1 0 7268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1357_
timestamp 1639504043
transform -1 0 9476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1358_
timestamp 1639504043
transform -1 0 9752 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1810_
timestamp 1639504043
transform 1 0 9752 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A1
timestamp 1639504043
transform 1 0 12880 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__B1
timestamp 1639504043
transform -1 0 13248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_115
timestamp 1639504043
transform 1 0 11684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_119
timestamp 1639504043
transform 1 0 12052 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_123
timestamp 1639504043
transform 1 0 12420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_127
timestamp 1639504043
transform 1 0 12788 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0949_
timestamp 1639504043
transform -1 0 12420 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__B1
timestamp 1639504043
transform -1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_132
timestamp 1639504043
transform 1 0 13248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_136
timestamp 1639504043
transform 1 0 13616 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_144
timestamp 1639504043
transform 1 0 14352 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1639504043
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0955_
timestamp 1639504043
transform -1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0956_
timestamp 1639504043
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1144_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1843_
timestamp 1639504043
transform 1 0 15732 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1639504043
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1639504043
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1129_
timestamp 1639504043
transform 1 0 17296 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _1130_
timestamp 1639504043
transform 1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_214
timestamp 1639504043
transform 1 0 20792 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1850_
timestamp 1639504043
transform 1 0 19228 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_16_226
timestamp 1639504043
transform 1 0 21896 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_238
timestamp 1639504043
transform 1 0 23000 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1639504043
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1639504043
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1639504043
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1639504043
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1639504043
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1639504043
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_301
timestamp 1639504043
transform 1 0 28796 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1639504043
transform -1 0 29440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_21
timestamp 1639504043
transform 1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1639504043
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1639504043
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1625_
timestamp 1639504043
transform -1 0 3036 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1671_
timestamp 1639504043
transform 1 0 1932 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_32
timestamp 1639504043
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_43
timestamp 1639504043
transform 1 0 5060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_2  _1178_
timestamp 1639504043
transform 1 0 4232 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1618_
timestamp 1639504043
transform 1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp 1639504043
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1639504043
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1191_
timestamp 1639504043
transform -1 0 5704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1793_
timestamp 1639504043
transform 1 0 6348 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_17_74
timestamp 1639504043
transform 1 0 7912 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1639504043
transform 1 0 8648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clk_i
timestamp 1639504043
transform -1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_i_A
timestamp 1639504043
transform 1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_100
timestamp 1639504043
transform 1 0 10304 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_90
timestamp 1639504043
transform 1 0 9384 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_96
timestamp 1639504043
transform 1 0 9936 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1350_
timestamp 1639504043
transform 1 0 10028 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1351_
timestamp 1639504043
transform 1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1352_
timestamp 1639504043
transform -1 0 11408 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__B1
timestamp 1639504043
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1639504043
transform 1 0 11684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1639504043
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1639504043
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0957_
timestamp 1639504043
transform 1 0 12144 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1890_
timestamp 1639504043
transform 1 0 12880 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__B1
timestamp 1639504043
transform 1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_149
timestamp 1639504043
transform 1 0 14812 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1143_
timestamp 1639504043
transform 1 0 15088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1639504043
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1639504043
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 1639504043
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1639504043
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__B1
timestamp 1639504043
transform -1 0 18400 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_188
timestamp 1639504043
transform 1 0 18400 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_196
timestamp 1639504043
transform 1 0 19136 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1678_
timestamp 1639504043
transform 1 0 17388 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_208
timestamp 1639504043
transform 1 0 20240 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_216
timestamp 1639504043
transform 1 0 20976 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1699_
timestamp 1639504043
transform 1 0 19412 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__A1
timestamp 1639504043
transform -1 0 21620 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__B1
timestamp 1639504043
transform 1 0 21252 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1639504043
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1639504043
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1409_
timestamp 1639504043
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1828_
timestamp 1639504043
transform 1 0 22540 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_17_250
timestamp 1639504043
transform 1 0 24104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1777_
timestamp 1639504043
transform 1 0 24472 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_17_271
timestamp 1639504043
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1639504043
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1639504043
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1639504043
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1639504043
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1639504043
transform -1 0 29440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_20
timestamp 1639504043
transform 1 0 2944 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1639504043
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 3036 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1742_
timestamp 1639504043
transform 1 0 1380 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 1639504043
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1639504043
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1738_
timestamp 1639504043
transform 1 0 3864 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__A
timestamp 1639504043
transform 1 0 5888 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_50
timestamp 1639504043
transform 1 0 5704 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_59
timestamp 1639504043
transform 1 0 6532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1166_
timestamp 1639504043
transform 1 0 5428 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1395_
timestamp 1639504043
transform 1 0 6072 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1639504043
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1639504043
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1837_
timestamp 1639504043
transform 1 0 7268 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106
timestamp 1639504043
transform 1 0 10856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_94
timestamp 1639504043
transform 1 0 9752 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1344_
timestamp 1639504043
transform 1 0 11040 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1353_
timestamp 1639504043
transform 1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1354_
timestamp 1639504043
transform -1 0 9752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__A1
timestamp 1639504043
transform -1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__B1
timestamp 1639504043
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_111
timestamp 1639504043
transform 1 0 11316 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_115
timestamp 1639504043
transform 1 0 11684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0947_
timestamp 1639504043
transform 1 0 12604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1342_
timestamp 1639504043
transform 1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1345_
timestamp 1639504043
transform 1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__B1
timestamp 1639504043
transform -1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_132
timestamp 1639504043
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_144
timestamp 1639504043
transform 1 0 14352 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1639504043
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0959_
timestamp 1639504043
transform -1 0 14352 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1142_
timestamp 1639504043
transform 1 0 14812 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1844_
timestamp 1639504043
transform 1 0 15640 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__B1
timestamp 1639504043
transform -1 0 17756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_175
timestamp 1639504043
transform 1 0 17204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1639504043
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1639504043
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1128_
timestamp 1639504043
transform 1 0 17756 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1639504043
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1812_
timestamp 1639504043
transform 1 0 19412 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_18_240
timestamp 1639504043
transform 1 0 23184 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1407_
timestamp 1639504043
transform -1 0 23184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1784_
timestamp 1639504043
transform -1 0 22908 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A1
timestamp 1639504043
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1639504043
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1413_
timestamp 1639504043
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1416_
timestamp 1639504043
transform 1 0 23552 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1779_
timestamp 1639504043
transform 1 0 24564 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_18_272
timestamp 1639504043
transform 1 0 26128 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_284
timestamp 1639504043
transform 1 0 27232 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_296
timestamp 1639504043
transform 1 0 28336 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_304
timestamp 1639504043
transform 1 0 29072 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1639504043
transform -1 0 29440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_18
timestamp 1639504043
transform 1 0 2760 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1639504043
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 1639504043
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1639504043
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1639504043
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1639504043
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1639504043
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1624_
timestamp 1639504043
transform -1 0 2760 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1647_
timestamp 1639504043
transform 1 0 2208 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_26
timestamp 1639504043
transform 1 0 3496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1639504043
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1639504043
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1639504043
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1639504043
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1639504043
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1667_
timestamp 1639504043
transform -1 0 4508 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_45
timestamp 1639504043
transform 1 0 5244 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1639504043
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_clk_i
timestamp 1639504043
transform -1 0 7084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1192_
timestamp 1639504043
transform -1 0 6716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1639504043
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_65
timestamp 1639504043
transform 1 0 7084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1639504043
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1639504043
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1839_
timestamp 1639504043
transform 1 0 6900 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1804_
timestamp 1639504043
transform 1 0 5336 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_19_75
timestamp 1639504043
transform 1 0 8004 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1639504043
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1639504043
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1639504043
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_2  _1194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 7268 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1809_
timestamp 1639504043
transform -1 0 10488 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1639504043
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1639504043
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1811_
timestamp 1639504043
transform -1 0 11316 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_clk_i
timestamp 1639504043
transform 1 0 10488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _1355_
timestamp 1639504043
transform -1 0 12236 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1349_
timestamp 1639504043
transform -1 0 12052 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0960_
timestamp 1639504043
transform 1 0 12144 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1639504043
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_119
timestamp 1639504043
transform 1 0 12052 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_130
timestamp 1639504043
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__B1
timestamp 1639504043
transform -1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__B1
timestamp 1639504043
transform -1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B1
timestamp 1639504043
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1889_
timestamp 1639504043
transform 1 0 12604 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__B1
timestamp 1639504043
transform -1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1639504043
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1639504043
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1639504043
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1639504043
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0958_
timestamp 1639504043
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1146_
timestamp 1639504043
transform 1 0 14812 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__B1
timestamp 1639504043
transform 1 0 17112 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1639504043
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1639504043
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1639504043
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_161
timestamp 1639504043
transform 1 0 15916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_173
timestamp 1639504043
transform 1 0 17020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1639504043
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1141_
timestamp 1639504043
transform -1 0 15916 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1639504043
transform 1 0 17388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_188
timestamp 1639504043
transform 1 0 18400 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1639504043
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1639504043
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1639504043
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1132_
timestamp 1639504043
transform -1 0 18124 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1705_
timestamp 1639504043
transform 1 0 17572 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1852_
timestamp 1639504043
transform -1 0 20056 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_clk_i
timestamp 1639504043
transform -1 0 18492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1639504043
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1639504043
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_i_A
timestamp 1639504043
transform 1 0 19872 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_clk_i
timestamp 1639504043
transform 1 0 20700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clk_i
timestamp 1639504043
transform 1 0 20056 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1341_
timestamp 1639504043
transform -1 0 20792 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_212
timestamp 1639504043
transform 1 0 20608 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_206
timestamp 1639504043
transform 1 0 20056 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1639504043
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_210
timestamp 1639504043
transform 1 0 20424 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1412_
timestamp 1639504043
transform 1 0 21068 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1410_
timestamp 1639504043
transform 1 0 21804 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1408_
timestamp 1639504043
transform -1 0 22080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1639504043
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1639504043
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1414_
timestamp 1639504043
transform 1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_232
timestamp 1639504043
transform 1 0 22448 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__B1
timestamp 1639504043
transform 1 0 22264 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A1
timestamp 1639504043
transform 1 0 22724 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__B1
timestamp 1639504043
transform 1 0 22080 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A1
timestamp 1639504043
transform 1 0 22540 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_237
timestamp 1639504043
transform 1 0 22908 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1639504043
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__A1
timestamp 1639504043
transform 1 0 23092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _1418_
timestamp 1639504043
transform 1 0 23920 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1417_
timestamp 1639504043
transform 1 0 23276 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_249
timestamp 1639504043
transform 1 0 24012 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_245
timestamp 1639504043
transform 1 0 23644 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__B1
timestamp 1639504043
transform 1 0 23736 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__B1
timestamp 1639504043
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _1415_
timestamp 1639504043
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1639504043
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__A1
timestamp 1639504043
transform 1 0 24840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__B1
timestamp 1639504043
transform 1 0 24656 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A1
timestamp 1639504043
transform 1 0 25116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_260
timestamp 1639504043
transform 1 0 25024 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__B1
timestamp 1639504043
transform 1 0 25300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1639504043
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1639504043
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1639504043
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1639504043
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1639504043
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1639504043
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1639504043
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_301
timestamp 1639504043
transform 1 0 28796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1639504043
transform -1 0 29440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1639504043
transform -1 0 29440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_11
timestamp 1639504043
transform 1 0 2116 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1639504043
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1639504043
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1462_
timestamp 1639504043
transform 1 0 2852 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _1464_
timestamp 1639504043
transform 1 0 2208 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1463_
timestamp 1639504043
transform 1 0 3312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1739_
timestamp 1639504043
transform 1 0 3588 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1639504043
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1639504043
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1639504043
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1153_
timestamp 1639504043
transform -1 0 7360 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _1457_
timestamp 1639504043
transform -1 0 5888 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A1
timestamp 1639504043
transform 1 0 7360 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_70
timestamp 1639504043
transform 1 0 7544 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1831_
timestamp 1639504043
transform 1 0 7912 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A
timestamp 1639504043
transform -1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1639504043
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_91
timestamp 1639504043
transform 1 0 9476 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1346_
timestamp 1639504043
transform -1 0 10396 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1347_
timestamp 1639504043
transform 1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1348_
timestamp 1639504043
transform -1 0 10672 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__B1
timestamp 1639504043
transform 1 0 12512 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1639504043
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_126
timestamp 1639504043
transform 1 0 12696 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1639504043
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0954_
timestamp 1639504043
transform 1 0 11776 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_132
timestamp 1639504043
transform 1 0 13248 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1639504043
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_144
timestamp 1639504043
transform 1 0 14352 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_150
timestamp 1639504043
transform 1 0 14904 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0951_
timestamp 1639504043
transform -1 0 14076 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0952_
timestamp 1639504043
transform 1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0966_
timestamp 1639504043
transform -1 0 14352 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1841_
timestamp 1639504043
transform 1 0 14996 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1639504043
transform 1 0 16928 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1639504043
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1140_
timestamp 1639504043
transform -1 0 16928 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1849_
timestamp 1639504043
transform 1 0 17112 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1635_
timestamp 1639504043
transform 1 0 18676 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1639504043
transform 1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1847_
timestamp 1639504043
transform -1 0 21252 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1639504043
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1639504043
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1639504043
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1781_
timestamp 1639504043
transform 1 0 21804 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1778_
timestamp 1639504043
transform 1 0 23368 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1780_
timestamp 1639504043
transform 1 0 24932 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1639504043
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1639504043
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1639504043
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1639504043
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1639504043
transform -1 0 29440 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1639504043
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1639504043
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1466_
timestamp 1639504043
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1639504043
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1639504043
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1639504043
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1465_
timestamp 1639504043
transform 1 0 3220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1645_
timestamp 1639504043
transform 1 0 4508 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_51
timestamp 1639504043
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1152_
timestamp 1639504043
transform -1 0 7176 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1456_
timestamp 1639504043
transform 1 0 5336 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A
timestamp 1639504043
transform 1 0 7912 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_66
timestamp 1639504043
transform 1 0 7176 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1639504043
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1639504043
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1639504043
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1215_
timestamp 1639504043
transform -1 0 8556 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A
timestamp 1639504043
transform 1 0 11040 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_104
timestamp 1639504043
transform 1 0 10672 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1639504043
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0976_
timestamp 1639504043
transform -1 0 11040 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1361_
timestamp 1639504043
transform 1 0 10396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_110
timestamp 1639504043
transform 1 0 11224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_114
timestamp 1639504043
transform 1 0 11592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1891_
timestamp 1639504043
transform -1 0 13616 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1639504043
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1639504043
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 1639504043
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1639504043
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0953_
timestamp 1639504043
transform -1 0 13892 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1145_
timestamp 1639504043
transform -1 0 15180 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1639504043
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_171
timestamp 1639504043
transform 1 0 16836 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1133_
timestamp 1639504043
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1134_
timestamp 1639504043
transform 1 0 16560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__B1
timestamp 1639504043
transform -1 0 18308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1639504043
transform 1 0 17940 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1639504043
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1126_
timestamp 1639504043
transform -1 0 17940 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1127_
timestamp 1639504043
transform 1 0 17388 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1137_
timestamp 1639504043
transform 1 0 18308 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__B1
timestamp 1639504043
transform -1 0 20240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_208
timestamp 1639504043
transform 1 0 20240 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _1136_
timestamp 1639504043
transform 1 0 19228 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__A1
timestamp 1639504043
transform 1 0 22172 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__B1
timestamp 1639504043
transform 1 0 22356 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_220
timestamp 1639504043
transform 1 0 21344 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1639504043
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _1411_
timestamp 1639504043
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1639504043
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1639504043
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_253
timestamp 1639504043
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_261
timestamp 1639504043
transform 1 0 25116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1639504043
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_267
timestamp 1639504043
transform 1 0 25668 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_279
timestamp 1639504043
transform 1 0 26772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0934_
timestamp 1639504043
transform 1 0 25392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_291
timestamp 1639504043
transform 1 0 27876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_303
timestamp 1639504043
transform 1 0 28980 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1639504043
transform -1 0 29440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1639504043
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1648_
timestamp 1639504043
transform 1 0 2944 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1743_
timestamp 1639504043
transform 1 0 1380 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_23_29
timestamp 1639504043
transform 1 0 3772 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_43
timestamp 1639504043
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1620_
timestamp 1639504043
transform -1 0 5060 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1668_
timestamp 1639504043
transform 1 0 3956 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1639504043
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1639504043
transform 1 0 6624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1639504043
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1639504043
transform -1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1737_
timestamp 1639504043
transform 1 0 6716 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1639504043
transform 1 0 7636 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_70
timestamp 1639504043
transform 1 0 7544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1149_
timestamp 1639504043
transform -1 0 9384 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1150_
timestamp 1639504043
transform 1 0 7820 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _1214_
timestamp 1639504043
transform 1 0 8372 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_102
timestamp 1639504043
transform 1 0 10488 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1639504043
transform 1 0 10856 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_90
timestamp 1639504043
transform 1 0 9384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_98
timestamp 1639504043
transform 1 0 10120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0977_
timestamp 1639504043
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1068_
timestamp 1639504043
transform 1 0 9476 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1373_
timestamp 1639504043
transform 1 0 11040 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A1
timestamp 1639504043
transform -1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1639504043
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_116
timestamp 1639504043
transform 1 0 11776 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_122
timestamp 1639504043
transform 1 0 12328 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1639504043
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0950_
timestamp 1639504043
transform 1 0 12420 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1374_
timestamp 1639504043
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1892_
timestamp 1639504043
transform 1 0 13340 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__B1
timestamp 1639504043
transform -1 0 16560 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_160
timestamp 1639504043
transform 1 0 15824 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1639504043
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0943_
timestamp 1639504043
transform -1 0 15548 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1138_
timestamp 1639504043
transform 1 0 15548 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1139_
timestamp 1639504043
transform 1 0 16652 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B1
timestamp 1639504043
transform -1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_180
timestamp 1639504043
transform 1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1848_
timestamp 1639504043
transform 1 0 17848 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_23_199
timestamp 1639504043
transform 1 0 19412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1846_
timestamp 1639504043
transform -1 0 21252 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1639504043
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1639504043
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1639504043
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_231
timestamp 1639504043
transform 1 0 22356 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1639504043
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1783_
timestamp 1639504043
transform 1 0 22448 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B1
timestamp 1639504043
transform 1 0 24288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0933_
timestamp 1639504043
transform 1 0 24472 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0942_
timestamp 1639504043
transform -1 0 24288 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1895_
timestamp 1639504043
transform 1 0 24748 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1639504043
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1639504043
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1639504043
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1639504043
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1639504043
transform -1 0 29440 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_14
timestamp 1639504043
transform 1 0 2392 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1639504043
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1639504043
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1165_
timestamp 1639504043
transform 1 0 2760 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1627_
timestamp 1639504043
transform -1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1639504043
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1639504043
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_37
timestamp 1639504043
transform 1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1639504043
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _1619_
timestamp 1639504043
transform 1 0 3864 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _1148_
timestamp 1639504043
transform -1 0 7636 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1840_
timestamp 1639504043
transform -1 0 6808 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__B
timestamp 1639504043
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1639504043
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1639504043
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1070_
timestamp 1639504043
transform -1 0 8648 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 7636 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1884_
timestamp 1639504043
transform 1 0 9016 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1803_
timestamp 1639504043
transform 1 0 10948 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 1639504043
transform 1 0 12880 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__B1
timestamp 1639504043
transform 1 0 13340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_132
timestamp 1639504043
transform 1 0 13248 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1639504043
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1639504043
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_141
timestamp 1639504043
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_150
timestamp 1639504043
transform 1 0 14904 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1639504043
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1392_
timestamp 1639504043
transform -1 0 14904 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_162
timestamp 1639504043
transform 1 0 16008 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1845_
timestamp 1639504043
transform 1 0 16100 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1639504043
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1639504043
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1124_
timestamp 1639504043
transform -1 0 18768 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1135_
timestamp 1639504043
transform 1 0 17664 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1639504043
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_205
timestamp 1639504043
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1853_
timestamp 1639504043
transform -1 0 21712 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1782_
timestamp 1639504043
transform 1 0 21712 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_24_241
timestamp 1639504043
transform 1 0 23276 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_256
timestamp 1639504043
transform 1 0 24656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1639504043
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0931_
timestamp 1639504043
transform 1 0 24748 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0932_
timestamp 1639504043
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0935_
timestamp 1639504043
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B1
timestamp 1639504043
transform 1 0 25484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_267
timestamp 1639504043
transform 1 0 25668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_279
timestamp 1639504043
transform 1 0 26772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_291
timestamp 1639504043
transform 1 0 27876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_303
timestamp 1639504043
transform 1 0 28980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1639504043
transform -1 0 29440 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1639504043
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1639504043
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1626_
timestamp 1639504043
transform -1 0 3220 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1672_
timestamp 1639504043
transform 1 0 1748 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_23
timestamp 1639504043
transform 1 0 3220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1639504043
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_36
timestamp 1639504043
transform 1 0 4416 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1179_
timestamp 1639504043
transform 1 0 3404 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1459_
timestamp 1639504043
transform 1 0 4508 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A1
timestamp 1639504043
transform 1 0 6624 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1639504043
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1639504043
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1639504043
transform 1 0 6808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1639504043
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_2  _1616_
timestamp 1639504043
transform 1 0 5244 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__C
timestamp 1639504043
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A
timestamp 1639504043
transform 1 0 7636 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1639504043
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__or3_2  _1003_
timestamp 1639504043
transform 1 0 8004 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1004_
timestamp 1639504043
transform 1 0 8556 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1076_
timestamp 1639504043
transform -1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__C1
timestamp 1639504043
transform 1 0 9568 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1639504043
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_88
timestamp 1639504043
transform 1 0 9200 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_94
timestamp 1639504043
transform 1 0 9752 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1639504043
transform -1 0 9568 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1639504043
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_125
timestamp 1639504043
transform 1 0 12604 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1639504043
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1795_
timestamp 1639504043
transform -1 0 15088 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_25_152
timestamp 1639504043
transform 1 0 15088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_156
timestamp 1639504043
transform 1 0 15456 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_160
timestamp 1639504043
transform 1 0 15824 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1639504043
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1639504043
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1639504043
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1387_
timestamp 1639504043
transform 1 0 15916 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1391_
timestamp 1639504043
transform -1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_184
timestamp 1639504043
transform 1 0 18032 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1131_
timestamp 1639504043
transform -1 0 18032 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1684_
timestamp 1639504043
transform 1 0 18952 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1702_
timestamp 1639504043
transform 1 0 18124 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__B1
timestamp 1639504043
transform -1 0 20976 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__B1
timestamp 1639504043
transform -1 0 21160 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_203
timestamp 1639504043
transform 1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1639504043
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _1125_
timestamp 1639504043
transform 1 0 19964 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1639504043
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1639504043
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1639504043
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_249
timestamp 1639504043
transform 1 0 24012 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_257
timestamp 1639504043
transform 1 0 24748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1896_
timestamp 1639504043
transform 1 0 24932 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1639504043
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1639504043
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1639504043
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1639504043
transform -1 0 29440 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1639504043
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1639504043
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1639504043
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1651_
timestamp 1639504043
transform 1 0 2208 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _1461_
timestamp 1639504043
transform 1 0 3036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1460_
timestamp 1639504043
transform -1 0 3036 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_27_11
timestamp 1639504043
transform 1 0 2116 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1639504043
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_15
timestamp 1639504043
transform 1 0 2484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1639504043
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1639504043
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1639504043
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_33
timestamp 1639504043
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_43
timestamp 1639504043
transform 1 0 5060 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1639504043
transform 1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1639504043
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1458_
timestamp 1639504043
transform -1 0 5244 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1652_
timestamp 1639504043
transform 1 0 4232 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1669_
timestamp 1639504043
transform 1 0 3772 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B2
timestamp 1639504043
transform 1 0 6900 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_65
timestamp 1639504043
transform 1 0 7084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1639504043
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1639504043
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1639504043
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_2  _1071_
timestamp 1639504043
transform 1 0 6992 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _1077_
timestamp 1639504043
transform 1 0 6348 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1874_
timestamp 1639504043
transform 1 0 5336 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_2  _1072_
timestamp 1639504043
transform 1 0 8004 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1066_
timestamp 1639504043
transform -1 0 8464 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1639504043
transform -1 0 7452 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1874__CLK
timestamp 1639504043
transform 1 0 7452 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A2
timestamp 1639504043
transform 1 0 7636 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A
timestamp 1639504043
transform -1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1639504043
transform -1 0 9384 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _1067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 9108 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1639504043
transform -1 0 8740 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1639504043
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1639504043
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1639504043
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__a221oi_2  _1075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 10120 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_106
timestamp 1639504043
transform 1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_98
timestamp 1639504043
transform 1 0 10120 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1639504043
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_2  _1467_
timestamp 1639504043
transform -1 0 12052 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_2  _1875_
timestamp 1639504043
transform 1 0 9384 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1277_
timestamp 1639504043
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1639504043
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_116
timestamp 1639504043
transform 1 0 11776 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1639504043
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_119
timestamp 1639504043
transform 1 0 12052 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1438_
timestamp 1639504043
transform -1 0 13708 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or3_2  _1428_
timestamp 1639504043
transform -1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0946_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 12328 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1639504043
transform -1 0 12788 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_127
timestamp 1639504043
transform 1 0 12788 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1639504043
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1639504043
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_150
timestamp 1639504043
transform 1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1639504043
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1639504043
transform 1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1427_
timestamp 1639504043
transform 1 0 13432 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1436_
timestamp 1639504043
transform -1 0 14904 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1797_
timestamp 1639504043
transform 1 0 15088 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 13708 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1639504043
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1639504043
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1639504043
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1013_
timestamp 1639504043
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_2  _1473_
timestamp 1639504043
transform 1 0 15548 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1119_
timestamp 1639504043
transform -1 0 17664 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1118_
timestamp 1639504043
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1117_
timestamp 1639504043
transform -1 0 18032 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1107_
timestamp 1639504043
transform 1 0 17480 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0916_
timestamp 1639504043
transform -1 0 17480 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1639504043
transform 1 0 18032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1639504043
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1120_
timestamp 1639504043
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1639504043
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1639504043
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1855_
timestamp 1639504043
transform 1 0 18216 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__B1
timestamp 1639504043
transform -1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1639504043
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_203
timestamp 1639504043
transform 1 0 19780 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_215
timestamp 1639504043
transform 1 0 20884 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1639504043
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _1121_
timestamp 1639504043
transform 1 0 19964 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1856_
timestamp 1639504043
transform -1 0 22356 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A1
timestamp 1639504043
transform 1 0 22632 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_231
timestamp 1639504043
transform 1 0 22356 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1639504043
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1639504043
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0938_
timestamp 1639504043
transform 1 0 22816 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1894_
timestamp 1639504043
transform -1 0 24472 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _0937_
timestamp 1639504043
transform -1 0 24104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0936_
timestamp 1639504043
transform 1 0 23552 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0941_
timestamp 1639504043
transform 1 0 24472 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0917_
timestamp 1639504043
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1639504043
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_256
timestamp 1639504043
transform 1 0 24656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B1
timestamp 1639504043
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0939_
timestamp 1639504043
transform 1 0 24932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_262
timestamp 1639504043
transform 1 0 25208 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_262
timestamp 1639504043
transform 1 0 25208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0940_
timestamp 1639504043
transform 1 0 25300 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0928_
timestamp 1639504043
transform 1 0 26036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0927_
timestamp 1639504043
transform 1 0 25668 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_270
timestamp 1639504043
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_270
timestamp 1639504043
transform 1 0 25944 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_266
timestamp 1639504043
transform 1 0 25576 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__B1
timestamp 1639504043
transform 1 0 25760 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A1
timestamp 1639504043
transform -1 0 25760 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1639504043
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1639504043
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1639504043
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_274
timestamp 1639504043
transform 1 0 26312 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_286
timestamp 1639504043
transform 1 0 27416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_298
timestamp 1639504043
transform 1 0 28520 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_304
timestamp 1639504043
transform 1 0 29072 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1639504043
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1639504043
transform -1 0 29440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1639504043
transform -1 0 29440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1741__CLK
timestamp 1639504043
transform 1 0 2944 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1639504043
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1741_
timestamp 1639504043
transform 1 0 1380 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_28_22
timestamp 1639504043
transform 1 0 3128 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_29
timestamp 1639504043
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1639504043
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1740_
timestamp 1639504043
transform 1 0 3864 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B1
timestamp 1639504043
transform 1 0 6992 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_47
timestamp 1639504043
transform 1 0 5428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_2  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 6164 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_28_66
timestamp 1639504043
transform 1 0 7176 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_72
timestamp 1639504043
transform 1 0 7728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1639504043
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp 1639504043
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1639504043
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1080_
timestamp 1639504043
transform 1 0 7820 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1875__CLK
timestamp 1639504043
transform 1 0 9200 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_103
timestamp 1639504043
transform 1 0 10580 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1639504043
transform 1 0 9384 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1639504043
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1639504043
transform 1 0 11132 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1083_
timestamp 1639504043
transform 1 0 9568 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1285_
timestamp 1639504043
transform 1 0 10672 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_28_112
timestamp 1639504043
transform 1 0 11408 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_127
timestamp 1639504043
transform 1 0 12788 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1014_
timestamp 1639504043
transform -1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1017_
timestamp 1639504043
transform 1 0 11500 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1278_
timestamp 1639504043
transform -1 0 12788 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1420_
timestamp 1639504043
transform 1 0 11776 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_i_A
timestamp 1639504043
transform -1 0 13708 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_134
timestamp 1639504043
transform 1 0 13432 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1639504043
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_144
timestamp 1639504043
transform 1 0 14352 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1639504043
transform 1 0 15088 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1639504043
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1639504043
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_165
timestamp 1639504043
transform 1 0 16284 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_171
timestamp 1639504043
transform 1 0 16836 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1639504043
transform -1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _0945_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 16008 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1388_
timestamp 1639504043
transform 1 0 16008 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__B1
timestamp 1639504043
transform 1 0 17848 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_178
timestamp 1639504043
transform 1 0 17480 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1639504043
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1639504043
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1122_
timestamp 1639504043
transform -1 0 18860 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1314_
timestamp 1639504043
transform 1 0 17204 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp 1639504043
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1123_
timestamp 1639504043
transform 1 0 20148 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1675_
timestamp 1639504043
transform -1 0 20148 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1854_
timestamp 1639504043
transform -1 0 22540 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_28_233
timestamp 1639504043
transform 1 0 22540 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0929_
timestamp 1639504043
transform 1 0 22908 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0930_
timestamp 1639504043
transform 1 0 23184 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_243
timestamp 1639504043
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1639504043
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1639504043
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1639504043
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1893_
timestamp 1639504043
transform 1 0 24564 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1639504043
transform 1 0 26496 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_288
timestamp 1639504043
transform 1 0 27600 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_300
timestamp 1639504043
transform 1 0 28704 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_304
timestamp 1639504043
transform 1 0 29072 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1639504043
transform -1 0 29440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_13
timestamp 1639504043
transform 1 0 2300 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1639504043
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1639504043
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1621_
timestamp 1639504043
transform -1 0 2852 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1622_
timestamp 1639504043
transform 1 0 2852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1670_
timestamp 1639504043
transform 1 0 1472 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1639504043
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1180_
timestamp 1639504043
transform -1 0 4692 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1657_
timestamp 1639504043
transform 1 0 3588 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1639504043
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1639504043
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_65
timestamp 1639504043
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1639504043
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1372_
timestamp 1639504043
transform -1 0 6072 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1873__CLK
timestamp 1639504043
transform 1 0 7360 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _1065_
timestamp 1639504043
transform 1 0 7544 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _1826_
timestamp 1639504043
transform 1 0 8004 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1826__CLK
timestamp 1639504043
transform 1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_106
timestamp 1639504043
transform 1 0 10856 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_98
timestamp 1639504043
transform 1 0 10120 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1011_
timestamp 1639504043
transform -1 0 11408 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_29_116
timestamp 1639504043
transform 1 0 11776 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_131
timestamp 1639504043
transform 1 0 13156 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1639504043
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1274_
timestamp 1639504043
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_2  _1424_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 13156 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_144
timestamp 1639504043
transform 1 0 14352 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1423_
timestamp 1639504043
transform -1 0 15364 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_2  _1437_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 13432 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1639504043
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1639504043
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0871_
timestamp 1639504043
transform 1 0 15364 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0910_
timestamp 1639504043
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_175
timestamp 1639504043
transform 1 0 17204 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_187
timestamp 1639504043
transform 1 0 18308 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1639504043
transform 1 0 18952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1115_
timestamp 1639504043
transform 1 0 18676 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__B1
timestamp 1639504043
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_207
timestamp 1639504043
transform 1 0 20148 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1639504043
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1696_
timestamp 1639504043
transform 1 0 19320 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1639504043
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1639504043
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_233
timestamp 1639504043
transform 1 0 22540 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 1639504043
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1639504043
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1639504043
transform 1 0 22632 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1898_
timestamp 1639504043
transform 1 0 23092 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_29_260
timestamp 1639504043
transform 1 0 25024 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1639504043
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1639504043
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1639504043
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1639504043
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1639504043
transform -1 0 29440 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1623__A2
timestamp 1639504043
transform 1 0 2668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_19
timestamp 1639504043
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1639504043
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1639504043
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1639504043
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _1623_
timestamp 1639504043
transform 1 0 1840 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1622__B1
timestamp 1639504043
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1639504043
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_31
timestamp 1639504043
transform 1 0 3956 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_43
timestamp 1639504043
transform 1 0 5060 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1639504043
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1639504043
transform 1 0 5152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _1082_
timestamp 1639504043
transform 1 0 5336 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1873_
timestamp 1639504043
transform 1 0 5796 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1639504043
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1639504043
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1639504043
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1639504043
transform -1 0 8464 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_2  _1081_
timestamp 1639504043
transform 1 0 7360 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_104
timestamp 1639504043
transform 1 0 10672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1639504043
transform 1 0 10396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1281_
timestamp 1639504043
transform 1 0 10856 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_2  _1282_
timestamp 1639504043
transform 1 0 9476 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__A2
timestamp 1639504043
transform 1 0 12328 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1639504043
transform 1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_2  _1279_
timestamp 1639504043
transform 1 0 11500 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_2  _1430_
timestamp 1639504043
transform 1 0 12512 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_136
timestamp 1639504043
transform 1 0 13616 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp 1639504043
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1639504043
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1639504043
transform -1 0 15272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1275_
timestamp 1639504043
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1425_
timestamp 1639504043
transform 1 0 14168 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0872_
timestamp 1639504043
transform -1 0 15548 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1426_
timestamp 1639504043
transform 1 0 15548 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dfrtp_2  _1796_
timestamp 1639504043
transform 1 0 16468 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_30_188
timestamp 1639504043
transform 1 0 18400 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1639504043
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1108_
timestamp 1639504043
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_clk_i
timestamp 1639504043
transform -1 0 18860 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _1116_
timestamp 1639504043
transform 1 0 20056 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1700_
timestamp 1639504043
transform -1 0 20056 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1857_
timestamp 1639504043
transform 1 0 20884 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_30_232
timestamp 1639504043
transform 1 0 22448 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0913_
timestamp 1639504043
transform -1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0923_
timestamp 1639504043
transform 1 0 22816 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A1
timestamp 1639504043
transform -1 0 24012 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__B1
timestamp 1639504043
transform -1 0 24196 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1639504043
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_253
timestamp 1639504043
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_262
timestamp 1639504043
transform 1 0 25208 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1639504043
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0911_
timestamp 1639504043
transform 1 0 23552 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0921_
timestamp 1639504043
transform 1 0 24656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0922_
timestamp 1639504043
transform -1 0 25208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_266
timestamp 1639504043
transform 1 0 25576 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_271
timestamp 1639504043
transform 1 0 26036 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_283
timestamp 1639504043
transform 1 0 27140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0918_
timestamp 1639504043
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0919_
timestamp 1639504043
transform 1 0 25760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_295
timestamp 1639504043
transform 1 0 28244 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_303
timestamp 1639504043
transform 1 0 28980 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1639504043
transform -1 0 29440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_11
timestamp 1639504043
transform 1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1639504043
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1639504043
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1653_
timestamp 1639504043
transform 1 0 2392 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_23
timestamp 1639504043
transform 1 0 3220 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_31
timestamp 1639504043
transform 1 0 3956 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1614_
timestamp 1639504043
transform -1 0 5612 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1644_
timestamp 1639504043
transform -1 0 4876 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1614__B2
timestamp 1639504043
transform 1 0 5612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1639504043
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1639504043
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_60
timestamp 1639504043
transform 1 0 6624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1639504043
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1455_
timestamp 1639504043
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_72
timestamp 1639504043
transform 1 0 7728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_79
timestamp 1639504043
transform 1 0 8372 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_84
timestamp 1639504043
transform 1 0 8832 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1272_
timestamp 1639504043
transform 1 0 8096 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1273_
timestamp 1639504043
transform 1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1639504043
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_2  _1286_
timestamp 1639504043
transform 1 0 10580 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1343_
timestamp 1639504043
transform -1 0 10580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_116
timestamp 1639504043
transform 1 0 11776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_121
timestamp 1639504043
transform 1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1639504043
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1276_
timestamp 1639504043
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1419_
timestamp 1639504043
transform -1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _1429_
timestamp 1639504043
transform -1 0 13340 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_31_133
timestamp 1639504043
transform 1 0 13340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1639504043
transform 1 0 14444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_150
timestamp 1639504043
transform 1 0 14904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1422_
timestamp 1639504043
transform -1 0 14904 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1639504043
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_172
timestamp 1639504043
transform 1 0 16928 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1639504043
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1389_
timestamp 1639504043
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1390_
timestamp 1639504043
transform 1 0 17112 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_177
timestamp 1639504043
transform 1 0 17388 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_184
timestamp 1639504043
transform 1 0 18032 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_196
timestamp 1639504043
transform 1 0 19136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1639504043
transform 1 0 17756 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1636_
timestamp 1639504043
transform 1 0 18308 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _1114_
timestamp 1639504043
transform 1 0 19320 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1858_
timestamp 1639504043
transform 1 0 20148 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1639504043
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1639504043
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1639504043
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_249
timestamp 1639504043
transform 1 0 24012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_253
timestamp 1639504043
transform 1 0 24380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0924_
timestamp 1639504043
transform 1 0 24472 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1899_
timestamp 1639504043
transform 1 0 24748 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1639504043
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1639504043
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1639504043
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1639504043
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1639504043
transform -1 0 29440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1639504043
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1639504043
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _1182_
timestamp 1639504043
transform 1 0 2760 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1189_
timestamp 1639504043
transform -1 0 2760 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1639504043
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1639504043
transform 1 0 4048 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_36
timestamp 1639504043
transform 1 0 4416 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1639504043
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1639504043
transform -1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 1639504043
transform -1 0 5336 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__A
timestamp 1639504043
transform 1 0 6256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_46
timestamp 1639504043
transform 1 0 5336 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_54
timestamp 1639504043
transform 1 0 6072 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_63
timestamp 1639504043
transform 1 0 6900 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1371_
timestamp 1639504043
transform -1 0 6900 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1825__CLK
timestamp 1639504043
transform 1 0 9016 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_71
timestamp 1639504043
transform 1 0 7636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_75
timestamp 1639504043
transform 1 0 8004 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1639504043
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1639504043
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1639504043
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1283_
timestamp 1639504043
transform 1 0 7728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_clk_i
timestamp 1639504043
transform -1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_100
timestamp 1639504043
transform 1 0 10304 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_88
timestamp 1639504043
transform 1 0 9200 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _1015_
timestamp 1639504043
transform -1 0 11684 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_115
timestamp 1639504043
transform 1 0 11684 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_123
timestamp 1639504043
transform 1 0 12420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_130
timestamp 1639504043
transform 1 0 13064 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1009_
timestamp 1639504043
transform -1 0 13064 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1280_
timestamp 1639504043
transform -1 0 13616 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1639504043
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1639504043
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1639504043
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_152
timestamp 1639504043
transform 1 0 15088 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1639504043
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1434_
timestamp 1639504043
transform 1 0 14536 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_161
timestamp 1639504043
transform 1 0 15916 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_172
timestamp 1639504043
transform 1 0 16928 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0909_
timestamp 1639504043
transform -1 0 16928 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1471_
timestamp 1639504043
transform 1 0 15364 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_32_180
timestamp 1639504043
transform 1 0 17664 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1639504043
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1639504043
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1639504043
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1085_
timestamp 1639504043
transform 1 0 17940 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1087_
timestamp 1639504043
transform 1 0 18216 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B1
timestamp 1639504043
transform -1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1639504043
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1639504043
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1639504043
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B1
timestamp 1639504043
transform 1 0 22448 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_221
timestamp 1639504043
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0907_
timestamp 1639504043
transform 1 0 22172 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0914_
timestamp 1639504043
transform 1 0 22632 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__B1
timestamp 1639504043
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_242
timestamp 1639504043
transform 1 0 23368 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_255
timestamp 1639504043
transform 1 0 24564 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_262
timestamp 1639504043
transform 1 0 25208 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1639504043
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0920_
timestamp 1639504043
transform 1 0 23552 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0925_
timestamp 1639504043
transform 1 0 24932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_274
timestamp 1639504043
transform 1 0 26312 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_286
timestamp 1639504043
transform 1 0 27416 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_298
timestamp 1639504043
transform 1 0 28520 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_304
timestamp 1639504043
transform 1 0 29072 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1639504043
transform -1 0 29440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__B1
timestamp 1639504043
transform 1 0 1656 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_17
timestamp 1639504043
transform 1 0 2668 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1639504043
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1639504043
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1639504043
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1405_
timestamp 1639504043
transform -1 0 3404 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _1406_
timestamp 1639504043
transform 1 0 1840 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1785_
timestamp 1639504043
transform -1 0 2944 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_33_32
timestamp 1639504043
transform 1 0 4048 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_37
timestamp 1639504043
transform 1 0 4508 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1639504043
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1156_
timestamp 1639504043
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_
timestamp 1639504043
transform -1 0 4508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _1615_
timestamp 1639504043
transform -1 0 4600 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1666_
timestamp 1639504043
transform -1 0 5428 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1674_
timestamp 1639504043
transform -1 0 4048 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1744_
timestamp 1639504043
transform 1 0 4692 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A
timestamp 1639504043
transform 1 0 6624 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_52
timestamp 1639504043
transform 1 0 5888 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_64
timestamp 1639504043
transform 1 0 6992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1639504043
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1639504043
transform -1 0 6624 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1639504043
transform 1 0 6808 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1613_
timestamp 1639504043
transform 1 0 5428 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _1825_
timestamp 1639504043
transform 1 0 7084 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _1288_
timestamp 1639504043
transform -1 0 7820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1284_
timestamp 1639504043
transform 1 0 7912 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0980_
timestamp 1639504043
transform 1 0 7176 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_73
timestamp 1639504043
transform 1 0 7820 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_69
timestamp 1639504043
transform 1 0 7452 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1639504043
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_85
timestamp 1639504043
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1639504043
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1639504043
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _1287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 9016 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__B
timestamp 1639504043
transform 1 0 9660 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_107
timestamp 1639504043
transform 1 0 10948 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_107
timestamp 1639504043
transform 1 0 10948 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_95
timestamp 1639504043
transform 1 0 9844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1639504043
transform 1 0 10672 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1021_
timestamp 1639504043
transform 1 0 9200 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1569_
timestamp 1639504043
transform -1 0 11316 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1649_
timestamp 1639504043
transform 1 0 9844 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1639504043
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_119
timestamp 1639504043
transform 1 0 12052 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_131
timestamp 1639504043
transform 1 0 13156 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1639504043
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1008_
timestamp 1639504043
transform 1 0 12604 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _1019_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 12604 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o2111ai_2  _1026_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_2  _1575_
timestamp 1639504043
transform 1 0 13708 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1018_
timestamp 1639504043
transform 1 0 13616 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1639504043
transform -1 0 13616 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1639504043
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1639504043
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1639504043
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1639504043
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_2  _1433_
timestamp 1639504043
transform 1 0 14536 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1016_
timestamp 1639504043
transform -1 0 14904 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_34_150
timestamp 1639504043
transform 1 0 14904 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__o22ai_2  _1472_
timestamp 1639504043
transform 1 0 15548 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _1309_
timestamp 1639504043
transform 1 0 16100 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1308_
timestamp 1639504043
transform 1 0 15272 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_162
timestamp 1639504043
transform 1 0 16008 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_153
timestamp 1639504043
transform 1 0 15180 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0873_
timestamp 1639504043
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1639504043
transform -1 0 16836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1639504043
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_171
timestamp 1639504043
transform 1 0 16836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1639504043
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1706_
timestamp 1639504043
transform 1 0 17296 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1679_
timestamp 1639504043
transform 1 0 17296 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_175
timestamp 1639504043
transform 1 0 17204 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_175
timestamp 1639504043
transform 1 0 17204 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1113_
timestamp 1639504043
transform 1 0 18308 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1111_
timestamp 1639504043
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1110_
timestamp 1639504043
transform 1 0 18584 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_189
timestamp 1639504043
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_185
timestamp 1639504043
transform 1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__B1
timestamp 1639504043
transform 1 0 18124 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1639504043
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_196
timestamp 1639504043
transform 1 0 19136 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__B1
timestamp 1639504043
transform -1 0 20792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_202
timestamp 1639504043
transform 1 0 19688 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_214
timestamp 1639504043
transform 1 0 20792 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _1112_
timestamp 1639504043
transform 1 0 19780 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1859_
timestamp 1639504043
transform -1 0 20792 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1860_
timestamp 1639504043
transform -1 0 22356 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__B1
timestamp 1639504043
transform 1 0 23000 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__B1
timestamp 1639504043
transform 1 0 23184 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1639504043
transform 1 0 22632 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1639504043
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0906_
timestamp 1639504043
transform -1 0 22632 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1900_
timestamp 1639504043
transform -1 0 23736 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_clk_i
timestamp 1639504043
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A1
timestamp 1639504043
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_246
timestamp 1639504043
transform 1 0 23736 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1639504043
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1639504043
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0926_
timestamp 1639504043
transform 1 0 23368 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1897_
timestamp 1639504043
transform 1 0 23828 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_33_268
timestamp 1639504043
transform 1 0 25760 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1639504043
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1639504043
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1639504043
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1639504043
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1639504043
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1639504043
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_301
timestamp 1639504043
transform 1 0 28796 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1639504043
transform -1 0 29440 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1639504043
transform -1 0 29440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_15
timestamp 1639504043
transform 1 0 2484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1639504043
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1639504043
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_23
timestamp 1639504043
transform 1 0 3220 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_33
timestamp 1639504043
transform 1 0 4140 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1157_
timestamp 1639504043
transform -1 0 4876 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1160_
timestamp 1639504043
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _1183_
timestamp 1639504043
transform 1 0 3404 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_44
timestamp 1639504043
transform 1 0 5152 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_50
timestamp 1639504043
transform 1 0 5704 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1639504043
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0978_
timestamp 1639504043
transform 1 0 6348 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1154_
timestamp 1639504043
transform 1 0 6808 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1155_
timestamp 1639504043
transform -1 0 6256 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_35_77
timestamp 1639504043
transform 1 0 8188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_85
timestamp 1639504043
transform 1 0 8924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0879_
timestamp 1639504043
transform 1 0 7636 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0995_
timestamp 1639504043
transform -1 0 9476 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1210_
timestamp 1639504043
transform -1 0 8188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_clk_i
timestamp 1639504043
transform -1 0 7636 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1639504043
transform -1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0991_
timestamp 1639504043
transform -1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_2  _0996_
timestamp 1639504043
transform 1 0 9476 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1006_
timestamp 1639504043
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B
timestamp 1639504043
transform -1 0 11684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_115
timestamp 1639504043
transform 1 0 11684 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1639504043
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_127
timestamp 1639504043
transform 1 0 12788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_131
timestamp 1639504043
transform 1 0 13156 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1639504043
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_2  _1421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 12144 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1800__CLK
timestamp 1639504043
transform 1 0 13248 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1800_
timestamp 1639504043
transform 1 0 13432 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_35_161
timestamp 1639504043
transform 1 0 15916 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1639504043
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_172
timestamp 1639504043
transform 1 0 16928 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1639504043
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0880_
timestamp 1639504043
transform 1 0 15364 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0915_
timestamp 1639504043
transform 1 0 15640 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1385_
timestamp 1639504043
transform 1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1386_
timestamp 1639504043
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1639504043
transform 1 0 18032 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_196
timestamp 1639504043
transform 1 0 19136 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_i_A
timestamp 1639504043
transform 1 0 19412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_205
timestamp 1639504043
transform 1 0 19964 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_213
timestamp 1639504043
transform 1 0 20700 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1639504043
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0896_
timestamp 1639504043
transform 1 0 20884 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clk_i
timestamp 1639504043
transform -1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A1
timestamp 1639504043
transform -1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1639504043
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0897_
timestamp 1639504043
transform 1 0 23000 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0903_
timestamp 1639504043
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0905_
timestamp 1639504043
transform -1 0 22816 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_262
timestamp 1639504043
transform 1 0 25208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _1903_
timestamp 1639504043
transform 1 0 23276 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_35_274
timestamp 1639504043
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1639504043
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1639504043
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1639504043
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1639504043
transform -1 0 29440 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_15
timestamp 1639504043
transform 1 0 2484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1639504043
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1639504043
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1190_
timestamp 1639504043
transform 1 0 2852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_22
timestamp 1639504043
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_35
timestamp 1639504043
transform 1 0 4324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1639504043
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1158_
timestamp 1639504043
transform -1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1196_
timestamp 1639504043
transform 1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1745_
timestamp 1639504043
transform 1 0 4876 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_58
timestamp 1639504043
transform 1 0 6440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_62
timestamp 1639504043
transform 1 0 6808 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1832_
timestamp 1639504043
transform 1 0 6900 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1639504043
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_2  _1213_
timestamp 1639504043
transform 1 0 8924 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_i_A
timestamp 1639504043
transform 1 0 10948 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_109
timestamp 1639504043
transform 1 0 11132 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_98
timestamp 1639504043
transform 1 0 10120 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0989_
timestamp 1639504043
transform -1 0 10672 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1639504043
transform 1 0 10672 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clk_i
timestamp 1639504043
transform -1 0 10120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1801__CLK
timestamp 1639504043
transform 1 0 11684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1801_
timestamp 1639504043
transform 1 0 11868 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1639504043
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1639504043
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1639504043
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0883_
timestamp 1639504043
transform -1 0 15364 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0997_
timestamp 1639504043
transform -1 0 15088 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_155
timestamp 1639504043
transform 1 0 15364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1798_
timestamp 1639504043
transform 1 0 15548 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_36_178
timestamp 1639504043
transform 1 0 17480 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1639504043
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1639504043
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1703_
timestamp 1639504043
transform 1 0 18032 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__B1
timestamp 1639504043
transform -1 0 20240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_208
timestamp 1639504043
transform 1 0 20240 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _1105_
timestamp 1639504043
transform 1 0 19228 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1901_
timestamp 1639504043
transform 1 0 20976 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_2  _0899_
timestamp 1639504043
transform 1 0 22908 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A1
timestamp 1639504043
transform -1 0 23828 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B1
timestamp 1639504043
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1639504043
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1639504043
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0898_
timestamp 1639504043
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1639504043
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1639504043
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1639504043
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_301
timestamp 1639504043
transform 1 0 28796 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1639504043
transform -1 0 29440 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1639504043
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1404_
timestamp 1639504043
transform -1 0 3404 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1835_
timestamp 1639504043
transform 1 0 1380 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_37_25
timestamp 1639504043
transform 1 0 3404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_42
timestamp 1639504043
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_2  _1162_
timestamp 1639504043
transform -1 0 4140 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1163_
timestamp 1639504043
transform -1 0 4968 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1198_
timestamp 1639504043
transform 1 0 4140 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1639504043
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1639504043
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_65
timestamp 1639504043
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1639504043
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_72
timestamp 1639504043
transform 1 0 7728 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_80
timestamp 1639504043
transform 1 0 8464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1211_
timestamp 1639504043
transform 1 0 7452 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1212_
timestamp 1639504043
transform 1 0 7912 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1289_
timestamp 1639504043
transform -1 0 8464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1290_
timestamp 1639504043
transform -1 0 7452 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1295_
timestamp 1639504043
transform -1 0 9476 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__B1
timestamp 1639504043
transform 1 0 10212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_101
timestamp 1639504043
transform 1 0 10396 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_91
timestamp 1639504043
transform 1 0 9476 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_2  _0992_
timestamp 1639504043
transform -1 0 10212 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1470_
timestamp 1639504043
transform -1 0 11408 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_123
timestamp 1639504043
transform 1 0 12420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_129
timestamp 1639504043
transform 1 0 12972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1639504043
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__a31oi_2  _1025_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 12420 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1378_
timestamp 1639504043
transform 1 0 13064 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_136
timestamp 1639504043
transform 1 0 13616 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_144
timestamp 1639504043
transform 1 0 14352 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_151
timestamp 1639504043
transform 1 0 14996 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1379_
timestamp 1639504043
transform -1 0 13616 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1380_
timestamp 1639504043
transform 1 0 14444 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1381_
timestamp 1639504043
transform -1 0 14996 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1639504043
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1639504043
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1639504043
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1639504043
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0884_
timestamp 1639504043
transform 1 0 15548 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1384_
timestamp 1639504043
transform 1 0 15824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1861_
timestamp 1639504043
transform 1 0 17020 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__o221a_2  _1109_
timestamp 1639504043
transform -1 0 19412 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_37_199
timestamp 1639504043
transform 1 0 19412 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0881_
timestamp 1639504043
transform 1 0 21068 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1863_
timestamp 1639504043
transform -1 0 21068 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1639504043
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_231
timestamp 1639504043
transform 1 0 22356 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_239
timestamp 1639504043
transform 1 0 23092 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1639504043
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0876_
timestamp 1639504043
transform -1 0 23092 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0893_
timestamp 1639504043
transform 1 0 22540 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0900_
timestamp 1639504043
transform -1 0 22080 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0904_
timestamp 1639504043
transform 1 0 22080 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_247
timestamp 1639504043
transform 1 0 23828 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1907_
timestamp 1639504043
transform 1 0 23920 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1639504043
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1639504043
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1639504043
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1639504043
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1639504043
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1639504043
transform -1 0 29440 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_10
timestamp 1639504043
transform 1 0 2024 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1639504043
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1639504043
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1205_
timestamp 1639504043
transform -1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1639504043
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_36
timestamp 1639504043
transform 1 0 4416 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1639504043
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_2  _1197_
timestamp 1639504043
transform -1 0 4416 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1786_
timestamp 1639504043
transform -1 0 6164 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_38_55
timestamp 1639504043
transform 1 0 6164 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1824_
timestamp 1639504043
transform -1 0 8280 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1824__CLK
timestamp 1639504043
transform -1 0 8464 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1639504043
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1639504043
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1639504043
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1022_
timestamp 1639504043
transform 1 0 10856 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _1023_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 9292 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _1024_
timestamp 1639504043
transform -1 0 10856 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_38_116
timestamp 1639504043
transform 1 0 11776 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1431_
timestamp 1639504043
transform 1 0 12880 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1469_
timestamp 1639504043
transform -1 0 11776 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1639504043
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_141
timestamp 1639504043
transform 1 0 14076 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_145
timestamp 1639504043
transform 1 0 14444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_149
timestamp 1639504043
transform 1 0 14812 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1639504043
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1375_
timestamp 1639504043
transform -1 0 15180 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1382_
timestamp 1639504043
transform 1 0 14168 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1432_
timestamp 1639504043
transform 1 0 13340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_153
timestamp 1639504043
transform 1 0 15180 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_2  _1794_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 15272 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__B1
timestamp 1639504043
transform -1 0 18860 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_175
timestamp 1639504043
transform 1 0 17204 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_187
timestamp 1639504043
transform 1 0 18308 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1639504043
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1639504043
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1102_
timestamp 1639504043
transform 1 0 18400 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_206
timestamp 1639504043
transform 1 0 20056 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_214
timestamp 1639504043
transform 1 0 20792 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1697_
timestamp 1639504043
transform 1 0 19228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1902_
timestamp 1639504043
transform -1 0 22816 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_38_236
timestamp 1639504043
transform 1 0 22816 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0874_
timestamp 1639504043
transform 1 0 22908 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1639504043
transform 1 0 23184 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A1
timestamp 1639504043
transform -1 0 24564 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__B1
timestamp 1639504043
transform -1 0 24748 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1639504043
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_257
timestamp 1639504043
transform 1 0 24748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1639504043
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0882_
timestamp 1639504043
transform 1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_269
timestamp 1639504043
transform 1 0 25852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_281
timestamp 1639504043
transform 1 0 26956 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_293
timestamp 1639504043
transform 1 0 28060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1639504043
transform -1 0 29440 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1639504043
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1639504043
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1639504043
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1161_
timestamp 1639504043
transform 1 0 2760 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _1202_
timestamp 1639504043
transform -1 0 3680 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _1207_
timestamp 1639504043
transform 1 0 1932 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1834_
timestamp 1639504043
transform 1 0 1380 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__o32a_2  _1204_
timestamp 1639504043
transform 1 0 3772 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1639504043
transform -1 0 3496 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1639504043
transform -1 0 3772 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1639504043
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_29
timestamp 1639504043
transform 1 0 3772 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _1403_
timestamp 1639504043
transform 1 0 4508 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1185_
timestamp 1639504043
transform -1 0 4416 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1639504043
transform -1 0 4876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_41
timestamp 1639504043
transform 1 0 4876 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_36
timestamp 1639504043
transform 1 0 4416 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1787_
timestamp 1639504043
transform 1 0 5060 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_39_45
timestamp 1639504043
transform 1 0 5244 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1639504043
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_60
timestamp 1639504043
transform 1 0 6624 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1639504043
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1402_
timestamp 1639504043
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1714_
timestamp 1639504043
transform 1 0 6348 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1876_
timestamp 1639504043
transform 1 0 6900 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_39_66
timestamp 1639504043
transform 1 0 7176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_71
timestamp 1639504043
transform 1 0 7636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_83
timestamp 1639504043
transform 1 0 8740 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1639504043
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _1060_
timestamp 1639504043
transform 1 0 8924 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1061_
timestamp 1639504043
transform -1 0 7636 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clk_i
timestamp 1639504043
transform -1 0 10120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_94
timestamp 1639504043
transform 1 0 9752 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_91
timestamp 1639504043
transform 1 0 9476 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1639504043
transform 1 0 10120 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0985_
timestamp 1639504043
transform 1 0 10028 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_39_103
timestamp 1639504043
transform 1 0 10580 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_i_A
timestamp 1639504043
transform 1 0 10396 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_108
timestamp 1639504043
transform 1 0 11040 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1639504043
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A2
timestamp 1639504043
transform 1 0 10856 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__C_N
timestamp 1639504043
transform 1 0 10856 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B
timestamp 1639504043
transform 1 0 10672 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_120
timestamp 1639504043
transform 1 0 12144 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1639504043
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__or3b_2  _1291_
timestamp 1639504043
transform -1 0 12144 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1376_
timestamp 1639504043
transform -1 0 13248 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1377_
timestamp 1639504043
transform -1 0 12972 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1802_
timestamp 1639504043
transform 1 0 11408 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_39_132
timestamp 1639504043
transform 1 0 13248 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1639504043
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1639504043
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1639504043
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_147
timestamp 1639504043
transform 1 0 14628 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1639504043
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1383_
timestamp 1639504043
transform 1 0 14352 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _1799_
timestamp 1639504043
transform 1 0 13340 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _1435_
timestamp 1639504043
transform 1 0 15272 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1092_
timestamp 1639504043
transform 1 0 15824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_163
timestamp 1639504043
transform 1 0 16100 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_157
timestamp 1639504043
transform 1 0 15548 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1394_
timestamp 1639504043
transform -1 0 16928 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1393_
timestamp 1639504043
transform 1 0 16192 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1639504043
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_172
timestamp 1639504043
transform 1 0 16928 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1639504043
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1864_
timestamp 1639504043
transform 1 0 16836 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_40_159
timestamp 1639504043
transform 1 0 15732 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__B1
timestamp 1639504043
transform -1 0 17664 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_i_A
timestamp 1639504043
transform -1 0 19136 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_192
timestamp 1639504043
transform 1 0 18768 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_188
timestamp 1639504043
transform 1 0 18400 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1639504043
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1103_
timestamp 1639504043
transform -1 0 18768 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1104_
timestamp 1639504043
transform -1 0 18492 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B1
timestamp 1639504043
transform 1 0 20148 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_209
timestamp 1639504043
transform 1 0 20332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_218
timestamp 1639504043
transform 1 0 21160 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _1106_
timestamp 1639504043
transform 1 0 19320 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1862_
timestamp 1639504043
transform -1 0 21160 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clk_i
timestamp 1639504043
transform -1 0 19596 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0902_
timestamp 1639504043
transform 1 0 21896 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0901_
timestamp 1639504043
transform -1 0 22080 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1639504043
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1639504043
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0894_
timestamp 1639504043
transform -1 0 22816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_236
timestamp 1639504043
transform 1 0 22816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_236
timestamp 1639504043
transform 1 0 22816 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_232
timestamp 1639504043
transform 1 0 22448 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_228
timestamp 1639504043
transform 1 0 22080 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__B1
timestamp 1639504043
transform 1 0 22632 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__B1
timestamp 1639504043
transform 1 0 23092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_242
timestamp 1639504043
transform 1 0 23368 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1639504043
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_256
timestamp 1639504043
transform 1 0 24656 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1639504043
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0877_
timestamp 1639504043
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1628_
timestamp 1639504043
transform 1 0 23460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1629_
timestamp 1639504043
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1908_
timestamp 1639504043
transform 1 0 23736 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_39_267
timestamp 1639504043
transform 1 0 25668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1639504043
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1639504043
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_264
timestamp 1639504043
transform 1 0 25392 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1639504043
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1815_
timestamp 1639504043
transform 1 0 25484 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1639504043
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_286
timestamp 1639504043
transform 1 0 27416 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_298
timestamp 1639504043
transform 1 0 28520 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_304
timestamp 1639504043
transform 1 0 29072 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1639504043
transform -1 0 29440 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1639504043
transform -1 0 29440 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_11
timestamp 1639504043
transform 1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_21
timestamp 1639504043
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1639504043
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1639504043
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1206_
timestamp 1639504043
transform 1 0 2392 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_41_33
timestamp 1639504043
transform 1 0 4140 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_37
timestamp 1639504043
transform 1 0 4508 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_41
timestamp 1639504043
transform 1 0 4876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1195_
timestamp 1639504043
transform -1 0 4508 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1203_
timestamp 1639504043
transform -1 0 4876 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1639504043
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_57
timestamp 1639504043
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1639504043
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1059_
timestamp 1639504043
transform 1 0 6900 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1058_
timestamp 1639504043
transform -1 0 7452 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1877_
timestamp 1639504043
transform 1 0 7452 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__or3b_2  _0984_
timestamp 1639504043
transform 1 0 10672 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1468_
timestamp 1639504043
transform -1 0 9844 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1640_
timestamp 1639504043
transform 1 0 9844 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1292_
timestamp 1639504043
transform -1 0 12236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1639504043
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_117
timestamp 1639504043
transform 1 0 11868 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1639504043
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__C_N
timestamp 1639504043
transform 1 0 11684 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1639504043
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1294_
timestamp 1639504043
transform 1 0 12696 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 1639504043
transform 1 0 12236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_129
timestamp 1639504043
transform 1 0 12972 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A
timestamp 1639504043
transform 1 0 12512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1821_
timestamp 1639504043
transform 1 0 13064 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_2  _1571_
timestamp 1639504043
transform 1 0 14996 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1571__B1
timestamp 1639504043
transform 1 0 15732 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1639504043
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1639504043
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1639504043
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1639504043
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_181
timestamp 1639504043
transform 1 0 17756 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_185
timestamp 1639504043
transform 1 0 18124 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_195
timestamp 1639504043
transform 1 0 19044 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1100_
timestamp 1639504043
transform 1 0 17848 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1685_
timestamp 1639504043
transform 1 0 18216 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_207
timestamp 1639504043
transform 1 0 20148 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_214
timestamp 1639504043
transform 1 0 20792 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1340_
timestamp 1639504043
transform 1 0 20516 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1676_
timestamp 1639504043
transform 1 0 19320 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_clk_i
timestamp 1639504043
transform 1 0 20976 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1639504043
transform 1 0 22080 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1639504043
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_230
timestamp 1639504043
transform 1 0 22264 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_238
timestamp 1639504043
transform 1 0 23000 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1639504043
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0891_
timestamp 1639504043
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1814_
timestamp 1639504043
transform -1 0 25116 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_41_261
timestamp 1639504043
transform 1 0 25116 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1333_
timestamp 1639504043
transform 1 0 25208 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A1
timestamp 1639504043
transform 1 0 26588 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__B1
timestamp 1639504043
transform -1 0 27140 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_270
timestamp 1639504043
transform 1 0 25944 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1639504043
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_283
timestamp 1639504043
transform 1 0 27140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1639504043
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1331_
timestamp 1639504043
transform 1 0 26036 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1332_
timestamp 1639504043
transform 1 0 26312 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_295
timestamp 1639504043
transform 1 0 28244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_303
timestamp 1639504043
transform 1 0 28980 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1639504043
transform -1 0 29440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_15
timestamp 1639504043
transform 1 0 2484 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1639504043
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1639504043
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1209_
timestamp 1639504043
transform 1 0 2576 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1639504043
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_37
timestamp 1639504043
transform 1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1639504043
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1199_
timestamp 1639504043
transform -1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1713_
timestamp 1639504043
transform 1 0 6808 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1788_
timestamp 1639504043
transform 1 0 5244 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_42_71
timestamp 1639504043
transform 1 0 7636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_75
timestamp 1639504043
transform 1 0 8004 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1639504043
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1639504043
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1054_
timestamp 1639504043
transform 1 0 8464 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1055_
timestamp 1639504043
transform -1 0 9200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_clk_i
timestamp 1639504043
transform -1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_105
timestamp 1639504043
transform 1 0 10764 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_88
timestamp 1639504043
transform 1 0 9200 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1641_
timestamp 1639504043
transform 1 0 9936 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__C_N
timestamp 1639504043
transform 1 0 11408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_111
timestamp 1639504043
transform 1 0 11316 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_127
timestamp 1639504043
transform 1 0 12788 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0983_
timestamp 1639504043
transform 1 0 12236 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _1020_
timestamp 1639504043
transform 1 0 11592 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1305_
timestamp 1639504043
transform 1 0 12880 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__A1
timestamp 1639504043
transform -1 0 14260 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__B1
timestamp 1639504043
transform -1 0 14444 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_136
timestamp 1639504043
transform 1 0 13616 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_145
timestamp 1639504043
transform 1 0 14444 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1639504043
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1570_
timestamp 1639504043
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1572_
timestamp 1639504043
transform -1 0 15456 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__B1
timestamp 1639504043
transform 1 0 15456 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_158
timestamp 1639504043
transform 1 0 15640 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_164
timestamp 1639504043
transform 1 0 16192 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1093_
timestamp 1639504043
transform -1 0 16560 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1680_
timestamp 1639504043
transform 1 0 16560 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_177
timestamp 1639504043
transform 1 0 17388 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_181
timestamp 1639504043
transform 1 0 17756 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1639504043
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1639504043
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1639504043
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1637_
timestamp 1639504043
transform 1 0 17848 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A
timestamp 1639504043
transform 1 0 20240 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_206
timestamp 1639504043
transform 1 0 20056 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_213
timestamp 1639504043
transform 1 0 20700 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1330_
timestamp 1639504043
transform 1 0 20424 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1701_
timestamp 1639504043
transform 1 0 19228 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1904_
timestamp 1639504043
transform 1 0 20792 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_2  _0895_
timestamp 1639504043
transform 1 0 22724 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__B1
timestamp 1639504043
transform -1 0 25116 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1639504043
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1639504043
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1334_
timestamp 1639504043
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1335_
timestamp 1639504043
transform -1 0 24932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1336_
timestamp 1639504043
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1339_
timestamp 1639504043
transform -1 0 25852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__B1
timestamp 1639504043
transform -1 0 26312 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_274
timestamp 1639504043
transform 1 0 26312 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1337_
timestamp 1639504043
transform 1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_286
timestamp 1639504043
transform 1 0 27416 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_298
timestamp 1639504043
transform 1 0 28520 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_304
timestamp 1639504043
transform 1 0 29072 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1639504043
transform -1 0 29440 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1639504043
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1639504043
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1833_
timestamp 1639504043
transform 1 0 1748 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_43_24
timestamp 1639504043
transform 1 0 3312 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1836_
timestamp 1639504043
transform 1 0 3588 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1639504043
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1639504043
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_65
timestamp 1639504043
transform 1 0 7084 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1639504043
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1397_
timestamp 1639504043
transform 1 0 5152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1401_
timestamp 1639504043
transform -1 0 7084 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_80
timestamp 1639504043
transform 1 0 8464 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1056_
timestamp 1639504043
transform 1 0 8832 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1057_
timestamp 1639504043
transform -1 0 8464 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_93
timestamp 1639504043
transform 1 0 9660 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1642_
timestamp 1639504043
transform 1 0 10212 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_clk_i
timestamp 1639504043
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A
timestamp 1639504043
transform 1 0 12420 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1639504043
transform 1 0 12696 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B
timestamp 1639504043
transform 1 0 12880 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__C
timestamp 1639504043
transform 1 0 13064 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_125
timestamp 1639504043
transform 1 0 12604 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1639504043
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1639504043
transform -1 0 12420 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0982_
timestamp 1639504043
transform 1 0 11500 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1639504043
transform 1 0 13248 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_134
timestamp 1639504043
transform 1 0 13432 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_142
timestamp 1639504043
transform 1 0 14168 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_147
timestamp 1639504043
transform 1 0 14628 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1304_
timestamp 1639504043
transform -1 0 14628 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1573_
timestamp 1639504043
transform -1 0 15456 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B1
timestamp 1639504043
transform -1 0 15732 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_156
timestamp 1639504043
transform 1 0 15456 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1639504043
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1098_
timestamp 1639504043
transform 1 0 15732 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1867_
timestamp 1639504043
transform -1 0 18216 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_43_186
timestamp 1639504043
transform 1 0 18216 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1099_
timestamp 1639504043
transform 1 0 18492 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_43_215
timestamp 1639504043
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1866_
timestamp 1639504043
transform -1 0 20884 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1639504043
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_228
timestamp 1639504043
transform 1 0 22080 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_240
timestamp 1639504043
transform 1 0 23184 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1639504043
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0892_
timestamp 1639504043
transform -1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__B1
timestamp 1639504043
transform 1 0 23460 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A1
timestamp 1639504043
transform -1 0 23460 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_245
timestamp 1639504043
transform 1 0 23644 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_257
timestamp 1639504043
transform 1 0 24748 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1813_
timestamp 1639504043
transform 1 0 24932 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1639504043
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1338_
timestamp 1639504043
transform -1 0 27232 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_284
timestamp 1639504043
transform 1 0 27232 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_296
timestamp 1639504043
transform 1 0 28336 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_304
timestamp 1639504043
transform 1 0 29072 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1639504043
transform -1 0 29440 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_15
timestamp 1639504043
transform 1 0 2484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_19
timestamp 1639504043
transform 1 0 2852 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1639504043
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1639504043
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1208_
timestamp 1639504043
transform 1 0 2944 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1639504043
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_29
timestamp 1639504043
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_35
timestamp 1639504043
transform 1 0 4324 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_43
timestamp 1639504043
transform 1 0 5060 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1639504043
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1187_
timestamp 1639504043
transform -1 0 4324 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_62
timestamp 1639504043
transform 1 0 6808 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1789_
timestamp 1639504043
transform 1 0 5244 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_44_70
timestamp 1639504043
transform 1 0 7544 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_79
timestamp 1639504043
transform 1 0 8372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1639504043
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1639504043
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1639504043
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1044_
timestamp 1639504043
transform -1 0 8096 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1050_
timestamp 1639504043
transform 1 0 8096 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_103
timestamp 1639504043
transform 1 0 10580 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_97
timestamp 1639504043
transform 1 0 10028 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1027_
timestamp 1639504043
transform -1 0 10580 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1643_
timestamp 1639504043
transform 1 0 10764 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__D
timestamp 1639504043
transform 1 0 12144 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1643__A1
timestamp 1639504043
transform -1 0 11776 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1639504043
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_122
timestamp 1639504043
transform 1 0 12328 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _1052_
timestamp 1639504043
transform 1 0 12604 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__B1
timestamp 1639504043
transform 1 0 13524 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1639504043
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_141
timestamp 1639504043
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1639504043
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1303_
timestamp 1639504043
transform -1 0 15180 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1574_
timestamp 1639504043
transform -1 0 14904 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1573__B1
timestamp 1639504043
transform 1 0 15456 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__B1
timestamp 1639504043
transform 1 0 15180 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_155
timestamp 1639504043
transform 1 0 15364 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_158
timestamp 1639504043
transform 1 0 15640 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1707_
timestamp 1639504043
transform 1 0 16376 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_44_175
timestamp 1639504043
transform 1 0 17204 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_187
timestamp 1639504043
transform 1 0 18308 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1639504043
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1095_
timestamp 1639504043
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 1639504043
transform 1 0 17480 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_clk_i
timestamp 1639504043
transform -1 0 18860 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__B1
timestamp 1639504043
transform -1 0 19688 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__B1
timestamp 1639504043
transform -1 0 19964 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_202
timestamp 1639504043
transform 1 0 19688 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_205
timestamp 1639504043
transform 1 0 19964 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_217
timestamp 1639504043
transform 1 0 21068 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1096_
timestamp 1639504043
transform -1 0 19504 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1639504043
transform -1 0 22448 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B1
timestamp 1639504043
transform 1 0 23000 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1639504043
transform -1 0 21620 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_226
timestamp 1639504043
transform 1 0 21896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_232
timestamp 1639504043
transform 1 0 22448 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0885_
timestamp 1639504043
transform 1 0 21988 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0887_
timestamp 1639504043
transform 1 0 23184 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0888_
timestamp 1639504043
transform -1 0 21896 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1639504043
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1639504043
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1639504043
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1639504043
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1639504043
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1639504043
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_301
timestamp 1639504043
transform 1 0 28796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1639504043
transform -1 0 29440 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_15
timestamp 1639504043
transform 1 0 2484 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1639504043
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1639504043
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1838_
timestamp 1639504043
transform 1 0 2760 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _1159_
timestamp 1639504043
transform -1 0 4876 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1186_
timestamp 1639504043
transform 1 0 4876 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_44
timestamp 1639504043
transform 1 0 5152 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_57
timestamp 1639504043
transform 1 0 6348 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1639504043
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1400_
timestamp 1639504043
transform 1 0 5520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1712_
timestamp 1639504043
transform 1 0 6440 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1878_
timestamp 1639504043
transform -1 0 9200 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_45_103
timestamp 1639504043
transform 1 0 10580 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0998_
timestamp 1639504043
transform -1 0 11408 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1047_
timestamp 1639504043
transform -1 0 10580 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_2  _1053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 9200 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1639504043
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_127
timestamp 1639504043
transform 1 0 12788 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1639504043
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2ai_2  _1031_
timestamp 1639504043
transform 1 0 11684 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_138
timestamp 1639504043
transform 1 0 13800 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1029_
timestamp 1639504043
transform 1 0 13524 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _1042_
timestamp 1639504043
transform 1 0 14352 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__B1
timestamp 1639504043
transform 1 0 15548 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__B1
timestamp 1639504043
transform -1 0 16560 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_159
timestamp 1639504043
transform 1 0 15732 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_165
timestamp 1639504043
transform 1 0 16284 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1639504043
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1097_
timestamp 1639504043
transform -1 0 17480 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1296_
timestamp 1639504043
transform 1 0 15272 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_178
timestamp 1639504043
transform 1 0 17480 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_184
timestamp 1639504043
transform 1 0 18032 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1101_
timestamp 1639504043
transform 1 0 18952 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1698_
timestamp 1639504043
transform 1 0 18124 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1865_
timestamp 1639504043
transform -1 0 21344 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_45_220
timestamp 1639504043
transform 1 0 21344 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1639504043
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0889_
timestamp 1639504043
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1905_
timestamp 1639504043
transform -1 0 23736 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1906_
timestamp 1639504043
transform -1 0 25668 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_45_270
timestamp 1639504043
transform 1 0 25944 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1639504043
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1639504043
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1639504043
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1326_
timestamp 1639504043
transform 1 0 25668 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1639504043
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1639504043
transform -1 0 29440 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1639504043
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1639504043
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1639504043
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1639504043
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1639504043
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1639504043
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1639504043
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_37
timestamp 1639504043
transform 1 0 4508 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_27
timestamp 1639504043
transform 1 0 3588 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_35
timestamp 1639504043
transform 1 0 4324 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1639504043
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1188_
timestamp 1639504043
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1708_
timestamp 1639504043
transform 1 0 4416 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_46_49
timestamp 1639504043
transform 1 0 5612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_61
timestamp 1639504043
transform 1 0 6716 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_45
timestamp 1639504043
transform 1 0 5244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1639504043
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1639504043
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1639504043
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1711_
timestamp 1639504043
transform 1 0 6532 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_46_73
timestamp 1639504043
transform 1 0 7820 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1639504043
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_68
timestamp 1639504043
transform 1 0 7360 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1639504043
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1045_
timestamp 1639504043
transform 1 0 7912 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_2  _1049_
timestamp 1639504043
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1051_
timestamp 1639504043
transform -1 0 8464 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1879_
timestamp 1639504043
transform -1 0 9384 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_46_107
timestamp 1639504043
transform 1 0 10948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_97
timestamp 1639504043
transform 1 0 10028 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_90
timestamp 1639504043
transform 1 0 9384 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _1034_
timestamp 1639504043
transform 1 0 10120 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1882_
timestamp 1639504043
transform 1 0 9476 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_47_113
timestamp 1639504043
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_121
timestamp 1639504043
transform 1 0 12236 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_126
timestamp 1639504043
transform 1 0 12696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1639504043
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0999_
timestamp 1639504043
transform 1 0 11500 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1000_
timestamp 1639504043
transform 1 0 12420 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1883_
timestamp 1639504043
transform -1 0 13708 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B1
timestamp 1639504043
transform 1 0 14996 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1639504043
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_138
timestamp 1639504043
transform 1 0 13800 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_144
timestamp 1639504043
transform 1 0 14352 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1639504043
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_2  _1030_
timestamp 1639504043
transform 1 0 14076 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__a22oi_2  _1048_
timestamp 1639504043
transform 1 0 14444 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__B1
timestamp 1639504043
transform 1 0 15364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_153
timestamp 1639504043
transform 1 0 15180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_157
timestamp 1639504043
transform 1 0 15548 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_157
timestamp 1639504043
transform 1 0 15548 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_165
timestamp 1639504043
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_169
timestamp 1639504043
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1639504043
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1868_
timestamp 1639504043
transform 1 0 15640 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1704_
timestamp 1639504043
transform 1 0 17572 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1686_
timestamp 1639504043
transform 1 0 17572 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_177
timestamp 1639504043
transform 1 0 17388 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_175
timestamp 1639504043
transform 1 0 17204 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1088_
timestamp 1639504043
transform -1 0 18952 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1086_
timestamp 1639504043
transform -1 0 18676 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1639504043
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_188
timestamp 1639504043
transform 1 0 18400 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1639504043
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1869_
timestamp 1639504043
transform -1 0 20332 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__B1
timestamp 1639504043
transform -1 0 20240 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A
timestamp 1639504043
transform -1 0 20424 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_213
timestamp 1639504043
transform 1 0 20700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_209
timestamp 1639504043
transform 1 0 20332 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_215
timestamp 1639504043
transform 1 0 20884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _1094_
timestamp 1639504043
transform -1 0 20056 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1307_
timestamp 1639504043
transform 1 0 20608 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1315_
timestamp 1639504043
transform 1 0 20424 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1639504043
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_225
timestamp 1639504043
transform 1 0 21804 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1639504043
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_225
timestamp 1639504043
transform 1 0 21804 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__B1
timestamp 1639504043
transform 1 0 21896 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1312_
timestamp 1639504043
transform 1 0 22264 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1311_
timestamp 1639504043
transform -1 0 23092 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1310_
timestamp 1639504043
transform -1 0 22816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0890_
timestamp 1639504043
transform 1 0 22724 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_228
timestamp 1639504043
transform 1 0 22080 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_233
timestamp 1639504043
transform 1 0 22540 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_239
timestamp 1639504043
transform 1 0 23092 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1327_
timestamp 1639504043
transform 1 0 23460 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0886_
timestamp 1639504043
transform 1 0 23828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_246
timestamp 1639504043
transform 1 0 23736 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__B1
timestamp 1639504043
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _1329_
timestamp 1639504043
transform 1 0 25208 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1325_
timestamp 1639504043
transform 1 0 24748 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1639504043
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1639504043
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1817_
timestamp 1639504043
transform 1 0 23276 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1816_
timestamp 1639504043
transform 1 0 25024 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__B1
timestamp 1639504043
transform 1 0 25944 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_281
timestamp 1639504043
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_272
timestamp 1639504043
transform 1 0 26128 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1639504043
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1639504043
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_293
timestamp 1639504043
transform 1 0 28060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1639504043
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1639504043
transform -1 0 29440 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1639504043
transform -1 0 29440 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1639504043
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1639504043
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1639504043
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1639504043
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_29
timestamp 1639504043
transform 1 0 3772 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_38
timestamp 1639504043
transform 1 0 4600 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1639504043
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1396_
timestamp 1639504043
transform 1 0 3864 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _1399_
timestamp 1639504043
transform 1 0 6716 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1790_
timestamp 1639504043
transform 1 0 5152 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_48_69
timestamp 1639504043
transform 1 0 7452 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_77
timestamp 1639504043
transform 1 0 8188 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1639504043
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1639504043
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1639504043
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1046_
timestamp 1639504043
transform -1 0 8648 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_100
timestamp 1639504043
transform 1 0 10304 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1032_
timestamp 1639504043
transform 1 0 10856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1033_
timestamp 1639504043
transform -1 0 11408 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1035_
timestamp 1639504043
transform -1 0 10304 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_112
timestamp 1639504043
transform 1 0 11408 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_124
timestamp 1639504043
transform 1 0 12512 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_130
timestamp 1639504043
transform 1 0 13064 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1299_
timestamp 1639504043
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__B1
timestamp 1639504043
transform -1 0 14260 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1639504043
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_143
timestamp 1639504043
transform 1 0 14260 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1639504043
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1297_
timestamp 1639504043
transform 1 0 15088 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1300_
timestamp 1639504043
transform -1 0 15088 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_155
timestamp 1639504043
transform 1 0 15364 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_162
timestamp 1639504043
transform 1 0 16008 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_174
timestamp 1639504043
transform 1 0 17112 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1306_
timestamp 1639504043
transform 1 0 15732 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__B1
timestamp 1639504043
transform 1 0 17204 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_186
timestamp 1639504043
transform 1 0 18216 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1639504043
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1639504043
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1091_
timestamp 1639504043
transform -1 0 18216 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1639504043
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_205
timestamp 1639504043
transform 1 0 19964 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1820_
timestamp 1639504043
transform -1 0 22080 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_2  _1313_
timestamp 1639504043
transform -1 0 22816 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1324_
timestamp 1639504043
transform 1 0 22816 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__B1
timestamp 1639504043
transform -1 0 24012 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1639504043
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_259
timestamp 1639504043
transform 1 0 24932 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1639504043
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1322_
timestamp 1639504043
transform 1 0 24380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1323_
timestamp 1639504043
transform -1 0 24932 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1328_
timestamp 1639504043
transform 1 0 23552 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_271
timestamp 1639504043
transform 1 0 26036 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_283
timestamp 1639504043
transform 1 0 27140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_295
timestamp 1639504043
transform 1 0 28244 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_303
timestamp 1639504043
transform 1 0 28980 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1639504043
transform -1 0 29440 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_15
timestamp 1639504043
transform 1 0 2484 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1639504043
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1639504043
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_23
timestamp 1639504043
transform 1 0 3220 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_42
timestamp 1639504043
transform 1 0 4968 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1792_
timestamp 1639504043
transform 1 0 3404 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1639504043
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_61
timestamp 1639504043
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1639504043
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1398_
timestamp 1639504043
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1709_
timestamp 1639504043
transform 1 0 6808 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_49_71
timestamp 1639504043
transform 1 0 7636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_83
timestamp 1639504043
transform 1 0 8740 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_101
timestamp 1639504043
transform 1 0 10396 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_105
timestamp 1639504043
transform 1 0 10764 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1028_
timestamp 1639504043
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1037_
timestamp 1639504043
transform -1 0 10764 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1038_
timestamp 1639504043
transform 1 0 9568 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1039_
timestamp 1639504043
transform -1 0 9568 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_113
timestamp 1639504043
transform 1 0 11500 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_126
timestamp 1639504043
transform 1 0 12696 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1639504043
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2ai_2  _1043_
timestamp 1639504043
transform 1 0 11592 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _1302_
timestamp 1639504043
transform 1 0 12880 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__B1
timestamp 1639504043
transform 1 0 13616 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1823_
timestamp 1639504043
transform 1 0 13800 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1639504043
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1639504043
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1298_
timestamp 1639504043
transform -1 0 16008 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1870_
timestamp 1639504043
transform 1 0 16652 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_49_186
timestamp 1639504043
transform 1 0 18216 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1871_
timestamp 1639504043
transform -1 0 20056 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_49_206
timestamp 1639504043
transform 1 0 20056 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_210
timestamp 1639504043
transform 1 0 20424 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_214
timestamp 1639504043
transform 1 0 20792 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1319_
timestamp 1639504043
transform -1 0 20792 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A1
timestamp 1639504043
transform -1 0 23092 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__B1
timestamp 1639504043
transform 1 0 23092 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1639504043
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_233
timestamp 1639504043
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1639504043
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1316_
timestamp 1639504043
transform 1 0 22632 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1318_
timestamp 1639504043
transform -1 0 22540 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_241
timestamp 1639504043
transform 1 0 23276 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_253
timestamp 1639504043
transform 1 0 24380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_265
timestamp 1639504043
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1639504043
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1639504043
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1639504043
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1639504043
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1639504043
transform -1 0 29440 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_15
timestamp 1639504043
transform 1 0 2484 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_21
timestamp 1639504043
transform 1 0 3036 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1639504043
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1639504043
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_25
timestamp 1639504043
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_29
timestamp 1639504043
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_37
timestamp 1639504043
transform 1 0 4508 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_41
timestamp 1639504043
transform 1 0 4876 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1639504043
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1631_
timestamp 1639504043
transform -1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1633_
timestamp 1639504043
transform 1 0 4600 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_47
timestamp 1639504043
transform 1 0 5428 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1710_
timestamp 1639504043
transform 1 0 7084 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1791_
timestamp 1639504043
transform 1 0 5520 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_50_74
timestamp 1639504043
transform 1 0 7912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1639504043
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_85
timestamp 1639504043
transform 1 0 8924 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1639504043
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1881_
timestamp 1639504043
transform 1 0 9016 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _1036_
timestamp 1639504043
transform -1 0 11224 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_110
timestamp 1639504043
transform 1 0 11224 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1880_
timestamp 1639504043
transform -1 0 13340 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1639504043
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1639504043
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1639504043
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1822_
timestamp 1639504043
transform -1 0 16008 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_50_162
timestamp 1639504043
transform 1 0 16008 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_168
timestamp 1639504043
transform 1 0 16560 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1872_
timestamp 1639504043
transform 1 0 16652 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1639504043
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1639504043
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1089_
timestamp 1639504043
transform -1 0 19044 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__B1
timestamp 1639504043
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_199
timestamp 1639504043
transform 1 0 19412 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1818_
timestamp 1639504043
transform -1 0 21436 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 1639504043
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1819_
timestamp 1639504043
transform 1 0 21804 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1639504043
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1639504043
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1639504043
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1639504043
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1639504043
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1639504043
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_301
timestamp 1639504043
transform 1 0 28796 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1639504043
transform -1 0 29440 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1639504043
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1639504043
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1639504043
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_27
timestamp 1639504043
transform 1 0 3588 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_29
timestamp 1639504043
transform 1 0 3772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_41
timestamp 1639504043
transform 1 0 4876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1639504043
transform 1 0 3680 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1639504043
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1639504043
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1639504043
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1639504043
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_81
timestamp 1639504043
transform 1 0 8556 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_85
timestamp 1639504043
transform 1 0 8924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1639504043
transform 1 0 8832 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_109
timestamp 1639504043
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_97
timestamp 1639504043
transform 1 0 10028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1639504043
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_119
timestamp 1639504043
transform 1 0 12052 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1639504043
transform 1 0 12420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1639504043
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1040_
timestamp 1639504043
transform 1 0 11776 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1041_
timestamp 1639504043
transform -1 0 12420 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_135
timestamp 1639504043
transform 1 0 13524 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_139
timestamp 1639504043
transform 1 0 13892 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_141
timestamp 1639504043
transform 1 0 14076 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_147
timestamp 1639504043
transform 1 0 14628 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_151
timestamp 1639504043
transform 1 0 14996 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1639504043
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1301_
timestamp 1639504043
transform -1 0 14996 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_163
timestamp 1639504043
transform 1 0 16100 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1639504043
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1639504043
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1639504043
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1639504043
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_193
timestamp 1639504043
transform 1 0 18860 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1639504043
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__B1
timestamp 1639504043
transform 1 0 20056 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_208
timestamp 1639504043
transform 1 0 20240 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1639504043
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _1090_
timestamp 1639504043
transform -1 0 20056 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1320_
timestamp 1639504043
transform -1 0 20792 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__A1
timestamp 1639504043
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__B1
timestamp 1639504043
transform 1 0 22540 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_235
timestamp 1639504043
transform 1 0 22724 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_239
timestamp 1639504043
transform 1 0 23092 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1639504043
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1317_
timestamp 1639504043
transform 1 0 22816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1321_
timestamp 1639504043
transform -1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_251
timestamp 1639504043
transform 1 0 24196 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_253
timestamp 1639504043
transform 1 0 24380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1639504043
transform 1 0 24288 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_265
timestamp 1639504043
transform 1 0 25484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1639504043
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1639504043
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1639504043
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1639504043
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1639504043
transform -1 0 29440 0 -1 30464
box -38 -48 314 592
<< labels >>
rlabel metal2 s 570 0 626 800 6 clk_i
port 0 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 data_addr_o[0]
port 1 nsew signal tristate
rlabel metal2 s 13910 31889 13966 32689 6 data_addr_o[10]
port 2 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 data_addr_o[11]
port 3 nsew signal tristate
rlabel metal2 s 5446 0 5502 800 6 data_addr_o[1]
port 4 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 data_addr_o[2]
port 5 nsew signal tristate
rlabel metal2 s 9034 0 9090 800 6 data_addr_o[3]
port 6 nsew signal tristate
rlabel metal3 s 0 12928 800 13048 6 data_addr_o[4]
port 7 nsew signal tristate
rlabel metal2 s 11518 0 11574 800 6 data_addr_o[5]
port 8 nsew signal tristate
rlabel metal3 s 0 15648 800 15768 6 data_addr_o[6]
port 9 nsew signal tristate
rlabel metal3 s 29745 10480 30545 10600 6 data_addr_o[7]
port 10 nsew signal tristate
rlabel metal2 s 14002 0 14058 800 6 data_addr_o[8]
port 11 nsew signal tristate
rlabel metal2 s 12530 31889 12586 32689 6 data_addr_o[9]
port 12 nsew signal tristate
rlabel metal2 s 2962 0 3018 800 6 data_be_o[0]
port 13 nsew signal tristate
rlabel metal2 s 3238 31889 3294 32689 6 data_be_o[1]
port 14 nsew signal tristate
rlabel metal2 s 7838 0 7894 800 6 data_be_o[2]
port 15 nsew signal tristate
rlabel metal2 s 4618 31889 4674 32689 6 data_be_o[3]
port 16 nsew signal tristate
rlabel metal2 s 662 31889 718 32689 6 data_gnt_i
port 17 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 data_rdata_i[0]
port 18 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 data_rdata_i[10]
port 19 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 data_rdata_i[11]
port 20 nsew signal input
rlabel metal3 s 29745 16192 30545 16312 6 data_rdata_i[12]
port 21 nsew signal input
rlabel metal3 s 29745 18232 30545 18352 6 data_rdata_i[13]
port 22 nsew signal input
rlabel metal2 s 16578 31889 16634 32689 6 data_rdata_i[14]
port 23 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 data_rdata_i[15]
port 24 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 data_rdata_i[16]
port 25 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 data_rdata_i[17]
port 26 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 data_rdata_i[18]
port 27 nsew signal input
rlabel metal2 s 20534 31889 20590 32689 6 data_rdata_i[19]
port 28 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 data_rdata_i[1]
port 29 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 data_rdata_i[20]
port 30 nsew signal input
rlabel metal3 s 29745 22040 30545 22160 6 data_rdata_i[21]
port 31 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 data_rdata_i[22]
port 32 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 data_rdata_i[23]
port 33 nsew signal input
rlabel metal2 s 25870 31889 25926 32689 6 data_rdata_i[24]
port 34 nsew signal input
rlabel metal3 s 29745 25848 30545 25968 6 data_rdata_i[25]
port 35 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 data_rdata_i[26]
port 36 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 data_rdata_i[27]
port 37 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 data_rdata_i[28]
port 38 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 data_rdata_i[29]
port 39 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 data_rdata_i[2]
port 40 nsew signal input
rlabel metal3 s 29745 29656 30545 29776 6 data_rdata_i[30]
port 41 nsew signal input
rlabel metal3 s 29745 31560 30545 31680 6 data_rdata_i[31]
port 42 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 data_rdata_i[3]
port 43 nsew signal input
rlabel metal2 s 5906 31889 5962 32689 6 data_rdata_i[4]
port 44 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 data_rdata_i[5]
port 45 nsew signal input
rlabel metal3 s 29745 8576 30545 8696 6 data_rdata_i[6]
port 46 nsew signal input
rlabel metal2 s 7286 31889 7342 32689 6 data_rdata_i[7]
port 47 nsew signal input
rlabel metal2 s 9954 31889 10010 32689 6 data_rdata_i[8]
port 48 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 data_rdata_i[9]
port 49 nsew signal input
rlabel metal3 s 0 688 800 808 6 data_req_o
port 50 nsew signal tristate
rlabel metal3 s 29745 960 30545 1080 6 data_rvalid_i
port 51 nsew signal input
rlabel metal3 s 29745 2864 30545 2984 6 data_wdata_o[0]
port 52 nsew signal tristate
rlabel metal3 s 29745 12384 30545 12504 6 data_wdata_o[10]
port 53 nsew signal tristate
rlabel metal3 s 29745 14288 30545 14408 6 data_wdata_o[11]
port 54 nsew signal tristate
rlabel metal2 s 15198 31889 15254 32689 6 data_wdata_o[12]
port 55 nsew signal tristate
rlabel metal2 s 18878 0 18934 800 6 data_wdata_o[13]
port 56 nsew signal tristate
rlabel metal3 s 29745 20136 30545 20256 6 data_wdata_o[14]
port 57 nsew signal tristate
rlabel metal2 s 17866 31889 17922 32689 6 data_wdata_o[15]
port 58 nsew signal tristate
rlabel metal2 s 22558 0 22614 800 6 data_wdata_o[16]
port 59 nsew signal tristate
rlabel metal2 s 19246 31889 19302 32689 6 data_wdata_o[17]
port 60 nsew signal tristate
rlabel metal2 s 24950 0 25006 800 6 data_wdata_o[18]
port 61 nsew signal tristate
rlabel metal2 s 21822 31889 21878 32689 6 data_wdata_o[19]
port 62 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 data_wdata_o[1]
port 63 nsew signal tristate
rlabel metal2 s 23202 31889 23258 32689 6 data_wdata_o[20]
port 64 nsew signal tristate
rlabel metal2 s 24490 31889 24546 32689 6 data_wdata_o[21]
port 65 nsew signal tristate
rlabel metal2 s 27434 0 27490 800 6 data_wdata_o[22]
port 66 nsew signal tristate
rlabel metal3 s 29745 23944 30545 24064 6 data_wdata_o[23]
port 67 nsew signal tristate
rlabel metal2 s 27158 31889 27214 32689 6 data_wdata_o[24]
port 68 nsew signal tristate
rlabel metal3 s 0 25168 800 25288 6 data_wdata_o[25]
port 69 nsew signal tristate
rlabel metal2 s 28630 0 28686 800 6 data_wdata_o[26]
port 70 nsew signal tristate
rlabel metal3 s 29745 27752 30545 27872 6 data_wdata_o[27]
port 71 nsew signal tristate
rlabel metal2 s 28538 31889 28594 32689 6 data_wdata_o[28]
port 72 nsew signal tristate
rlabel metal3 s 0 30608 800 30728 6 data_wdata_o[29]
port 73 nsew signal tristate
rlabel metal3 s 29745 4768 30545 4888 6 data_wdata_o[2]
port 74 nsew signal tristate
rlabel metal3 s 0 31968 800 32088 6 data_wdata_o[30]
port 75 nsew signal tristate
rlabel metal2 s 29826 31889 29882 32689 6 data_wdata_o[31]
port 76 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 data_wdata_o[3]
port 77 nsew signal tristate
rlabel metal3 s 0 14288 800 14408 6 data_wdata_o[4]
port 78 nsew signal tristate
rlabel metal3 s 29745 6672 30545 6792 6 data_wdata_o[5]
port 79 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 data_wdata_o[6]
port 80 nsew signal tristate
rlabel metal2 s 8574 31889 8630 32689 6 data_wdata_o[7]
port 81 nsew signal tristate
rlabel metal2 s 11242 31889 11298 32689 6 data_wdata_o[8]
port 82 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 data_wdata_o[9]
port 83 nsew signal tristate
rlabel metal2 s 1950 31889 2006 32689 6 data_we_o
port 84 nsew signal tristate
rlabel metal2 s 1766 0 1822 800 6 rst_i
port 85 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 rx_i
port 86 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 tx_o
port 87 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 uart_error
port 88 nsew signal tristate
rlabel metal4 s 5667 2128 5987 30512 6 vccd1
port 89 nsew power input
rlabel metal4 s 15112 2128 15432 30512 6 vccd1
port 89 nsew power input
rlabel metal4 s 24557 2128 24877 30512 6 vccd1
port 89 nsew power input
rlabel metal4 s 10389 2128 10709 30512 6 vssd1
port 90 nsew ground input
rlabel metal4 s 19834 2128 20154 30512 6 vssd1
port 90 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 30545 32689
<< end >>
