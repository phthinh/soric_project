magic
tech sky130A
magscale 1 2
timestamp 1640365532
<< obsli1 >>
rect 1104 1717 238987 237745
<< obsm1 >>
rect 14 1300 238999 237776
<< metal2 >>
rect 1214 239200 1270 240000
rect 3606 239200 3662 240000
rect 5998 239200 6054 240000
rect 8390 239200 8446 240000
rect 10782 239200 10838 240000
rect 13174 239200 13230 240000
rect 15566 239200 15622 240000
rect 17958 239200 18014 240000
rect 20350 239200 20406 240000
rect 22742 239200 22798 240000
rect 25134 239200 25190 240000
rect 27526 239200 27582 240000
rect 30010 239200 30066 240000
rect 32402 239200 32458 240000
rect 34794 239200 34850 240000
rect 37186 239200 37242 240000
rect 39578 239200 39634 240000
rect 41970 239200 42026 240000
rect 44362 239200 44418 240000
rect 46754 239200 46810 240000
rect 49146 239200 49202 240000
rect 51538 239200 51594 240000
rect 53930 239200 53986 240000
rect 56414 239200 56470 240000
rect 58806 239200 58862 240000
rect 61198 239200 61254 240000
rect 63590 239200 63646 240000
rect 65982 239200 66038 240000
rect 68374 239200 68430 240000
rect 70766 239200 70822 240000
rect 73158 239200 73214 240000
rect 75550 239200 75606 240000
rect 77942 239200 77998 240000
rect 80334 239200 80390 240000
rect 82818 239200 82874 240000
rect 85210 239200 85266 240000
rect 87602 239200 87658 240000
rect 89994 239200 90050 240000
rect 92386 239200 92442 240000
rect 94778 239200 94834 240000
rect 97170 239200 97226 240000
rect 99562 239200 99618 240000
rect 101954 239200 102010 240000
rect 104346 239200 104402 240000
rect 106738 239200 106794 240000
rect 109222 239200 109278 240000
rect 111614 239200 111670 240000
rect 114006 239200 114062 240000
rect 116398 239200 116454 240000
rect 118790 239200 118846 240000
rect 121182 239200 121238 240000
rect 123574 239200 123630 240000
rect 125966 239200 126022 240000
rect 128358 239200 128414 240000
rect 130750 239200 130806 240000
rect 133142 239200 133198 240000
rect 135626 239200 135682 240000
rect 138018 239200 138074 240000
rect 140410 239200 140466 240000
rect 142802 239200 142858 240000
rect 145194 239200 145250 240000
rect 147586 239200 147642 240000
rect 149978 239200 150034 240000
rect 152370 239200 152426 240000
rect 154762 239200 154818 240000
rect 157154 239200 157210 240000
rect 159546 239200 159602 240000
rect 162030 239200 162086 240000
rect 164422 239200 164478 240000
rect 166814 239200 166870 240000
rect 169206 239200 169262 240000
rect 171598 239200 171654 240000
rect 173990 239200 174046 240000
rect 176382 239200 176438 240000
rect 178774 239200 178830 240000
rect 181166 239200 181222 240000
rect 183558 239200 183614 240000
rect 185950 239200 186006 240000
rect 188434 239200 188490 240000
rect 190826 239200 190882 240000
rect 193218 239200 193274 240000
rect 195610 239200 195666 240000
rect 198002 239200 198058 240000
rect 200394 239200 200450 240000
rect 202786 239200 202842 240000
rect 205178 239200 205234 240000
rect 207570 239200 207626 240000
rect 209962 239200 210018 240000
rect 212354 239200 212410 240000
rect 214838 239200 214894 240000
rect 217230 239200 217286 240000
rect 219622 239200 219678 240000
rect 222014 239200 222070 240000
rect 224406 239200 224462 240000
rect 226798 239200 226854 240000
rect 229190 239200 229246 240000
rect 231582 239200 231638 240000
rect 233974 239200 234030 240000
rect 236366 239200 236422 240000
rect 238758 239200 238814 240000
rect 1122 0 1178 800
rect 3330 0 3386 800
rect 5630 0 5686 800
rect 7930 0 7986 800
rect 10230 0 10286 800
rect 12530 0 12586 800
rect 14830 0 14886 800
rect 17038 0 17094 800
rect 19338 0 19394 800
rect 21638 0 21694 800
rect 23938 0 23994 800
rect 26238 0 26294 800
rect 28538 0 28594 800
rect 30838 0 30894 800
rect 33046 0 33102 800
rect 35346 0 35402 800
rect 37646 0 37702 800
rect 39946 0 40002 800
rect 42246 0 42302 800
rect 44546 0 44602 800
rect 46754 0 46810 800
rect 49054 0 49110 800
rect 51354 0 51410 800
rect 53654 0 53710 800
rect 55954 0 56010 800
rect 58254 0 58310 800
rect 60554 0 60610 800
rect 62762 0 62818 800
rect 65062 0 65118 800
rect 67362 0 67418 800
rect 69662 0 69718 800
rect 71962 0 72018 800
rect 74262 0 74318 800
rect 76470 0 76526 800
rect 78770 0 78826 800
rect 81070 0 81126 800
rect 83370 0 83426 800
rect 85670 0 85726 800
rect 87970 0 88026 800
rect 90270 0 90326 800
rect 92478 0 92534 800
rect 94778 0 94834 800
rect 97078 0 97134 800
rect 99378 0 99434 800
rect 101678 0 101734 800
rect 103978 0 104034 800
rect 106186 0 106242 800
rect 108486 0 108542 800
rect 110786 0 110842 800
rect 113086 0 113142 800
rect 115386 0 115442 800
rect 117686 0 117742 800
rect 119986 0 120042 800
rect 122194 0 122250 800
rect 124494 0 124550 800
rect 126794 0 126850 800
rect 129094 0 129150 800
rect 131394 0 131450 800
rect 133694 0 133750 800
rect 135994 0 136050 800
rect 138202 0 138258 800
rect 140502 0 140558 800
rect 142802 0 142858 800
rect 145102 0 145158 800
rect 147402 0 147458 800
rect 149702 0 149758 800
rect 151910 0 151966 800
rect 154210 0 154266 800
rect 156510 0 156566 800
rect 158810 0 158866 800
rect 161110 0 161166 800
rect 163410 0 163466 800
rect 165710 0 165766 800
rect 167918 0 167974 800
rect 170218 0 170274 800
rect 172518 0 172574 800
rect 174818 0 174874 800
rect 177118 0 177174 800
rect 179418 0 179474 800
rect 181626 0 181682 800
rect 183926 0 183982 800
rect 186226 0 186282 800
rect 188526 0 188582 800
rect 190826 0 190882 800
rect 193126 0 193182 800
rect 195426 0 195482 800
rect 197634 0 197690 800
rect 199934 0 199990 800
rect 202234 0 202290 800
rect 204534 0 204590 800
rect 206834 0 206890 800
rect 209134 0 209190 800
rect 211342 0 211398 800
rect 213642 0 213698 800
rect 215942 0 215998 800
rect 218242 0 218298 800
rect 220542 0 220598 800
rect 222842 0 222898 800
rect 225142 0 225198 800
rect 227350 0 227406 800
rect 229650 0 229706 800
rect 231950 0 232006 800
rect 234250 0 234306 800
rect 236550 0 236606 800
rect 238850 0 238906 800
<< obsm2 >>
rect 20 239144 1158 239306
rect 1326 239144 3550 239306
rect 3718 239144 5942 239306
rect 6110 239144 8334 239306
rect 8502 239144 10726 239306
rect 10894 239144 13118 239306
rect 13286 239144 15510 239306
rect 15678 239144 17902 239306
rect 18070 239144 20294 239306
rect 20462 239144 22686 239306
rect 22854 239144 25078 239306
rect 25246 239144 27470 239306
rect 27638 239144 29954 239306
rect 30122 239144 32346 239306
rect 32514 239144 34738 239306
rect 34906 239144 37130 239306
rect 37298 239144 39522 239306
rect 39690 239144 41914 239306
rect 42082 239144 44306 239306
rect 44474 239144 46698 239306
rect 46866 239144 49090 239306
rect 49258 239144 51482 239306
rect 51650 239144 53874 239306
rect 54042 239144 56358 239306
rect 56526 239144 58750 239306
rect 58918 239144 61142 239306
rect 61310 239144 63534 239306
rect 63702 239144 65926 239306
rect 66094 239144 68318 239306
rect 68486 239144 70710 239306
rect 70878 239144 73102 239306
rect 73270 239144 75494 239306
rect 75662 239144 77886 239306
rect 78054 239144 80278 239306
rect 80446 239144 82762 239306
rect 82930 239144 85154 239306
rect 85322 239144 87546 239306
rect 87714 239144 89938 239306
rect 90106 239144 92330 239306
rect 92498 239144 94722 239306
rect 94890 239144 97114 239306
rect 97282 239144 99506 239306
rect 99674 239144 101898 239306
rect 102066 239144 104290 239306
rect 104458 239144 106682 239306
rect 106850 239144 109166 239306
rect 109334 239144 111558 239306
rect 111726 239144 113950 239306
rect 114118 239144 116342 239306
rect 116510 239144 118734 239306
rect 118902 239144 121126 239306
rect 121294 239144 123518 239306
rect 123686 239144 125910 239306
rect 126078 239144 128302 239306
rect 128470 239144 130694 239306
rect 130862 239144 133086 239306
rect 133254 239144 135570 239306
rect 135738 239144 137962 239306
rect 138130 239144 140354 239306
rect 140522 239144 142746 239306
rect 142914 239144 145138 239306
rect 145306 239144 147530 239306
rect 147698 239144 149922 239306
rect 150090 239144 152314 239306
rect 152482 239144 154706 239306
rect 154874 239144 157098 239306
rect 157266 239144 159490 239306
rect 159658 239144 161974 239306
rect 162142 239144 164366 239306
rect 164534 239144 166758 239306
rect 166926 239144 169150 239306
rect 169318 239144 171542 239306
rect 171710 239144 173934 239306
rect 174102 239144 176326 239306
rect 176494 239144 178718 239306
rect 178886 239144 181110 239306
rect 181278 239144 183502 239306
rect 183670 239144 185894 239306
rect 186062 239144 188378 239306
rect 188546 239144 190770 239306
rect 190938 239144 193162 239306
rect 193330 239144 195554 239306
rect 195722 239144 197946 239306
rect 198114 239144 200338 239306
rect 200506 239144 202730 239306
rect 202898 239144 205122 239306
rect 205290 239144 207514 239306
rect 207682 239144 209906 239306
rect 210074 239144 212298 239306
rect 212466 239144 214782 239306
rect 214950 239144 217174 239306
rect 217342 239144 219566 239306
rect 219734 239144 221958 239306
rect 222126 239144 224350 239306
rect 224518 239144 226742 239306
rect 226910 239144 229134 239306
rect 229302 239144 231526 239306
rect 231694 239144 233918 239306
rect 234086 239144 236310 239306
rect 236478 239144 238702 239306
rect 238870 239144 238904 239306
rect 20 856 238904 239144
rect 20 734 1066 856
rect 1234 734 3274 856
rect 3442 734 5574 856
rect 5742 734 7874 856
rect 8042 734 10174 856
rect 10342 734 12474 856
rect 12642 734 14774 856
rect 14942 734 16982 856
rect 17150 734 19282 856
rect 19450 734 21582 856
rect 21750 734 23882 856
rect 24050 734 26182 856
rect 26350 734 28482 856
rect 28650 734 30782 856
rect 30950 734 32990 856
rect 33158 734 35290 856
rect 35458 734 37590 856
rect 37758 734 39890 856
rect 40058 734 42190 856
rect 42358 734 44490 856
rect 44658 734 46698 856
rect 46866 734 48998 856
rect 49166 734 51298 856
rect 51466 734 53598 856
rect 53766 734 55898 856
rect 56066 734 58198 856
rect 58366 734 60498 856
rect 60666 734 62706 856
rect 62874 734 65006 856
rect 65174 734 67306 856
rect 67474 734 69606 856
rect 69774 734 71906 856
rect 72074 734 74206 856
rect 74374 734 76414 856
rect 76582 734 78714 856
rect 78882 734 81014 856
rect 81182 734 83314 856
rect 83482 734 85614 856
rect 85782 734 87914 856
rect 88082 734 90214 856
rect 90382 734 92422 856
rect 92590 734 94722 856
rect 94890 734 97022 856
rect 97190 734 99322 856
rect 99490 734 101622 856
rect 101790 734 103922 856
rect 104090 734 106130 856
rect 106298 734 108430 856
rect 108598 734 110730 856
rect 110898 734 113030 856
rect 113198 734 115330 856
rect 115498 734 117630 856
rect 117798 734 119930 856
rect 120098 734 122138 856
rect 122306 734 124438 856
rect 124606 734 126738 856
rect 126906 734 129038 856
rect 129206 734 131338 856
rect 131506 734 133638 856
rect 133806 734 135938 856
rect 136106 734 138146 856
rect 138314 734 140446 856
rect 140614 734 142746 856
rect 142914 734 145046 856
rect 145214 734 147346 856
rect 147514 734 149646 856
rect 149814 734 151854 856
rect 152022 734 154154 856
rect 154322 734 156454 856
rect 156622 734 158754 856
rect 158922 734 161054 856
rect 161222 734 163354 856
rect 163522 734 165654 856
rect 165822 734 167862 856
rect 168030 734 170162 856
rect 170330 734 172462 856
rect 172630 734 174762 856
rect 174930 734 177062 856
rect 177230 734 179362 856
rect 179530 734 181570 856
rect 181738 734 183870 856
rect 184038 734 186170 856
rect 186338 734 188470 856
rect 188638 734 190770 856
rect 190938 734 193070 856
rect 193238 734 195370 856
rect 195538 734 197578 856
rect 197746 734 199878 856
rect 200046 734 202178 856
rect 202346 734 204478 856
rect 204646 734 206778 856
rect 206946 734 209078 856
rect 209246 734 211286 856
rect 211454 734 213586 856
rect 213754 734 215886 856
rect 216054 734 218186 856
rect 218354 734 220486 856
rect 220654 734 222786 856
rect 222954 734 225086 856
rect 225254 734 227294 856
rect 227462 734 229594 856
rect 229762 734 231894 856
rect 232062 734 234194 856
rect 234362 734 236494 856
rect 236662 734 238794 856
<< metal3 >>
rect 239200 238824 240000 238944
rect 0 238552 800 238672
rect 239200 236512 240000 236632
rect 0 235968 800 236088
rect 239200 234200 240000 234320
rect 0 233384 800 233504
rect 239200 231888 240000 232008
rect 0 230800 800 230920
rect 239200 229576 240000 229696
rect 0 228216 800 228336
rect 239200 227264 240000 227384
rect 0 225496 800 225616
rect 239200 224952 240000 225072
rect 0 222912 800 223032
rect 239200 222640 240000 222760
rect 0 220328 800 220448
rect 239200 220328 240000 220448
rect 239200 218016 240000 218136
rect 0 217744 800 217864
rect 239200 215704 240000 215824
rect 0 215160 800 215280
rect 239200 213392 240000 213512
rect 0 212440 800 212560
rect 239200 211080 240000 211200
rect 0 209856 800 209976
rect 239200 208768 240000 208888
rect 0 207272 800 207392
rect 239200 206456 240000 206576
rect 0 204688 800 204808
rect 239200 204144 240000 204264
rect 0 202104 800 202224
rect 239200 201832 240000 201952
rect 0 199520 800 199640
rect 239200 199520 240000 199640
rect 239200 197208 240000 197328
rect 0 196800 800 196920
rect 239200 194896 240000 195016
rect 0 194216 800 194336
rect 239200 192584 240000 192704
rect 0 191632 800 191752
rect 239200 190272 240000 190392
rect 0 189048 800 189168
rect 239200 187960 240000 188080
rect 0 186464 800 186584
rect 239200 185648 240000 185768
rect 0 183744 800 183864
rect 239200 183336 240000 183456
rect 0 181160 800 181280
rect 239200 181024 240000 181144
rect 0 178576 800 178696
rect 239200 178712 240000 178832
rect 239200 176400 240000 176520
rect 0 175992 800 176112
rect 239200 174088 240000 174208
rect 0 173408 800 173528
rect 239200 171776 240000 171896
rect 0 170824 800 170944
rect 239200 169464 240000 169584
rect 0 168104 800 168224
rect 239200 167152 240000 167272
rect 0 165520 800 165640
rect 239200 164840 240000 164960
rect 0 162936 800 163056
rect 239200 162528 240000 162648
rect 0 160352 800 160472
rect 239200 160352 240000 160472
rect 239200 158040 240000 158160
rect 0 157768 800 157888
rect 239200 155728 240000 155848
rect 0 155048 800 155168
rect 239200 153416 240000 153536
rect 0 152464 800 152584
rect 239200 151104 240000 151224
rect 0 149880 800 150000
rect 239200 148792 240000 148912
rect 0 147296 800 147416
rect 239200 146480 240000 146600
rect 0 144712 800 144832
rect 239200 144168 240000 144288
rect 0 141992 800 142112
rect 239200 141856 240000 141976
rect 0 139408 800 139528
rect 239200 139544 240000 139664
rect 239200 137232 240000 137352
rect 0 136824 800 136944
rect 239200 134920 240000 135040
rect 0 134240 800 134360
rect 239200 132608 240000 132728
rect 0 131656 800 131776
rect 239200 130296 240000 130416
rect 0 129072 800 129192
rect 239200 127984 240000 128104
rect 0 126352 800 126472
rect 239200 125672 240000 125792
rect 0 123768 800 123888
rect 239200 123360 240000 123480
rect 0 121184 800 121304
rect 239200 121048 240000 121168
rect 0 118600 800 118720
rect 239200 118736 240000 118856
rect 239200 116424 240000 116544
rect 0 116016 800 116136
rect 239200 114112 240000 114232
rect 0 113296 800 113416
rect 239200 111800 240000 111920
rect 0 110712 800 110832
rect 239200 109488 240000 109608
rect 0 108128 800 108248
rect 239200 107176 240000 107296
rect 0 105544 800 105664
rect 239200 104864 240000 104984
rect 0 102960 800 103080
rect 239200 102552 240000 102672
rect 0 100376 800 100496
rect 239200 100240 240000 100360
rect 239200 97928 240000 98048
rect 0 97656 800 97776
rect 239200 95616 240000 95736
rect 0 95072 800 95192
rect 239200 93304 240000 93424
rect 0 92488 800 92608
rect 239200 90992 240000 91112
rect 0 89904 800 90024
rect 239200 88680 240000 88800
rect 0 87320 800 87440
rect 239200 86368 240000 86488
rect 0 84600 800 84720
rect 239200 84056 240000 84176
rect 0 82016 800 82136
rect 239200 81744 240000 81864
rect 0 79432 800 79552
rect 239200 79568 240000 79688
rect 239200 77256 240000 77376
rect 0 76848 800 76968
rect 239200 74944 240000 75064
rect 0 74264 800 74384
rect 239200 72632 240000 72752
rect 0 71544 800 71664
rect 239200 70320 240000 70440
rect 0 68960 800 69080
rect 239200 68008 240000 68128
rect 0 66376 800 66496
rect 239200 65696 240000 65816
rect 0 63792 800 63912
rect 239200 63384 240000 63504
rect 0 61208 800 61328
rect 239200 61072 240000 61192
rect 0 58624 800 58744
rect 239200 58760 240000 58880
rect 239200 56448 240000 56568
rect 0 55904 800 56024
rect 239200 54136 240000 54256
rect 0 53320 800 53440
rect 239200 51824 240000 51944
rect 0 50736 800 50856
rect 239200 49512 240000 49632
rect 0 48152 800 48272
rect 239200 47200 240000 47320
rect 0 45568 800 45688
rect 239200 44888 240000 45008
rect 0 42848 800 42968
rect 239200 42576 240000 42696
rect 0 40264 800 40384
rect 239200 40264 240000 40384
rect 239200 37952 240000 38072
rect 0 37680 800 37800
rect 239200 35640 240000 35760
rect 0 35096 800 35216
rect 239200 33328 240000 33448
rect 0 32512 800 32632
rect 239200 31016 240000 31136
rect 0 29928 800 30048
rect 239200 28704 240000 28824
rect 0 27208 800 27328
rect 239200 26392 240000 26512
rect 0 24624 800 24744
rect 239200 24080 240000 24200
rect 0 22040 800 22160
rect 239200 21768 240000 21888
rect 0 19456 800 19576
rect 239200 19456 240000 19576
rect 239200 17144 240000 17264
rect 0 16872 800 16992
rect 239200 14832 240000 14952
rect 0 14152 800 14272
rect 239200 12520 240000 12640
rect 0 11568 800 11688
rect 239200 10208 240000 10328
rect 0 8984 800 9104
rect 239200 7896 240000 8016
rect 0 6400 800 6520
rect 239200 5584 240000 5704
rect 0 3816 800 3936
rect 239200 3272 240000 3392
rect 0 1232 800 1352
rect 239200 1096 240000 1216
<< obsm3 >>
rect 800 238752 239120 238917
rect 880 238744 239120 238752
rect 880 238472 239322 238744
rect 800 236712 239322 238472
rect 800 236432 239120 236712
rect 800 236168 239322 236432
rect 880 235888 239322 236168
rect 800 234400 239322 235888
rect 800 234120 239120 234400
rect 800 233584 239322 234120
rect 880 233304 239322 233584
rect 800 232088 239322 233304
rect 800 231808 239120 232088
rect 800 231000 239322 231808
rect 880 230720 239322 231000
rect 800 229776 239322 230720
rect 800 229496 239120 229776
rect 800 228416 239322 229496
rect 880 228136 239322 228416
rect 800 227464 239322 228136
rect 800 227184 239120 227464
rect 800 225696 239322 227184
rect 880 225416 239322 225696
rect 800 225152 239322 225416
rect 800 224872 239120 225152
rect 800 223112 239322 224872
rect 880 222840 239322 223112
rect 880 222832 239120 222840
rect 800 222560 239120 222832
rect 800 220528 239322 222560
rect 880 220248 239120 220528
rect 800 218216 239322 220248
rect 800 217944 239120 218216
rect 880 217936 239120 217944
rect 880 217664 239322 217936
rect 800 215904 239322 217664
rect 800 215624 239120 215904
rect 800 215360 239322 215624
rect 880 215080 239322 215360
rect 800 213592 239322 215080
rect 800 213312 239120 213592
rect 800 212640 239322 213312
rect 880 212360 239322 212640
rect 800 211280 239322 212360
rect 800 211000 239120 211280
rect 800 210056 239322 211000
rect 880 209776 239322 210056
rect 800 208968 239322 209776
rect 800 208688 239120 208968
rect 800 207472 239322 208688
rect 880 207192 239322 207472
rect 800 206656 239322 207192
rect 800 206376 239120 206656
rect 800 204888 239322 206376
rect 880 204608 239322 204888
rect 800 204344 239322 204608
rect 800 204064 239120 204344
rect 800 202304 239322 204064
rect 880 202032 239322 202304
rect 880 202024 239120 202032
rect 800 201752 239120 202024
rect 800 199720 239322 201752
rect 880 199440 239120 199720
rect 800 197408 239322 199440
rect 800 197128 239120 197408
rect 800 197000 239322 197128
rect 880 196720 239322 197000
rect 800 195096 239322 196720
rect 800 194816 239120 195096
rect 800 194416 239322 194816
rect 880 194136 239322 194416
rect 800 192784 239322 194136
rect 800 192504 239120 192784
rect 800 191832 239322 192504
rect 880 191552 239322 191832
rect 800 190472 239322 191552
rect 800 190192 239120 190472
rect 800 189248 239322 190192
rect 880 188968 239322 189248
rect 800 188160 239322 188968
rect 800 187880 239120 188160
rect 800 186664 239322 187880
rect 880 186384 239322 186664
rect 800 185848 239322 186384
rect 800 185568 239120 185848
rect 800 183944 239322 185568
rect 880 183664 239322 183944
rect 800 183536 239322 183664
rect 800 183256 239120 183536
rect 800 181360 239322 183256
rect 880 181224 239322 181360
rect 880 181080 239120 181224
rect 800 180944 239120 181080
rect 800 178912 239322 180944
rect 800 178776 239120 178912
rect 880 178632 239120 178776
rect 880 178496 239322 178632
rect 800 176600 239322 178496
rect 800 176320 239120 176600
rect 800 176192 239322 176320
rect 880 175912 239322 176192
rect 800 174288 239322 175912
rect 800 174008 239120 174288
rect 800 173608 239322 174008
rect 880 173328 239322 173608
rect 800 171976 239322 173328
rect 800 171696 239120 171976
rect 800 171024 239322 171696
rect 880 170744 239322 171024
rect 800 169664 239322 170744
rect 800 169384 239120 169664
rect 800 168304 239322 169384
rect 880 168024 239322 168304
rect 800 167352 239322 168024
rect 800 167072 239120 167352
rect 800 165720 239322 167072
rect 880 165440 239322 165720
rect 800 165040 239322 165440
rect 800 164760 239120 165040
rect 800 163136 239322 164760
rect 880 162856 239322 163136
rect 800 162728 239322 162856
rect 800 162448 239120 162728
rect 800 160552 239322 162448
rect 880 160272 239120 160552
rect 800 158240 239322 160272
rect 800 157968 239120 158240
rect 880 157960 239120 157968
rect 880 157688 239322 157960
rect 800 155928 239322 157688
rect 800 155648 239120 155928
rect 800 155248 239322 155648
rect 880 154968 239322 155248
rect 800 153616 239322 154968
rect 800 153336 239120 153616
rect 800 152664 239322 153336
rect 880 152384 239322 152664
rect 800 151304 239322 152384
rect 800 151024 239120 151304
rect 800 150080 239322 151024
rect 880 149800 239322 150080
rect 800 148992 239322 149800
rect 800 148712 239120 148992
rect 800 147496 239322 148712
rect 880 147216 239322 147496
rect 800 146680 239322 147216
rect 800 146400 239120 146680
rect 800 144912 239322 146400
rect 880 144632 239322 144912
rect 800 144368 239322 144632
rect 800 144088 239120 144368
rect 800 142192 239322 144088
rect 880 142056 239322 142192
rect 880 141912 239120 142056
rect 800 141776 239120 141912
rect 800 139744 239322 141776
rect 800 139608 239120 139744
rect 880 139464 239120 139608
rect 880 139328 239322 139464
rect 800 137432 239322 139328
rect 800 137152 239120 137432
rect 800 137024 239322 137152
rect 880 136744 239322 137024
rect 800 135120 239322 136744
rect 800 134840 239120 135120
rect 800 134440 239322 134840
rect 880 134160 239322 134440
rect 800 132808 239322 134160
rect 800 132528 239120 132808
rect 800 131856 239322 132528
rect 880 131576 239322 131856
rect 800 130496 239322 131576
rect 800 130216 239120 130496
rect 800 129272 239322 130216
rect 880 128992 239322 129272
rect 800 128184 239322 128992
rect 800 127904 239120 128184
rect 800 126552 239322 127904
rect 880 126272 239322 126552
rect 800 125872 239322 126272
rect 800 125592 239120 125872
rect 800 123968 239322 125592
rect 880 123688 239322 123968
rect 800 123560 239322 123688
rect 800 123280 239120 123560
rect 800 121384 239322 123280
rect 880 121248 239322 121384
rect 880 121104 239120 121248
rect 800 120968 239120 121104
rect 800 118936 239322 120968
rect 800 118800 239120 118936
rect 880 118656 239120 118800
rect 880 118520 239322 118656
rect 800 116624 239322 118520
rect 800 116344 239120 116624
rect 800 116216 239322 116344
rect 880 115936 239322 116216
rect 800 114312 239322 115936
rect 800 114032 239120 114312
rect 800 113496 239322 114032
rect 880 113216 239322 113496
rect 800 112000 239322 113216
rect 800 111720 239120 112000
rect 800 110912 239322 111720
rect 880 110632 239322 110912
rect 800 109688 239322 110632
rect 800 109408 239120 109688
rect 800 108328 239322 109408
rect 880 108048 239322 108328
rect 800 107376 239322 108048
rect 800 107096 239120 107376
rect 800 105744 239322 107096
rect 880 105464 239322 105744
rect 800 105064 239322 105464
rect 800 104784 239120 105064
rect 800 103160 239322 104784
rect 880 102880 239322 103160
rect 800 102752 239322 102880
rect 800 102472 239120 102752
rect 800 100576 239322 102472
rect 880 100440 239322 100576
rect 880 100296 239120 100440
rect 800 100160 239120 100296
rect 800 98128 239322 100160
rect 800 97856 239120 98128
rect 880 97848 239120 97856
rect 880 97576 239322 97848
rect 800 95816 239322 97576
rect 800 95536 239120 95816
rect 800 95272 239322 95536
rect 880 94992 239322 95272
rect 800 93504 239322 94992
rect 800 93224 239120 93504
rect 800 92688 239322 93224
rect 880 92408 239322 92688
rect 800 91192 239322 92408
rect 800 90912 239120 91192
rect 800 90104 239322 90912
rect 880 89824 239322 90104
rect 800 88880 239322 89824
rect 800 88600 239120 88880
rect 800 87520 239322 88600
rect 880 87240 239322 87520
rect 800 86568 239322 87240
rect 800 86288 239120 86568
rect 800 84800 239322 86288
rect 880 84520 239322 84800
rect 800 84256 239322 84520
rect 800 83976 239120 84256
rect 800 82216 239322 83976
rect 880 81944 239322 82216
rect 880 81936 239120 81944
rect 800 81664 239120 81936
rect 800 79768 239322 81664
rect 800 79632 239120 79768
rect 880 79488 239120 79632
rect 880 79352 239322 79488
rect 800 77456 239322 79352
rect 800 77176 239120 77456
rect 800 77048 239322 77176
rect 880 76768 239322 77048
rect 800 75144 239322 76768
rect 800 74864 239120 75144
rect 800 74464 239322 74864
rect 880 74184 239322 74464
rect 800 72832 239322 74184
rect 800 72552 239120 72832
rect 800 71744 239322 72552
rect 880 71464 239322 71744
rect 800 70520 239322 71464
rect 800 70240 239120 70520
rect 800 69160 239322 70240
rect 880 68880 239322 69160
rect 800 68208 239322 68880
rect 800 67928 239120 68208
rect 800 66576 239322 67928
rect 880 66296 239322 66576
rect 800 65896 239322 66296
rect 800 65616 239120 65896
rect 800 63992 239322 65616
rect 880 63712 239322 63992
rect 800 63584 239322 63712
rect 800 63304 239120 63584
rect 800 61408 239322 63304
rect 880 61272 239322 61408
rect 880 61128 239120 61272
rect 800 60992 239120 61128
rect 800 58960 239322 60992
rect 800 58824 239120 58960
rect 880 58680 239120 58824
rect 880 58544 239322 58680
rect 800 56648 239322 58544
rect 800 56368 239120 56648
rect 800 56104 239322 56368
rect 880 55824 239322 56104
rect 800 54336 239322 55824
rect 800 54056 239120 54336
rect 800 53520 239322 54056
rect 880 53240 239322 53520
rect 800 52024 239322 53240
rect 800 51744 239120 52024
rect 800 50936 239322 51744
rect 880 50656 239322 50936
rect 800 49712 239322 50656
rect 800 49432 239120 49712
rect 800 48352 239322 49432
rect 880 48072 239322 48352
rect 800 47400 239322 48072
rect 800 47120 239120 47400
rect 800 45768 239322 47120
rect 880 45488 239322 45768
rect 800 45088 239322 45488
rect 800 44808 239120 45088
rect 800 43048 239322 44808
rect 880 42776 239322 43048
rect 880 42768 239120 42776
rect 800 42496 239120 42768
rect 800 40464 239322 42496
rect 880 40184 239120 40464
rect 800 38152 239322 40184
rect 800 37880 239120 38152
rect 880 37872 239120 37880
rect 880 37600 239322 37872
rect 800 35840 239322 37600
rect 800 35560 239120 35840
rect 800 35296 239322 35560
rect 880 35016 239322 35296
rect 800 33528 239322 35016
rect 800 33248 239120 33528
rect 800 32712 239322 33248
rect 880 32432 239322 32712
rect 800 31216 239322 32432
rect 800 30936 239120 31216
rect 800 30128 239322 30936
rect 880 29848 239322 30128
rect 800 28904 239322 29848
rect 800 28624 239120 28904
rect 800 27408 239322 28624
rect 880 27128 239322 27408
rect 800 26592 239322 27128
rect 800 26312 239120 26592
rect 800 24824 239322 26312
rect 880 24544 239322 24824
rect 800 24280 239322 24544
rect 800 24000 239120 24280
rect 800 22240 239322 24000
rect 880 21968 239322 22240
rect 880 21960 239120 21968
rect 800 21688 239120 21960
rect 800 19656 239322 21688
rect 880 19376 239120 19656
rect 800 17344 239322 19376
rect 800 17072 239120 17344
rect 880 17064 239120 17072
rect 880 16792 239322 17064
rect 800 15032 239322 16792
rect 800 14752 239120 15032
rect 800 14352 239322 14752
rect 880 14072 239322 14352
rect 800 12720 239322 14072
rect 800 12440 239120 12720
rect 800 11768 239322 12440
rect 880 11488 239322 11768
rect 800 10408 239322 11488
rect 800 10128 239120 10408
rect 800 9184 239322 10128
rect 880 8904 239322 9184
rect 800 8096 239322 8904
rect 800 7816 239120 8096
rect 800 6600 239322 7816
rect 880 6320 239322 6600
rect 800 5784 239322 6320
rect 800 5504 239120 5784
rect 800 4016 239322 5504
rect 880 3736 239322 4016
rect 800 3472 239322 3736
rect 800 3192 239120 3472
rect 800 1432 239322 3192
rect 880 1296 239322 1432
rect 880 1152 239120 1296
rect 800 1123 239120 1152
<< metal4 >>
rect 4208 2128 4528 237776
rect 9208 2128 9528 237776
rect 14208 2128 14528 237776
rect 19208 2128 19528 237776
rect 24208 2128 24528 237776
rect 29208 2128 29528 237776
rect 34208 2128 34528 237776
rect 39208 2128 39528 237776
rect 44208 2128 44528 237776
rect 49208 2128 49528 237776
rect 54208 2128 54528 237776
rect 59208 2128 59528 237776
rect 64208 2128 64528 237776
rect 69208 2128 69528 237776
rect 74208 2128 74528 237776
rect 79208 2128 79528 237776
rect 84208 2128 84528 237776
rect 89208 2128 89528 237776
rect 94208 2128 94528 237776
rect 99208 2128 99528 237776
rect 104208 2128 104528 237776
rect 109208 2128 109528 237776
rect 114208 2128 114528 237776
rect 119208 2128 119528 237776
rect 124208 2128 124528 237776
rect 129208 2128 129528 237776
rect 134208 2128 134528 237776
rect 139208 2128 139528 237776
rect 144208 2128 144528 237776
rect 149208 2128 149528 237776
rect 154208 2128 154528 237776
rect 159208 2128 159528 237776
rect 164208 2128 164528 237776
rect 169208 2128 169528 237776
rect 174208 2128 174528 237776
rect 179208 2128 179528 237776
rect 184208 2128 184528 237776
rect 189208 2128 189528 237776
rect 194208 2128 194528 237776
rect 199208 2128 199528 237776
rect 204208 2128 204528 237776
rect 209208 2128 209528 237776
rect 214208 2128 214528 237776
rect 219208 2128 219528 237776
rect 224208 2128 224528 237776
rect 229208 2128 229528 237776
rect 234208 2128 234528 237776
<< obsm4 >>
rect 35571 25467 39128 206957
rect 39608 25467 44128 206957
rect 44608 25467 49128 206957
rect 49608 25467 54128 206957
rect 54608 25467 59128 206957
rect 59608 25467 64128 206957
rect 64608 25467 69128 206957
rect 69608 25467 74128 206957
rect 74608 25467 79128 206957
rect 79608 25467 84128 206957
rect 84608 25467 89128 206957
rect 89608 25467 94128 206957
rect 94608 25467 99128 206957
rect 99608 25467 104128 206957
rect 104608 25467 109128 206957
rect 109608 25467 114128 206957
rect 114608 25467 119128 206957
rect 119608 25467 124128 206957
rect 124608 25467 129128 206957
rect 129608 25467 134128 206957
rect 134608 25467 139128 206957
rect 139608 25467 144128 206957
rect 144608 25467 149128 206957
rect 149608 25467 154128 206957
rect 154608 25467 159128 206957
rect 159608 25467 163885 206957
<< labels >>
rlabel metal3 s 239200 14832 240000 14952 6 boot_addr_i[0]
port 1 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 boot_addr_i[10]
port 2 nsew signal input
rlabel metal2 s 85210 239200 85266 240000 6 boot_addr_i[11]
port 3 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 boot_addr_i[12]
port 4 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 boot_addr_i[13]
port 5 nsew signal input
rlabel metal2 s 109222 239200 109278 240000 6 boot_addr_i[14]
port 6 nsew signal input
rlabel metal3 s 239200 121048 240000 121168 6 boot_addr_i[15]
port 7 nsew signal input
rlabel metal2 s 135626 239200 135682 240000 6 boot_addr_i[16]
port 8 nsew signal input
rlabel metal3 s 239200 134920 240000 135040 6 boot_addr_i[17]
port 9 nsew signal input
rlabel metal2 s 142802 239200 142858 240000 6 boot_addr_i[18]
port 10 nsew signal input
rlabel metal3 s 0 144712 800 144832 6 boot_addr_i[19]
port 11 nsew signal input
rlabel metal3 s 239200 26392 240000 26512 6 boot_addr_i[1]
port 12 nsew signal input
rlabel metal2 s 177118 0 177174 800 6 boot_addr_i[20]
port 13 nsew signal input
rlabel metal2 s 164422 239200 164478 240000 6 boot_addr_i[21]
port 14 nsew signal input
rlabel metal3 s 0 162936 800 163056 6 boot_addr_i[22]
port 15 nsew signal input
rlabel metal2 s 181166 239200 181222 240000 6 boot_addr_i[23]
port 16 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 boot_addr_i[24]
port 17 nsew signal input
rlabel metal2 s 193218 239200 193274 240000 6 boot_addr_i[25]
port 18 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 boot_addr_i[26]
port 19 nsew signal input
rlabel metal3 s 239200 208768 240000 208888 6 boot_addr_i[27]
port 20 nsew signal input
rlabel metal3 s 0 217744 800 217864 6 boot_addr_i[28]
port 21 nsew signal input
rlabel metal3 s 0 228216 800 228336 6 boot_addr_i[29]
port 22 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 boot_addr_i[2]
port 23 nsew signal input
rlabel metal2 s 229650 0 229706 800 6 boot_addr_i[30]
port 24 nsew signal input
rlabel metal2 s 226798 239200 226854 240000 6 boot_addr_i[31]
port 25 nsew signal input
rlabel metal3 s 239200 35640 240000 35760 6 boot_addr_i[3]
port 26 nsew signal input
rlabel metal3 s 239200 49512 240000 49632 6 boot_addr_i[4]
port 27 nsew signal input
rlabel metal2 s 49146 239200 49202 240000 6 boot_addr_i[5]
port 28 nsew signal input
rlabel metal3 s 239200 68008 240000 68128 6 boot_addr_i[6]
port 29 nsew signal input
rlabel metal3 s 239200 79568 240000 79688 6 boot_addr_i[7]
port 30 nsew signal input
rlabel metal2 s 80334 239200 80390 240000 6 boot_addr_i[8]
port 31 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 boot_addr_i[9]
port 32 nsew signal input
rlabel metal3 s 239200 1096 240000 1216 6 clk_i
port 33 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 cluster_id_i[0]
port 34 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 cluster_id_i[1]
port 35 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 cluster_id_i[2]
port 36 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 cluster_id_i[3]
port 37 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 cluster_id_i[4]
port 38 nsew signal input
rlabel metal2 s 51538 239200 51594 240000 6 cluster_id_i[5]
port 39 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 core_id_i[0]
port 40 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 core_id_i[1]
port 41 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 core_id_i[2]
port 42 nsew signal input
rlabel metal2 s 37186 239200 37242 240000 6 core_id_i[3]
port 43 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 data_addr_o[0]
port 44 nsew signal output
rlabel metal2 s 82818 239200 82874 240000 6 data_addr_o[10]
port 45 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 data_addr_o[11]
port 46 nsew signal output
rlabel metal2 s 92386 239200 92442 240000 6 data_addr_o[12]
port 47 nsew signal output
rlabel metal2 s 99562 239200 99618 240000 6 data_addr_o[13]
port 48 nsew signal output
rlabel metal3 s 239200 116424 240000 116544 6 data_addr_o[14]
port 49 nsew signal output
rlabel metal2 s 123574 239200 123630 240000 6 data_addr_o[15]
port 50 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 data_addr_o[16]
port 51 nsew signal output
rlabel metal2 s 158810 0 158866 800 6 data_addr_o[17]
port 52 nsew signal output
rlabel metal2 s 145194 239200 145250 240000 6 data_addr_o[18]
port 53 nsew signal output
rlabel metal3 s 0 147296 800 147416 6 data_addr_o[19]
port 54 nsew signal output
rlabel metal2 s 15566 239200 15622 240000 6 data_addr_o[1]
port 55 nsew signal output
rlabel metal2 s 157154 239200 157210 240000 6 data_addr_o[20]
port 56 nsew signal output
rlabel metal3 s 239200 162528 240000 162648 6 data_addr_o[21]
port 57 nsew signal output
rlabel metal2 s 171598 239200 171654 240000 6 data_addr_o[22]
port 58 nsew signal output
rlabel metal3 s 0 173408 800 173528 6 data_addr_o[23]
port 59 nsew signal output
rlabel metal2 s 190826 239200 190882 240000 6 data_addr_o[24]
port 60 nsew signal output
rlabel metal3 s 239200 197208 240000 197328 6 data_addr_o[25]
port 61 nsew signal output
rlabel metal3 s 0 202104 800 202224 6 data_addr_o[26]
port 62 nsew signal output
rlabel metal3 s 239200 211080 240000 211200 6 data_addr_o[27]
port 63 nsew signal output
rlabel metal3 s 0 220328 800 220448 6 data_addr_o[28]
port 64 nsew signal output
rlabel metal2 s 218242 0 218298 800 6 data_addr_o[29]
port 65 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 data_addr_o[2]
port 66 nsew signal output
rlabel metal3 s 0 230800 800 230920 6 data_addr_o[30]
port 67 nsew signal output
rlabel metal3 s 239200 234200 240000 234320 6 data_addr_o[31]
port 68 nsew signal output
rlabel metal3 s 239200 37952 240000 38072 6 data_addr_o[3]
port 69 nsew signal output
rlabel metal3 s 239200 51824 240000 51944 6 data_addr_o[4]
port 70 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 data_addr_o[5]
port 71 nsew signal output
rlabel metal2 s 63590 239200 63646 240000 6 data_addr_o[6]
port 72 nsew signal output
rlabel metal3 s 239200 81744 240000 81864 6 data_addr_o[7]
port 73 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 data_addr_o[8]
port 74 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 data_addr_o[9]
port 75 nsew signal output
rlabel metal2 s 8390 239200 8446 240000 6 data_be_o[0]
port 76 nsew signal output
rlabel metal2 s 17958 239200 18014 240000 6 data_be_o[1]
port 77 nsew signal output
rlabel metal2 s 27526 239200 27582 240000 6 data_be_o[2]
port 78 nsew signal output
rlabel metal3 s 239200 40264 240000 40384 6 data_be_o[3]
port 79 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 data_err_i
port 80 nsew signal input
rlabel metal3 s 0 1232 800 1352 6 data_gnt_i
port 81 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 data_rdata_i[0]
port 82 nsew signal input
rlabel metal3 s 239200 102552 240000 102672 6 data_rdata_i[10]
port 83 nsew signal input
rlabel metal3 s 239200 107176 240000 107296 6 data_rdata_i[11]
port 84 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 data_rdata_i[12]
port 85 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 data_rdata_i[13]
port 86 nsew signal input
rlabel metal2 s 111614 239200 111670 240000 6 data_rdata_i[14]
port 87 nsew signal input
rlabel metal2 s 125966 239200 126022 240000 6 data_rdata_i[15]
port 88 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 data_rdata_i[16]
port 89 nsew signal input
rlabel metal3 s 239200 137232 240000 137352 6 data_rdata_i[17]
port 90 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 data_rdata_i[18]
port 91 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 data_rdata_i[19]
port 92 nsew signal input
rlabel metal2 s 20350 239200 20406 240000 6 data_rdata_i[1]
port 93 nsew signal input
rlabel metal3 s 0 155048 800 155168 6 data_rdata_i[20]
port 94 nsew signal input
rlabel metal2 s 166814 239200 166870 240000 6 data_rdata_i[21]
port 95 nsew signal input
rlabel metal3 s 239200 178712 240000 178832 6 data_rdata_i[22]
port 96 nsew signal input
rlabel metal3 s 0 175992 800 176112 6 data_rdata_i[23]
port 97 nsew signal input
rlabel metal3 s 0 186464 800 186584 6 data_rdata_i[24]
port 98 nsew signal input
rlabel metal3 s 239200 199520 240000 199640 6 data_rdata_i[25]
port 99 nsew signal input
rlabel metal3 s 0 204688 800 204808 6 data_rdata_i[26]
port 100 nsew signal input
rlabel metal3 s 0 215160 800 215280 6 data_rdata_i[27]
port 101 nsew signal input
rlabel metal3 s 239200 218016 240000 218136 6 data_rdata_i[28]
port 102 nsew signal input
rlabel metal2 s 212354 239200 212410 240000 6 data_rdata_i[29]
port 103 nsew signal input
rlabel metal2 s 30010 239200 30066 240000 6 data_rdata_i[2]
port 104 nsew signal input
rlabel metal2 s 219622 239200 219678 240000 6 data_rdata_i[30]
port 105 nsew signal input
rlabel metal3 s 239200 236512 240000 236632 6 data_rdata_i[31]
port 106 nsew signal input
rlabel metal3 s 239200 42576 240000 42696 6 data_rdata_i[3]
port 107 nsew signal input
rlabel metal3 s 239200 54136 240000 54256 6 data_rdata_i[4]
port 108 nsew signal input
rlabel metal2 s 53930 239200 53986 240000 6 data_rdata_i[5]
port 109 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 data_rdata_i[6]
port 110 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 data_rdata_i[7]
port 111 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 data_rdata_i[8]
port 112 nsew signal input
rlabel metal3 s 239200 93304 240000 93424 6 data_rdata_i[9]
port 113 nsew signal input
rlabel metal3 s 239200 3272 240000 3392 6 data_req_o
port 114 nsew signal output
rlabel metal3 s 239200 5584 240000 5704 6 data_rvalid_i
port 115 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 data_wdata_o[0]
port 116 nsew signal output
rlabel metal2 s 126794 0 126850 800 6 data_wdata_o[10]
port 117 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 data_wdata_o[11]
port 118 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 data_wdata_o[12]
port 119 nsew signal output
rlabel metal2 s 101954 239200 102010 240000 6 data_wdata_o[13]
port 120 nsew signal output
rlabel metal2 s 114006 239200 114062 240000 6 data_wdata_o[14]
port 121 nsew signal output
rlabel metal2 s 128358 239200 128414 240000 6 data_wdata_o[15]
port 122 nsew signal output
rlabel metal3 s 239200 125672 240000 125792 6 data_wdata_o[16]
port 123 nsew signal output
rlabel metal3 s 239200 139544 240000 139664 6 data_wdata_o[17]
port 124 nsew signal output
rlabel metal2 s 163410 0 163466 800 6 data_wdata_o[18]
port 125 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 data_wdata_o[19]
port 126 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 data_wdata_o[1]
port 127 nsew signal output
rlabel metal2 s 159546 239200 159602 240000 6 data_wdata_o[20]
port 128 nsew signal output
rlabel metal3 s 239200 164840 240000 164960 6 data_wdata_o[21]
port 129 nsew signal output
rlabel metal2 s 173990 239200 174046 240000 6 data_wdata_o[22]
port 130 nsew signal output
rlabel metal2 s 183558 239200 183614 240000 6 data_wdata_o[23]
port 131 nsew signal output
rlabel metal3 s 0 189048 800 189168 6 data_wdata_o[24]
port 132 nsew signal output
rlabel metal2 s 193126 0 193182 800 6 data_wdata_o[25]
port 133 nsew signal output
rlabel metal3 s 0 207272 800 207392 6 data_wdata_o[26]
port 134 nsew signal output
rlabel metal2 s 209134 0 209190 800 6 data_wdata_o[27]
port 135 nsew signal output
rlabel metal3 s 0 222912 800 223032 6 data_wdata_o[28]
port 136 nsew signal output
rlabel metal2 s 220542 0 220598 800 6 data_wdata_o[29]
port 137 nsew signal output
rlabel metal2 s 32402 239200 32458 240000 6 data_wdata_o[2]
port 138 nsew signal output
rlabel metal2 s 231950 0 232006 800 6 data_wdata_o[30]
port 139 nsew signal output
rlabel metal2 s 229190 239200 229246 240000 6 data_wdata_o[31]
port 140 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 data_wdata_o[3]
port 141 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 data_wdata_o[4]
port 142 nsew signal output
rlabel metal2 s 56414 239200 56470 240000 6 data_wdata_o[5]
port 143 nsew signal output
rlabel metal3 s 0 55904 800 56024 6 data_wdata_o[6]
port 144 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 data_wdata_o[7]
port 145 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 data_wdata_o[8]
port 146 nsew signal output
rlabel metal2 s 113086 0 113142 800 6 data_wdata_o[9]
port 147 nsew signal output
rlabel metal2 s 1214 239200 1270 240000 6 data_we_o
port 148 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 debug_req_i
port 149 nsew signal input
rlabel metal2 s 10782 239200 10838 240000 6 eFPGA_delay_o[0]
port 150 nsew signal output
rlabel metal2 s 22742 239200 22798 240000 6 eFPGA_delay_o[1]
port 151 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 eFPGA_delay_o[2]
port 152 nsew signal output
rlabel metal2 s 39578 239200 39634 240000 6 eFPGA_delay_o[3]
port 153 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 eFPGA_en_o
port 154 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 eFPGA_fpga_done_i
port 155 nsew signal input
rlabel metal3 s 239200 17144 240000 17264 6 eFPGA_operand_a_o[0]
port 156 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 eFPGA_operand_a_o[10]
port 157 nsew signal output
rlabel metal3 s 239200 109488 240000 109608 6 eFPGA_operand_a_o[11]
port 158 nsew signal output
rlabel metal2 s 142802 0 142858 800 6 eFPGA_operand_a_o[12]
port 159 nsew signal output
rlabel metal3 s 0 102960 800 103080 6 eFPGA_operand_a_o[13]
port 160 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 eFPGA_operand_a_o[14]
port 161 nsew signal output
rlabel metal3 s 0 118600 800 118720 6 eFPGA_operand_a_o[15]
port 162 nsew signal output
rlabel metal2 s 138018 239200 138074 240000 6 eFPGA_operand_a_o[16]
port 163 nsew signal output
rlabel metal3 s 239200 141856 240000 141976 6 eFPGA_operand_a_o[17]
port 164 nsew signal output
rlabel metal3 s 0 141992 800 142112 6 eFPGA_operand_a_o[18]
port 165 nsew signal output
rlabel metal3 s 239200 153416 240000 153536 6 eFPGA_operand_a_o[19]
port 166 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 eFPGA_operand_a_o[1]
port 167 nsew signal output
rlabel metal2 s 179418 0 179474 800 6 eFPGA_operand_a_o[20]
port 168 nsew signal output
rlabel metal3 s 239200 167152 240000 167272 6 eFPGA_operand_a_o[21]
port 169 nsew signal output
rlabel metal3 s 0 165520 800 165640 6 eFPGA_operand_a_o[22]
port 170 nsew signal output
rlabel metal3 s 239200 185648 240000 185768 6 eFPGA_operand_a_o[23]
port 171 nsew signal output
rlabel metal3 s 239200 187960 240000 188080 6 eFPGA_operand_a_o[24]
port 172 nsew signal output
rlabel metal2 s 195426 0 195482 800 6 eFPGA_operand_a_o[25]
port 173 nsew signal output
rlabel metal3 s 0 209856 800 209976 6 eFPGA_operand_a_o[26]
port 174 nsew signal output
rlabel metal3 s 239200 213392 240000 213512 6 eFPGA_operand_a_o[27]
port 175 nsew signal output
rlabel metal2 s 207570 239200 207626 240000 6 eFPGA_operand_a_o[28]
port 176 nsew signal output
rlabel metal2 s 214838 239200 214894 240000 6 eFPGA_operand_a_o[29]
port 177 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 eFPGA_operand_a_o[2]
port 178 nsew signal output
rlabel metal2 s 234250 0 234306 800 6 eFPGA_operand_a_o[30]
port 179 nsew signal output
rlabel metal3 s 0 235968 800 236088 6 eFPGA_operand_a_o[31]
port 180 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 eFPGA_operand_a_o[3]
port 181 nsew signal output
rlabel metal3 s 239200 56448 240000 56568 6 eFPGA_operand_a_o[4]
port 182 nsew signal output
rlabel metal3 s 239200 65696 240000 65816 6 eFPGA_operand_a_o[5]
port 183 nsew signal output
rlabel metal2 s 65982 239200 66038 240000 6 eFPGA_operand_a_o[6]
port 184 nsew signal output
rlabel metal3 s 0 63792 800 63912 6 eFPGA_operand_a_o[7]
port 185 nsew signal output
rlabel metal3 s 239200 88680 240000 88800 6 eFPGA_operand_a_o[8]
port 186 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 eFPGA_operand_a_o[9]
port 187 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 eFPGA_operand_b_o[0]
port 188 nsew signal output
rlabel metal3 s 239200 104864 240000 104984 6 eFPGA_operand_b_o[10]
port 189 nsew signal output
rlabel metal2 s 87602 239200 87658 240000 6 eFPGA_operand_b_o[11]
port 190 nsew signal output
rlabel metal3 s 239200 114112 240000 114232 6 eFPGA_operand_b_o[12]
port 191 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 eFPGA_operand_b_o[13]
port 192 nsew signal output
rlabel metal3 s 239200 118736 240000 118856 6 eFPGA_operand_b_o[14]
port 193 nsew signal output
rlabel metal3 s 239200 123360 240000 123480 6 eFPGA_operand_b_o[15]
port 194 nsew signal output
rlabel metal2 s 140410 239200 140466 240000 6 eFPGA_operand_b_o[16]
port 195 nsew signal output
rlabel metal3 s 0 131656 800 131776 6 eFPGA_operand_b_o[17]
port 196 nsew signal output
rlabel metal3 s 239200 148792 240000 148912 6 eFPGA_operand_b_o[18]
port 197 nsew signal output
rlabel metal2 s 152370 239200 152426 240000 6 eFPGA_operand_b_o[19]
port 198 nsew signal output
rlabel metal2 s 25134 239200 25190 240000 6 eFPGA_operand_b_o[1]
port 199 nsew signal output
rlabel metal3 s 239200 158040 240000 158160 6 eFPGA_operand_b_o[20]
port 200 nsew signal output
rlabel metal3 s 239200 169464 240000 169584 6 eFPGA_operand_b_o[21]
port 201 nsew signal output
rlabel metal3 s 0 168104 800 168224 6 eFPGA_operand_b_o[22]
port 202 nsew signal output
rlabel metal2 s 185950 239200 186006 240000 6 eFPGA_operand_b_o[23]
port 203 nsew signal output
rlabel metal3 s 0 191632 800 191752 6 eFPGA_operand_b_o[24]
port 204 nsew signal output
rlabel metal3 s 0 196800 800 196920 6 eFPGA_operand_b_o[25]
port 205 nsew signal output
rlabel metal3 s 0 212440 800 212560 6 eFPGA_operand_b_o[26]
port 206 nsew signal output
rlabel metal2 s 200394 239200 200450 240000 6 eFPGA_operand_b_o[27]
port 207 nsew signal output
rlabel metal3 s 239200 220328 240000 220448 6 eFPGA_operand_b_o[28]
port 208 nsew signal output
rlabel metal2 s 222842 0 222898 800 6 eFPGA_operand_b_o[29]
port 209 nsew signal output
rlabel metal3 s 239200 33328 240000 33448 6 eFPGA_operand_b_o[2]
port 210 nsew signal output
rlabel metal2 s 236550 0 236606 800 6 eFPGA_operand_b_o[30]
port 211 nsew signal output
rlabel metal3 s 239200 238824 240000 238944 6 eFPGA_operand_b_o[31]
port 212 nsew signal output
rlabel metal3 s 239200 44888 240000 45008 6 eFPGA_operand_b_o[3]
port 213 nsew signal output
rlabel metal2 s 44362 239200 44418 240000 6 eFPGA_operand_b_o[4]
port 214 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 eFPGA_operand_b_o[5]
port 215 nsew signal output
rlabel metal3 s 239200 70320 240000 70440 6 eFPGA_operand_b_o[6]
port 216 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 eFPGA_operand_b_o[7]
port 217 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 eFPGA_operand_b_o[8]
port 218 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 eFPGA_operand_b_o[9]
port 219 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 eFPGA_operator_o[0]
port 220 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 eFPGA_operator_o[1]
port 221 nsew signal output
rlabel metal3 s 239200 19456 240000 19576 6 eFPGA_result_a_i[0]
port 222 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 eFPGA_result_a_i[10]
port 223 nsew signal input
rlabel metal2 s 89994 239200 90050 240000 6 eFPGA_result_a_i[11]
port 224 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 eFPGA_result_a_i[12]
port 225 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 eFPGA_result_a_i[13]
port 226 nsew signal input
rlabel metal2 s 116398 239200 116454 240000 6 eFPGA_result_a_i[14]
port 227 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 eFPGA_result_a_i[15]
port 228 nsew signal input
rlabel metal3 s 239200 127984 240000 128104 6 eFPGA_result_a_i[16]
port 229 nsew signal input
rlabel metal3 s 0 134240 800 134360 6 eFPGA_result_a_i[17]
port 230 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 eFPGA_result_a_i[18]
port 231 nsew signal input
rlabel metal3 s 0 149880 800 150000 6 eFPGA_result_a_i[19]
port 232 nsew signal input
rlabel metal3 s 239200 28704 240000 28824 6 eFPGA_result_a_i[1]
port 233 nsew signal input
rlabel metal2 s 181626 0 181682 800 6 eFPGA_result_a_i[20]
port 234 nsew signal input
rlabel metal3 s 239200 171776 240000 171896 6 eFPGA_result_a_i[21]
port 235 nsew signal input
rlabel metal3 s 239200 181024 240000 181144 6 eFPGA_result_a_i[22]
port 236 nsew signal input
rlabel metal2 s 188434 239200 188490 240000 6 eFPGA_result_a_i[23]
port 237 nsew signal input
rlabel metal3 s 239200 190272 240000 190392 6 eFPGA_result_a_i[24]
port 238 nsew signal input
rlabel metal3 s 239200 201832 240000 201952 6 eFPGA_result_a_i[25]
port 239 nsew signal input
rlabel metal3 s 239200 206456 240000 206576 6 eFPGA_result_a_i[26]
port 240 nsew signal input
rlabel metal2 s 211342 0 211398 800 6 eFPGA_result_a_i[27]
port 241 nsew signal input
rlabel metal3 s 0 225496 800 225616 6 eFPGA_result_a_i[28]
port 242 nsew signal input
rlabel metal3 s 239200 227264 240000 227384 6 eFPGA_result_a_i[29]
port 243 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 eFPGA_result_a_i[2]
port 244 nsew signal input
rlabel metal2 s 222014 239200 222070 240000 6 eFPGA_result_a_i[30]
port 245 nsew signal input
rlabel metal2 s 231582 239200 231638 240000 6 eFPGA_result_a_i[31]
port 246 nsew signal input
rlabel metal3 s 239200 47200 240000 47320 6 eFPGA_result_a_i[3]
port 247 nsew signal input
rlabel metal3 s 239200 58760 240000 58880 6 eFPGA_result_a_i[4]
port 248 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 eFPGA_result_a_i[5]
port 249 nsew signal input
rlabel metal2 s 68374 239200 68430 240000 6 eFPGA_result_a_i[6]
port 250 nsew signal input
rlabel metal3 s 239200 84056 240000 84176 6 eFPGA_result_a_i[7]
port 251 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 eFPGA_result_a_i[8]
port 252 nsew signal input
rlabel metal3 s 239200 95616 240000 95736 6 eFPGA_result_a_i[9]
port 253 nsew signal input
rlabel metal2 s 13174 239200 13230 240000 6 eFPGA_result_b_i[0]
port 254 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 eFPGA_result_b_i[10]
port 255 nsew signal input
rlabel metal3 s 239200 111800 240000 111920 6 eFPGA_result_b_i[11]
port 256 nsew signal input
rlabel metal3 s 0 95072 800 95192 6 eFPGA_result_b_i[12]
port 257 nsew signal input
rlabel metal3 s 0 110712 800 110832 6 eFPGA_result_b_i[13]
port 258 nsew signal input
rlabel metal2 s 118790 239200 118846 240000 6 eFPGA_result_b_i[14]
port 259 nsew signal input
rlabel metal2 s 130750 239200 130806 240000 6 eFPGA_result_b_i[15]
port 260 nsew signal input
rlabel metal3 s 239200 130296 240000 130416 6 eFPGA_result_b_i[16]
port 261 nsew signal input
rlabel metal3 s 239200 144168 240000 144288 6 eFPGA_result_b_i[17]
port 262 nsew signal input
rlabel metal2 s 147586 239200 147642 240000 6 eFPGA_result_b_i[18]
port 263 nsew signal input
rlabel metal2 s 154762 239200 154818 240000 6 eFPGA_result_b_i[19]
port 264 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 eFPGA_result_b_i[1]
port 265 nsew signal input
rlabel metal3 s 239200 160352 240000 160472 6 eFPGA_result_b_i[20]
port 266 nsew signal input
rlabel metal3 s 0 160352 800 160472 6 eFPGA_result_b_i[21]
port 267 nsew signal input
rlabel metal3 s 0 170824 800 170944 6 eFPGA_result_b_i[22]
port 268 nsew signal input
rlabel metal3 s 0 178576 800 178696 6 eFPGA_result_b_i[23]
port 269 nsew signal input
rlabel metal3 s 239200 192584 240000 192704 6 eFPGA_result_b_i[24]
port 270 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 eFPGA_result_b_i[25]
port 271 nsew signal input
rlabel metal2 s 198002 239200 198058 240000 6 eFPGA_result_b_i[26]
port 272 nsew signal input
rlabel metal3 s 239200 215704 240000 215824 6 eFPGA_result_b_i[27]
port 273 nsew signal input
rlabel metal3 s 239200 222640 240000 222760 6 eFPGA_result_b_i[28]
port 274 nsew signal input
rlabel metal3 s 239200 229576 240000 229696 6 eFPGA_result_b_i[29]
port 275 nsew signal input
rlabel metal2 s 34794 239200 34850 240000 6 eFPGA_result_b_i[2]
port 276 nsew signal input
rlabel metal2 s 224406 239200 224462 240000 6 eFPGA_result_b_i[30]
port 277 nsew signal input
rlabel metal3 s 0 238552 800 238672 6 eFPGA_result_b_i[31]
port 278 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 eFPGA_result_b_i[3]
port 279 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 eFPGA_result_b_i[4]
port 280 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 eFPGA_result_b_i[5]
port 281 nsew signal input
rlabel metal2 s 70766 239200 70822 240000 6 eFPGA_result_b_i[6]
port 282 nsew signal input
rlabel metal2 s 73158 239200 73214 240000 6 eFPGA_result_b_i[7]
port 283 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 eFPGA_result_b_i[8]
port 284 nsew signal input
rlabel metal3 s 239200 97928 240000 98048 6 eFPGA_result_b_i[9]
port 285 nsew signal input
rlabel metal3 s 239200 21768 240000 21888 6 eFPGA_result_c_i[0]
port 286 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 eFPGA_result_c_i[10]
port 287 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 eFPGA_result_c_i[11]
port 288 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 eFPGA_result_c_i[12]
port 289 nsew signal input
rlabel metal2 s 104346 239200 104402 240000 6 eFPGA_result_c_i[13]
port 290 nsew signal input
rlabel metal3 s 0 116016 800 116136 6 eFPGA_result_c_i[14]
port 291 nsew signal input
rlabel metal3 s 0 121184 800 121304 6 eFPGA_result_c_i[15]
port 292 nsew signal input
rlabel metal3 s 0 126352 800 126472 6 eFPGA_result_c_i[16]
port 293 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 eFPGA_result_c_i[17]
port 294 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 eFPGA_result_c_i[18]
port 295 nsew signal input
rlabel metal2 s 174818 0 174874 800 6 eFPGA_result_c_i[19]
port 296 nsew signal input
rlabel metal3 s 239200 31016 240000 31136 6 eFPGA_result_c_i[1]
port 297 nsew signal input
rlabel metal2 s 162030 239200 162086 240000 6 eFPGA_result_c_i[20]
port 298 nsew signal input
rlabel metal3 s 239200 174088 240000 174208 6 eFPGA_result_c_i[21]
port 299 nsew signal input
rlabel metal2 s 176382 239200 176438 240000 6 eFPGA_result_c_i[22]
port 300 nsew signal input
rlabel metal2 s 186226 0 186282 800 6 eFPGA_result_c_i[23]
port 301 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 eFPGA_result_c_i[24]
port 302 nsew signal input
rlabel metal3 s 0 199520 800 199640 6 eFPGA_result_c_i[25]
port 303 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 eFPGA_result_c_i[26]
port 304 nsew signal input
rlabel metal2 s 202786 239200 202842 240000 6 eFPGA_result_c_i[27]
port 305 nsew signal input
rlabel metal2 s 215942 0 215998 800 6 eFPGA_result_c_i[28]
port 306 nsew signal input
rlabel metal2 s 225142 0 225198 800 6 eFPGA_result_c_i[29]
port 307 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 eFPGA_result_c_i[2]
port 308 nsew signal input
rlabel metal3 s 239200 231888 240000 232008 6 eFPGA_result_c_i[30]
port 309 nsew signal input
rlabel metal2 s 233974 239200 234030 240000 6 eFPGA_result_c_i[31]
port 310 nsew signal input
rlabel metal2 s 41970 239200 42026 240000 6 eFPGA_result_c_i[3]
port 311 nsew signal input
rlabel metal3 s 239200 61072 240000 61192 6 eFPGA_result_c_i[4]
port 312 nsew signal input
rlabel metal3 s 0 50736 800 50856 6 eFPGA_result_c_i[5]
port 313 nsew signal input
rlabel metal3 s 239200 72632 240000 72752 6 eFPGA_result_c_i[6]
port 314 nsew signal input
rlabel metal2 s 75550 239200 75606 240000 6 eFPGA_result_c_i[7]
port 315 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 eFPGA_result_c_i[8]
port 316 nsew signal input
rlabel metal3 s 239200 100240 240000 100360 6 eFPGA_result_c_i[9]
port 317 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 eFPGA_write_strobe_o
port 318 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 ext_perf_counters_i
port 319 nsew signal input
rlabel metal3 s 239200 7896 240000 8016 6 fetch_enable_i
port 320 nsew signal input
rlabel metal3 s 239200 24080 240000 24200 6 instr_addr_o[0]
port 321 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 instr_addr_o[10]
port 322 nsew signal output
rlabel metal3 s 0 82016 800 82136 6 instr_addr_o[11]
port 323 nsew signal output
rlabel metal2 s 94778 239200 94834 240000 6 instr_addr_o[12]
port 324 nsew signal output
rlabel metal2 s 106738 239200 106794 240000 6 instr_addr_o[13]
port 325 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 instr_addr_o[14]
port 326 nsew signal output
rlabel metal2 s 133142 239200 133198 240000 6 instr_addr_o[15]
port 327 nsew signal output
rlabel metal3 s 0 129072 800 129192 6 instr_addr_o[16]
port 328 nsew signal output
rlabel metal3 s 239200 146480 240000 146600 6 instr_addr_o[17]
port 329 nsew signal output
rlabel metal2 s 149978 239200 150034 240000 6 instr_addr_o[18]
port 330 nsew signal output
rlabel metal3 s 0 152464 800 152584 6 instr_addr_o[19]
port 331 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 instr_addr_o[1]
port 332 nsew signal output
rlabel metal3 s 0 157768 800 157888 6 instr_addr_o[20]
port 333 nsew signal output
rlabel metal3 s 239200 176400 240000 176520 6 instr_addr_o[21]
port 334 nsew signal output
rlabel metal2 s 178774 239200 178830 240000 6 instr_addr_o[22]
port 335 nsew signal output
rlabel metal3 s 0 181160 800 181280 6 instr_addr_o[23]
port 336 nsew signal output
rlabel metal3 s 239200 194896 240000 195016 6 instr_addr_o[24]
port 337 nsew signal output
rlabel metal2 s 195610 239200 195666 240000 6 instr_addr_o[25]
port 338 nsew signal output
rlabel metal2 s 204534 0 204590 800 6 instr_addr_o[26]
port 339 nsew signal output
rlabel metal2 s 213642 0 213698 800 6 instr_addr_o[27]
port 340 nsew signal output
rlabel metal2 s 209962 239200 210018 240000 6 instr_addr_o[28]
port 341 nsew signal output
rlabel metal2 s 217230 239200 217286 240000 6 instr_addr_o[29]
port 342 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 instr_addr_o[2]
port 343 nsew signal output
rlabel metal3 s 0 233384 800 233504 6 instr_addr_o[30]
port 344 nsew signal output
rlabel metal2 s 236366 239200 236422 240000 6 instr_addr_o[31]
port 345 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 instr_addr_o[3]
port 346 nsew signal output
rlabel metal2 s 46754 239200 46810 240000 6 instr_addr_o[4]
port 347 nsew signal output
rlabel metal2 s 58806 239200 58862 240000 6 instr_addr_o[5]
port 348 nsew signal output
rlabel metal3 s 239200 74944 240000 75064 6 instr_addr_o[6]
port 349 nsew signal output
rlabel metal2 s 77942 239200 77998 240000 6 instr_addr_o[7]
port 350 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 instr_addr_o[8]
port 351 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 instr_addr_o[9]
port 352 nsew signal output
rlabel metal3 s 239200 10208 240000 10328 6 instr_gnt_i
port 353 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 instr_rdata_i[0]
port 354 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 instr_rdata_i[10]
port 355 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 instr_rdata_i[11]
port 356 nsew signal input
rlabel metal2 s 97170 239200 97226 240000 6 instr_rdata_i[12]
port 357 nsew signal input
rlabel metal3 s 0 113296 800 113416 6 instr_rdata_i[13]
port 358 nsew signal input
rlabel metal2 s 121182 239200 121238 240000 6 instr_rdata_i[14]
port 359 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 instr_rdata_i[15]
port 360 nsew signal input
rlabel metal3 s 239200 132608 240000 132728 6 instr_rdata_i[16]
port 361 nsew signal input
rlabel metal3 s 0 136824 800 136944 6 instr_rdata_i[17]
port 362 nsew signal input
rlabel metal3 s 239200 151104 240000 151224 6 instr_rdata_i[18]
port 363 nsew signal input
rlabel metal3 s 239200 155728 240000 155848 6 instr_rdata_i[19]
port 364 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 instr_rdata_i[1]
port 365 nsew signal input
rlabel metal2 s 183926 0 183982 800 6 instr_rdata_i[20]
port 366 nsew signal input
rlabel metal2 s 169206 239200 169262 240000 6 instr_rdata_i[21]
port 367 nsew signal input
rlabel metal3 s 239200 183336 240000 183456 6 instr_rdata_i[22]
port 368 nsew signal input
rlabel metal3 s 0 183744 800 183864 6 instr_rdata_i[23]
port 369 nsew signal input
rlabel metal3 s 0 194216 800 194336 6 instr_rdata_i[24]
port 370 nsew signal input
rlabel metal3 s 239200 204144 240000 204264 6 instr_rdata_i[25]
port 371 nsew signal input
rlabel metal2 s 206834 0 206890 800 6 instr_rdata_i[26]
port 372 nsew signal input
rlabel metal2 s 205178 239200 205234 240000 6 instr_rdata_i[27]
port 373 nsew signal input
rlabel metal3 s 239200 224952 240000 225072 6 instr_rdata_i[28]
port 374 nsew signal input
rlabel metal2 s 227350 0 227406 800 6 instr_rdata_i[29]
port 375 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 instr_rdata_i[2]
port 376 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 instr_rdata_i[30]
port 377 nsew signal input
rlabel metal2 s 238758 239200 238814 240000 6 instr_rdata_i[31]
port 378 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 instr_rdata_i[3]
port 379 nsew signal input
rlabel metal3 s 239200 63384 240000 63504 6 instr_rdata_i[4]
port 380 nsew signal input
rlabel metal2 s 61198 239200 61254 240000 6 instr_rdata_i[5]
port 381 nsew signal input
rlabel metal3 s 239200 77256 240000 77376 6 instr_rdata_i[6]
port 382 nsew signal input
rlabel metal3 s 239200 86368 240000 86488 6 instr_rdata_i[7]
port 383 nsew signal input
rlabel metal3 s 239200 90992 240000 91112 6 instr_rdata_i[8]
port 384 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 instr_rdata_i[9]
port 385 nsew signal input
rlabel metal3 s 239200 12520 240000 12640 6 instr_req_o
port 386 nsew signal output
rlabel metal2 s 3606 239200 3662 240000 6 instr_rvalid_i
port 387 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 irq_ack_o
port 388 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 irq_i
port 389 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 irq_id_i[0]
port 390 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 irq_id_i[1]
port 391 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 irq_id_i[2]
port 392 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 irq_id_i[3]
port 393 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 irq_id_i[4]
port 394 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 irq_id_o[0]
port 395 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 irq_id_o[1]
port 396 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 irq_id_o[2]
port 397 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 irq_id_o[3]
port 398 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 irq_id_o[4]
port 399 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 rst_ni
port 400 nsew signal input
rlabel metal2 s 5998 239200 6054 240000 6 test_en_i
port 401 nsew signal input
rlabel metal4 s 4208 2128 4528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 14208 2128 14528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 24208 2128 24528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 34208 2128 34528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 44208 2128 44528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 54208 2128 54528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 64208 2128 64528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 74208 2128 74528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 84208 2128 84528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 94208 2128 94528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 104208 2128 104528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 114208 2128 114528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 124208 2128 124528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 134208 2128 134528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 144208 2128 144528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 154208 2128 154528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 164208 2128 164528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 174208 2128 174528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 184208 2128 184528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 194208 2128 194528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 204208 2128 204528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 214208 2128 214528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 224208 2128 224528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 234208 2128 234528 237776 6 vccd1
port 402 nsew power input
rlabel metal4 s 9208 2128 9528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 19208 2128 19528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 29208 2128 29528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 39208 2128 39528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 49208 2128 49528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 59208 2128 59528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 69208 2128 69528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 79208 2128 79528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 89208 2128 89528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 99208 2128 99528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 109208 2128 109528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 119208 2128 119528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 129208 2128 129528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 139208 2128 139528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 149208 2128 149528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 159208 2128 159528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 169208 2128 169528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 179208 2128 179528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 189208 2128 189528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 199208 2128 199528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 209208 2128 209528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 219208 2128 219528 237776 6 vssd1
port 403 nsew ground input
rlabel metal4 s 229208 2128 229528 237776 6 vssd1
port 403 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 240000 240000
string LEFview TRUE
string GDS_FILE /project/openlane/flexbex_ibex_core/runs/flexbex_ibex_core/results/magic/flexbex_ibex_core.gds
string GDS_END 100766730
string GDS_START 571538
<< end >>

