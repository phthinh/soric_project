VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO soric_soc
  CLASS BLOCK ;
  FOREIGN soric_soc ;
  ORIGIN 0.000 0.000 ;
  SIZE 1700.000 BY 300.000 ;
  PIN error_uart_to_mem
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 269.320 1700.000 269.920 ;
    END
  END error_uart_to_mem
  PIN master_data_addr_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 296.000 1.290 300.000 ;
    END
  END master_data_addr_to_inter_i[0]
  PIN master_data_addr_to_inter_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 296.000 160.450 300.000 ;
    END
  END master_data_addr_to_inter_i[10]
  PIN master_data_addr_to_inter_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 296.000 171.490 300.000 ;
    END
  END master_data_addr_to_inter_i[11]
  PIN master_data_addr_to_inter_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 296.000 182.530 300.000 ;
    END
  END master_data_addr_to_inter_i[12]
  PIN master_data_addr_to_inter_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 296.000 193.570 300.000 ;
    END
  END master_data_addr_to_inter_i[13]
  PIN master_data_addr_to_inter_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 296.000 204.610 300.000 ;
    END
  END master_data_addr_to_inter_i[14]
  PIN master_data_addr_to_inter_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 296.000 215.650 300.000 ;
    END
  END master_data_addr_to_inter_i[15]
  PIN master_data_addr_to_inter_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 296.000 226.690 300.000 ;
    END
  END master_data_addr_to_inter_i[16]
  PIN master_data_addr_to_inter_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 296.000 237.730 300.000 ;
    END
  END master_data_addr_to_inter_i[17]
  PIN master_data_addr_to_inter_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 296.000 249.230 300.000 ;
    END
  END master_data_addr_to_inter_i[18]
  PIN master_data_addr_to_inter_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 296.000 260.270 300.000 ;
    END
  END master_data_addr_to_inter_i[19]
  PIN master_data_addr_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 296.000 29.810 300.000 ;
    END
  END master_data_addr_to_inter_i[1]
  PIN master_data_addr_to_inter_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 296.000 271.310 300.000 ;
    END
  END master_data_addr_to_inter_i[20]
  PIN master_data_addr_to_inter_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 296.000 282.350 300.000 ;
    END
  END master_data_addr_to_inter_i[21]
  PIN master_data_addr_to_inter_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 296.000 293.390 300.000 ;
    END
  END master_data_addr_to_inter_i[22]
  PIN master_data_addr_to_inter_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 296.000 304.430 300.000 ;
    END
  END master_data_addr_to_inter_i[23]
  PIN master_data_addr_to_inter_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 296.000 315.470 300.000 ;
    END
  END master_data_addr_to_inter_i[24]
  PIN master_data_addr_to_inter_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 296.000 326.510 300.000 ;
    END
  END master_data_addr_to_inter_i[25]
  PIN master_data_addr_to_inter_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 296.000 337.550 300.000 ;
    END
  END master_data_addr_to_inter_i[26]
  PIN master_data_addr_to_inter_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 296.000 346.290 300.000 ;
    END
  END master_data_addr_to_inter_i[27]
  PIN master_data_addr_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 296.000 58.790 300.000 ;
    END
  END master_data_addr_to_inter_i[2]
  PIN master_data_addr_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 296.000 72.130 300.000 ;
    END
  END master_data_addr_to_inter_i[3]
  PIN master_data_addr_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 296.000 85.010 300.000 ;
    END
  END master_data_addr_to_inter_i[4]
  PIN master_data_addr_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 296.000 98.350 300.000 ;
    END
  END master_data_addr_to_inter_i[5]
  PIN master_data_addr_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 296.000 111.690 300.000 ;
    END
  END master_data_addr_to_inter_i[6]
  PIN master_data_addr_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 296.000 125.030 300.000 ;
    END
  END master_data_addr_to_inter_i[7]
  PIN master_data_addr_to_inter_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 296.000 138.370 300.000 ;
    END
  END master_data_addr_to_inter_i[8]
  PIN master_data_addr_to_inter_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 296.000 149.410 300.000 ;
    END
  END master_data_addr_to_inter_i[9]
  PIN master_data_addr_to_inter_ro_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 296.000 3.130 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[0]
  PIN master_data_addr_to_inter_ro_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 296.000 162.750 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[10]
  PIN master_data_addr_to_inter_ro_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 296.000 173.790 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[11]
  PIN master_data_addr_to_inter_ro_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 296.000 184.830 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[12]
  PIN master_data_addr_to_inter_ro_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 296.000 195.870 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[13]
  PIN master_data_addr_to_inter_ro_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 296.000 206.910 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[14]
  PIN master_data_addr_to_inter_ro_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 296.000 217.950 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[15]
  PIN master_data_addr_to_inter_ro_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 296.000 228.990 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[16]
  PIN master_data_addr_to_inter_ro_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 296.000 240.030 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[17]
  PIN master_data_addr_to_inter_ro_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 296.000 251.070 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[18]
  PIN master_data_addr_to_inter_ro_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 296.000 262.110 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[19]
  PIN master_data_addr_to_inter_ro_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 296.000 32.110 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[1]
  PIN master_data_addr_to_inter_ro_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 296.000 273.150 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[20]
  PIN master_data_addr_to_inter_ro_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 296.000 284.650 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[21]
  PIN master_data_addr_to_inter_ro_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 296.000 295.690 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[22]
  PIN master_data_addr_to_inter_ro_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 296.000 306.730 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[23]
  PIN master_data_addr_to_inter_ro_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 296.000 317.770 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[24]
  PIN master_data_addr_to_inter_ro_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 296.000 328.810 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[25]
  PIN master_data_addr_to_inter_ro_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 296.000 60.630 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[2]
  PIN master_data_addr_to_inter_ro_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 296.000 73.970 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[3]
  PIN master_data_addr_to_inter_ro_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 296.000 87.310 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[4]
  PIN master_data_addr_to_inter_ro_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 296.000 100.650 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[5]
  PIN master_data_addr_to_inter_ro_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 296.000 113.990 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[6]
  PIN master_data_addr_to_inter_ro_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 296.000 127.330 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[7]
  PIN master_data_addr_to_inter_ro_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 296.000 140.670 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[8]
  PIN master_data_addr_to_inter_ro_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 296.000 151.710 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[9]
  PIN master_data_be_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 296.000 5.430 300.000 ;
    END
  END master_data_be_to_inter_i[0]
  PIN master_data_be_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 296.000 34.410 300.000 ;
    END
  END master_data_be_to_inter_i[1]
  PIN master_data_be_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 296.000 62.930 300.000 ;
    END
  END master_data_be_to_inter_i[2]
  PIN master_data_be_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 296.000 76.270 300.000 ;
    END
  END master_data_be_to_inter_i[3]
  PIN master_data_be_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 296.000 89.610 300.000 ;
    END
  END master_data_be_to_inter_i[4]
  PIN master_data_be_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 296.000 102.950 300.000 ;
    END
  END master_data_be_to_inter_i[5]
  PIN master_data_be_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 296.000 116.290 300.000 ;
    END
  END master_data_be_to_inter_i[6]
  PIN master_data_be_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 296.000 129.630 300.000 ;
    END
  END master_data_be_to_inter_i[7]
  PIN master_data_gnt_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 296.000 7.730 300.000 ;
    END
  END master_data_gnt_to_inter_o[0]
  PIN master_data_gnt_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 296.000 36.710 300.000 ;
    END
  END master_data_gnt_to_inter_o[1]
  PIN master_data_gnt_to_inter_ro_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 296.000 10.030 300.000 ;
    END
  END master_data_gnt_to_inter_ro_o[0]
  PIN master_data_gnt_to_inter_ro_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 296.000 38.550 300.000 ;
    END
  END master_data_gnt_to_inter_ro_o[1]
  PIN master_data_rdata_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 296.000 12.330 300.000 ;
    END
  END master_data_rdata_to_inter_o[0]
  PIN master_data_rdata_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 296.000 165.050 300.000 ;
    END
  END master_data_rdata_to_inter_o[10]
  PIN master_data_rdata_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 296.000 176.090 300.000 ;
    END
  END master_data_rdata_to_inter_o[11]
  PIN master_data_rdata_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 296.000 187.130 300.000 ;
    END
  END master_data_rdata_to_inter_o[12]
  PIN master_data_rdata_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 296.000 198.170 300.000 ;
    END
  END master_data_rdata_to_inter_o[13]
  PIN master_data_rdata_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 296.000 209.210 300.000 ;
    END
  END master_data_rdata_to_inter_o[14]
  PIN master_data_rdata_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 296.000 220.250 300.000 ;
    END
  END master_data_rdata_to_inter_o[15]
  PIN master_data_rdata_to_inter_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 296.000 231.290 300.000 ;
    END
  END master_data_rdata_to_inter_o[16]
  PIN master_data_rdata_to_inter_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 296.000 242.330 300.000 ;
    END
  END master_data_rdata_to_inter_o[17]
  PIN master_data_rdata_to_inter_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 296.000 253.370 300.000 ;
    END
  END master_data_rdata_to_inter_o[18]
  PIN master_data_rdata_to_inter_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 296.000 264.410 300.000 ;
    END
  END master_data_rdata_to_inter_o[19]
  PIN master_data_rdata_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 296.000 40.850 300.000 ;
    END
  END master_data_rdata_to_inter_o[1]
  PIN master_data_rdata_to_inter_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 296.000 275.450 300.000 ;
    END
  END master_data_rdata_to_inter_o[20]
  PIN master_data_rdata_to_inter_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 296.000 286.490 300.000 ;
    END
  END master_data_rdata_to_inter_o[21]
  PIN master_data_rdata_to_inter_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 296.000 297.530 300.000 ;
    END
  END master_data_rdata_to_inter_o[22]
  PIN master_data_rdata_to_inter_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 296.000 308.570 300.000 ;
    END
  END master_data_rdata_to_inter_o[23]
  PIN master_data_rdata_to_inter_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 296.000 320.070 300.000 ;
    END
  END master_data_rdata_to_inter_o[24]
  PIN master_data_rdata_to_inter_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 296.000 331.110 300.000 ;
    END
  END master_data_rdata_to_inter_o[25]
  PIN master_data_rdata_to_inter_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 296.000 339.850 300.000 ;
    END
  END master_data_rdata_to_inter_o[26]
  PIN master_data_rdata_to_inter_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 296.000 348.590 300.000 ;
    END
  END master_data_rdata_to_inter_o[27]
  PIN master_data_rdata_to_inter_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 296.000 355.490 300.000 ;
    END
  END master_data_rdata_to_inter_o[28]
  PIN master_data_rdata_to_inter_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 296.000 361.930 300.000 ;
    END
  END master_data_rdata_to_inter_o[29]
  PIN master_data_rdata_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 296.000 65.230 300.000 ;
    END
  END master_data_rdata_to_inter_o[2]
  PIN master_data_rdata_to_inter_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 296.000 368.370 300.000 ;
    END
  END master_data_rdata_to_inter_o[30]
  PIN master_data_rdata_to_inter_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 296.000 375.270 300.000 ;
    END
  END master_data_rdata_to_inter_o[31]
  PIN master_data_rdata_to_inter_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 296.000 381.710 300.000 ;
    END
  END master_data_rdata_to_inter_o[32]
  PIN master_data_rdata_to_inter_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 296.000 388.610 300.000 ;
    END
  END master_data_rdata_to_inter_o[33]
  PIN master_data_rdata_to_inter_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 296.000 395.050 300.000 ;
    END
  END master_data_rdata_to_inter_o[34]
  PIN master_data_rdata_to_inter_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 296.000 401.950 300.000 ;
    END
  END master_data_rdata_to_inter_o[35]
  PIN master_data_rdata_to_inter_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 296.000 408.390 300.000 ;
    END
  END master_data_rdata_to_inter_o[36]
  PIN master_data_rdata_to_inter_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 296.000 414.830 300.000 ;
    END
  END master_data_rdata_to_inter_o[37]
  PIN master_data_rdata_to_inter_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 296.000 421.730 300.000 ;
    END
  END master_data_rdata_to_inter_o[38]
  PIN master_data_rdata_to_inter_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 296.000 428.170 300.000 ;
    END
  END master_data_rdata_to_inter_o[39]
  PIN master_data_rdata_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 296.000 78.570 300.000 ;
    END
  END master_data_rdata_to_inter_o[3]
  PIN master_data_rdata_to_inter_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 296.000 435.070 300.000 ;
    END
  END master_data_rdata_to_inter_o[40]
  PIN master_data_rdata_to_inter_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 296.000 441.510 300.000 ;
    END
  END master_data_rdata_to_inter_o[41]
  PIN master_data_rdata_to_inter_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 296.000 448.410 300.000 ;
    END
  END master_data_rdata_to_inter_o[42]
  PIN master_data_rdata_to_inter_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 296.000 454.850 300.000 ;
    END
  END master_data_rdata_to_inter_o[43]
  PIN master_data_rdata_to_inter_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 296.000 461.750 300.000 ;
    END
  END master_data_rdata_to_inter_o[44]
  PIN master_data_rdata_to_inter_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 296.000 468.190 300.000 ;
    END
  END master_data_rdata_to_inter_o[45]
  PIN master_data_rdata_to_inter_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 296.000 474.630 300.000 ;
    END
  END master_data_rdata_to_inter_o[46]
  PIN master_data_rdata_to_inter_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 296.000 481.530 300.000 ;
    END
  END master_data_rdata_to_inter_o[47]
  PIN master_data_rdata_to_inter_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 296.000 487.970 300.000 ;
    END
  END master_data_rdata_to_inter_o[48]
  PIN master_data_rdata_to_inter_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 296.000 494.870 300.000 ;
    END
  END master_data_rdata_to_inter_o[49]
  PIN master_data_rdata_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 296.000 91.910 300.000 ;
    END
  END master_data_rdata_to_inter_o[4]
  PIN master_data_rdata_to_inter_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 296.000 501.310 300.000 ;
    END
  END master_data_rdata_to_inter_o[50]
  PIN master_data_rdata_to_inter_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 296.000 508.210 300.000 ;
    END
  END master_data_rdata_to_inter_o[51]
  PIN master_data_rdata_to_inter_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 296.000 514.650 300.000 ;
    END
  END master_data_rdata_to_inter_o[52]
  PIN master_data_rdata_to_inter_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 296.000 521.090 300.000 ;
    END
  END master_data_rdata_to_inter_o[53]
  PIN master_data_rdata_to_inter_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 296.000 527.990 300.000 ;
    END
  END master_data_rdata_to_inter_o[54]
  PIN master_data_rdata_to_inter_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 296.000 534.430 300.000 ;
    END
  END master_data_rdata_to_inter_o[55]
  PIN master_data_rdata_to_inter_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 296.000 541.330 300.000 ;
    END
  END master_data_rdata_to_inter_o[56]
  PIN master_data_rdata_to_inter_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 296.000 547.770 300.000 ;
    END
  END master_data_rdata_to_inter_o[57]
  PIN master_data_rdata_to_inter_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 296.000 554.670 300.000 ;
    END
  END master_data_rdata_to_inter_o[58]
  PIN master_data_rdata_to_inter_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 296.000 561.110 300.000 ;
    END
  END master_data_rdata_to_inter_o[59]
  PIN master_data_rdata_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 296.000 105.250 300.000 ;
    END
  END master_data_rdata_to_inter_o[5]
  PIN master_data_rdata_to_inter_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 296.000 568.010 300.000 ;
    END
  END master_data_rdata_to_inter_o[60]
  PIN master_data_rdata_to_inter_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 296.000 574.450 300.000 ;
    END
  END master_data_rdata_to_inter_o[61]
  PIN master_data_rdata_to_inter_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 296.000 580.890 300.000 ;
    END
  END master_data_rdata_to_inter_o[62]
  PIN master_data_rdata_to_inter_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 296.000 587.790 300.000 ;
    END
  END master_data_rdata_to_inter_o[63]
  PIN master_data_rdata_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 296.000 118.590 300.000 ;
    END
  END master_data_rdata_to_inter_o[6]
  PIN master_data_rdata_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 296.000 131.470 300.000 ;
    END
  END master_data_rdata_to_inter_o[7]
  PIN master_data_rdata_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 296.000 142.970 300.000 ;
    END
  END master_data_rdata_to_inter_o[8]
  PIN master_data_rdata_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 296.000 154.010 300.000 ;
    END
  END master_data_rdata_to_inter_o[9]
  PIN master_data_rdata_to_inter_ro_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 296.000 14.170 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[0]
  PIN master_data_rdata_to_inter_ro_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 296.000 166.890 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[10]
  PIN master_data_rdata_to_inter_ro_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 296.000 178.390 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[11]
  PIN master_data_rdata_to_inter_ro_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 296.000 189.430 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[12]
  PIN master_data_rdata_to_inter_ro_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 296.000 200.470 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[13]
  PIN master_data_rdata_to_inter_ro_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 296.000 211.510 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[14]
  PIN master_data_rdata_to_inter_ro_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 296.000 222.550 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[15]
  PIN master_data_rdata_to_inter_ro_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 296.000 233.590 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[16]
  PIN master_data_rdata_to_inter_ro_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 296.000 244.630 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[17]
  PIN master_data_rdata_to_inter_ro_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 296.000 255.670 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[18]
  PIN master_data_rdata_to_inter_ro_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 296.000 266.710 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[19]
  PIN master_data_rdata_to_inter_ro_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 296.000 43.150 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[1]
  PIN master_data_rdata_to_inter_ro_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 296.000 277.750 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[20]
  PIN master_data_rdata_to_inter_ro_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 296.000 288.790 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[21]
  PIN master_data_rdata_to_inter_ro_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 296.000 299.830 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[22]
  PIN master_data_rdata_to_inter_ro_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 296.000 310.870 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[23]
  PIN master_data_rdata_to_inter_ro_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 296.000 321.910 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[24]
  PIN master_data_rdata_to_inter_ro_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 296.000 332.950 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[25]
  PIN master_data_rdata_to_inter_ro_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 296.000 342.150 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[26]
  PIN master_data_rdata_to_inter_ro_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 296.000 350.890 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[27]
  PIN master_data_rdata_to_inter_ro_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 296.000 357.330 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[28]
  PIN master_data_rdata_to_inter_ro_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 296.000 364.230 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[29]
  PIN master_data_rdata_to_inter_ro_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 296.000 67.530 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[2]
  PIN master_data_rdata_to_inter_ro_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 296.000 370.670 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[30]
  PIN master_data_rdata_to_inter_ro_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 296.000 377.570 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[31]
  PIN master_data_rdata_to_inter_ro_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 296.000 384.010 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[32]
  PIN master_data_rdata_to_inter_ro_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 296.000 390.910 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[33]
  PIN master_data_rdata_to_inter_ro_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 296.000 397.350 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[34]
  PIN master_data_rdata_to_inter_ro_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 296.000 403.790 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[35]
  PIN master_data_rdata_to_inter_ro_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 296.000 410.690 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[36]
  PIN master_data_rdata_to_inter_ro_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 296.000 417.130 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[37]
  PIN master_data_rdata_to_inter_ro_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 296.000 424.030 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[38]
  PIN master_data_rdata_to_inter_ro_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 296.000 430.470 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[39]
  PIN master_data_rdata_to_inter_ro_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 296.000 80.870 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[3]
  PIN master_data_rdata_to_inter_ro_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 296.000 437.370 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[40]
  PIN master_data_rdata_to_inter_ro_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 296.000 443.810 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[41]
  PIN master_data_rdata_to_inter_ro_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 296.000 450.250 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[42]
  PIN master_data_rdata_to_inter_ro_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 296.000 457.150 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[43]
  PIN master_data_rdata_to_inter_ro_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 296.000 463.590 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[44]
  PIN master_data_rdata_to_inter_ro_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 296.000 470.490 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[45]
  PIN master_data_rdata_to_inter_ro_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 296.000 476.930 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[46]
  PIN master_data_rdata_to_inter_ro_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 296.000 483.830 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[47]
  PIN master_data_rdata_to_inter_ro_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 296.000 490.270 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[48]
  PIN master_data_rdata_to_inter_ro_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 296.000 497.170 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[49]
  PIN master_data_rdata_to_inter_ro_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 296.000 94.210 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[4]
  PIN master_data_rdata_to_inter_ro_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 296.000 503.610 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[50]
  PIN master_data_rdata_to_inter_ro_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 296.000 510.050 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[51]
  PIN master_data_rdata_to_inter_ro_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 296.000 516.950 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[52]
  PIN master_data_rdata_to_inter_ro_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 296.000 523.390 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[53]
  PIN master_data_rdata_to_inter_ro_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 296.000 530.290 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[54]
  PIN master_data_rdata_to_inter_ro_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 296.000 536.730 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[55]
  PIN master_data_rdata_to_inter_ro_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 296.000 543.630 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[56]
  PIN master_data_rdata_to_inter_ro_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 296.000 550.070 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[57]
  PIN master_data_rdata_to_inter_ro_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 296.000 556.510 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[58]
  PIN master_data_rdata_to_inter_ro_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 296.000 563.410 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[59]
  PIN master_data_rdata_to_inter_ro_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 296.000 107.550 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[5]
  PIN master_data_rdata_to_inter_ro_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 296.000 569.850 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[60]
  PIN master_data_rdata_to_inter_ro_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 296.000 576.750 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[61]
  PIN master_data_rdata_to_inter_ro_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 296.000 583.190 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[62]
  PIN master_data_rdata_to_inter_ro_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 296.000 590.090 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[63]
  PIN master_data_rdata_to_inter_ro_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 296.000 120.430 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[6]
  PIN master_data_rdata_to_inter_ro_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 296.000 133.770 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[7]
  PIN master_data_rdata_to_inter_ro_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 296.000 144.810 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[8]
  PIN master_data_rdata_to_inter_ro_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 296.000 155.850 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[9]
  PIN master_data_req_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 296.000 16.470 300.000 ;
    END
  END master_data_req_to_inter_i[0]
  PIN master_data_req_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 296.000 45.450 300.000 ;
    END
  END master_data_req_to_inter_i[1]
  PIN master_data_req_to_inter_ro_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 296.000 18.770 300.000 ;
    END
  END master_data_req_to_inter_ro_i[0]
  PIN master_data_req_to_inter_ro_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 296.000 47.750 300.000 ;
    END
  END master_data_req_to_inter_ro_i[1]
  PIN master_data_rvalid_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 296.000 21.070 300.000 ;
    END
  END master_data_rvalid_to_inter_o[0]
  PIN master_data_rvalid_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 296.000 49.590 300.000 ;
    END
  END master_data_rvalid_to_inter_o[1]
  PIN master_data_rvalid_to_inter_ro_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 296.000 23.370 300.000 ;
    END
  END master_data_rvalid_to_inter_ro_o[0]
  PIN master_data_rvalid_to_inter_ro_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 296.000 51.890 300.000 ;
    END
  END master_data_rvalid_to_inter_ro_o[1]
  PIN master_data_wdata_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 296.000 25.210 300.000 ;
    END
  END master_data_wdata_to_inter_i[0]
  PIN master_data_wdata_to_inter_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 296.000 169.190 300.000 ;
    END
  END master_data_wdata_to_inter_i[10]
  PIN master_data_wdata_to_inter_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 296.000 180.230 300.000 ;
    END
  END master_data_wdata_to_inter_i[11]
  PIN master_data_wdata_to_inter_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 296.000 191.270 300.000 ;
    END
  END master_data_wdata_to_inter_i[12]
  PIN master_data_wdata_to_inter_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 296.000 202.310 300.000 ;
    END
  END master_data_wdata_to_inter_i[13]
  PIN master_data_wdata_to_inter_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 296.000 213.810 300.000 ;
    END
  END master_data_wdata_to_inter_i[14]
  PIN master_data_wdata_to_inter_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 296.000 224.850 300.000 ;
    END
  END master_data_wdata_to_inter_i[15]
  PIN master_data_wdata_to_inter_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 296.000 235.890 300.000 ;
    END
  END master_data_wdata_to_inter_i[16]
  PIN master_data_wdata_to_inter_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 296.000 246.930 300.000 ;
    END
  END master_data_wdata_to_inter_i[17]
  PIN master_data_wdata_to_inter_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 296.000 257.970 300.000 ;
    END
  END master_data_wdata_to_inter_i[18]
  PIN master_data_wdata_to_inter_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 296.000 269.010 300.000 ;
    END
  END master_data_wdata_to_inter_i[19]
  PIN master_data_wdata_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 296.000 54.190 300.000 ;
    END
  END master_data_wdata_to_inter_i[1]
  PIN master_data_wdata_to_inter_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 296.000 280.050 300.000 ;
    END
  END master_data_wdata_to_inter_i[20]
  PIN master_data_wdata_to_inter_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 296.000 291.090 300.000 ;
    END
  END master_data_wdata_to_inter_i[21]
  PIN master_data_wdata_to_inter_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 296.000 302.130 300.000 ;
    END
  END master_data_wdata_to_inter_i[22]
  PIN master_data_wdata_to_inter_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 296.000 313.170 300.000 ;
    END
  END master_data_wdata_to_inter_i[23]
  PIN master_data_wdata_to_inter_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 296.000 324.210 300.000 ;
    END
  END master_data_wdata_to_inter_i[24]
  PIN master_data_wdata_to_inter_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 296.000 335.250 300.000 ;
    END
  END master_data_wdata_to_inter_i[25]
  PIN master_data_wdata_to_inter_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 296.000 343.990 300.000 ;
    END
  END master_data_wdata_to_inter_i[26]
  PIN master_data_wdata_to_inter_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 296.000 353.190 300.000 ;
    END
  END master_data_wdata_to_inter_i[27]
  PIN master_data_wdata_to_inter_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 296.000 359.630 300.000 ;
    END
  END master_data_wdata_to_inter_i[28]
  PIN master_data_wdata_to_inter_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 296.000 366.530 300.000 ;
    END
  END master_data_wdata_to_inter_i[29]
  PIN master_data_wdata_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 296.000 69.830 300.000 ;
    END
  END master_data_wdata_to_inter_i[2]
  PIN master_data_wdata_to_inter_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 296.000 372.970 300.000 ;
    END
  END master_data_wdata_to_inter_i[30]
  PIN master_data_wdata_to_inter_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 296.000 379.410 300.000 ;
    END
  END master_data_wdata_to_inter_i[31]
  PIN master_data_wdata_to_inter_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 296.000 386.310 300.000 ;
    END
  END master_data_wdata_to_inter_i[32]
  PIN master_data_wdata_to_inter_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 296.000 392.750 300.000 ;
    END
  END master_data_wdata_to_inter_i[33]
  PIN master_data_wdata_to_inter_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 296.000 399.650 300.000 ;
    END
  END master_data_wdata_to_inter_i[34]
  PIN master_data_wdata_to_inter_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 296.000 406.090 300.000 ;
    END
  END master_data_wdata_to_inter_i[35]
  PIN master_data_wdata_to_inter_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 296.000 412.990 300.000 ;
    END
  END master_data_wdata_to_inter_i[36]
  PIN master_data_wdata_to_inter_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 296.000 419.430 300.000 ;
    END
  END master_data_wdata_to_inter_i[37]
  PIN master_data_wdata_to_inter_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 296.000 426.330 300.000 ;
    END
  END master_data_wdata_to_inter_i[38]
  PIN master_data_wdata_to_inter_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 296.000 432.770 300.000 ;
    END
  END master_data_wdata_to_inter_i[39]
  PIN master_data_wdata_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 296.000 83.170 300.000 ;
    END
  END master_data_wdata_to_inter_i[3]
  PIN master_data_wdata_to_inter_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 296.000 439.210 300.000 ;
    END
  END master_data_wdata_to_inter_i[40]
  PIN master_data_wdata_to_inter_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 296.000 446.110 300.000 ;
    END
  END master_data_wdata_to_inter_i[41]
  PIN master_data_wdata_to_inter_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 296.000 452.550 300.000 ;
    END
  END master_data_wdata_to_inter_i[42]
  PIN master_data_wdata_to_inter_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 296.000 459.450 300.000 ;
    END
  END master_data_wdata_to_inter_i[43]
  PIN master_data_wdata_to_inter_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 296.000 465.890 300.000 ;
    END
  END master_data_wdata_to_inter_i[44]
  PIN master_data_wdata_to_inter_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 296.000 472.790 300.000 ;
    END
  END master_data_wdata_to_inter_i[45]
  PIN master_data_wdata_to_inter_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 296.000 479.230 300.000 ;
    END
  END master_data_wdata_to_inter_i[46]
  PIN master_data_wdata_to_inter_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 296.000 485.670 300.000 ;
    END
  END master_data_wdata_to_inter_i[47]
  PIN master_data_wdata_to_inter_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 296.000 492.570 300.000 ;
    END
  END master_data_wdata_to_inter_i[48]
  PIN master_data_wdata_to_inter_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 296.000 499.010 300.000 ;
    END
  END master_data_wdata_to_inter_i[49]
  PIN master_data_wdata_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 296.000 96.050 300.000 ;
    END
  END master_data_wdata_to_inter_i[4]
  PIN master_data_wdata_to_inter_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 296.000 505.910 300.000 ;
    END
  END master_data_wdata_to_inter_i[50]
  PIN master_data_wdata_to_inter_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 296.000 512.350 300.000 ;
    END
  END master_data_wdata_to_inter_i[51]
  PIN master_data_wdata_to_inter_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 296.000 519.250 300.000 ;
    END
  END master_data_wdata_to_inter_i[52]
  PIN master_data_wdata_to_inter_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 296.000 525.690 300.000 ;
    END
  END master_data_wdata_to_inter_i[53]
  PIN master_data_wdata_to_inter_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 296.000 532.590 300.000 ;
    END
  END master_data_wdata_to_inter_i[54]
  PIN master_data_wdata_to_inter_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 296.000 539.030 300.000 ;
    END
  END master_data_wdata_to_inter_i[55]
  PIN master_data_wdata_to_inter_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 296.000 545.470 300.000 ;
    END
  END master_data_wdata_to_inter_i[56]
  PIN master_data_wdata_to_inter_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 296.000 552.370 300.000 ;
    END
  END master_data_wdata_to_inter_i[57]
  PIN master_data_wdata_to_inter_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 296.000 558.810 300.000 ;
    END
  END master_data_wdata_to_inter_i[58]
  PIN master_data_wdata_to_inter_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 296.000 565.710 300.000 ;
    END
  END master_data_wdata_to_inter_i[59]
  PIN master_data_wdata_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 296.000 109.390 300.000 ;
    END
  END master_data_wdata_to_inter_i[5]
  PIN master_data_wdata_to_inter_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 296.000 572.150 300.000 ;
    END
  END master_data_wdata_to_inter_i[60]
  PIN master_data_wdata_to_inter_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 296.000 579.050 300.000 ;
    END
  END master_data_wdata_to_inter_i[61]
  PIN master_data_wdata_to_inter_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 296.000 585.490 300.000 ;
    END
  END master_data_wdata_to_inter_i[62]
  PIN master_data_wdata_to_inter_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 296.000 591.930 300.000 ;
    END
  END master_data_wdata_to_inter_i[63]
  PIN master_data_wdata_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 296.000 122.730 300.000 ;
    END
  END master_data_wdata_to_inter_i[6]
  PIN master_data_wdata_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 296.000 136.070 300.000 ;
    END
  END master_data_wdata_to_inter_i[7]
  PIN master_data_wdata_to_inter_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 296.000 147.110 300.000 ;
    END
  END master_data_wdata_to_inter_i[8]
  PIN master_data_wdata_to_inter_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 296.000 158.150 300.000 ;
    END
  END master_data_wdata_to_inter_i[9]
  PIN master_data_we_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 296.000 27.510 300.000 ;
    END
  END master_data_we_to_inter_i[0]
  PIN master_data_we_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 296.000 56.490 300.000 ;
    END
  END master_data_we_to_inter_i[1]
  PIN rxd_uart
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 29.960 1700.000 30.560 ;
    END
  END rxd_uart
  PIN rxd_uart_to_mem
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 89.800 1700.000 90.400 ;
    END
  END rxd_uart_to_mem
  PIN slave_data_addr_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 296.000 594.230 300.000 ;
    END
  END slave_data_addr_to_inter_o[0]
  PIN slave_data_addr_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 296.000 753.850 300.000 ;
    END
  END slave_data_addr_to_inter_o[10]
  PIN slave_data_addr_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 296.000 767.190 300.000 ;
    END
  END slave_data_addr_to_inter_o[11]
  PIN slave_data_addr_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 296.000 780.530 300.000 ;
    END
  END slave_data_addr_to_inter_o[12]
  PIN slave_data_addr_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 296.000 793.410 300.000 ;
    END
  END slave_data_addr_to_inter_o[13]
  PIN slave_data_addr_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 296.000 806.750 300.000 ;
    END
  END slave_data_addr_to_inter_o[14]
  PIN slave_data_addr_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 296.000 820.090 300.000 ;
    END
  END slave_data_addr_to_inter_o[15]
  PIN slave_data_addr_to_inter_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 296.000 833.430 300.000 ;
    END
  END slave_data_addr_to_inter_o[16]
  PIN slave_data_addr_to_inter_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 296.000 844.470 300.000 ;
    END
  END slave_data_addr_to_inter_o[17]
  PIN slave_data_addr_to_inter_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.230 296.000 855.510 300.000 ;
    END
  END slave_data_addr_to_inter_o[18]
  PIN slave_data_addr_to_inter_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 296.000 866.550 300.000 ;
    END
  END slave_data_addr_to_inter_o[19]
  PIN slave_data_addr_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 296.000 614.470 300.000 ;
    END
  END slave_data_addr_to_inter_o[1]
  PIN slave_data_addr_to_inter_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 296.000 877.590 300.000 ;
    END
  END slave_data_addr_to_inter_o[20]
  PIN slave_data_addr_to_inter_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 296.000 888.630 300.000 ;
    END
  END slave_data_addr_to_inter_o[21]
  PIN slave_data_addr_to_inter_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 296.000 899.670 300.000 ;
    END
  END slave_data_addr_to_inter_o[22]
  PIN slave_data_addr_to_inter_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.430 296.000 910.710 300.000 ;
    END
  END slave_data_addr_to_inter_o[23]
  PIN slave_data_addr_to_inter_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 296.000 922.210 300.000 ;
    END
  END slave_data_addr_to_inter_o[24]
  PIN slave_data_addr_to_inter_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.970 296.000 933.250 300.000 ;
    END
  END slave_data_addr_to_inter_o[25]
  PIN slave_data_addr_to_inter_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 296.000 944.290 300.000 ;
    END
  END slave_data_addr_to_inter_o[26]
  PIN slave_data_addr_to_inter_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 296.000 955.330 300.000 ;
    END
  END slave_data_addr_to_inter_o[27]
  PIN slave_data_addr_to_inter_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 296.000 966.370 300.000 ;
    END
  END slave_data_addr_to_inter_o[28]
  PIN slave_data_addr_to_inter_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 296.000 977.410 300.000 ;
    END
  END slave_data_addr_to_inter_o[29]
  PIN slave_data_addr_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 296.000 634.250 300.000 ;
    END
  END slave_data_addr_to_inter_o[2]
  PIN slave_data_addr_to_inter_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 296.000 988.450 300.000 ;
    END
  END slave_data_addr_to_inter_o[30]
  PIN slave_data_addr_to_inter_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.210 296.000 999.490 300.000 ;
    END
  END slave_data_addr_to_inter_o[31]
  PIN slave_data_addr_to_inter_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 296.000 1010.530 300.000 ;
    END
  END slave_data_addr_to_inter_o[32]
  PIN slave_data_addr_to_inter_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.290 296.000 1021.570 300.000 ;
    END
  END slave_data_addr_to_inter_o[33]
  PIN slave_data_addr_to_inter_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 296.000 1032.610 300.000 ;
    END
  END slave_data_addr_to_inter_o[34]
  PIN slave_data_addr_to_inter_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 296.000 1043.650 300.000 ;
    END
  END slave_data_addr_to_inter_o[35]
  PIN slave_data_addr_to_inter_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 296.000 1054.690 300.000 ;
    END
  END slave_data_addr_to_inter_o[36]
  PIN slave_data_addr_to_inter_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 296.000 1065.730 300.000 ;
    END
  END slave_data_addr_to_inter_o[37]
  PIN slave_data_addr_to_inter_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 296.000 1076.770 300.000 ;
    END
  END slave_data_addr_to_inter_o[38]
  PIN slave_data_addr_to_inter_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 296.000 1087.810 300.000 ;
    END
  END slave_data_addr_to_inter_o[39]
  PIN slave_data_addr_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 296.000 654.030 300.000 ;
    END
  END slave_data_addr_to_inter_o[3]
  PIN slave_data_addr_to_inter_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 296.000 1099.310 300.000 ;
    END
  END slave_data_addr_to_inter_o[40]
  PIN slave_data_addr_to_inter_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 296.000 1110.350 300.000 ;
    END
  END slave_data_addr_to_inter_o[41]
  PIN slave_data_addr_to_inter_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 296.000 1121.390 300.000 ;
    END
  END slave_data_addr_to_inter_o[42]
  PIN slave_data_addr_to_inter_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.150 296.000 1132.430 300.000 ;
    END
  END slave_data_addr_to_inter_o[43]
  PIN slave_data_addr_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 296.000 674.270 300.000 ;
    END
  END slave_data_addr_to_inter_o[4]
  PIN slave_data_addr_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 296.000 687.150 300.000 ;
    END
  END slave_data_addr_to_inter_o[5]
  PIN slave_data_addr_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 296.000 700.490 300.000 ;
    END
  END slave_data_addr_to_inter_o[6]
  PIN slave_data_addr_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 296.000 713.830 300.000 ;
    END
  END slave_data_addr_to_inter_o[7]
  PIN slave_data_addr_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 296.000 727.170 300.000 ;
    END
  END slave_data_addr_to_inter_o[8]
  PIN slave_data_addr_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 296.000 740.510 300.000 ;
    END
  END slave_data_addr_to_inter_o[9]
  PIN slave_data_addr_to_inter_ro_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 296.000 596.530 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[0]
  PIN slave_data_addr_to_inter_ro_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 296.000 756.150 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[10]
  PIN slave_data_addr_to_inter_ro_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 296.000 769.030 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[11]
  PIN slave_data_addr_to_inter_ro_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 296.000 782.370 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[12]
  PIN slave_data_addr_to_inter_ro_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 296.000 795.710 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[13]
  PIN slave_data_addr_to_inter_ro_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 296.000 809.050 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[14]
  PIN slave_data_addr_to_inter_ro_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 296.000 822.390 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[15]
  PIN slave_data_addr_to_inter_ro_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 296.000 835.730 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[16]
  PIN slave_data_addr_to_inter_ro_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 296.000 846.770 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[17]
  PIN slave_data_addr_to_inter_ro_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.530 296.000 857.810 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[18]
  PIN slave_data_addr_to_inter_ro_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 296.000 868.850 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[19]
  PIN slave_data_addr_to_inter_ro_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 296.000 616.310 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[1]
  PIN slave_data_addr_to_inter_ro_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 296.000 879.890 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[20]
  PIN slave_data_addr_to_inter_ro_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.650 296.000 890.930 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[21]
  PIN slave_data_addr_to_inter_ro_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 296.000 901.970 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[22]
  PIN slave_data_addr_to_inter_ro_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.730 296.000 913.010 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[23]
  PIN slave_data_addr_to_inter_ro_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 296.000 924.050 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[24]
  PIN slave_data_addr_to_inter_ro_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 296.000 935.090 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[25]
  PIN slave_data_addr_to_inter_ro_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.850 296.000 946.130 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[26]
  PIN slave_data_addr_to_inter_ro_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 296.000 957.630 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[27]
  PIN slave_data_addr_to_inter_ro_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 296.000 968.670 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[28]
  PIN slave_data_addr_to_inter_ro_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 296.000 979.710 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[29]
  PIN slave_data_addr_to_inter_ro_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 296.000 636.550 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[2]
  PIN slave_data_addr_to_inter_ro_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 296.000 990.750 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[30]
  PIN slave_data_addr_to_inter_ro_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 296.000 1001.790 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[31]
  PIN slave_data_addr_to_inter_ro_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 296.000 1012.830 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[32]
  PIN slave_data_addr_to_inter_ro_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.590 296.000 1023.870 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[33]
  PIN slave_data_addr_to_inter_ro_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.630 296.000 1034.910 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[34]
  PIN slave_data_addr_to_inter_ro_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.670 296.000 1045.950 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[35]
  PIN slave_data_addr_to_inter_ro_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 296.000 1056.990 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[36]
  PIN slave_data_addr_to_inter_ro_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.750 296.000 1068.030 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[37]
  PIN slave_data_addr_to_inter_ro_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 296.000 1079.070 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[38]
  PIN slave_data_addr_to_inter_ro_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.830 296.000 1090.110 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[39]
  PIN slave_data_addr_to_inter_ro_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 296.000 656.330 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[3]
  PIN slave_data_addr_to_inter_ro_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.870 296.000 1101.150 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[40]
  PIN slave_data_addr_to_inter_ro_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 296.000 1112.190 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[41]
  PIN slave_data_addr_to_inter_ro_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.950 296.000 1123.230 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[42]
  PIN slave_data_addr_to_inter_ro_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 296.000 1134.730 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[43]
  PIN slave_data_addr_to_inter_ro_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 296.000 676.110 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[4]
  PIN slave_data_addr_to_inter_ro_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 296.000 689.450 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[5]
  PIN slave_data_addr_to_inter_ro_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 296.000 702.790 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[6]
  PIN slave_data_addr_to_inter_ro_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 296.000 716.130 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[7]
  PIN slave_data_addr_to_inter_ro_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 296.000 729.470 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[8]
  PIN slave_data_addr_to_inter_ro_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 296.000 742.810 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[9]
  PIN slave_data_be_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 296.000 598.830 300.000 ;
    END
  END slave_data_be_to_inter_o[0]
  PIN slave_data_be_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 296.000 757.990 300.000 ;
    END
  END slave_data_be_to_inter_o[10]
  PIN slave_data_be_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 296.000 771.330 300.000 ;
    END
  END slave_data_be_to_inter_o[11]
  PIN slave_data_be_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 296.000 784.670 300.000 ;
    END
  END slave_data_be_to_inter_o[12]
  PIN slave_data_be_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 296.000 798.010 300.000 ;
    END
  END slave_data_be_to_inter_o[13]
  PIN slave_data_be_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 296.000 811.350 300.000 ;
    END
  END slave_data_be_to_inter_o[14]
  PIN slave_data_be_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 296.000 824.690 300.000 ;
    END
  END slave_data_be_to_inter_o[15]
  PIN slave_data_be_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 296.000 618.610 300.000 ;
    END
  END slave_data_be_to_inter_o[1]
  PIN slave_data_be_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 296.000 638.850 300.000 ;
    END
  END slave_data_be_to_inter_o[2]
  PIN slave_data_be_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 296.000 658.630 300.000 ;
    END
  END slave_data_be_to_inter_o[3]
  PIN slave_data_be_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 296.000 678.410 300.000 ;
    END
  END slave_data_be_to_inter_o[4]
  PIN slave_data_be_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 296.000 691.750 300.000 ;
    END
  END slave_data_be_to_inter_o[5]
  PIN slave_data_be_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 296.000 705.090 300.000 ;
    END
  END slave_data_be_to_inter_o[6]
  PIN slave_data_be_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 296.000 718.430 300.000 ;
    END
  END slave_data_be_to_inter_o[7]
  PIN slave_data_be_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 296.000 731.770 300.000 ;
    END
  END slave_data_be_to_inter_o[8]
  PIN slave_data_be_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 296.000 745.110 300.000 ;
    END
  END slave_data_be_to_inter_o[9]
  PIN slave_data_rdata_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 296.000 601.130 300.000 ;
    END
  END slave_data_rdata_to_inter_i[0]
  PIN slave_data_rdata_to_inter_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.870 296.000 1515.150 300.000 ;
    END
  END slave_data_rdata_to_inter_i[100]
  PIN slave_data_rdata_to_inter_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.770 296.000 1522.050 300.000 ;
    END
  END slave_data_rdata_to_inter_i[101]
  PIN slave_data_rdata_to_inter_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.210 296.000 1528.490 300.000 ;
    END
  END slave_data_rdata_to_inter_i[102]
  PIN slave_data_rdata_to_inter_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.110 296.000 1535.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[103]
  PIN slave_data_rdata_to_inter_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.550 296.000 1541.830 300.000 ;
    END
  END slave_data_rdata_to_inter_i[104]
  PIN slave_data_rdata_to_inter_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.990 296.000 1548.270 300.000 ;
    END
  END slave_data_rdata_to_inter_i[105]
  PIN slave_data_rdata_to_inter_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.890 296.000 1555.170 300.000 ;
    END
  END slave_data_rdata_to_inter_i[106]
  PIN slave_data_rdata_to_inter_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.330 296.000 1561.610 300.000 ;
    END
  END slave_data_rdata_to_inter_i[107]
  PIN slave_data_rdata_to_inter_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 296.000 1568.510 300.000 ;
    END
  END slave_data_rdata_to_inter_i[108]
  PIN slave_data_rdata_to_inter_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.670 296.000 1574.950 300.000 ;
    END
  END slave_data_rdata_to_inter_i[109]
  PIN slave_data_rdata_to_inter_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 296.000 760.290 300.000 ;
    END
  END slave_data_rdata_to_inter_i[10]
  PIN slave_data_rdata_to_inter_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.570 296.000 1581.850 300.000 ;
    END
  END slave_data_rdata_to_inter_i[110]
  PIN slave_data_rdata_to_inter_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.010 296.000 1588.290 300.000 ;
    END
  END slave_data_rdata_to_inter_i[111]
  PIN slave_data_rdata_to_inter_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.910 296.000 1595.190 300.000 ;
    END
  END slave_data_rdata_to_inter_i[112]
  PIN slave_data_rdata_to_inter_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1601.350 296.000 1601.630 300.000 ;
    END
  END slave_data_rdata_to_inter_i[113]
  PIN slave_data_rdata_to_inter_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.790 296.000 1608.070 300.000 ;
    END
  END slave_data_rdata_to_inter_i[114]
  PIN slave_data_rdata_to_inter_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.690 296.000 1614.970 300.000 ;
    END
  END slave_data_rdata_to_inter_i[115]
  PIN slave_data_rdata_to_inter_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.130 296.000 1621.410 300.000 ;
    END
  END slave_data_rdata_to_inter_i[116]
  PIN slave_data_rdata_to_inter_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.030 296.000 1628.310 300.000 ;
    END
  END slave_data_rdata_to_inter_i[117]
  PIN slave_data_rdata_to_inter_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.470 296.000 1634.750 300.000 ;
    END
  END slave_data_rdata_to_inter_i[118]
  PIN slave_data_rdata_to_inter_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.370 296.000 1641.650 300.000 ;
    END
  END slave_data_rdata_to_inter_i[119]
  PIN slave_data_rdata_to_inter_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 296.000 773.630 300.000 ;
    END
  END slave_data_rdata_to_inter_i[11]
  PIN slave_data_rdata_to_inter_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.810 296.000 1648.090 300.000 ;
    END
  END slave_data_rdata_to_inter_i[120]
  PIN slave_data_rdata_to_inter_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.250 296.000 1654.530 300.000 ;
    END
  END slave_data_rdata_to_inter_i[121]
  PIN slave_data_rdata_to_inter_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.150 296.000 1661.430 300.000 ;
    END
  END slave_data_rdata_to_inter_i[122]
  PIN slave_data_rdata_to_inter_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.590 296.000 1667.870 300.000 ;
    END
  END slave_data_rdata_to_inter_i[123]
  PIN slave_data_rdata_to_inter_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 296.000 1674.770 300.000 ;
    END
  END slave_data_rdata_to_inter_i[124]
  PIN slave_data_rdata_to_inter_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.930 296.000 1681.210 300.000 ;
    END
  END slave_data_rdata_to_inter_i[125]
  PIN slave_data_rdata_to_inter_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.830 296.000 1688.110 300.000 ;
    END
  END slave_data_rdata_to_inter_i[126]
  PIN slave_data_rdata_to_inter_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.270 296.000 1694.550 300.000 ;
    END
  END slave_data_rdata_to_inter_i[127]
  PIN slave_data_rdata_to_inter_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 296.000 786.970 300.000 ;
    END
  END slave_data_rdata_to_inter_i[12]
  PIN slave_data_rdata_to_inter_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 296.000 800.310 300.000 ;
    END
  END slave_data_rdata_to_inter_i[13]
  PIN slave_data_rdata_to_inter_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 296.000 813.650 300.000 ;
    END
  END slave_data_rdata_to_inter_i[14]
  PIN slave_data_rdata_to_inter_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 296.000 826.990 300.000 ;
    END
  END slave_data_rdata_to_inter_i[15]
  PIN slave_data_rdata_to_inter_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 296.000 838.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[16]
  PIN slave_data_rdata_to_inter_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 296.000 849.070 300.000 ;
    END
  END slave_data_rdata_to_inter_i[17]
  PIN slave_data_rdata_to_inter_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 296.000 860.110 300.000 ;
    END
  END slave_data_rdata_to_inter_i[18]
  PIN slave_data_rdata_to_inter_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 296.000 871.150 300.000 ;
    END
  END slave_data_rdata_to_inter_i[19]
  PIN slave_data_rdata_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 296.000 620.910 300.000 ;
    END
  END slave_data_rdata_to_inter_i[1]
  PIN slave_data_rdata_to_inter_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.910 296.000 882.190 300.000 ;
    END
  END slave_data_rdata_to_inter_i[20]
  PIN slave_data_rdata_to_inter_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 296.000 893.230 300.000 ;
    END
  END slave_data_rdata_to_inter_i[21]
  PIN slave_data_rdata_to_inter_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 296.000 904.270 300.000 ;
    END
  END slave_data_rdata_to_inter_i[22]
  PIN slave_data_rdata_to_inter_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 296.000 915.310 300.000 ;
    END
  END slave_data_rdata_to_inter_i[23]
  PIN slave_data_rdata_to_inter_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 296.000 926.350 300.000 ;
    END
  END slave_data_rdata_to_inter_i[24]
  PIN slave_data_rdata_to_inter_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 296.000 937.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[25]
  PIN slave_data_rdata_to_inter_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 296.000 948.430 300.000 ;
    END
  END slave_data_rdata_to_inter_i[26]
  PIN slave_data_rdata_to_inter_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 296.000 959.470 300.000 ;
    END
  END slave_data_rdata_to_inter_i[27]
  PIN slave_data_rdata_to_inter_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 296.000 970.510 300.000 ;
    END
  END slave_data_rdata_to_inter_i[28]
  PIN slave_data_rdata_to_inter_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 296.000 981.550 300.000 ;
    END
  END slave_data_rdata_to_inter_i[29]
  PIN slave_data_rdata_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 296.000 640.690 300.000 ;
    END
  END slave_data_rdata_to_inter_i[2]
  PIN slave_data_rdata_to_inter_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.770 296.000 993.050 300.000 ;
    END
  END slave_data_rdata_to_inter_i[30]
  PIN slave_data_rdata_to_inter_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.810 296.000 1004.090 300.000 ;
    END
  END slave_data_rdata_to_inter_i[31]
  PIN slave_data_rdata_to_inter_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.850 296.000 1015.130 300.000 ;
    END
  END slave_data_rdata_to_inter_i[32]
  PIN slave_data_rdata_to_inter_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.890 296.000 1026.170 300.000 ;
    END
  END slave_data_rdata_to_inter_i[33]
  PIN slave_data_rdata_to_inter_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 296.000 1037.210 300.000 ;
    END
  END slave_data_rdata_to_inter_i[34]
  PIN slave_data_rdata_to_inter_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.970 296.000 1048.250 300.000 ;
    END
  END slave_data_rdata_to_inter_i[35]
  PIN slave_data_rdata_to_inter_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 296.000 1059.290 300.000 ;
    END
  END slave_data_rdata_to_inter_i[36]
  PIN slave_data_rdata_to_inter_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 296.000 1070.330 300.000 ;
    END
  END slave_data_rdata_to_inter_i[37]
  PIN slave_data_rdata_to_inter_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.090 296.000 1081.370 300.000 ;
    END
  END slave_data_rdata_to_inter_i[38]
  PIN slave_data_rdata_to_inter_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.130 296.000 1092.410 300.000 ;
    END
  END slave_data_rdata_to_inter_i[39]
  PIN slave_data_rdata_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 296.000 660.930 300.000 ;
    END
  END slave_data_rdata_to_inter_i[3]
  PIN slave_data_rdata_to_inter_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.170 296.000 1103.450 300.000 ;
    END
  END slave_data_rdata_to_inter_i[40]
  PIN slave_data_rdata_to_inter_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 296.000 1114.490 300.000 ;
    END
  END slave_data_rdata_to_inter_i[41]
  PIN slave_data_rdata_to_inter_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.250 296.000 1125.530 300.000 ;
    END
  END slave_data_rdata_to_inter_i[42]
  PIN slave_data_rdata_to_inter_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.290 296.000 1136.570 300.000 ;
    END
  END slave_data_rdata_to_inter_i[43]
  PIN slave_data_rdata_to_inter_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 296.000 1143.470 300.000 ;
    END
  END slave_data_rdata_to_inter_i[44]
  PIN slave_data_rdata_to_inter_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 296.000 1149.910 300.000 ;
    END
  END slave_data_rdata_to_inter_i[45]
  PIN slave_data_rdata_to_inter_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.530 296.000 1156.810 300.000 ;
    END
  END slave_data_rdata_to_inter_i[46]
  PIN slave_data_rdata_to_inter_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.970 296.000 1163.250 300.000 ;
    END
  END slave_data_rdata_to_inter_i[47]
  PIN slave_data_rdata_to_inter_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 296.000 1170.150 300.000 ;
    END
  END slave_data_rdata_to_inter_i[48]
  PIN slave_data_rdata_to_inter_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.310 296.000 1176.590 300.000 ;
    END
  END slave_data_rdata_to_inter_i[49]
  PIN slave_data_rdata_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 296.000 680.710 300.000 ;
    END
  END slave_data_rdata_to_inter_i[4]
  PIN slave_data_rdata_to_inter_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.750 296.000 1183.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[50]
  PIN slave_data_rdata_to_inter_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.650 296.000 1189.930 300.000 ;
    END
  END slave_data_rdata_to_inter_i[51]
  PIN slave_data_rdata_to_inter_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.090 296.000 1196.370 300.000 ;
    END
  END slave_data_rdata_to_inter_i[52]
  PIN slave_data_rdata_to_inter_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.990 296.000 1203.270 300.000 ;
    END
  END slave_data_rdata_to_inter_i[53]
  PIN slave_data_rdata_to_inter_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.430 296.000 1209.710 300.000 ;
    END
  END slave_data_rdata_to_inter_i[54]
  PIN slave_data_rdata_to_inter_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.330 296.000 1216.610 300.000 ;
    END
  END slave_data_rdata_to_inter_i[55]
  PIN slave_data_rdata_to_inter_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1222.770 296.000 1223.050 300.000 ;
    END
  END slave_data_rdata_to_inter_i[56]
  PIN slave_data_rdata_to_inter_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.210 296.000 1229.490 300.000 ;
    END
  END slave_data_rdata_to_inter_i[57]
  PIN slave_data_rdata_to_inter_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.110 296.000 1236.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[58]
  PIN slave_data_rdata_to_inter_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 296.000 1242.830 300.000 ;
    END
  END slave_data_rdata_to_inter_i[59]
  PIN slave_data_rdata_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 296.000 694.050 300.000 ;
    END
  END slave_data_rdata_to_inter_i[5]
  PIN slave_data_rdata_to_inter_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 296.000 1249.730 300.000 ;
    END
  END slave_data_rdata_to_inter_i[60]
  PIN slave_data_rdata_to_inter_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 296.000 1256.170 300.000 ;
    END
  END slave_data_rdata_to_inter_i[61]
  PIN slave_data_rdata_to_inter_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.790 296.000 1263.070 300.000 ;
    END
  END slave_data_rdata_to_inter_i[62]
  PIN slave_data_rdata_to_inter_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.230 296.000 1269.510 300.000 ;
    END
  END slave_data_rdata_to_inter_i[63]
  PIN slave_data_rdata_to_inter_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.130 296.000 1276.410 300.000 ;
    END
  END slave_data_rdata_to_inter_i[64]
  PIN slave_data_rdata_to_inter_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.570 296.000 1282.850 300.000 ;
    END
  END slave_data_rdata_to_inter_i[65]
  PIN slave_data_rdata_to_inter_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 296.000 1289.290 300.000 ;
    END
  END slave_data_rdata_to_inter_i[66]
  PIN slave_data_rdata_to_inter_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.910 296.000 1296.190 300.000 ;
    END
  END slave_data_rdata_to_inter_i[67]
  PIN slave_data_rdata_to_inter_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.350 296.000 1302.630 300.000 ;
    END
  END slave_data_rdata_to_inter_i[68]
  PIN slave_data_rdata_to_inter_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.250 296.000 1309.530 300.000 ;
    END
  END slave_data_rdata_to_inter_i[69]
  PIN slave_data_rdata_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 296.000 707.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[6]
  PIN slave_data_rdata_to_inter_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.690 296.000 1315.970 300.000 ;
    END
  END slave_data_rdata_to_inter_i[70]
  PIN slave_data_rdata_to_inter_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.590 296.000 1322.870 300.000 ;
    END
  END slave_data_rdata_to_inter_i[71]
  PIN slave_data_rdata_to_inter_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.030 296.000 1329.310 300.000 ;
    END
  END slave_data_rdata_to_inter_i[72]
  PIN slave_data_rdata_to_inter_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 296.000 1335.750 300.000 ;
    END
  END slave_data_rdata_to_inter_i[73]
  PIN slave_data_rdata_to_inter_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 296.000 1342.650 300.000 ;
    END
  END slave_data_rdata_to_inter_i[74]
  PIN slave_data_rdata_to_inter_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.810 296.000 1349.090 300.000 ;
    END
  END slave_data_rdata_to_inter_i[75]
  PIN slave_data_rdata_to_inter_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 296.000 1355.990 300.000 ;
    END
  END slave_data_rdata_to_inter_i[76]
  PIN slave_data_rdata_to_inter_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 296.000 1362.430 300.000 ;
    END
  END slave_data_rdata_to_inter_i[77]
  PIN slave_data_rdata_to_inter_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.050 296.000 1369.330 300.000 ;
    END
  END slave_data_rdata_to_inter_i[78]
  PIN slave_data_rdata_to_inter_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.490 296.000 1375.770 300.000 ;
    END
  END slave_data_rdata_to_inter_i[79]
  PIN slave_data_rdata_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 296.000 720.730 300.000 ;
    END
  END slave_data_rdata_to_inter_i[7]
  PIN slave_data_rdata_to_inter_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.390 296.000 1382.670 300.000 ;
    END
  END slave_data_rdata_to_inter_i[80]
  PIN slave_data_rdata_to_inter_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.830 296.000 1389.110 300.000 ;
    END
  END slave_data_rdata_to_inter_i[81]
  PIN slave_data_rdata_to_inter_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.270 296.000 1395.550 300.000 ;
    END
  END slave_data_rdata_to_inter_i[82]
  PIN slave_data_rdata_to_inter_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.170 296.000 1402.450 300.000 ;
    END
  END slave_data_rdata_to_inter_i[83]
  PIN slave_data_rdata_to_inter_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.610 296.000 1408.890 300.000 ;
    END
  END slave_data_rdata_to_inter_i[84]
  PIN slave_data_rdata_to_inter_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.510 296.000 1415.790 300.000 ;
    END
  END slave_data_rdata_to_inter_i[85]
  PIN slave_data_rdata_to_inter_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.950 296.000 1422.230 300.000 ;
    END
  END slave_data_rdata_to_inter_i[86]
  PIN slave_data_rdata_to_inter_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.850 296.000 1429.130 300.000 ;
    END
  END slave_data_rdata_to_inter_i[87]
  PIN slave_data_rdata_to_inter_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 296.000 1435.570 300.000 ;
    END
  END slave_data_rdata_to_inter_i[88]
  PIN slave_data_rdata_to_inter_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.730 296.000 1442.010 300.000 ;
    END
  END slave_data_rdata_to_inter_i[89]
  PIN slave_data_rdata_to_inter_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 296.000 733.610 300.000 ;
    END
  END slave_data_rdata_to_inter_i[8]
  PIN slave_data_rdata_to_inter_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.630 296.000 1448.910 300.000 ;
    END
  END slave_data_rdata_to_inter_i[90]
  PIN slave_data_rdata_to_inter_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.070 296.000 1455.350 300.000 ;
    END
  END slave_data_rdata_to_inter_i[91]
  PIN slave_data_rdata_to_inter_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 296.000 1462.250 300.000 ;
    END
  END slave_data_rdata_to_inter_i[92]
  PIN slave_data_rdata_to_inter_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 296.000 1468.690 300.000 ;
    END
  END slave_data_rdata_to_inter_i[93]
  PIN slave_data_rdata_to_inter_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 296.000 1475.590 300.000 ;
    END
  END slave_data_rdata_to_inter_i[94]
  PIN slave_data_rdata_to_inter_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.750 296.000 1482.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[95]
  PIN slave_data_rdata_to_inter_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.650 296.000 1488.930 300.000 ;
    END
  END slave_data_rdata_to_inter_i[96]
  PIN slave_data_rdata_to_inter_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.090 296.000 1495.370 300.000 ;
    END
  END slave_data_rdata_to_inter_i[97]
  PIN slave_data_rdata_to_inter_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.530 296.000 1501.810 300.000 ;
    END
  END slave_data_rdata_to_inter_i[98]
  PIN slave_data_rdata_to_inter_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.430 296.000 1508.710 300.000 ;
    END
  END slave_data_rdata_to_inter_i[99]
  PIN slave_data_rdata_to_inter_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 296.000 746.950 300.000 ;
    END
  END slave_data_rdata_to_inter_i[9]
  PIN slave_data_rdata_to_inter_ro_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 296.000 603.430 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[0]
  PIN slave_data_rdata_to_inter_ro_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.170 296.000 1517.450 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[100]
  PIN slave_data_rdata_to_inter_ro_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.070 296.000 1524.350 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[101]
  PIN slave_data_rdata_to_inter_ro_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.510 296.000 1530.790 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[102]
  PIN slave_data_rdata_to_inter_ro_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.950 296.000 1537.230 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[103]
  PIN slave_data_rdata_to_inter_ro_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1543.850 296.000 1544.130 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[104]
  PIN slave_data_rdata_to_inter_ro_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.290 296.000 1550.570 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[105]
  PIN slave_data_rdata_to_inter_ro_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 296.000 1557.470 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[106]
  PIN slave_data_rdata_to_inter_ro_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.630 296.000 1563.910 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[107]
  PIN slave_data_rdata_to_inter_ro_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.530 296.000 1570.810 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[108]
  PIN slave_data_rdata_to_inter_ro_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.970 296.000 1577.250 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[109]
  PIN slave_data_rdata_to_inter_ro_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 296.000 762.590 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[10]
  PIN slave_data_rdata_to_inter_ro_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.410 296.000 1583.690 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[110]
  PIN slave_data_rdata_to_inter_ro_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.310 296.000 1590.590 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[111]
  PIN slave_data_rdata_to_inter_ro_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.750 296.000 1597.030 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[112]
  PIN slave_data_rdata_to_inter_ro_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 296.000 1603.930 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[113]
  PIN slave_data_rdata_to_inter_ro_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 296.000 1610.370 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[114]
  PIN slave_data_rdata_to_inter_ro_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.990 296.000 1617.270 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[115]
  PIN slave_data_rdata_to_inter_ro_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.430 296.000 1623.710 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[116]
  PIN slave_data_rdata_to_inter_ro_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.330 296.000 1630.610 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[117]
  PIN slave_data_rdata_to_inter_ro_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.770 296.000 1637.050 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[118]
  PIN slave_data_rdata_to_inter_ro_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.210 296.000 1643.490 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[119]
  PIN slave_data_rdata_to_inter_ro_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 296.000 775.930 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[11]
  PIN slave_data_rdata_to_inter_ro_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.110 296.000 1650.390 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[120]
  PIN slave_data_rdata_to_inter_ro_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.550 296.000 1656.830 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[121]
  PIN slave_data_rdata_to_inter_ro_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.450 296.000 1663.730 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[122]
  PIN slave_data_rdata_to_inter_ro_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.890 296.000 1670.170 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[123]
  PIN slave_data_rdata_to_inter_ro_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.790 296.000 1677.070 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[124]
  PIN slave_data_rdata_to_inter_ro_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.230 296.000 1683.510 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[125]
  PIN slave_data_rdata_to_inter_ro_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.670 296.000 1689.950 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[126]
  PIN slave_data_rdata_to_inter_ro_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.570 296.000 1696.850 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[127]
  PIN slave_data_rdata_to_inter_ro_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 296.000 789.270 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[12]
  PIN slave_data_rdata_to_inter_ro_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 296.000 802.610 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[13]
  PIN slave_data_rdata_to_inter_ro_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 296.000 815.950 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[14]
  PIN slave_data_rdata_to_inter_ro_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 296.000 828.830 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[15]
  PIN slave_data_rdata_to_inter_ro_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 296.000 839.870 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[16]
  PIN slave_data_rdata_to_inter_ro_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 296.000 851.370 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[17]
  PIN slave_data_rdata_to_inter_ro_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 296.000 862.410 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[18]
  PIN slave_data_rdata_to_inter_ro_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 296.000 873.450 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[19]
  PIN slave_data_rdata_to_inter_ro_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 296.000 623.210 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[1]
  PIN slave_data_rdata_to_inter_ro_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 296.000 884.490 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[20]
  PIN slave_data_rdata_to_inter_ro_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 296.000 895.530 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[21]
  PIN slave_data_rdata_to_inter_ro_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.290 296.000 906.570 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[22]
  PIN slave_data_rdata_to_inter_ro_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.330 296.000 917.610 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[23]
  PIN slave_data_rdata_to_inter_ro_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.370 296.000 928.650 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[24]
  PIN slave_data_rdata_to_inter_ro_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.410 296.000 939.690 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[25]
  PIN slave_data_rdata_to_inter_ro_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.450 296.000 950.730 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[26]
  PIN slave_data_rdata_to_inter_ro_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 296.000 961.770 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[27]
  PIN slave_data_rdata_to_inter_ro_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 296.000 972.810 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[28]
  PIN slave_data_rdata_to_inter_ro_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 296.000 983.850 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[29]
  PIN slave_data_rdata_to_inter_ro_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 296.000 642.990 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[2]
  PIN slave_data_rdata_to_inter_ro_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.610 296.000 994.890 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[30]
  PIN slave_data_rdata_to_inter_ro_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.650 296.000 1005.930 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[31]
  PIN slave_data_rdata_to_inter_ro_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 296.000 1016.970 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[32]
  PIN slave_data_rdata_to_inter_ro_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.190 296.000 1028.470 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[33]
  PIN slave_data_rdata_to_inter_ro_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.230 296.000 1039.510 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[34]
  PIN slave_data_rdata_to_inter_ro_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 296.000 1050.550 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[35]
  PIN slave_data_rdata_to_inter_ro_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.310 296.000 1061.590 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[36]
  PIN slave_data_rdata_to_inter_ro_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 296.000 1072.630 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[37]
  PIN slave_data_rdata_to_inter_ro_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.390 296.000 1083.670 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[38]
  PIN slave_data_rdata_to_inter_ro_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.430 296.000 1094.710 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[39]
  PIN slave_data_rdata_to_inter_ro_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 296.000 662.770 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[3]
  PIN slave_data_rdata_to_inter_ro_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.470 296.000 1105.750 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[40]
  PIN slave_data_rdata_to_inter_ro_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.510 296.000 1116.790 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[41]
  PIN slave_data_rdata_to_inter_ro_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.550 296.000 1127.830 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[42]
  PIN slave_data_rdata_to_inter_ro_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.590 296.000 1138.870 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[43]
  PIN slave_data_rdata_to_inter_ro_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.490 296.000 1145.770 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[44]
  PIN slave_data_rdata_to_inter_ro_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.930 296.000 1152.210 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[45]
  PIN slave_data_rdata_to_inter_ro_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.370 296.000 1158.650 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[46]
  PIN slave_data_rdata_to_inter_ro_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.270 296.000 1165.550 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[47]
  PIN slave_data_rdata_to_inter_ro_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.710 296.000 1171.990 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[48]
  PIN slave_data_rdata_to_inter_ro_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 296.000 1178.890 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[49]
  PIN slave_data_rdata_to_inter_ro_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 296.000 683.010 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[4]
  PIN slave_data_rdata_to_inter_ro_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 296.000 1185.330 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[50]
  PIN slave_data_rdata_to_inter_ro_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 296.000 1192.230 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[51]
  PIN slave_data_rdata_to_inter_ro_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.390 296.000 1198.670 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[52]
  PIN slave_data_rdata_to_inter_ro_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.290 296.000 1205.570 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[53]
  PIN slave_data_rdata_to_inter_ro_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.730 296.000 1212.010 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[54]
  PIN slave_data_rdata_to_inter_ro_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 296.000 1218.450 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[55]
  PIN slave_data_rdata_to_inter_ro_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.070 296.000 1225.350 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[56]
  PIN slave_data_rdata_to_inter_ro_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.510 296.000 1231.790 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[57]
  PIN slave_data_rdata_to_inter_ro_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.410 296.000 1238.690 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[58]
  PIN slave_data_rdata_to_inter_ro_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.850 296.000 1245.130 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[59]
  PIN slave_data_rdata_to_inter_ro_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 296.000 696.350 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[5]
  PIN slave_data_rdata_to_inter_ro_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.750 296.000 1252.030 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[60]
  PIN slave_data_rdata_to_inter_ro_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.190 296.000 1258.470 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[61]
  PIN slave_data_rdata_to_inter_ro_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.630 296.000 1264.910 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[62]
  PIN slave_data_rdata_to_inter_ro_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.530 296.000 1271.810 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[63]
  PIN slave_data_rdata_to_inter_ro_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.970 296.000 1278.250 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[64]
  PIN slave_data_rdata_to_inter_ro_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 296.000 1285.150 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[65]
  PIN slave_data_rdata_to_inter_ro_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 296.000 1291.590 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[66]
  PIN slave_data_rdata_to_inter_ro_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 296.000 1298.490 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[67]
  PIN slave_data_rdata_to_inter_ro_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.650 296.000 1304.930 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[68]
  PIN slave_data_rdata_to_inter_ro_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.550 296.000 1311.830 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[69]
  PIN slave_data_rdata_to_inter_ro_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 296.000 709.690 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[6]
  PIN slave_data_rdata_to_inter_ro_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.990 296.000 1318.270 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[70]
  PIN slave_data_rdata_to_inter_ro_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.430 296.000 1324.710 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[71]
  PIN slave_data_rdata_to_inter_ro_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.330 296.000 1331.610 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[72]
  PIN slave_data_rdata_to_inter_ro_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.770 296.000 1338.050 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[73]
  PIN slave_data_rdata_to_inter_ro_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.670 296.000 1344.950 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[74]
  PIN slave_data_rdata_to_inter_ro_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.110 296.000 1351.390 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[75]
  PIN slave_data_rdata_to_inter_ro_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.010 296.000 1358.290 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[76]
  PIN slave_data_rdata_to_inter_ro_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.450 296.000 1364.730 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[77]
  PIN slave_data_rdata_to_inter_ro_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.890 296.000 1371.170 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[78]
  PIN slave_data_rdata_to_inter_ro_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.790 296.000 1378.070 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[79]
  PIN slave_data_rdata_to_inter_ro_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 296.000 722.570 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[7]
  PIN slave_data_rdata_to_inter_ro_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.230 296.000 1384.510 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[80]
  PIN slave_data_rdata_to_inter_ro_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 296.000 1391.410 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[81]
  PIN slave_data_rdata_to_inter_ro_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 296.000 1397.850 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[82]
  PIN slave_data_rdata_to_inter_ro_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.470 296.000 1404.750 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[83]
  PIN slave_data_rdata_to_inter_ro_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 296.000 1411.190 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[84]
  PIN slave_data_rdata_to_inter_ro_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.810 296.000 1418.090 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[85]
  PIN slave_data_rdata_to_inter_ro_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.250 296.000 1424.530 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[86]
  PIN slave_data_rdata_to_inter_ro_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1430.690 296.000 1430.970 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[87]
  PIN slave_data_rdata_to_inter_ro_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.590 296.000 1437.870 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[88]
  PIN slave_data_rdata_to_inter_ro_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.030 296.000 1444.310 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[89]
  PIN slave_data_rdata_to_inter_ro_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 296.000 735.910 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[8]
  PIN slave_data_rdata_to_inter_ro_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.930 296.000 1451.210 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[90]
  PIN slave_data_rdata_to_inter_ro_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.370 296.000 1457.650 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[91]
  PIN slave_data_rdata_to_inter_ro_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.270 296.000 1464.550 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[92]
  PIN slave_data_rdata_to_inter_ro_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.710 296.000 1470.990 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[93]
  PIN slave_data_rdata_to_inter_ro_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.150 296.000 1477.430 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[94]
  PIN slave_data_rdata_to_inter_ro_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.050 296.000 1484.330 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[95]
  PIN slave_data_rdata_to_inter_ro_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 296.000 1490.770 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[96]
  PIN slave_data_rdata_to_inter_ro_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 296.000 1497.670 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[97]
  PIN slave_data_rdata_to_inter_ro_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 296.000 1504.110 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[98]
  PIN slave_data_rdata_to_inter_ro_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.730 296.000 1511.010 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[99]
  PIN slave_data_rdata_to_inter_ro_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 296.000 749.250 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[9]
  PIN slave_data_req_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 296.000 605.270 300.000 ;
    END
  END slave_data_req_to_inter_o[0]
  PIN slave_data_req_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 296.000 625.510 300.000 ;
    END
  END slave_data_req_to_inter_o[1]
  PIN slave_data_req_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 296.000 645.290 300.000 ;
    END
  END slave_data_req_to_inter_o[2]
  PIN slave_data_req_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 296.000 665.070 300.000 ;
    END
  END slave_data_req_to_inter_o[3]
  PIN slave_data_req_to_inter_ro_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 296.000 607.570 300.000 ;
    END
  END slave_data_req_to_inter_ro_o[0]
  PIN slave_data_req_to_inter_ro_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 296.000 627.350 300.000 ;
    END
  END slave_data_req_to_inter_ro_o[1]
  PIN slave_data_req_to_inter_ro_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 296.000 647.590 300.000 ;
    END
  END slave_data_req_to_inter_ro_o[2]
  PIN slave_data_req_to_inter_ro_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 296.000 667.370 300.000 ;
    END
  END slave_data_req_to_inter_ro_o[3]
  PIN slave_data_wdata_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 296.000 609.870 300.000 ;
    END
  END slave_data_wdata_to_inter_o[0]
  PIN slave_data_wdata_to_inter_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.470 296.000 1519.750 300.000 ;
    END
  END slave_data_wdata_to_inter_o[100]
  PIN slave_data_wdata_to_inter_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.910 296.000 1526.190 300.000 ;
    END
  END slave_data_wdata_to_inter_o[101]
  PIN slave_data_wdata_to_inter_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 296.000 1533.090 300.000 ;
    END
  END slave_data_wdata_to_inter_o[102]
  PIN slave_data_wdata_to_inter_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 296.000 1539.530 300.000 ;
    END
  END slave_data_wdata_to_inter_o[103]
  PIN slave_data_wdata_to_inter_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.150 296.000 1546.430 300.000 ;
    END
  END slave_data_wdata_to_inter_o[104]
  PIN slave_data_wdata_to_inter_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.590 296.000 1552.870 300.000 ;
    END
  END slave_data_wdata_to_inter_o[105]
  PIN slave_data_wdata_to_inter_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.490 296.000 1559.770 300.000 ;
    END
  END slave_data_wdata_to_inter_o[106]
  PIN slave_data_wdata_to_inter_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.930 296.000 1566.210 300.000 ;
    END
  END slave_data_wdata_to_inter_o[107]
  PIN slave_data_wdata_to_inter_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.370 296.000 1572.650 300.000 ;
    END
  END slave_data_wdata_to_inter_o[108]
  PIN slave_data_wdata_to_inter_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.270 296.000 1579.550 300.000 ;
    END
  END slave_data_wdata_to_inter_o[109]
  PIN slave_data_wdata_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 296.000 764.890 300.000 ;
    END
  END slave_data_wdata_to_inter_o[10]
  PIN slave_data_wdata_to_inter_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.710 296.000 1585.990 300.000 ;
    END
  END slave_data_wdata_to_inter_o[110]
  PIN slave_data_wdata_to_inter_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.610 296.000 1592.890 300.000 ;
    END
  END slave_data_wdata_to_inter_o[111]
  PIN slave_data_wdata_to_inter_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.050 296.000 1599.330 300.000 ;
    END
  END slave_data_wdata_to_inter_o[112]
  PIN slave_data_wdata_to_inter_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.950 296.000 1606.230 300.000 ;
    END
  END slave_data_wdata_to_inter_o[113]
  PIN slave_data_wdata_to_inter_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.390 296.000 1612.670 300.000 ;
    END
  END slave_data_wdata_to_inter_o[114]
  PIN slave_data_wdata_to_inter_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.830 296.000 1619.110 300.000 ;
    END
  END slave_data_wdata_to_inter_o[115]
  PIN slave_data_wdata_to_inter_o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 296.000 1626.010 300.000 ;
    END
  END slave_data_wdata_to_inter_o[116]
  PIN slave_data_wdata_to_inter_o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.170 296.000 1632.450 300.000 ;
    END
  END slave_data_wdata_to_inter_o[117]
  PIN slave_data_wdata_to_inter_o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 296.000 1639.350 300.000 ;
    END
  END slave_data_wdata_to_inter_o[118]
  PIN slave_data_wdata_to_inter_o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 296.000 1645.790 300.000 ;
    END
  END slave_data_wdata_to_inter_o[119]
  PIN slave_data_wdata_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 296.000 778.230 300.000 ;
    END
  END slave_data_wdata_to_inter_o[11]
  PIN slave_data_wdata_to_inter_o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.410 296.000 1652.690 300.000 ;
    END
  END slave_data_wdata_to_inter_o[120]
  PIN slave_data_wdata_to_inter_o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 296.000 1659.130 300.000 ;
    END
  END slave_data_wdata_to_inter_o[121]
  PIN slave_data_wdata_to_inter_o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.750 296.000 1666.030 300.000 ;
    END
  END slave_data_wdata_to_inter_o[122]
  PIN slave_data_wdata_to_inter_o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 296.000 1672.470 300.000 ;
    END
  END slave_data_wdata_to_inter_o[123]
  PIN slave_data_wdata_to_inter_o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.630 296.000 1678.910 300.000 ;
    END
  END slave_data_wdata_to_inter_o[124]
  PIN slave_data_wdata_to_inter_o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.530 296.000 1685.810 300.000 ;
    END
  END slave_data_wdata_to_inter_o[125]
  PIN slave_data_wdata_to_inter_o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 296.000 1692.250 300.000 ;
    END
  END slave_data_wdata_to_inter_o[126]
  PIN slave_data_wdata_to_inter_o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.870 296.000 1699.150 300.000 ;
    END
  END slave_data_wdata_to_inter_o[127]
  PIN slave_data_wdata_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 296.000 791.570 300.000 ;
    END
  END slave_data_wdata_to_inter_o[12]
  PIN slave_data_wdata_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 296.000 804.450 300.000 ;
    END
  END slave_data_wdata_to_inter_o[13]
  PIN slave_data_wdata_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 296.000 817.790 300.000 ;
    END
  END slave_data_wdata_to_inter_o[14]
  PIN slave_data_wdata_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 296.000 831.130 300.000 ;
    END
  END slave_data_wdata_to_inter_o[15]
  PIN slave_data_wdata_to_inter_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 296.000 842.170 300.000 ;
    END
  END slave_data_wdata_to_inter_o[16]
  PIN slave_data_wdata_to_inter_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 296.000 853.210 300.000 ;
    END
  END slave_data_wdata_to_inter_o[17]
  PIN slave_data_wdata_to_inter_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 296.000 864.250 300.000 ;
    END
  END slave_data_wdata_to_inter_o[18]
  PIN slave_data_wdata_to_inter_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 296.000 875.290 300.000 ;
    END
  END slave_data_wdata_to_inter_o[19]
  PIN slave_data_wdata_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 296.000 629.650 300.000 ;
    END
  END slave_data_wdata_to_inter_o[1]
  PIN slave_data_wdata_to_inter_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 296.000 886.790 300.000 ;
    END
  END slave_data_wdata_to_inter_o[20]
  PIN slave_data_wdata_to_inter_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 296.000 897.830 300.000 ;
    END
  END slave_data_wdata_to_inter_o[21]
  PIN slave_data_wdata_to_inter_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 296.000 908.870 300.000 ;
    END
  END slave_data_wdata_to_inter_o[22]
  PIN slave_data_wdata_to_inter_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.630 296.000 919.910 300.000 ;
    END
  END slave_data_wdata_to_inter_o[23]
  PIN slave_data_wdata_to_inter_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 296.000 930.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[24]
  PIN slave_data_wdata_to_inter_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.710 296.000 941.990 300.000 ;
    END
  END slave_data_wdata_to_inter_o[25]
  PIN slave_data_wdata_to_inter_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 296.000 953.030 300.000 ;
    END
  END slave_data_wdata_to_inter_o[26]
  PIN slave_data_wdata_to_inter_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 296.000 964.070 300.000 ;
    END
  END slave_data_wdata_to_inter_o[27]
  PIN slave_data_wdata_to_inter_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.830 296.000 975.110 300.000 ;
    END
  END slave_data_wdata_to_inter_o[28]
  PIN slave_data_wdata_to_inter_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.870 296.000 986.150 300.000 ;
    END
  END slave_data_wdata_to_inter_o[29]
  PIN slave_data_wdata_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 296.000 649.890 300.000 ;
    END
  END slave_data_wdata_to_inter_o[2]
  PIN slave_data_wdata_to_inter_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 296.000 997.190 300.000 ;
    END
  END slave_data_wdata_to_inter_o[30]
  PIN slave_data_wdata_to_inter_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 296.000 1008.230 300.000 ;
    END
  END slave_data_wdata_to_inter_o[31]
  PIN slave_data_wdata_to_inter_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 296.000 1019.270 300.000 ;
    END
  END slave_data_wdata_to_inter_o[32]
  PIN slave_data_wdata_to_inter_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.030 296.000 1030.310 300.000 ;
    END
  END slave_data_wdata_to_inter_o[33]
  PIN slave_data_wdata_to_inter_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.070 296.000 1041.350 300.000 ;
    END
  END slave_data_wdata_to_inter_o[34]
  PIN slave_data_wdata_to_inter_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.110 296.000 1052.390 300.000 ;
    END
  END slave_data_wdata_to_inter_o[35]
  PIN slave_data_wdata_to_inter_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.610 296.000 1063.890 300.000 ;
    END
  END slave_data_wdata_to_inter_o[36]
  PIN slave_data_wdata_to_inter_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.650 296.000 1074.930 300.000 ;
    END
  END slave_data_wdata_to_inter_o[37]
  PIN slave_data_wdata_to_inter_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.690 296.000 1085.970 300.000 ;
    END
  END slave_data_wdata_to_inter_o[38]
  PIN slave_data_wdata_to_inter_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.730 296.000 1097.010 300.000 ;
    END
  END slave_data_wdata_to_inter_o[39]
  PIN slave_data_wdata_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 296.000 669.670 300.000 ;
    END
  END slave_data_wdata_to_inter_o[3]
  PIN slave_data_wdata_to_inter_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 296.000 1108.050 300.000 ;
    END
  END slave_data_wdata_to_inter_o[40]
  PIN slave_data_wdata_to_inter_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.810 296.000 1119.090 300.000 ;
    END
  END slave_data_wdata_to_inter_o[41]
  PIN slave_data_wdata_to_inter_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.850 296.000 1130.130 300.000 ;
    END
  END slave_data_wdata_to_inter_o[42]
  PIN slave_data_wdata_to_inter_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.890 296.000 1141.170 300.000 ;
    END
  END slave_data_wdata_to_inter_o[43]
  PIN slave_data_wdata_to_inter_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.330 296.000 1147.610 300.000 ;
    END
  END slave_data_wdata_to_inter_o[44]
  PIN slave_data_wdata_to_inter_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.230 296.000 1154.510 300.000 ;
    END
  END slave_data_wdata_to_inter_o[45]
  PIN slave_data_wdata_to_inter_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.670 296.000 1160.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[46]
  PIN slave_data_wdata_to_inter_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.570 296.000 1167.850 300.000 ;
    END
  END slave_data_wdata_to_inter_o[47]
  PIN slave_data_wdata_to_inter_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.010 296.000 1174.290 300.000 ;
    END
  END slave_data_wdata_to_inter_o[48]
  PIN slave_data_wdata_to_inter_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.910 296.000 1181.190 300.000 ;
    END
  END slave_data_wdata_to_inter_o[49]
  PIN slave_data_wdata_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 296.000 685.310 300.000 ;
    END
  END slave_data_wdata_to_inter_o[4]
  PIN slave_data_wdata_to_inter_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.350 296.000 1187.630 300.000 ;
    END
  END slave_data_wdata_to_inter_o[50]
  PIN slave_data_wdata_to_inter_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.790 296.000 1194.070 300.000 ;
    END
  END slave_data_wdata_to_inter_o[51]
  PIN slave_data_wdata_to_inter_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.690 296.000 1200.970 300.000 ;
    END
  END slave_data_wdata_to_inter_o[52]
  PIN slave_data_wdata_to_inter_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.130 296.000 1207.410 300.000 ;
    END
  END slave_data_wdata_to_inter_o[53]
  PIN slave_data_wdata_to_inter_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 296.000 1214.310 300.000 ;
    END
  END slave_data_wdata_to_inter_o[54]
  PIN slave_data_wdata_to_inter_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 296.000 1220.750 300.000 ;
    END
  END slave_data_wdata_to_inter_o[55]
  PIN slave_data_wdata_to_inter_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 296.000 1227.650 300.000 ;
    END
  END slave_data_wdata_to_inter_o[56]
  PIN slave_data_wdata_to_inter_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 296.000 1234.090 300.000 ;
    END
  END slave_data_wdata_to_inter_o[57]
  PIN slave_data_wdata_to_inter_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.710 296.000 1240.990 300.000 ;
    END
  END slave_data_wdata_to_inter_o[58]
  PIN slave_data_wdata_to_inter_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.150 296.000 1247.430 300.000 ;
    END
  END slave_data_wdata_to_inter_o[59]
  PIN slave_data_wdata_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 296.000 698.190 300.000 ;
    END
  END slave_data_wdata_to_inter_o[5]
  PIN slave_data_wdata_to_inter_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.590 296.000 1253.870 300.000 ;
    END
  END slave_data_wdata_to_inter_o[60]
  PIN slave_data_wdata_to_inter_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.490 296.000 1260.770 300.000 ;
    END
  END slave_data_wdata_to_inter_o[61]
  PIN slave_data_wdata_to_inter_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 296.000 1267.210 300.000 ;
    END
  END slave_data_wdata_to_inter_o[62]
  PIN slave_data_wdata_to_inter_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 296.000 1274.110 300.000 ;
    END
  END slave_data_wdata_to_inter_o[63]
  PIN slave_data_wdata_to_inter_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 296.000 1280.550 300.000 ;
    END
  END slave_data_wdata_to_inter_o[64]
  PIN slave_data_wdata_to_inter_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.170 296.000 1287.450 300.000 ;
    END
  END slave_data_wdata_to_inter_o[65]
  PIN slave_data_wdata_to_inter_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.610 296.000 1293.890 300.000 ;
    END
  END slave_data_wdata_to_inter_o[66]
  PIN slave_data_wdata_to_inter_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.050 296.000 1300.330 300.000 ;
    END
  END slave_data_wdata_to_inter_o[67]
  PIN slave_data_wdata_to_inter_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.950 296.000 1307.230 300.000 ;
    END
  END slave_data_wdata_to_inter_o[68]
  PIN slave_data_wdata_to_inter_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.390 296.000 1313.670 300.000 ;
    END
  END slave_data_wdata_to_inter_o[69]
  PIN slave_data_wdata_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 296.000 711.530 300.000 ;
    END
  END slave_data_wdata_to_inter_o[6]
  PIN slave_data_wdata_to_inter_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.290 296.000 1320.570 300.000 ;
    END
  END slave_data_wdata_to_inter_o[70]
  PIN slave_data_wdata_to_inter_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 296.000 1327.010 300.000 ;
    END
  END slave_data_wdata_to_inter_o[71]
  PIN slave_data_wdata_to_inter_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 296.000 1333.910 300.000 ;
    END
  END slave_data_wdata_to_inter_o[72]
  PIN slave_data_wdata_to_inter_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.070 296.000 1340.350 300.000 ;
    END
  END slave_data_wdata_to_inter_o[73]
  PIN slave_data_wdata_to_inter_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.970 296.000 1347.250 300.000 ;
    END
  END slave_data_wdata_to_inter_o[74]
  PIN slave_data_wdata_to_inter_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.410 296.000 1353.690 300.000 ;
    END
  END slave_data_wdata_to_inter_o[75]
  PIN slave_data_wdata_to_inter_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.850 296.000 1360.130 300.000 ;
    END
  END slave_data_wdata_to_inter_o[76]
  PIN slave_data_wdata_to_inter_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.750 296.000 1367.030 300.000 ;
    END
  END slave_data_wdata_to_inter_o[77]
  PIN slave_data_wdata_to_inter_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.190 296.000 1373.470 300.000 ;
    END
  END slave_data_wdata_to_inter_o[78]
  PIN slave_data_wdata_to_inter_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 296.000 1380.370 300.000 ;
    END
  END slave_data_wdata_to_inter_o[79]
  PIN slave_data_wdata_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 296.000 724.870 300.000 ;
    END
  END slave_data_wdata_to_inter_o[7]
  PIN slave_data_wdata_to_inter_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.530 296.000 1386.810 300.000 ;
    END
  END slave_data_wdata_to_inter_o[80]
  PIN slave_data_wdata_to_inter_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.430 296.000 1393.710 300.000 ;
    END
  END slave_data_wdata_to_inter_o[81]
  PIN slave_data_wdata_to_inter_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.870 296.000 1400.150 300.000 ;
    END
  END slave_data_wdata_to_inter_o[82]
  PIN slave_data_wdata_to_inter_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.310 296.000 1406.590 300.000 ;
    END
  END slave_data_wdata_to_inter_o[83]
  PIN slave_data_wdata_to_inter_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.210 296.000 1413.490 300.000 ;
    END
  END slave_data_wdata_to_inter_o[84]
  PIN slave_data_wdata_to_inter_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.650 296.000 1419.930 300.000 ;
    END
  END slave_data_wdata_to_inter_o[85]
  PIN slave_data_wdata_to_inter_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 296.000 1426.830 300.000 ;
    END
  END slave_data_wdata_to_inter_o[86]
  PIN slave_data_wdata_to_inter_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 296.000 1433.270 300.000 ;
    END
  END slave_data_wdata_to_inter_o[87]
  PIN slave_data_wdata_to_inter_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 296.000 1440.170 300.000 ;
    END
  END slave_data_wdata_to_inter_o[88]
  PIN slave_data_wdata_to_inter_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 296.000 1446.610 300.000 ;
    END
  END slave_data_wdata_to_inter_o[89]
  PIN slave_data_wdata_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 296.000 738.210 300.000 ;
    END
  END slave_data_wdata_to_inter_o[8]
  PIN slave_data_wdata_to_inter_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.230 296.000 1453.510 300.000 ;
    END
  END slave_data_wdata_to_inter_o[90]
  PIN slave_data_wdata_to_inter_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.670 296.000 1459.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[91]
  PIN slave_data_wdata_to_inter_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.110 296.000 1466.390 300.000 ;
    END
  END slave_data_wdata_to_inter_o[92]
  PIN slave_data_wdata_to_inter_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.010 296.000 1473.290 300.000 ;
    END
  END slave_data_wdata_to_inter_o[93]
  PIN slave_data_wdata_to_inter_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.450 296.000 1479.730 300.000 ;
    END
  END slave_data_wdata_to_inter_o[94]
  PIN slave_data_wdata_to_inter_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.350 296.000 1486.630 300.000 ;
    END
  END slave_data_wdata_to_inter_o[95]
  PIN slave_data_wdata_to_inter_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 296.000 1493.070 300.000 ;
    END
  END slave_data_wdata_to_inter_o[96]
  PIN slave_data_wdata_to_inter_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 296.000 1499.970 300.000 ;
    END
  END slave_data_wdata_to_inter_o[97]
  PIN slave_data_wdata_to_inter_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.130 296.000 1506.410 300.000 ;
    END
  END slave_data_wdata_to_inter_o[98]
  PIN slave_data_wdata_to_inter_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.570 296.000 1512.850 300.000 ;
    END
  END slave_data_wdata_to_inter_o[99]
  PIN slave_data_wdata_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 296.000 751.550 300.000 ;
    END
  END slave_data_wdata_to_inter_o[9]
  PIN slave_data_we_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 296.000 612.170 300.000 ;
    END
  END slave_data_we_to_inter_o[0]
  PIN slave_data_we_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 296.000 631.950 300.000 ;
    END
  END slave_data_we_to_inter_o[1]
  PIN slave_data_we_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 296.000 651.730 300.000 ;
    END
  END slave_data_we_to_inter_o[2]
  PIN slave_data_we_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 296.000 671.970 300.000 ;
    END
  END slave_data_we_to_inter_o[3]
  PIN txd_uart
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 149.640 1700.000 150.240 ;
    END
  END txd_uart
  PIN txd_uart_to_mem
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 209.480 1700.000 210.080 ;
    END
  END txd_uart_to_mem
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.870 0.000 1676.150 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 0.000 1692.250 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 0.000 858.270 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.830 0.000 906.110 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 0.000 954.410 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 0.000 1002.250 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 0.000 1050.550 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 0.000 1194.990 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 0.000 1242.830 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.850 0.000 1291.130 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.150 0.000 1339.430 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.990 0.000 1387.270 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 0.000 1435.570 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.130 0.000 1483.410 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.430 0.000 1531.710 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.730 0.000 1580.010 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.570 0.000 1627.850 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 0.000 681.630 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 0.000 826.070 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 0.000 873.910 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 0.000 922.210 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 0.000 970.510 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.070 0.000 1018.350 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 0.000 1066.650 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.650 0.000 1258.930 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.950 0.000 1307.230 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.790 0.000 1355.070 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.090 0.000 1403.370 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.390 0.000 1451.670 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.230 0.000 1499.510 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.530 0.000 1547.810 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.370 0.000 1595.650 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.670 0.000 1643.950 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 0.000 890.010 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 0.000 938.310 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.870 0.000 986.150 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 0.000 1034.450 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.470 0.000 1082.750 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.450 0.000 1226.730 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.750 0.000 1275.030 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 0.000 1323.330 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.890 0.000 1371.170 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.190 0.000 1419.470 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.030 0.000 1467.310 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.330 0.000 1515.610 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.630 0.000 1563.910 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.470 0.000 1611.750 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1659.770 0.000 1660.050 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1694.180 288.405 ;
      LAYER met1 ;
        RECT 0.990 10.240 1699.170 299.840 ;
      LAYER met2 ;
        RECT 1.570 295.720 2.570 299.870 ;
        RECT 3.410 295.720 4.870 299.870 ;
        RECT 5.710 295.720 7.170 299.870 ;
        RECT 8.010 295.720 9.470 299.870 ;
        RECT 10.310 295.720 11.770 299.870 ;
        RECT 12.610 295.720 13.610 299.870 ;
        RECT 14.450 295.720 15.910 299.870 ;
        RECT 16.750 295.720 18.210 299.870 ;
        RECT 19.050 295.720 20.510 299.870 ;
        RECT 21.350 295.720 22.810 299.870 ;
        RECT 23.650 295.720 24.650 299.870 ;
        RECT 25.490 295.720 26.950 299.870 ;
        RECT 27.790 295.720 29.250 299.870 ;
        RECT 30.090 295.720 31.550 299.870 ;
        RECT 32.390 295.720 33.850 299.870 ;
        RECT 34.690 295.720 36.150 299.870 ;
        RECT 36.990 295.720 37.990 299.870 ;
        RECT 38.830 295.720 40.290 299.870 ;
        RECT 41.130 295.720 42.590 299.870 ;
        RECT 43.430 295.720 44.890 299.870 ;
        RECT 45.730 295.720 47.190 299.870 ;
        RECT 48.030 295.720 49.030 299.870 ;
        RECT 49.870 295.720 51.330 299.870 ;
        RECT 52.170 295.720 53.630 299.870 ;
        RECT 54.470 295.720 55.930 299.870 ;
        RECT 56.770 295.720 58.230 299.870 ;
        RECT 59.070 295.720 60.070 299.870 ;
        RECT 60.910 295.720 62.370 299.870 ;
        RECT 63.210 295.720 64.670 299.870 ;
        RECT 65.510 295.720 66.970 299.870 ;
        RECT 67.810 295.720 69.270 299.870 ;
        RECT 70.110 295.720 71.570 299.870 ;
        RECT 72.410 295.720 73.410 299.870 ;
        RECT 74.250 295.720 75.710 299.870 ;
        RECT 76.550 295.720 78.010 299.870 ;
        RECT 78.850 295.720 80.310 299.870 ;
        RECT 81.150 295.720 82.610 299.870 ;
        RECT 83.450 295.720 84.450 299.870 ;
        RECT 85.290 295.720 86.750 299.870 ;
        RECT 87.590 295.720 89.050 299.870 ;
        RECT 89.890 295.720 91.350 299.870 ;
        RECT 92.190 295.720 93.650 299.870 ;
        RECT 94.490 295.720 95.490 299.870 ;
        RECT 96.330 295.720 97.790 299.870 ;
        RECT 98.630 295.720 100.090 299.870 ;
        RECT 100.930 295.720 102.390 299.870 ;
        RECT 103.230 295.720 104.690 299.870 ;
        RECT 105.530 295.720 106.990 299.870 ;
        RECT 107.830 295.720 108.830 299.870 ;
        RECT 109.670 295.720 111.130 299.870 ;
        RECT 111.970 295.720 113.430 299.870 ;
        RECT 114.270 295.720 115.730 299.870 ;
        RECT 116.570 295.720 118.030 299.870 ;
        RECT 118.870 295.720 119.870 299.870 ;
        RECT 120.710 295.720 122.170 299.870 ;
        RECT 123.010 295.720 124.470 299.870 ;
        RECT 125.310 295.720 126.770 299.870 ;
        RECT 127.610 295.720 129.070 299.870 ;
        RECT 129.910 295.720 130.910 299.870 ;
        RECT 131.750 295.720 133.210 299.870 ;
        RECT 134.050 295.720 135.510 299.870 ;
        RECT 136.350 295.720 137.810 299.870 ;
        RECT 138.650 295.720 140.110 299.870 ;
        RECT 140.950 295.720 142.410 299.870 ;
        RECT 143.250 295.720 144.250 299.870 ;
        RECT 145.090 295.720 146.550 299.870 ;
        RECT 147.390 295.720 148.850 299.870 ;
        RECT 149.690 295.720 151.150 299.870 ;
        RECT 151.990 295.720 153.450 299.870 ;
        RECT 154.290 295.720 155.290 299.870 ;
        RECT 156.130 295.720 157.590 299.870 ;
        RECT 158.430 295.720 159.890 299.870 ;
        RECT 160.730 295.720 162.190 299.870 ;
        RECT 163.030 295.720 164.490 299.870 ;
        RECT 165.330 295.720 166.330 299.870 ;
        RECT 167.170 295.720 168.630 299.870 ;
        RECT 169.470 295.720 170.930 299.870 ;
        RECT 171.770 295.720 173.230 299.870 ;
        RECT 174.070 295.720 175.530 299.870 ;
        RECT 176.370 295.720 177.830 299.870 ;
        RECT 178.670 295.720 179.670 299.870 ;
        RECT 180.510 295.720 181.970 299.870 ;
        RECT 182.810 295.720 184.270 299.870 ;
        RECT 185.110 295.720 186.570 299.870 ;
        RECT 187.410 295.720 188.870 299.870 ;
        RECT 189.710 295.720 190.710 299.870 ;
        RECT 191.550 295.720 193.010 299.870 ;
        RECT 193.850 295.720 195.310 299.870 ;
        RECT 196.150 295.720 197.610 299.870 ;
        RECT 198.450 295.720 199.910 299.870 ;
        RECT 200.750 295.720 201.750 299.870 ;
        RECT 202.590 295.720 204.050 299.870 ;
        RECT 204.890 295.720 206.350 299.870 ;
        RECT 207.190 295.720 208.650 299.870 ;
        RECT 209.490 295.720 210.950 299.870 ;
        RECT 211.790 295.720 213.250 299.870 ;
        RECT 214.090 295.720 215.090 299.870 ;
        RECT 215.930 295.720 217.390 299.870 ;
        RECT 218.230 295.720 219.690 299.870 ;
        RECT 220.530 295.720 221.990 299.870 ;
        RECT 222.830 295.720 224.290 299.870 ;
        RECT 225.130 295.720 226.130 299.870 ;
        RECT 226.970 295.720 228.430 299.870 ;
        RECT 229.270 295.720 230.730 299.870 ;
        RECT 231.570 295.720 233.030 299.870 ;
        RECT 233.870 295.720 235.330 299.870 ;
        RECT 236.170 295.720 237.170 299.870 ;
        RECT 238.010 295.720 239.470 299.870 ;
        RECT 240.310 295.720 241.770 299.870 ;
        RECT 242.610 295.720 244.070 299.870 ;
        RECT 244.910 295.720 246.370 299.870 ;
        RECT 247.210 295.720 248.670 299.870 ;
        RECT 249.510 295.720 250.510 299.870 ;
        RECT 251.350 295.720 252.810 299.870 ;
        RECT 253.650 295.720 255.110 299.870 ;
        RECT 255.950 295.720 257.410 299.870 ;
        RECT 258.250 295.720 259.710 299.870 ;
        RECT 260.550 295.720 261.550 299.870 ;
        RECT 262.390 295.720 263.850 299.870 ;
        RECT 264.690 295.720 266.150 299.870 ;
        RECT 266.990 295.720 268.450 299.870 ;
        RECT 269.290 295.720 270.750 299.870 ;
        RECT 271.590 295.720 272.590 299.870 ;
        RECT 273.430 295.720 274.890 299.870 ;
        RECT 275.730 295.720 277.190 299.870 ;
        RECT 278.030 295.720 279.490 299.870 ;
        RECT 280.330 295.720 281.790 299.870 ;
        RECT 282.630 295.720 284.090 299.870 ;
        RECT 284.930 295.720 285.930 299.870 ;
        RECT 286.770 295.720 288.230 299.870 ;
        RECT 289.070 295.720 290.530 299.870 ;
        RECT 291.370 295.720 292.830 299.870 ;
        RECT 293.670 295.720 295.130 299.870 ;
        RECT 295.970 295.720 296.970 299.870 ;
        RECT 297.810 295.720 299.270 299.870 ;
        RECT 300.110 295.720 301.570 299.870 ;
        RECT 302.410 295.720 303.870 299.870 ;
        RECT 304.710 295.720 306.170 299.870 ;
        RECT 307.010 295.720 308.010 299.870 ;
        RECT 308.850 295.720 310.310 299.870 ;
        RECT 311.150 295.720 312.610 299.870 ;
        RECT 313.450 295.720 314.910 299.870 ;
        RECT 315.750 295.720 317.210 299.870 ;
        RECT 318.050 295.720 319.510 299.870 ;
        RECT 320.350 295.720 321.350 299.870 ;
        RECT 322.190 295.720 323.650 299.870 ;
        RECT 324.490 295.720 325.950 299.870 ;
        RECT 326.790 295.720 328.250 299.870 ;
        RECT 329.090 295.720 330.550 299.870 ;
        RECT 331.390 295.720 332.390 299.870 ;
        RECT 333.230 295.720 334.690 299.870 ;
        RECT 335.530 295.720 336.990 299.870 ;
        RECT 337.830 295.720 339.290 299.870 ;
        RECT 340.130 295.720 341.590 299.870 ;
        RECT 342.430 295.720 343.430 299.870 ;
        RECT 344.270 295.720 345.730 299.870 ;
        RECT 346.570 295.720 348.030 299.870 ;
        RECT 348.870 295.720 350.330 299.870 ;
        RECT 351.170 295.720 352.630 299.870 ;
        RECT 353.470 295.720 354.930 299.870 ;
        RECT 355.770 295.720 356.770 299.870 ;
        RECT 357.610 295.720 359.070 299.870 ;
        RECT 359.910 295.720 361.370 299.870 ;
        RECT 362.210 295.720 363.670 299.870 ;
        RECT 364.510 295.720 365.970 299.870 ;
        RECT 366.810 295.720 367.810 299.870 ;
        RECT 368.650 295.720 370.110 299.870 ;
        RECT 370.950 295.720 372.410 299.870 ;
        RECT 373.250 295.720 374.710 299.870 ;
        RECT 375.550 295.720 377.010 299.870 ;
        RECT 377.850 295.720 378.850 299.870 ;
        RECT 379.690 295.720 381.150 299.870 ;
        RECT 381.990 295.720 383.450 299.870 ;
        RECT 384.290 295.720 385.750 299.870 ;
        RECT 386.590 295.720 388.050 299.870 ;
        RECT 388.890 295.720 390.350 299.870 ;
        RECT 391.190 295.720 392.190 299.870 ;
        RECT 393.030 295.720 394.490 299.870 ;
        RECT 395.330 295.720 396.790 299.870 ;
        RECT 397.630 295.720 399.090 299.870 ;
        RECT 399.930 295.720 401.390 299.870 ;
        RECT 402.230 295.720 403.230 299.870 ;
        RECT 404.070 295.720 405.530 299.870 ;
        RECT 406.370 295.720 407.830 299.870 ;
        RECT 408.670 295.720 410.130 299.870 ;
        RECT 410.970 295.720 412.430 299.870 ;
        RECT 413.270 295.720 414.270 299.870 ;
        RECT 415.110 295.720 416.570 299.870 ;
        RECT 417.410 295.720 418.870 299.870 ;
        RECT 419.710 295.720 421.170 299.870 ;
        RECT 422.010 295.720 423.470 299.870 ;
        RECT 424.310 295.720 425.770 299.870 ;
        RECT 426.610 295.720 427.610 299.870 ;
        RECT 428.450 295.720 429.910 299.870 ;
        RECT 430.750 295.720 432.210 299.870 ;
        RECT 433.050 295.720 434.510 299.870 ;
        RECT 435.350 295.720 436.810 299.870 ;
        RECT 437.650 295.720 438.650 299.870 ;
        RECT 439.490 295.720 440.950 299.870 ;
        RECT 441.790 295.720 443.250 299.870 ;
        RECT 444.090 295.720 445.550 299.870 ;
        RECT 446.390 295.720 447.850 299.870 ;
        RECT 448.690 295.720 449.690 299.870 ;
        RECT 450.530 295.720 451.990 299.870 ;
        RECT 452.830 295.720 454.290 299.870 ;
        RECT 455.130 295.720 456.590 299.870 ;
        RECT 457.430 295.720 458.890 299.870 ;
        RECT 459.730 295.720 461.190 299.870 ;
        RECT 462.030 295.720 463.030 299.870 ;
        RECT 463.870 295.720 465.330 299.870 ;
        RECT 466.170 295.720 467.630 299.870 ;
        RECT 468.470 295.720 469.930 299.870 ;
        RECT 470.770 295.720 472.230 299.870 ;
        RECT 473.070 295.720 474.070 299.870 ;
        RECT 474.910 295.720 476.370 299.870 ;
        RECT 477.210 295.720 478.670 299.870 ;
        RECT 479.510 295.720 480.970 299.870 ;
        RECT 481.810 295.720 483.270 299.870 ;
        RECT 484.110 295.720 485.110 299.870 ;
        RECT 485.950 295.720 487.410 299.870 ;
        RECT 488.250 295.720 489.710 299.870 ;
        RECT 490.550 295.720 492.010 299.870 ;
        RECT 492.850 295.720 494.310 299.870 ;
        RECT 495.150 295.720 496.610 299.870 ;
        RECT 497.450 295.720 498.450 299.870 ;
        RECT 499.290 295.720 500.750 299.870 ;
        RECT 501.590 295.720 503.050 299.870 ;
        RECT 503.890 295.720 505.350 299.870 ;
        RECT 506.190 295.720 507.650 299.870 ;
        RECT 508.490 295.720 509.490 299.870 ;
        RECT 510.330 295.720 511.790 299.870 ;
        RECT 512.630 295.720 514.090 299.870 ;
        RECT 514.930 295.720 516.390 299.870 ;
        RECT 517.230 295.720 518.690 299.870 ;
        RECT 519.530 295.720 520.530 299.870 ;
        RECT 521.370 295.720 522.830 299.870 ;
        RECT 523.670 295.720 525.130 299.870 ;
        RECT 525.970 295.720 527.430 299.870 ;
        RECT 528.270 295.720 529.730 299.870 ;
        RECT 530.570 295.720 532.030 299.870 ;
        RECT 532.870 295.720 533.870 299.870 ;
        RECT 534.710 295.720 536.170 299.870 ;
        RECT 537.010 295.720 538.470 299.870 ;
        RECT 539.310 295.720 540.770 299.870 ;
        RECT 541.610 295.720 543.070 299.870 ;
        RECT 543.910 295.720 544.910 299.870 ;
        RECT 545.750 295.720 547.210 299.870 ;
        RECT 548.050 295.720 549.510 299.870 ;
        RECT 550.350 295.720 551.810 299.870 ;
        RECT 552.650 295.720 554.110 299.870 ;
        RECT 554.950 295.720 555.950 299.870 ;
        RECT 556.790 295.720 558.250 299.870 ;
        RECT 559.090 295.720 560.550 299.870 ;
        RECT 561.390 295.720 562.850 299.870 ;
        RECT 563.690 295.720 565.150 299.870 ;
        RECT 565.990 295.720 567.450 299.870 ;
        RECT 568.290 295.720 569.290 299.870 ;
        RECT 570.130 295.720 571.590 299.870 ;
        RECT 572.430 295.720 573.890 299.870 ;
        RECT 574.730 295.720 576.190 299.870 ;
        RECT 577.030 295.720 578.490 299.870 ;
        RECT 579.330 295.720 580.330 299.870 ;
        RECT 581.170 295.720 582.630 299.870 ;
        RECT 583.470 295.720 584.930 299.870 ;
        RECT 585.770 295.720 587.230 299.870 ;
        RECT 588.070 295.720 589.530 299.870 ;
        RECT 590.370 295.720 591.370 299.870 ;
        RECT 592.210 295.720 593.670 299.870 ;
        RECT 594.510 295.720 595.970 299.870 ;
        RECT 596.810 295.720 598.270 299.870 ;
        RECT 599.110 295.720 600.570 299.870 ;
        RECT 601.410 295.720 602.870 299.870 ;
        RECT 603.710 295.720 604.710 299.870 ;
        RECT 605.550 295.720 607.010 299.870 ;
        RECT 607.850 295.720 609.310 299.870 ;
        RECT 610.150 295.720 611.610 299.870 ;
        RECT 612.450 295.720 613.910 299.870 ;
        RECT 614.750 295.720 615.750 299.870 ;
        RECT 616.590 295.720 618.050 299.870 ;
        RECT 618.890 295.720 620.350 299.870 ;
        RECT 621.190 295.720 622.650 299.870 ;
        RECT 623.490 295.720 624.950 299.870 ;
        RECT 625.790 295.720 626.790 299.870 ;
        RECT 627.630 295.720 629.090 299.870 ;
        RECT 629.930 295.720 631.390 299.870 ;
        RECT 632.230 295.720 633.690 299.870 ;
        RECT 634.530 295.720 635.990 299.870 ;
        RECT 636.830 295.720 638.290 299.870 ;
        RECT 639.130 295.720 640.130 299.870 ;
        RECT 640.970 295.720 642.430 299.870 ;
        RECT 643.270 295.720 644.730 299.870 ;
        RECT 645.570 295.720 647.030 299.870 ;
        RECT 647.870 295.720 649.330 299.870 ;
        RECT 650.170 295.720 651.170 299.870 ;
        RECT 652.010 295.720 653.470 299.870 ;
        RECT 654.310 295.720 655.770 299.870 ;
        RECT 656.610 295.720 658.070 299.870 ;
        RECT 658.910 295.720 660.370 299.870 ;
        RECT 661.210 295.720 662.210 299.870 ;
        RECT 663.050 295.720 664.510 299.870 ;
        RECT 665.350 295.720 666.810 299.870 ;
        RECT 667.650 295.720 669.110 299.870 ;
        RECT 669.950 295.720 671.410 299.870 ;
        RECT 672.250 295.720 673.710 299.870 ;
        RECT 674.550 295.720 675.550 299.870 ;
        RECT 676.390 295.720 677.850 299.870 ;
        RECT 678.690 295.720 680.150 299.870 ;
        RECT 680.990 295.720 682.450 299.870 ;
        RECT 683.290 295.720 684.750 299.870 ;
        RECT 685.590 295.720 686.590 299.870 ;
        RECT 687.430 295.720 688.890 299.870 ;
        RECT 689.730 295.720 691.190 299.870 ;
        RECT 692.030 295.720 693.490 299.870 ;
        RECT 694.330 295.720 695.790 299.870 ;
        RECT 696.630 295.720 697.630 299.870 ;
        RECT 698.470 295.720 699.930 299.870 ;
        RECT 700.770 295.720 702.230 299.870 ;
        RECT 703.070 295.720 704.530 299.870 ;
        RECT 705.370 295.720 706.830 299.870 ;
        RECT 707.670 295.720 709.130 299.870 ;
        RECT 709.970 295.720 710.970 299.870 ;
        RECT 711.810 295.720 713.270 299.870 ;
        RECT 714.110 295.720 715.570 299.870 ;
        RECT 716.410 295.720 717.870 299.870 ;
        RECT 718.710 295.720 720.170 299.870 ;
        RECT 721.010 295.720 722.010 299.870 ;
        RECT 722.850 295.720 724.310 299.870 ;
        RECT 725.150 295.720 726.610 299.870 ;
        RECT 727.450 295.720 728.910 299.870 ;
        RECT 729.750 295.720 731.210 299.870 ;
        RECT 732.050 295.720 733.050 299.870 ;
        RECT 733.890 295.720 735.350 299.870 ;
        RECT 736.190 295.720 737.650 299.870 ;
        RECT 738.490 295.720 739.950 299.870 ;
        RECT 740.790 295.720 742.250 299.870 ;
        RECT 743.090 295.720 744.550 299.870 ;
        RECT 745.390 295.720 746.390 299.870 ;
        RECT 747.230 295.720 748.690 299.870 ;
        RECT 749.530 295.720 750.990 299.870 ;
        RECT 751.830 295.720 753.290 299.870 ;
        RECT 754.130 295.720 755.590 299.870 ;
        RECT 756.430 295.720 757.430 299.870 ;
        RECT 758.270 295.720 759.730 299.870 ;
        RECT 760.570 295.720 762.030 299.870 ;
        RECT 762.870 295.720 764.330 299.870 ;
        RECT 765.170 295.720 766.630 299.870 ;
        RECT 767.470 295.720 768.470 299.870 ;
        RECT 769.310 295.720 770.770 299.870 ;
        RECT 771.610 295.720 773.070 299.870 ;
        RECT 773.910 295.720 775.370 299.870 ;
        RECT 776.210 295.720 777.670 299.870 ;
        RECT 778.510 295.720 779.970 299.870 ;
        RECT 780.810 295.720 781.810 299.870 ;
        RECT 782.650 295.720 784.110 299.870 ;
        RECT 784.950 295.720 786.410 299.870 ;
        RECT 787.250 295.720 788.710 299.870 ;
        RECT 789.550 295.720 791.010 299.870 ;
        RECT 791.850 295.720 792.850 299.870 ;
        RECT 793.690 295.720 795.150 299.870 ;
        RECT 795.990 295.720 797.450 299.870 ;
        RECT 798.290 295.720 799.750 299.870 ;
        RECT 800.590 295.720 802.050 299.870 ;
        RECT 802.890 295.720 803.890 299.870 ;
        RECT 804.730 295.720 806.190 299.870 ;
        RECT 807.030 295.720 808.490 299.870 ;
        RECT 809.330 295.720 810.790 299.870 ;
        RECT 811.630 295.720 813.090 299.870 ;
        RECT 813.930 295.720 815.390 299.870 ;
        RECT 816.230 295.720 817.230 299.870 ;
        RECT 818.070 295.720 819.530 299.870 ;
        RECT 820.370 295.720 821.830 299.870 ;
        RECT 822.670 295.720 824.130 299.870 ;
        RECT 824.970 295.720 826.430 299.870 ;
        RECT 827.270 295.720 828.270 299.870 ;
        RECT 829.110 295.720 830.570 299.870 ;
        RECT 831.410 295.720 832.870 299.870 ;
        RECT 833.710 295.720 835.170 299.870 ;
        RECT 836.010 295.720 837.470 299.870 ;
        RECT 838.310 295.720 839.310 299.870 ;
        RECT 840.150 295.720 841.610 299.870 ;
        RECT 842.450 295.720 843.910 299.870 ;
        RECT 844.750 295.720 846.210 299.870 ;
        RECT 847.050 295.720 848.510 299.870 ;
        RECT 849.350 295.720 850.810 299.870 ;
        RECT 851.650 295.720 852.650 299.870 ;
        RECT 853.490 295.720 854.950 299.870 ;
        RECT 855.790 295.720 857.250 299.870 ;
        RECT 858.090 295.720 859.550 299.870 ;
        RECT 860.390 295.720 861.850 299.870 ;
        RECT 862.690 295.720 863.690 299.870 ;
        RECT 864.530 295.720 865.990 299.870 ;
        RECT 866.830 295.720 868.290 299.870 ;
        RECT 869.130 295.720 870.590 299.870 ;
        RECT 871.430 295.720 872.890 299.870 ;
        RECT 873.730 295.720 874.730 299.870 ;
        RECT 875.570 295.720 877.030 299.870 ;
        RECT 877.870 295.720 879.330 299.870 ;
        RECT 880.170 295.720 881.630 299.870 ;
        RECT 882.470 295.720 883.930 299.870 ;
        RECT 884.770 295.720 886.230 299.870 ;
        RECT 887.070 295.720 888.070 299.870 ;
        RECT 888.910 295.720 890.370 299.870 ;
        RECT 891.210 295.720 892.670 299.870 ;
        RECT 893.510 295.720 894.970 299.870 ;
        RECT 895.810 295.720 897.270 299.870 ;
        RECT 898.110 295.720 899.110 299.870 ;
        RECT 899.950 295.720 901.410 299.870 ;
        RECT 902.250 295.720 903.710 299.870 ;
        RECT 904.550 295.720 906.010 299.870 ;
        RECT 906.850 295.720 908.310 299.870 ;
        RECT 909.150 295.720 910.150 299.870 ;
        RECT 910.990 295.720 912.450 299.870 ;
        RECT 913.290 295.720 914.750 299.870 ;
        RECT 915.590 295.720 917.050 299.870 ;
        RECT 917.890 295.720 919.350 299.870 ;
        RECT 920.190 295.720 921.650 299.870 ;
        RECT 922.490 295.720 923.490 299.870 ;
        RECT 924.330 295.720 925.790 299.870 ;
        RECT 926.630 295.720 928.090 299.870 ;
        RECT 928.930 295.720 930.390 299.870 ;
        RECT 931.230 295.720 932.690 299.870 ;
        RECT 933.530 295.720 934.530 299.870 ;
        RECT 935.370 295.720 936.830 299.870 ;
        RECT 937.670 295.720 939.130 299.870 ;
        RECT 939.970 295.720 941.430 299.870 ;
        RECT 942.270 295.720 943.730 299.870 ;
        RECT 944.570 295.720 945.570 299.870 ;
        RECT 946.410 295.720 947.870 299.870 ;
        RECT 948.710 295.720 950.170 299.870 ;
        RECT 951.010 295.720 952.470 299.870 ;
        RECT 953.310 295.720 954.770 299.870 ;
        RECT 955.610 295.720 957.070 299.870 ;
        RECT 957.910 295.720 958.910 299.870 ;
        RECT 959.750 295.720 961.210 299.870 ;
        RECT 962.050 295.720 963.510 299.870 ;
        RECT 964.350 295.720 965.810 299.870 ;
        RECT 966.650 295.720 968.110 299.870 ;
        RECT 968.950 295.720 969.950 299.870 ;
        RECT 970.790 295.720 972.250 299.870 ;
        RECT 973.090 295.720 974.550 299.870 ;
        RECT 975.390 295.720 976.850 299.870 ;
        RECT 977.690 295.720 979.150 299.870 ;
        RECT 979.990 295.720 980.990 299.870 ;
        RECT 981.830 295.720 983.290 299.870 ;
        RECT 984.130 295.720 985.590 299.870 ;
        RECT 986.430 295.720 987.890 299.870 ;
        RECT 988.730 295.720 990.190 299.870 ;
        RECT 991.030 295.720 992.490 299.870 ;
        RECT 993.330 295.720 994.330 299.870 ;
        RECT 995.170 295.720 996.630 299.870 ;
        RECT 997.470 295.720 998.930 299.870 ;
        RECT 999.770 295.720 1001.230 299.870 ;
        RECT 1002.070 295.720 1003.530 299.870 ;
        RECT 1004.370 295.720 1005.370 299.870 ;
        RECT 1006.210 295.720 1007.670 299.870 ;
        RECT 1008.510 295.720 1009.970 299.870 ;
        RECT 1010.810 295.720 1012.270 299.870 ;
        RECT 1013.110 295.720 1014.570 299.870 ;
        RECT 1015.410 295.720 1016.410 299.870 ;
        RECT 1017.250 295.720 1018.710 299.870 ;
        RECT 1019.550 295.720 1021.010 299.870 ;
        RECT 1021.850 295.720 1023.310 299.870 ;
        RECT 1024.150 295.720 1025.610 299.870 ;
        RECT 1026.450 295.720 1027.910 299.870 ;
        RECT 1028.750 295.720 1029.750 299.870 ;
        RECT 1030.590 295.720 1032.050 299.870 ;
        RECT 1032.890 295.720 1034.350 299.870 ;
        RECT 1035.190 295.720 1036.650 299.870 ;
        RECT 1037.490 295.720 1038.950 299.870 ;
        RECT 1039.790 295.720 1040.790 299.870 ;
        RECT 1041.630 295.720 1043.090 299.870 ;
        RECT 1043.930 295.720 1045.390 299.870 ;
        RECT 1046.230 295.720 1047.690 299.870 ;
        RECT 1048.530 295.720 1049.990 299.870 ;
        RECT 1050.830 295.720 1051.830 299.870 ;
        RECT 1052.670 295.720 1054.130 299.870 ;
        RECT 1054.970 295.720 1056.430 299.870 ;
        RECT 1057.270 295.720 1058.730 299.870 ;
        RECT 1059.570 295.720 1061.030 299.870 ;
        RECT 1061.870 295.720 1063.330 299.870 ;
        RECT 1064.170 295.720 1065.170 299.870 ;
        RECT 1066.010 295.720 1067.470 299.870 ;
        RECT 1068.310 295.720 1069.770 299.870 ;
        RECT 1070.610 295.720 1072.070 299.870 ;
        RECT 1072.910 295.720 1074.370 299.870 ;
        RECT 1075.210 295.720 1076.210 299.870 ;
        RECT 1077.050 295.720 1078.510 299.870 ;
        RECT 1079.350 295.720 1080.810 299.870 ;
        RECT 1081.650 295.720 1083.110 299.870 ;
        RECT 1083.950 295.720 1085.410 299.870 ;
        RECT 1086.250 295.720 1087.250 299.870 ;
        RECT 1088.090 295.720 1089.550 299.870 ;
        RECT 1090.390 295.720 1091.850 299.870 ;
        RECT 1092.690 295.720 1094.150 299.870 ;
        RECT 1094.990 295.720 1096.450 299.870 ;
        RECT 1097.290 295.720 1098.750 299.870 ;
        RECT 1099.590 295.720 1100.590 299.870 ;
        RECT 1101.430 295.720 1102.890 299.870 ;
        RECT 1103.730 295.720 1105.190 299.870 ;
        RECT 1106.030 295.720 1107.490 299.870 ;
        RECT 1108.330 295.720 1109.790 299.870 ;
        RECT 1110.630 295.720 1111.630 299.870 ;
        RECT 1112.470 295.720 1113.930 299.870 ;
        RECT 1114.770 295.720 1116.230 299.870 ;
        RECT 1117.070 295.720 1118.530 299.870 ;
        RECT 1119.370 295.720 1120.830 299.870 ;
        RECT 1121.670 295.720 1122.670 299.870 ;
        RECT 1123.510 295.720 1124.970 299.870 ;
        RECT 1125.810 295.720 1127.270 299.870 ;
        RECT 1128.110 295.720 1129.570 299.870 ;
        RECT 1130.410 295.720 1131.870 299.870 ;
        RECT 1132.710 295.720 1134.170 299.870 ;
        RECT 1135.010 295.720 1136.010 299.870 ;
        RECT 1136.850 295.720 1138.310 299.870 ;
        RECT 1139.150 295.720 1140.610 299.870 ;
        RECT 1141.450 295.720 1142.910 299.870 ;
        RECT 1143.750 295.720 1145.210 299.870 ;
        RECT 1146.050 295.720 1147.050 299.870 ;
        RECT 1147.890 295.720 1149.350 299.870 ;
        RECT 1150.190 295.720 1151.650 299.870 ;
        RECT 1152.490 295.720 1153.950 299.870 ;
        RECT 1154.790 295.720 1156.250 299.870 ;
        RECT 1157.090 295.720 1158.090 299.870 ;
        RECT 1158.930 295.720 1160.390 299.870 ;
        RECT 1161.230 295.720 1162.690 299.870 ;
        RECT 1163.530 295.720 1164.990 299.870 ;
        RECT 1165.830 295.720 1167.290 299.870 ;
        RECT 1168.130 295.720 1169.590 299.870 ;
        RECT 1170.430 295.720 1171.430 299.870 ;
        RECT 1172.270 295.720 1173.730 299.870 ;
        RECT 1174.570 295.720 1176.030 299.870 ;
        RECT 1176.870 295.720 1178.330 299.870 ;
        RECT 1179.170 295.720 1180.630 299.870 ;
        RECT 1181.470 295.720 1182.470 299.870 ;
        RECT 1183.310 295.720 1184.770 299.870 ;
        RECT 1185.610 295.720 1187.070 299.870 ;
        RECT 1187.910 295.720 1189.370 299.870 ;
        RECT 1190.210 295.720 1191.670 299.870 ;
        RECT 1192.510 295.720 1193.510 299.870 ;
        RECT 1194.350 295.720 1195.810 299.870 ;
        RECT 1196.650 295.720 1198.110 299.870 ;
        RECT 1198.950 295.720 1200.410 299.870 ;
        RECT 1201.250 295.720 1202.710 299.870 ;
        RECT 1203.550 295.720 1205.010 299.870 ;
        RECT 1205.850 295.720 1206.850 299.870 ;
        RECT 1207.690 295.720 1209.150 299.870 ;
        RECT 1209.990 295.720 1211.450 299.870 ;
        RECT 1212.290 295.720 1213.750 299.870 ;
        RECT 1214.590 295.720 1216.050 299.870 ;
        RECT 1216.890 295.720 1217.890 299.870 ;
        RECT 1218.730 295.720 1220.190 299.870 ;
        RECT 1221.030 295.720 1222.490 299.870 ;
        RECT 1223.330 295.720 1224.790 299.870 ;
        RECT 1225.630 295.720 1227.090 299.870 ;
        RECT 1227.930 295.720 1228.930 299.870 ;
        RECT 1229.770 295.720 1231.230 299.870 ;
        RECT 1232.070 295.720 1233.530 299.870 ;
        RECT 1234.370 295.720 1235.830 299.870 ;
        RECT 1236.670 295.720 1238.130 299.870 ;
        RECT 1238.970 295.720 1240.430 299.870 ;
        RECT 1241.270 295.720 1242.270 299.870 ;
        RECT 1243.110 295.720 1244.570 299.870 ;
        RECT 1245.410 295.720 1246.870 299.870 ;
        RECT 1247.710 295.720 1249.170 299.870 ;
        RECT 1250.010 295.720 1251.470 299.870 ;
        RECT 1252.310 295.720 1253.310 299.870 ;
        RECT 1254.150 295.720 1255.610 299.870 ;
        RECT 1256.450 295.720 1257.910 299.870 ;
        RECT 1258.750 295.720 1260.210 299.870 ;
        RECT 1261.050 295.720 1262.510 299.870 ;
        RECT 1263.350 295.720 1264.350 299.870 ;
        RECT 1265.190 295.720 1266.650 299.870 ;
        RECT 1267.490 295.720 1268.950 299.870 ;
        RECT 1269.790 295.720 1271.250 299.870 ;
        RECT 1272.090 295.720 1273.550 299.870 ;
        RECT 1274.390 295.720 1275.850 299.870 ;
        RECT 1276.690 295.720 1277.690 299.870 ;
        RECT 1278.530 295.720 1279.990 299.870 ;
        RECT 1280.830 295.720 1282.290 299.870 ;
        RECT 1283.130 295.720 1284.590 299.870 ;
        RECT 1285.430 295.720 1286.890 299.870 ;
        RECT 1287.730 295.720 1288.730 299.870 ;
        RECT 1289.570 295.720 1291.030 299.870 ;
        RECT 1291.870 295.720 1293.330 299.870 ;
        RECT 1294.170 295.720 1295.630 299.870 ;
        RECT 1296.470 295.720 1297.930 299.870 ;
        RECT 1298.770 295.720 1299.770 299.870 ;
        RECT 1300.610 295.720 1302.070 299.870 ;
        RECT 1302.910 295.720 1304.370 299.870 ;
        RECT 1305.210 295.720 1306.670 299.870 ;
        RECT 1307.510 295.720 1308.970 299.870 ;
        RECT 1309.810 295.720 1311.270 299.870 ;
        RECT 1312.110 295.720 1313.110 299.870 ;
        RECT 1313.950 295.720 1315.410 299.870 ;
        RECT 1316.250 295.720 1317.710 299.870 ;
        RECT 1318.550 295.720 1320.010 299.870 ;
        RECT 1320.850 295.720 1322.310 299.870 ;
        RECT 1323.150 295.720 1324.150 299.870 ;
        RECT 1324.990 295.720 1326.450 299.870 ;
        RECT 1327.290 295.720 1328.750 299.870 ;
        RECT 1329.590 295.720 1331.050 299.870 ;
        RECT 1331.890 295.720 1333.350 299.870 ;
        RECT 1334.190 295.720 1335.190 299.870 ;
        RECT 1336.030 295.720 1337.490 299.870 ;
        RECT 1338.330 295.720 1339.790 299.870 ;
        RECT 1340.630 295.720 1342.090 299.870 ;
        RECT 1342.930 295.720 1344.390 299.870 ;
        RECT 1345.230 295.720 1346.690 299.870 ;
        RECT 1347.530 295.720 1348.530 299.870 ;
        RECT 1349.370 295.720 1350.830 299.870 ;
        RECT 1351.670 295.720 1353.130 299.870 ;
        RECT 1353.970 295.720 1355.430 299.870 ;
        RECT 1356.270 295.720 1357.730 299.870 ;
        RECT 1358.570 295.720 1359.570 299.870 ;
        RECT 1360.410 295.720 1361.870 299.870 ;
        RECT 1362.710 295.720 1364.170 299.870 ;
        RECT 1365.010 295.720 1366.470 299.870 ;
        RECT 1367.310 295.720 1368.770 299.870 ;
        RECT 1369.610 295.720 1370.610 299.870 ;
        RECT 1371.450 295.720 1372.910 299.870 ;
        RECT 1373.750 295.720 1375.210 299.870 ;
        RECT 1376.050 295.720 1377.510 299.870 ;
        RECT 1378.350 295.720 1379.810 299.870 ;
        RECT 1380.650 295.720 1382.110 299.870 ;
        RECT 1382.950 295.720 1383.950 299.870 ;
        RECT 1384.790 295.720 1386.250 299.870 ;
        RECT 1387.090 295.720 1388.550 299.870 ;
        RECT 1389.390 295.720 1390.850 299.870 ;
        RECT 1391.690 295.720 1393.150 299.870 ;
        RECT 1393.990 295.720 1394.990 299.870 ;
        RECT 1395.830 295.720 1397.290 299.870 ;
        RECT 1398.130 295.720 1399.590 299.870 ;
        RECT 1400.430 295.720 1401.890 299.870 ;
        RECT 1402.730 295.720 1404.190 299.870 ;
        RECT 1405.030 295.720 1406.030 299.870 ;
        RECT 1406.870 295.720 1408.330 299.870 ;
        RECT 1409.170 295.720 1410.630 299.870 ;
        RECT 1411.470 295.720 1412.930 299.870 ;
        RECT 1413.770 295.720 1415.230 299.870 ;
        RECT 1416.070 295.720 1417.530 299.870 ;
        RECT 1418.370 295.720 1419.370 299.870 ;
        RECT 1420.210 295.720 1421.670 299.870 ;
        RECT 1422.510 295.720 1423.970 299.870 ;
        RECT 1424.810 295.720 1426.270 299.870 ;
        RECT 1427.110 295.720 1428.570 299.870 ;
        RECT 1429.410 295.720 1430.410 299.870 ;
        RECT 1431.250 295.720 1432.710 299.870 ;
        RECT 1433.550 295.720 1435.010 299.870 ;
        RECT 1435.850 295.720 1437.310 299.870 ;
        RECT 1438.150 295.720 1439.610 299.870 ;
        RECT 1440.450 295.720 1441.450 299.870 ;
        RECT 1442.290 295.720 1443.750 299.870 ;
        RECT 1444.590 295.720 1446.050 299.870 ;
        RECT 1446.890 295.720 1448.350 299.870 ;
        RECT 1449.190 295.720 1450.650 299.870 ;
        RECT 1451.490 295.720 1452.950 299.870 ;
        RECT 1453.790 295.720 1454.790 299.870 ;
        RECT 1455.630 295.720 1457.090 299.870 ;
        RECT 1457.930 295.720 1459.390 299.870 ;
        RECT 1460.230 295.720 1461.690 299.870 ;
        RECT 1462.530 295.720 1463.990 299.870 ;
        RECT 1464.830 295.720 1465.830 299.870 ;
        RECT 1466.670 295.720 1468.130 299.870 ;
        RECT 1468.970 295.720 1470.430 299.870 ;
        RECT 1471.270 295.720 1472.730 299.870 ;
        RECT 1473.570 295.720 1475.030 299.870 ;
        RECT 1475.870 295.720 1476.870 299.870 ;
        RECT 1477.710 295.720 1479.170 299.870 ;
        RECT 1480.010 295.720 1481.470 299.870 ;
        RECT 1482.310 295.720 1483.770 299.870 ;
        RECT 1484.610 295.720 1486.070 299.870 ;
        RECT 1486.910 295.720 1488.370 299.870 ;
        RECT 1489.210 295.720 1490.210 299.870 ;
        RECT 1491.050 295.720 1492.510 299.870 ;
        RECT 1493.350 295.720 1494.810 299.870 ;
        RECT 1495.650 295.720 1497.110 299.870 ;
        RECT 1497.950 295.720 1499.410 299.870 ;
        RECT 1500.250 295.720 1501.250 299.870 ;
        RECT 1502.090 295.720 1503.550 299.870 ;
        RECT 1504.390 295.720 1505.850 299.870 ;
        RECT 1506.690 295.720 1508.150 299.870 ;
        RECT 1508.990 295.720 1510.450 299.870 ;
        RECT 1511.290 295.720 1512.290 299.870 ;
        RECT 1513.130 295.720 1514.590 299.870 ;
        RECT 1515.430 295.720 1516.890 299.870 ;
        RECT 1517.730 295.720 1519.190 299.870 ;
        RECT 1520.030 295.720 1521.490 299.870 ;
        RECT 1522.330 295.720 1523.790 299.870 ;
        RECT 1524.630 295.720 1525.630 299.870 ;
        RECT 1526.470 295.720 1527.930 299.870 ;
        RECT 1528.770 295.720 1530.230 299.870 ;
        RECT 1531.070 295.720 1532.530 299.870 ;
        RECT 1533.370 295.720 1534.830 299.870 ;
        RECT 1535.670 295.720 1536.670 299.870 ;
        RECT 1537.510 295.720 1538.970 299.870 ;
        RECT 1539.810 295.720 1541.270 299.870 ;
        RECT 1542.110 295.720 1543.570 299.870 ;
        RECT 1544.410 295.720 1545.870 299.870 ;
        RECT 1546.710 295.720 1547.710 299.870 ;
        RECT 1548.550 295.720 1550.010 299.870 ;
        RECT 1550.850 295.720 1552.310 299.870 ;
        RECT 1553.150 295.720 1554.610 299.870 ;
        RECT 1555.450 295.720 1556.910 299.870 ;
        RECT 1557.750 295.720 1559.210 299.870 ;
        RECT 1560.050 295.720 1561.050 299.870 ;
        RECT 1561.890 295.720 1563.350 299.870 ;
        RECT 1564.190 295.720 1565.650 299.870 ;
        RECT 1566.490 295.720 1567.950 299.870 ;
        RECT 1568.790 295.720 1570.250 299.870 ;
        RECT 1571.090 295.720 1572.090 299.870 ;
        RECT 1572.930 295.720 1574.390 299.870 ;
        RECT 1575.230 295.720 1576.690 299.870 ;
        RECT 1577.530 295.720 1578.990 299.870 ;
        RECT 1579.830 295.720 1581.290 299.870 ;
        RECT 1582.130 295.720 1583.130 299.870 ;
        RECT 1583.970 295.720 1585.430 299.870 ;
        RECT 1586.270 295.720 1587.730 299.870 ;
        RECT 1588.570 295.720 1590.030 299.870 ;
        RECT 1590.870 295.720 1592.330 299.870 ;
        RECT 1593.170 295.720 1594.630 299.870 ;
        RECT 1595.470 295.720 1596.470 299.870 ;
        RECT 1597.310 295.720 1598.770 299.870 ;
        RECT 1599.610 295.720 1601.070 299.870 ;
        RECT 1601.910 295.720 1603.370 299.870 ;
        RECT 1604.210 295.720 1605.670 299.870 ;
        RECT 1606.510 295.720 1607.510 299.870 ;
        RECT 1608.350 295.720 1609.810 299.870 ;
        RECT 1610.650 295.720 1612.110 299.870 ;
        RECT 1612.950 295.720 1614.410 299.870 ;
        RECT 1615.250 295.720 1616.710 299.870 ;
        RECT 1617.550 295.720 1618.550 299.870 ;
        RECT 1619.390 295.720 1620.850 299.870 ;
        RECT 1621.690 295.720 1623.150 299.870 ;
        RECT 1623.990 295.720 1625.450 299.870 ;
        RECT 1626.290 295.720 1627.750 299.870 ;
        RECT 1628.590 295.720 1630.050 299.870 ;
        RECT 1630.890 295.720 1631.890 299.870 ;
        RECT 1632.730 295.720 1634.190 299.870 ;
        RECT 1635.030 295.720 1636.490 299.870 ;
        RECT 1637.330 295.720 1638.790 299.870 ;
        RECT 1639.630 295.720 1641.090 299.870 ;
        RECT 1641.930 295.720 1642.930 299.870 ;
        RECT 1643.770 295.720 1645.230 299.870 ;
        RECT 1646.070 295.720 1647.530 299.870 ;
        RECT 1648.370 295.720 1649.830 299.870 ;
        RECT 1650.670 295.720 1652.130 299.870 ;
        RECT 1652.970 295.720 1653.970 299.870 ;
        RECT 1654.810 295.720 1656.270 299.870 ;
        RECT 1657.110 295.720 1658.570 299.870 ;
        RECT 1659.410 295.720 1660.870 299.870 ;
        RECT 1661.710 295.720 1663.170 299.870 ;
        RECT 1664.010 295.720 1665.470 299.870 ;
        RECT 1666.310 295.720 1667.310 299.870 ;
        RECT 1668.150 295.720 1669.610 299.870 ;
        RECT 1670.450 295.720 1671.910 299.870 ;
        RECT 1672.750 295.720 1674.210 299.870 ;
        RECT 1675.050 295.720 1676.510 299.870 ;
        RECT 1677.350 295.720 1678.350 299.870 ;
        RECT 1679.190 295.720 1680.650 299.870 ;
        RECT 1681.490 295.720 1682.950 299.870 ;
        RECT 1683.790 295.720 1685.250 299.870 ;
        RECT 1686.090 295.720 1687.550 299.870 ;
        RECT 1688.390 295.720 1689.390 299.870 ;
        RECT 1690.230 295.720 1691.690 299.870 ;
        RECT 1692.530 295.720 1693.990 299.870 ;
        RECT 1694.830 295.720 1696.290 299.870 ;
        RECT 1697.130 295.720 1698.590 299.870 ;
        RECT 1.020 4.280 1699.140 295.720 ;
        RECT 1.020 3.670 7.630 4.280 ;
        RECT 8.470 3.670 23.270 4.280 ;
        RECT 24.110 3.670 39.370 4.280 ;
        RECT 40.210 3.670 55.470 4.280 ;
        RECT 56.310 3.670 71.570 4.280 ;
        RECT 72.410 3.670 87.670 4.280 ;
        RECT 88.510 3.670 103.770 4.280 ;
        RECT 104.610 3.670 119.870 4.280 ;
        RECT 120.710 3.670 135.510 4.280 ;
        RECT 136.350 3.670 151.610 4.280 ;
        RECT 152.450 3.670 167.710 4.280 ;
        RECT 168.550 3.670 183.810 4.280 ;
        RECT 184.650 3.670 199.910 4.280 ;
        RECT 200.750 3.670 216.010 4.280 ;
        RECT 216.850 3.670 232.110 4.280 ;
        RECT 232.950 3.670 248.210 4.280 ;
        RECT 249.050 3.670 263.850 4.280 ;
        RECT 264.690 3.670 279.950 4.280 ;
        RECT 280.790 3.670 296.050 4.280 ;
        RECT 296.890 3.670 312.150 4.280 ;
        RECT 312.990 3.670 328.250 4.280 ;
        RECT 329.090 3.670 344.350 4.280 ;
        RECT 345.190 3.670 360.450 4.280 ;
        RECT 361.290 3.670 376.090 4.280 ;
        RECT 376.930 3.670 392.190 4.280 ;
        RECT 393.030 3.670 408.290 4.280 ;
        RECT 409.130 3.670 424.390 4.280 ;
        RECT 425.230 3.670 440.490 4.280 ;
        RECT 441.330 3.670 456.590 4.280 ;
        RECT 457.430 3.670 472.690 4.280 ;
        RECT 473.530 3.670 488.790 4.280 ;
        RECT 489.630 3.670 504.430 4.280 ;
        RECT 505.270 3.670 520.530 4.280 ;
        RECT 521.370 3.670 536.630 4.280 ;
        RECT 537.470 3.670 552.730 4.280 ;
        RECT 553.570 3.670 568.830 4.280 ;
        RECT 569.670 3.670 584.930 4.280 ;
        RECT 585.770 3.670 601.030 4.280 ;
        RECT 601.870 3.670 616.670 4.280 ;
        RECT 617.510 3.670 632.770 4.280 ;
        RECT 633.610 3.670 648.870 4.280 ;
        RECT 649.710 3.670 664.970 4.280 ;
        RECT 665.810 3.670 681.070 4.280 ;
        RECT 681.910 3.670 697.170 4.280 ;
        RECT 698.010 3.670 713.270 4.280 ;
        RECT 714.110 3.670 729.370 4.280 ;
        RECT 730.210 3.670 745.010 4.280 ;
        RECT 745.850 3.670 761.110 4.280 ;
        RECT 761.950 3.670 777.210 4.280 ;
        RECT 778.050 3.670 793.310 4.280 ;
        RECT 794.150 3.670 809.410 4.280 ;
        RECT 810.250 3.670 825.510 4.280 ;
        RECT 826.350 3.670 841.610 4.280 ;
        RECT 842.450 3.670 857.710 4.280 ;
        RECT 858.550 3.670 873.350 4.280 ;
        RECT 874.190 3.670 889.450 4.280 ;
        RECT 890.290 3.670 905.550 4.280 ;
        RECT 906.390 3.670 921.650 4.280 ;
        RECT 922.490 3.670 937.750 4.280 ;
        RECT 938.590 3.670 953.850 4.280 ;
        RECT 954.690 3.670 969.950 4.280 ;
        RECT 970.790 3.670 985.590 4.280 ;
        RECT 986.430 3.670 1001.690 4.280 ;
        RECT 1002.530 3.670 1017.790 4.280 ;
        RECT 1018.630 3.670 1033.890 4.280 ;
        RECT 1034.730 3.670 1049.990 4.280 ;
        RECT 1050.830 3.670 1066.090 4.280 ;
        RECT 1066.930 3.670 1082.190 4.280 ;
        RECT 1083.030 3.670 1098.290 4.280 ;
        RECT 1099.130 3.670 1113.930 4.280 ;
        RECT 1114.770 3.670 1130.030 4.280 ;
        RECT 1130.870 3.670 1146.130 4.280 ;
        RECT 1146.970 3.670 1162.230 4.280 ;
        RECT 1163.070 3.670 1178.330 4.280 ;
        RECT 1179.170 3.670 1194.430 4.280 ;
        RECT 1195.270 3.670 1210.530 4.280 ;
        RECT 1211.370 3.670 1226.170 4.280 ;
        RECT 1227.010 3.670 1242.270 4.280 ;
        RECT 1243.110 3.670 1258.370 4.280 ;
        RECT 1259.210 3.670 1274.470 4.280 ;
        RECT 1275.310 3.670 1290.570 4.280 ;
        RECT 1291.410 3.670 1306.670 4.280 ;
        RECT 1307.510 3.670 1322.770 4.280 ;
        RECT 1323.610 3.670 1338.870 4.280 ;
        RECT 1339.710 3.670 1354.510 4.280 ;
        RECT 1355.350 3.670 1370.610 4.280 ;
        RECT 1371.450 3.670 1386.710 4.280 ;
        RECT 1387.550 3.670 1402.810 4.280 ;
        RECT 1403.650 3.670 1418.910 4.280 ;
        RECT 1419.750 3.670 1435.010 4.280 ;
        RECT 1435.850 3.670 1451.110 4.280 ;
        RECT 1451.950 3.670 1466.750 4.280 ;
        RECT 1467.590 3.670 1482.850 4.280 ;
        RECT 1483.690 3.670 1498.950 4.280 ;
        RECT 1499.790 3.670 1515.050 4.280 ;
        RECT 1515.890 3.670 1531.150 4.280 ;
        RECT 1531.990 3.670 1547.250 4.280 ;
        RECT 1548.090 3.670 1563.350 4.280 ;
        RECT 1564.190 3.670 1579.450 4.280 ;
        RECT 1580.290 3.670 1595.090 4.280 ;
        RECT 1595.930 3.670 1611.190 4.280 ;
        RECT 1612.030 3.670 1627.290 4.280 ;
        RECT 1628.130 3.670 1643.390 4.280 ;
        RECT 1644.230 3.670 1659.490 4.280 ;
        RECT 1660.330 3.670 1675.590 4.280 ;
        RECT 1676.430 3.670 1691.690 4.280 ;
        RECT 1692.530 3.670 1699.140 4.280 ;
      LAYER met3 ;
        RECT 11.105 270.320 1696.000 294.945 ;
        RECT 11.105 268.920 1695.600 270.320 ;
        RECT 11.105 210.480 1696.000 268.920 ;
        RECT 11.105 209.080 1695.600 210.480 ;
        RECT 11.105 150.640 1696.000 209.080 ;
        RECT 11.105 149.240 1695.600 150.640 ;
        RECT 11.105 90.800 1696.000 149.240 ;
        RECT 11.105 89.400 1695.600 90.800 ;
        RECT 11.105 30.960 1696.000 89.400 ;
        RECT 11.105 29.560 1695.600 30.960 ;
        RECT 11.105 10.715 1696.000 29.560 ;
      LAYER met4 ;
        RECT 191.655 288.960 1539.785 294.265 ;
        RECT 191.655 17.175 251.040 288.960 ;
        RECT 253.440 17.175 327.840 288.960 ;
        RECT 330.240 17.175 404.640 288.960 ;
        RECT 407.040 17.175 481.440 288.960 ;
        RECT 483.840 17.175 558.240 288.960 ;
        RECT 560.640 17.175 635.040 288.960 ;
        RECT 637.440 17.175 711.840 288.960 ;
        RECT 714.240 17.175 788.640 288.960 ;
        RECT 791.040 17.175 865.440 288.960 ;
        RECT 867.840 17.175 942.240 288.960 ;
        RECT 944.640 17.175 1019.040 288.960 ;
        RECT 1021.440 17.175 1095.840 288.960 ;
        RECT 1098.240 17.175 1172.640 288.960 ;
        RECT 1175.040 17.175 1249.440 288.960 ;
        RECT 1251.840 17.175 1326.240 288.960 ;
        RECT 1328.640 17.175 1403.040 288.960 ;
        RECT 1405.440 17.175 1479.840 288.960 ;
        RECT 1482.240 17.175 1539.785 288.960 ;
  END
END soric_soc
END LIBRARY

