VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ibex_top
  CLASS BLOCK ;
  FOREIGN ibex_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN alert_major_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END alert_major_o
  PIN alert_minor_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 3.440 1200.000 4.040 ;
    END
  END alert_minor_o
  PIN boot_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END boot_addr_i[0]
  PIN boot_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 403.280 1200.000 403.880 ;
    END
  END boot_addr_i[10]
  PIN boot_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END boot_addr_i[11]
  PIN boot_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 454.280 1200.000 454.880 ;
    END
  END boot_addr_i[12]
  PIN boot_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 1196.000 414.370 1200.000 ;
    END
  END boot_addr_i[13]
  PIN boot_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END boot_addr_i[14]
  PIN boot_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 1196.000 461.750 1200.000 ;
    END
  END boot_addr_i[15]
  PIN boot_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END boot_addr_i[16]
  PIN boot_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END boot_addr_i[17]
  PIN boot_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 606.600 1200.000 607.200 ;
    END
  END boot_addr_i[18]
  PIN boot_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 635.840 1200.000 636.440 ;
    END
  END boot_addr_i[19]
  PIN boot_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END boot_addr_i[1]
  PIN boot_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 672.560 1200.000 673.160 ;
    END
  END boot_addr_i[20]
  PIN boot_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 0.000 762.590 4.000 ;
    END
  END boot_addr_i[21]
  PIN boot_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END boot_addr_i[22]
  PIN boot_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 752.120 1200.000 752.720 ;
    END
  END boot_addr_i[23]
  PIN boot_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.880 4.000 825.480 ;
    END
  END boot_addr_i[24]
  PIN boot_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.160 4.000 873.760 ;
    END
  END boot_addr_i[25]
  PIN boot_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 1196.000 776.390 1200.000 ;
    END
  END boot_addr_i[26]
  PIN boot_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 913.280 4.000 913.880 ;
    END
  END boot_addr_i[27]
  PIN boot_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.810 1196.000 843.090 1200.000 ;
    END
  END boot_addr_i[28]
  PIN boot_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 0.000 937.850 4.000 ;
    END
  END boot_addr_i[29]
  PIN boot_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END boot_addr_i[2]
  PIN boot_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.720 4.000 970.320 ;
    END
  END boot_addr_i[30]
  PIN boot_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 977.880 1200.000 978.480 ;
    END
  END boot_addr_i[31]
  PIN boot_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END boot_addr_i[3]
  PIN boot_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 1196.000 166.890 1200.000 ;
    END
  END boot_addr_i[4]
  PIN boot_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 1196.000 214.270 1200.000 ;
    END
  END boot_addr_i[5]
  PIN boot_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END boot_addr_i[6]
  PIN boot_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 323.040 1200.000 323.640 ;
    END
  END boot_addr_i[7]
  PIN boot_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 366.560 1200.000 367.160 ;
    END
  END boot_addr_i[8]
  PIN boot_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 1196.000 252.450 1200.000 ;
    END
  END boot_addr_i[9]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 10.240 1200.000 10.840 ;
    END
  END clk_i
  PIN core_sleep_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END core_sleep_o
  PIN crash_dump_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END crash_dump_o[0]
  PIN crash_dump_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.200 4.000 1147.800 ;
    END
  END crash_dump_o[100]
  PIN crash_dump_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1130.880 1200.000 1131.480 ;
    END
  END crash_dump_o[101]
  PIN crash_dump_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1154.680 4.000 1155.280 ;
    END
  END crash_dump_o[102]
  PIN crash_dump_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.230 0.000 1154.510 4.000 ;
    END
  END crash_dump_o[103]
  PIN crash_dump_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END crash_dump_o[104]
  PIN crash_dump_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END crash_dump_o[105]
  PIN crash_dump_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1171.000 4.000 1171.600 ;
    END
  END crash_dump_o[106]
  PIN crash_dump_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1137.680 1200.000 1138.280 ;
    END
  END crash_dump_o[107]
  PIN crash_dump_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.160 4.000 1179.760 ;
    END
  END crash_dump_o[108]
  PIN crash_dump_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1145.160 1200.000 1145.760 ;
    END
  END crash_dump_o[109]
  PIN crash_dump_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END crash_dump_o[10]
  PIN crash_dump_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1152.640 1200.000 1153.240 ;
    END
  END crash_dump_o[110]
  PIN crash_dump_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1159.440 1200.000 1160.040 ;
    END
  END crash_dump_o[111]
  PIN crash_dump_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1166.920 1200.000 1167.520 ;
    END
  END crash_dump_o[112]
  PIN crash_dump_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.790 0.000 1171.070 4.000 ;
    END
  END crash_dump_o[113]
  PIN crash_dump_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.070 0.000 1179.350 4.000 ;
    END
  END crash_dump_o[114]
  PIN crash_dump_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1174.400 1200.000 1175.000 ;
    END
  END crash_dump_o[115]
  PIN crash_dump_o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1181.200 1200.000 1181.800 ;
    END
  END crash_dump_o[116]
  PIN crash_dump_o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1187.320 4.000 1187.920 ;
    END
  END crash_dump_o[117]
  PIN crash_dump_o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.990 1196.000 1157.270 1200.000 ;
    END
  END crash_dump_o[118]
  PIN crash_dump_o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.350 0.000 1187.630 4.000 ;
    END
  END crash_dump_o[119]
  PIN crash_dump_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 432.520 1200.000 433.120 ;
    END
  END crash_dump_o[11]
  PIN crash_dump_o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1188.680 1200.000 1189.280 ;
    END
  END crash_dump_o[120]
  PIN crash_dump_o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.650 1196.000 1166.930 1200.000 ;
    END
  END crash_dump_o[121]
  PIN crash_dump_o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 1196.000 1176.130 1200.000 ;
    END
  END crash_dump_o[122]
  PIN crash_dump_o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1196.160 1200.000 1196.760 ;
    END
  END crash_dump_o[123]
  PIN crash_dump_o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.510 1196.000 1185.790 1200.000 ;
    END
  END crash_dump_o[124]
  PIN crash_dump_o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.630 0.000 1195.910 4.000 ;
    END
  END crash_dump_o[125]
  PIN crash_dump_o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1195.480 4.000 1196.080 ;
    END
  END crash_dump_o[126]
  PIN crash_dump_o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 1196.000 1195.450 1200.000 ;
    END
  END crash_dump_o[127]
  PIN crash_dump_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 1196.000 376.190 1200.000 ;
    END
  END crash_dump_o[12]
  PIN crash_dump_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END crash_dump_o[13]
  PIN crash_dump_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END crash_dump_o[14]
  PIN crash_dump_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 527.040 1200.000 527.640 ;
    END
  END crash_dump_o[15]
  PIN crash_dump_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 1196.000 481.070 1200.000 ;
    END
  END crash_dump_o[16]
  PIN crash_dump_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END crash_dump_o[17]
  PIN crash_dump_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 687.520 4.000 688.120 ;
    END
  END crash_dump_o[18]
  PIN crash_dump_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 643.320 1200.000 643.920 ;
    END
  END crash_dump_o[19]
  PIN crash_dump_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 1196.000 71.210 1200.000 ;
    END
  END crash_dump_o[1]
  PIN crash_dump_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 679.360 1200.000 679.960 ;
    END
  END crash_dump_o[20]
  PIN crash_dump_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 1196.000 623.670 1200.000 ;
    END
  END crash_dump_o[21]
  PIN crash_dump_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 1196.000 652.650 1200.000 ;
    END
  END crash_dump_o[22]
  PIN crash_dump_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 1196.000 690.370 1200.000 ;
    END
  END crash_dump_o[23]
  PIN crash_dump_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 1196.000 718.890 1200.000 ;
    END
  END crash_dump_o[24]
  PIN crash_dump_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 1196.000 747.870 1200.000 ;
    END
  END crash_dump_o[25]
  PIN crash_dump_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 1196.000 785.590 1200.000 ;
    END
  END crash_dump_o[26]
  PIN crash_dump_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END crash_dump_o[27]
  PIN crash_dump_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 1196.000 852.290 1200.000 ;
    END
  END crash_dump_o[28]
  PIN crash_dump_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 926.880 1200.000 927.480 ;
    END
  END crash_dump_o[29]
  PIN crash_dump_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 112.240 1200.000 112.840 ;
    END
  END crash_dump_o[2]
  PIN crash_dump_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 948.640 1200.000 949.240 ;
    END
  END crash_dump_o[30]
  PIN crash_dump_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END crash_dump_o[31]
  PIN crash_dump_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.160 4.000 1026.760 ;
    END
  END crash_dump_o[32]
  PIN crash_dump_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1007.120 1200.000 1007.720 ;
    END
  END crash_dump_o[33]
  PIN crash_dump_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 0.000 1029.390 4.000 ;
    END
  END crash_dump_o[34]
  PIN crash_dump_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.890 1196.000 957.170 1200.000 ;
    END
  END crash_dump_o[35]
  PIN crash_dump_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1013.920 1200.000 1014.520 ;
    END
  END crash_dump_o[36]
  PIN crash_dump_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 1196.000 966.830 1200.000 ;
    END
  END crash_dump_o[37]
  PIN crash_dump_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 1196.000 976.490 1200.000 ;
    END
  END crash_dump_o[38]
  PIN crash_dump_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1034.320 4.000 1034.920 ;
    END
  END crash_dump_o[39]
  PIN crash_dump_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END crash_dump_o[3]
  PIN crash_dump_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1021.400 1200.000 1022.000 ;
    END
  END crash_dump_o[40]
  PIN crash_dump_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END crash_dump_o[41]
  PIN crash_dump_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 1196.000 985.690 1200.000 ;
    END
  END crash_dump_o[42]
  PIN crash_dump_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1028.880 1200.000 1029.480 ;
    END
  END crash_dump_o[43]
  PIN crash_dump_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1042.480 4.000 1043.080 ;
    END
  END crash_dump_o[44]
  PIN crash_dump_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 1196.000 995.350 1200.000 ;
    END
  END crash_dump_o[45]
  PIN crash_dump_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.670 0.000 1045.950 4.000 ;
    END
  END crash_dump_o[46]
  PIN crash_dump_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 0.000 1054.230 4.000 ;
    END
  END crash_dump_o[47]
  PIN crash_dump_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 1196.000 1005.010 1200.000 ;
    END
  END crash_dump_o[48]
  PIN crash_dump_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.960 4.000 1050.560 ;
    END
  END crash_dump_o[49]
  PIN crash_dump_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END crash_dump_o[4]
  PIN crash_dump_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 1196.000 1014.210 1200.000 ;
    END
  END crash_dump_o[50]
  PIN crash_dump_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.590 1196.000 1023.870 1200.000 ;
    END
  END crash_dump_o[51]
  PIN crash_dump_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1058.120 4.000 1058.720 ;
    END
  END crash_dump_o[52]
  PIN crash_dump_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 1196.000 1033.530 1200.000 ;
    END
  END crash_dump_o[53]
  PIN crash_dump_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.230 0.000 1062.510 4.000 ;
    END
  END crash_dump_o[54]
  PIN crash_dump_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.280 4.000 1066.880 ;
    END
  END crash_dump_o[55]
  PIN crash_dump_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1035.680 1200.000 1036.280 ;
    END
  END crash_dump_o[56]
  PIN crash_dump_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.450 1196.000 1042.730 1200.000 ;
    END
  END crash_dump_o[57]
  PIN crash_dump_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END crash_dump_o[58]
  PIN crash_dump_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.110 1196.000 1052.390 1200.000 ;
    END
  END crash_dump_o[59]
  PIN crash_dump_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 221.040 1200.000 221.640 ;
    END
  END crash_dump_o[5]
  PIN crash_dump_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1043.160 1200.000 1043.760 ;
    END
  END crash_dump_o[60]
  PIN crash_dump_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.770 1196.000 1062.050 1200.000 ;
    END
  END crash_dump_o[61]
  PIN crash_dump_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.970 0.000 1071.250 4.000 ;
    END
  END crash_dump_o[62]
  PIN crash_dump_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1082.600 4.000 1083.200 ;
    END
  END crash_dump_o[63]
  PIN crash_dump_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1090.760 4.000 1091.360 ;
    END
  END crash_dump_o[64]
  PIN crash_dump_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 0.000 1079.530 4.000 ;
    END
  END crash_dump_o[65]
  PIN crash_dump_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1050.640 1200.000 1051.240 ;
    END
  END crash_dump_o[66]
  PIN crash_dump_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 1196.000 1071.710 1200.000 ;
    END
  END crash_dump_o[67]
  PIN crash_dump_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 1196.000 1080.910 1200.000 ;
    END
  END crash_dump_o[68]
  PIN crash_dump_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 1196.000 1090.570 1200.000 ;
    END
  END crash_dump_o[69]
  PIN crash_dump_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END crash_dump_o[6]
  PIN crash_dump_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.920 4.000 1099.520 ;
    END
  END crash_dump_o[70]
  PIN crash_dump_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1106.400 4.000 1107.000 ;
    END
  END crash_dump_o[71]
  PIN crash_dump_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 0.000 1087.810 4.000 ;
    END
  END crash_dump_o[72]
  PIN crash_dump_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1114.560 4.000 1115.160 ;
    END
  END crash_dump_o[73]
  PIN crash_dump_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.950 1196.000 1100.230 1200.000 ;
    END
  END crash_dump_o[74]
  PIN crash_dump_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1058.120 1200.000 1058.720 ;
    END
  END crash_dump_o[75]
  PIN crash_dump_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1064.920 1200.000 1065.520 ;
    END
  END crash_dump_o[76]
  PIN crash_dump_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1072.400 1200.000 1073.000 ;
    END
  END crash_dump_o[77]
  PIN crash_dump_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 1196.000 1109.430 1200.000 ;
    END
  END crash_dump_o[78]
  PIN crash_dump_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 0.000 1096.090 4.000 ;
    END
  END crash_dump_o[79]
  PIN crash_dump_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END crash_dump_o[7]
  PIN crash_dump_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1079.880 1200.000 1080.480 ;
    END
  END crash_dump_o[80]
  PIN crash_dump_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.810 1196.000 1119.090 1200.000 ;
    END
  END crash_dump_o[81]
  PIN crash_dump_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END crash_dump_o[82]
  PIN crash_dump_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1086.680 1200.000 1087.280 ;
    END
  END crash_dump_o[83]
  PIN crash_dump_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1094.160 1200.000 1094.760 ;
    END
  END crash_dump_o[84]
  PIN crash_dump_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 1196.000 1128.750 1200.000 ;
    END
  END crash_dump_o[85]
  PIN crash_dump_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.720 4.000 1123.320 ;
    END
  END crash_dump_o[86]
  PIN crash_dump_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.370 0.000 1112.650 4.000 ;
    END
  END crash_dump_o[87]
  PIN crash_dump_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1130.880 4.000 1131.480 ;
    END
  END crash_dump_o[88]
  PIN crash_dump_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END crash_dump_o[89]
  PIN crash_dump_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END crash_dump_o[8]
  PIN crash_dump_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1101.640 1200.000 1102.240 ;
    END
  END crash_dump_o[90]
  PIN crash_dump_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1108.440 1200.000 1109.040 ;
    END
  END crash_dump_o[91]
  PIN crash_dump_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1115.920 1200.000 1116.520 ;
    END
  END crash_dump_o[92]
  PIN crash_dump_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 1196.000 1138.410 1200.000 ;
    END
  END crash_dump_o[93]
  PIN crash_dump_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 4.000 ;
    END
  END crash_dump_o[94]
  PIN crash_dump_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1123.400 1200.000 1124.000 ;
    END
  END crash_dump_o[95]
  PIN crash_dump_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.330 1196.000 1147.610 1200.000 ;
    END
  END crash_dump_o[96]
  PIN crash_dump_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END crash_dump_o[97]
  PIN crash_dump_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.670 0.000 1137.950 4.000 ;
    END
  END crash_dump_o[98]
  PIN crash_dump_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 0.000 1146.230 4.000 ;
    END
  END crash_dump_o[99]
  PIN crash_dump_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 395.800 1200.000 396.400 ;
    END
  END crash_dump_o[9]
  PIN data_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END data_addr_o[0]
  PIN data_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 494.400 4.000 495.000 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 461.080 1200.000 461.680 ;
    END
  END data_addr_o[12]
  PIN data_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END data_addr_o[13]
  PIN data_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END data_addr_o[14]
  PIN data_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END data_addr_o[15]
  PIN data_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 1196.000 490.730 1200.000 ;
    END
  END data_addr_o[16]
  PIN data_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END data_addr_o[17]
  PIN data_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 1196.000 528.450 1200.000 ;
    END
  END data_addr_o[18]
  PIN data_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 0.000 712.910 4.000 ;
    END
  END data_addr_o[19]
  PIN data_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1196.000 80.870 1200.000 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 1196.000 585.950 1200.000 ;
    END
  END data_addr_o[20]
  PIN data_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 708.600 1200.000 709.200 ;
    END
  END data_addr_o[21]
  PIN data_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 4.000 ;
    END
  END data_addr_o[22]
  PIN data_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 1196.000 700.030 1200.000 ;
    END
  END data_addr_o[23]
  PIN data_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 1196.000 728.550 1200.000 ;
    END
  END data_addr_o[24]
  PIN data_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 810.600 1200.000 811.200 ;
    END
  END data_addr_o[25]
  PIN data_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 839.840 1200.000 840.440 ;
    END
  END data_addr_o[26]
  PIN data_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 1196.000 814.570 1200.000 ;
    END
  END data_addr_o[27]
  PIN data_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 0.000 912.550 4.000 ;
    END
  END data_addr_o[28]
  PIN data_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 953.400 4.000 954.000 ;
    END
  END data_addr_o[29]
  PIN data_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1196.000 100.190 1200.000 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END data_addr_o[30]
  PIN data_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.710 1196.000 918.990 1200.000 ;
    END
  END data_addr_o[31]
  PIN data_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 177.520 1200.000 178.120 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 199.280 1200.000 199.880 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 228.520 1200.000 229.120 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 374.040 1200.000 374.640 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END data_addr_o[9]
  PIN data_be_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 46.960 1200.000 47.560 ;
    END
  END data_be_o[0]
  PIN data_be_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END data_be_o[1]
  PIN data_be_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END data_be_o[2]
  PIN data_be_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 185.000 1200.000 185.600 ;
    END
  END data_be_o[3]
  PIN data_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END data_err_i
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END data_gnt_i
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END data_rdata_i[0]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 410.760 1200.000 411.360 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 439.320 1200.000 439.920 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 468.560 1200.000 469.160 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 1196.000 424.030 1200.000 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 1196.000 499.930 1200.000 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 570.560 1200.000 571.160 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.680 4.000 696.280 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1196.000 90.530 1200.000 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 686.840 1200.000 687.440 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 788.840 1200.000 789.440 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 1196.000 757.070 1200.000 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 0.000 862.870 4.000 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 0.000 887.710 4.000 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 905.120 1200.000 905.720 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 934.360 1200.000 934.960 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.880 4.000 978.480 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 330.520 1200.000 331.120 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END data_rdata_i[9]
  PIN data_rdata_intg_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END data_rdata_intg_i[0]
  PIN data_rdata_intg_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END data_rdata_intg_i[1]
  PIN data_rdata_intg_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 1196.000 109.390 1200.000 ;
    END
  END data_rdata_intg_i[2]
  PIN data_rdata_intg_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 1196.000 128.710 1200.000 ;
    END
  END data_rdata_intg_i[3]
  PIN data_rdata_intg_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 206.760 1200.000 207.360 ;
    END
  END data_rdata_intg_i[4]
  PIN data_rdata_intg_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END data_rdata_intg_i[5]
  PIN data_rdata_intg_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 265.240 1200.000 265.840 ;
    END
  END data_rdata_intg_i[6]
  PIN data_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END data_req_o
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 1196.000 4.970 1200.000 ;
    END
  END data_rvalid_i
  PIN data_wdata_intg_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END data_wdata_intg_o[0]
  PIN data_wdata_intg_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END data_wdata_intg_o[1]
  PIN data_wdata_intg_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 119.720 1200.000 120.320 ;
    END
  END data_wdata_intg_o[2]
  PIN data_wdata_intg_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 1196.000 137.910 1200.000 ;
    END
  END data_wdata_intg_o[3]
  PIN data_wdata_intg_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 1196.000 176.090 1200.000 ;
    END
  END data_wdata_intg_o[4]
  PIN data_wdata_intg_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 236.000 1200.000 236.600 ;
    END
  END data_wdata_intg_o[5]
  PIN data_wdata_intg_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 272.040 1200.000 272.640 ;
    END
  END data_wdata_intg_o[6]
  PIN data_wdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END data_wdata_o[0]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 1196.000 328.810 1200.000 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 1196.000 442.890 1200.000 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 533.840 1200.000 534.440 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 614.080 1200.000 614.680 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 1196.000 566.630 1200.000 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 68.720 1200.000 69.320 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 1196.000 595.150 1200.000 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 0.000 779.150 4.000 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 759.600 1200.000 760.200 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 0.000 829.290 4.000 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 818.080 1200.000 818.680 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.960 4.000 897.560 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 1196.000 861.950 1200.000 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.530 1196.000 880.810 1200.000 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 126.520 1200.000 127.120 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 985.360 1200.000 985.960 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 1196.000 223.930 1200.000 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 279.520 1200.000 280.120 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 338.000 1200.000 338.600 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END data_wdata_o[9]
  PIN data_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END data_we_o
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 1196.000 14.170 1200.000 ;
    END
  END debug_req_i
  PIN eFPGA_delay_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 1196.000 52.350 1200.000 ;
    END
  END eFPGA_delay_o[0]
  PIN eFPGA_delay_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END eFPGA_delay_o[1]
  PIN eFPGA_delay_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 134.000 1200.000 134.600 ;
    END
  END eFPGA_delay_o[2]
  PIN eFPGA_delay_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END eFPGA_delay_o[3]
  PIN eFPGA_en_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 17.720 1200.000 18.320 ;
    END
  END eFPGA_en_o
  PIN eFPGA_fpga_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 1196.000 23.830 1200.000 ;
    END
  END eFPGA_fpga_done_i
  PIN eFPGA_operand_a_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END eFPGA_operand_a_o[0]
  PIN eFPGA_operand_a_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 417.560 1200.000 418.160 ;
    END
  END eFPGA_operand_a_o[10]
  PIN eFPGA_operand_a_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 1196.000 338.010 1200.000 ;
    END
  END eFPGA_operand_a_o[11]
  PIN eFPGA_operand_a_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 476.040 1200.000 476.640 ;
    END
  END eFPGA_operand_a_o[12]
  PIN eFPGA_operand_a_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END eFPGA_operand_a_o[13]
  PIN eFPGA_operand_a_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END eFPGA_operand_a_o[14]
  PIN eFPGA_operand_a_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END eFPGA_operand_a_o[15]
  PIN eFPGA_operand_a_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 1196.000 509.590 1200.000 ;
    END
  END eFPGA_operand_a_o[16]
  PIN eFPGA_operand_a_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 578.040 1200.000 578.640 ;
    END
  END eFPGA_operand_a_o[17]
  PIN eFPGA_operand_a_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END eFPGA_operand_a_o[18]
  PIN eFPGA_operand_a_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 650.800 1200.000 651.400 ;
    END
  END eFPGA_operand_a_o[19]
  PIN eFPGA_operand_a_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END eFPGA_operand_a_o[1]
  PIN eFPGA_operand_a_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 694.320 1200.000 694.920 ;
    END
  END eFPGA_operand_a_o[20]
  PIN eFPGA_operand_a_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 0.000 787.890 4.000 ;
    END
  END eFPGA_operand_a_o[21]
  PIN eFPGA_operand_a_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 1196.000 661.850 1200.000 ;
    END
  END eFPGA_operand_a_o[22]
  PIN eFPGA_operand_a_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 767.080 1200.000 767.680 ;
    END
  END eFPGA_operand_a_o[23]
  PIN eFPGA_operand_a_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END eFPGA_operand_a_o[24]
  PIN eFPGA_operand_a_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END eFPGA_operand_a_o[25]
  PIN eFPGA_operand_a_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 846.640 1200.000 847.240 ;
    END
  END eFPGA_operand_a_o[26]
  PIN eFPGA_operand_a_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 875.880 1200.000 876.480 ;
    END
  END eFPGA_operand_a_o[27]
  PIN eFPGA_operand_a_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 929.600 4.000 930.200 ;
    END
  END eFPGA_operand_a_o[28]
  PIN eFPGA_operand_a_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 1196.000 890.470 1200.000 ;
    END
  END eFPGA_operand_a_o[29]
  PIN eFPGA_operand_a_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 141.480 1200.000 142.080 ;
    END
  END eFPGA_operand_a_o[2]
  PIN eFPGA_operand_a_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 1196.000 909.790 1200.000 ;
    END
  END eFPGA_operand_a_o[30]
  PIN eFPGA_operand_a_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 992.160 1200.000 992.760 ;
    END
  END eFPGA_operand_a_o[31]
  PIN eFPGA_operand_a_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 1196.000 147.570 1200.000 ;
    END
  END eFPGA_operand_a_o[3]
  PIN eFPGA_operand_a_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END eFPGA_operand_a_o[4]
  PIN eFPGA_operand_a_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 243.480 1200.000 244.080 ;
    END
  END eFPGA_operand_a_o[5]
  PIN eFPGA_operand_a_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 287.000 1200.000 287.600 ;
    END
  END eFPGA_operand_a_o[6]
  PIN eFPGA_operand_a_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END eFPGA_operand_a_o[7]
  PIN eFPGA_operand_a_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END eFPGA_operand_a_o[8]
  PIN eFPGA_operand_a_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 1196.000 262.110 1200.000 ;
    END
  END eFPGA_operand_a_o[9]
  PIN eFPGA_operand_b_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 53.760 1200.000 54.360 ;
    END
  END eFPGA_operand_b_o[0]
  PIN eFPGA_operand_b_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END eFPGA_operand_b_o[10]
  PIN eFPGA_operand_b_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 4.000 503.160 ;
    END
  END eFPGA_operand_b_o[11]
  PIN eFPGA_operand_b_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END eFPGA_operand_b_o[12]
  PIN eFPGA_operand_b_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 483.520 1200.000 484.120 ;
    END
  END eFPGA_operand_b_o[13]
  PIN eFPGA_operand_b_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 505.280 1200.000 505.880 ;
    END
  END eFPGA_operand_b_o[14]
  PIN eFPGA_operand_b_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END eFPGA_operand_b_o[15]
  PIN eFPGA_operand_b_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END eFPGA_operand_b_o[16]
  PIN eFPGA_operand_b_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 584.840 1200.000 585.440 ;
    END
  END eFPGA_operand_b_o[17]
  PIN eFPGA_operand_b_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 621.560 1200.000 622.160 ;
    END
  END eFPGA_operand_b_o[18]
  PIN eFPGA_operand_b_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.000 4.000 712.600 ;
    END
  END eFPGA_operand_b_o[19]
  PIN eFPGA_operand_b_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END eFPGA_operand_b_o[1]
  PIN eFPGA_operand_b_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 728.320 4.000 728.920 ;
    END
  END eFPGA_operand_b_o[20]
  PIN eFPGA_operand_b_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END eFPGA_operand_b_o[21]
  PIN eFPGA_operand_b_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END eFPGA_operand_b_o[22]
  PIN eFPGA_operand_b_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END eFPGA_operand_b_o[23]
  PIN eFPGA_operand_b_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END eFPGA_operand_b_o[24]
  PIN eFPGA_operand_b_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END eFPGA_operand_b_o[25]
  PIN eFPGA_operand_b_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 854.120 1200.000 854.720 ;
    END
  END eFPGA_operand_b_o[26]
  PIN eFPGA_operand_b_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END eFPGA_operand_b_o[27]
  PIN eFPGA_operand_b_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 0.000 920.830 4.000 ;
    END
  END eFPGA_operand_b_o[28]
  PIN eFPGA_operand_b_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.850 0.000 946.130 4.000 ;
    END
  END eFPGA_operand_b_o[29]
  PIN eFPGA_operand_b_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 148.280 1200.000 148.880 ;
    END
  END eFPGA_operand_b_o[2]
  PIN eFPGA_operand_b_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 0.000 996.270 4.000 ;
    END
  END eFPGA_operand_b_o[30]
  PIN eFPGA_operand_b_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.680 4.000 1002.280 ;
    END
  END eFPGA_operand_b_o[31]
  PIN eFPGA_operand_b_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END eFPGA_operand_b_o[3]
  PIN eFPGA_operand_b_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 1196.000 185.750 1200.000 ;
    END
  END eFPGA_operand_b_o[4]
  PIN eFPGA_operand_b_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END eFPGA_operand_b_o[5]
  PIN eFPGA_operand_b_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 293.800 1200.000 294.400 ;
    END
  END eFPGA_operand_b_o[6]
  PIN eFPGA_operand_b_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 344.800 1200.000 345.400 ;
    END
  END eFPGA_operand_b_o[7]
  PIN eFPGA_operand_b_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END eFPGA_operand_b_o[8]
  PIN eFPGA_operand_b_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 1196.000 271.310 1200.000 ;
    END
  END eFPGA_operand_b_o[9]
  PIN eFPGA_operator_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 1196.000 62.010 1200.000 ;
    END
  END eFPGA_operator_o[0]
  PIN eFPGA_operator_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 75.520 1200.000 76.120 ;
    END
  END eFPGA_operator_o[1]
  PIN eFPGA_result_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END eFPGA_result_a_i[0]
  PIN eFPGA_result_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END eFPGA_result_a_i[10]
  PIN eFPGA_result_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.720 4.000 511.320 ;
    END
  END eFPGA_result_a_i[11]
  PIN eFPGA_result_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END eFPGA_result_a_i[12]
  PIN eFPGA_result_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 490.320 1200.000 490.920 ;
    END
  END eFPGA_result_a_i[13]
  PIN eFPGA_result_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END eFPGA_result_a_i[14]
  PIN eFPGA_result_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.280 4.000 607.880 ;
    END
  END eFPGA_result_a_i[15]
  PIN eFPGA_result_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 563.080 1200.000 563.680 ;
    END
  END eFPGA_result_a_i[16]
  PIN eFPGA_result_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 4.000 664.320 ;
    END
  END eFPGA_result_a_i[17]
  PIN eFPGA_result_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 1196.000 538.110 1200.000 ;
    END
  END eFPGA_result_a_i[18]
  PIN eFPGA_result_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END eFPGA_result_a_i[19]
  PIN eFPGA_result_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 83.000 1200.000 83.600 ;
    END
  END eFPGA_result_a_i[1]
  PIN eFPGA_result_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END eFPGA_result_a_i[20]
  PIN eFPGA_result_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 716.080 1200.000 716.680 ;
    END
  END eFPGA_result_a_i[21]
  PIN eFPGA_result_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END eFPGA_result_a_i[22]
  PIN eFPGA_result_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 1196.000 709.690 1200.000 ;
    END
  END eFPGA_result_a_i[23]
  PIN eFPGA_result_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 795.640 1200.000 796.240 ;
    END
  END eFPGA_result_a_i[24]
  PIN eFPGA_result_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END eFPGA_result_a_i[25]
  PIN eFPGA_result_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 1196.000 795.250 1200.000 ;
    END
  END eFPGA_result_a_i[26]
  PIN eFPGA_result_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 883.360 1200.000 883.960 ;
    END
  END eFPGA_result_a_i[27]
  PIN eFPGA_result_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.330 1196.000 871.610 1200.000 ;
    END
  END eFPGA_result_a_i[28]
  PIN eFPGA_result_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 941.160 1200.000 941.760 ;
    END
  END eFPGA_result_a_i[29]
  PIN eFPGA_result_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 155.760 1200.000 156.360 ;
    END
  END eFPGA_result_a_i[2]
  PIN eFPGA_result_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.270 0.000 1004.550 4.000 ;
    END
  END eFPGA_result_a_i[30]
  PIN eFPGA_result_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.370 1196.000 928.650 1200.000 ;
    END
  END eFPGA_result_a_i[31]
  PIN eFPGA_result_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END eFPGA_result_a_i[3]
  PIN eFPGA_result_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END eFPGA_result_a_i[4]
  PIN eFPGA_result_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END eFPGA_result_a_i[5]
  PIN eFPGA_result_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 1196.000 233.130 1200.000 ;
    END
  END eFPGA_result_a_i[6]
  PIN eFPGA_result_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END eFPGA_result_a_i[7]
  PIN eFPGA_result_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 381.520 1200.000 382.120 ;
    END
  END eFPGA_result_a_i[8]
  PIN eFPGA_result_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END eFPGA_result_a_i[9]
  PIN eFPGA_result_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END eFPGA_result_b_i[0]
  PIN eFPGA_result_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 1196.000 290.630 1200.000 ;
    END
  END eFPGA_result_b_i[10]
  PIN eFPGA_result_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 1196.000 347.670 1200.000 ;
    END
  END eFPGA_result_b_i[11]
  PIN eFPGA_result_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 1196.000 385.850 1200.000 ;
    END
  END eFPGA_result_b_i[12]
  PIN eFPGA_result_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 1196.000 433.230 1200.000 ;
    END
  END eFPGA_result_b_i[13]
  PIN eFPGA_result_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 1196.000 452.550 1200.000 ;
    END
  END eFPGA_result_b_i[14]
  PIN eFPGA_result_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 541.320 1200.000 541.920 ;
    END
  END eFPGA_result_b_i[15]
  PIN eFPGA_result_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END eFPGA_result_b_i[16]
  PIN eFPGA_result_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END eFPGA_result_b_i[17]
  PIN eFPGA_result_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 1196.000 547.770 1200.000 ;
    END
  END eFPGA_result_b_i[18]
  PIN eFPGA_result_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 1196.000 576.290 1200.000 ;
    END
  END eFPGA_result_b_i[19]
  PIN eFPGA_result_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 90.480 1200.000 91.080 ;
    END
  END eFPGA_result_b_i[1]
  PIN eFPGA_result_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1196.000 604.810 1200.000 ;
    END
  END eFPGA_result_b_i[20]
  PIN eFPGA_result_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 1196.000 633.330 1200.000 ;
    END
  END eFPGA_result_b_i[21]
  PIN eFPGA_result_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 737.840 1200.000 738.440 ;
    END
  END eFPGA_result_b_i[22]
  PIN eFPGA_result_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 800.400 4.000 801.000 ;
    END
  END eFPGA_result_b_i[23]
  PIN eFPGA_result_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 803.120 1200.000 803.720 ;
    END
  END eFPGA_result_b_i[24]
  PIN eFPGA_result_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 824.880 1200.000 825.480 ;
    END
  END eFPGA_result_b_i[25]
  PIN eFPGA_result_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 1196.000 804.910 1200.000 ;
    END
  END eFPGA_result_b_i[26]
  PIN eFPGA_result_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 890.840 1200.000 891.440 ;
    END
  END eFPGA_result_b_i[27]
  PIN eFPGA_result_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.760 4.000 938.360 ;
    END
  END eFPGA_result_b_i[28]
  PIN eFPGA_result_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 0.000 954.410 4.000 ;
    END
  END eFPGA_result_b_i[29]
  PIN eFPGA_result_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 163.240 1200.000 163.840 ;
    END
  END eFPGA_result_b_i[2]
  PIN eFPGA_result_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END eFPGA_result_b_i[30]
  PIN eFPGA_result_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 1196.000 938.310 1200.000 ;
    END
  END eFPGA_result_b_i[31]
  PIN eFPGA_result_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 1196.000 157.230 1200.000 ;
    END
  END eFPGA_result_b_i[3]
  PIN eFPGA_result_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 1196.000 195.410 1200.000 ;
    END
  END eFPGA_result_b_i[4]
  PIN eFPGA_result_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END eFPGA_result_b_i[5]
  PIN eFPGA_result_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 301.280 1200.000 301.880 ;
    END
  END eFPGA_result_b_i[6]
  PIN eFPGA_result_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END eFPGA_result_b_i[7]
  PIN eFPGA_result_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.160 4.000 414.760 ;
    END
  END eFPGA_result_b_i[8]
  PIN eFPGA_result_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 1196.000 280.970 1200.000 ;
    END
  END eFPGA_result_b_i[9]
  PIN eFPGA_result_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END eFPGA_result_c_i[0]
  PIN eFPGA_result_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 425.040 1200.000 425.640 ;
    END
  END eFPGA_result_c_i[10]
  PIN eFPGA_result_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.880 4.000 519.480 ;
    END
  END eFPGA_result_c_i[11]
  PIN eFPGA_result_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 1196.000 395.050 1200.000 ;
    END
  END eFPGA_result_c_i[12]
  PIN eFPGA_result_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END eFPGA_result_c_i[13]
  PIN eFPGA_result_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END eFPGA_result_c_i[14]
  PIN eFPGA_result_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 548.800 1200.000 549.400 ;
    END
  END eFPGA_result_c_i[15]
  PIN eFPGA_result_c_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END eFPGA_result_c_i[16]
  PIN eFPGA_result_c_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 592.320 1200.000 592.920 ;
    END
  END eFPGA_result_c_i[17]
  PIN eFPGA_result_c_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END eFPGA_result_c_i[18]
  PIN eFPGA_result_c_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END eFPGA_result_c_i[19]
  PIN eFPGA_result_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END eFPGA_result_c_i[1]
  PIN eFPGA_result_c_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 701.120 1200.000 701.720 ;
    END
  END eFPGA_result_c_i[20]
  PIN eFPGA_result_c_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 723.560 1200.000 724.160 ;
    END
  END eFPGA_result_c_i[21]
  PIN eFPGA_result_c_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 1196.000 671.510 1200.000 ;
    END
  END eFPGA_result_c_i[22]
  PIN eFPGA_result_c_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 773.880 1200.000 774.480 ;
    END
  END eFPGA_result_c_i[23]
  PIN eFPGA_result_c_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.680 4.000 849.280 ;
    END
  END eFPGA_result_c_i[24]
  PIN eFPGA_result_c_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 889.480 4.000 890.080 ;
    END
  END eFPGA_result_c_i[25]
  PIN eFPGA_result_c_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 861.600 1200.000 862.200 ;
    END
  END eFPGA_result_c_i[26]
  PIN eFPGA_result_c_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 1196.000 823.770 1200.000 ;
    END
  END eFPGA_result_c_i[27]
  PIN eFPGA_result_c_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 912.600 1200.000 913.200 ;
    END
  END eFPGA_result_c_i[28]
  PIN eFPGA_result_c_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 0.000 962.690 4.000 ;
    END
  END eFPGA_result_c_i[29]
  PIN eFPGA_result_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 170.720 1200.000 171.320 ;
    END
  END eFPGA_result_c_i[2]
  PIN eFPGA_result_c_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 956.120 1200.000 956.720 ;
    END
  END eFPGA_result_c_i[30]
  PIN eFPGA_result_c_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END eFPGA_result_c_i[31]
  PIN eFPGA_result_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 192.480 1200.000 193.080 ;
    END
  END eFPGA_result_c_i[3]
  PIN eFPGA_result_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 214.240 1200.000 214.840 ;
    END
  END eFPGA_result_c_i[4]
  PIN eFPGA_result_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END eFPGA_result_c_i[5]
  PIN eFPGA_result_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END eFPGA_result_c_i[6]
  PIN eFPGA_result_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 352.280 1200.000 352.880 ;
    END
  END eFPGA_result_c_i[7]
  PIN eFPGA_result_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END eFPGA_result_c_i[8]
  PIN eFPGA_result_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END eFPGA_result_c_i[9]
  PIN eFPGA_write_strobe_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END eFPGA_write_strobe_o
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 1196.000 33.490 1200.000 ;
    END
  END fetch_enable_i
  PIN hart_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END hart_id_i[0]
  PIN hart_id_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1196.000 299.830 1200.000 ;
    END
  END hart_id_i[10]
  PIN hart_id_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 1196.000 357.330 1200.000 ;
    END
  END hart_id_i[11]
  PIN hart_id_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END hart_id_i[12]
  PIN hart_id_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END hart_id_i[13]
  PIN hart_id_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 512.080 1200.000 512.680 ;
    END
  END hart_id_i[14]
  PIN hart_id_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 555.600 1200.000 556.200 ;
    END
  END hart_id_i[15]
  PIN hart_id_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 1196.000 519.250 1200.000 ;
    END
  END hart_id_i[16]
  PIN hart_id_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 599.800 1200.000 600.400 ;
    END
  END hart_id_i[17]
  PIN hart_id_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END hart_id_i[18]
  PIN hart_id_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 657.600 1200.000 658.200 ;
    END
  END hart_id_i[19]
  PIN hart_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 97.960 1200.000 98.560 ;
    END
  END hart_id_i[1]
  PIN hart_id_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 0.000 746.030 4.000 ;
    END
  END hart_id_i[20]
  PIN hart_id_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END hart_id_i[21]
  PIN hart_id_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 745.320 1200.000 745.920 ;
    END
  END hart_id_i[22]
  PIN hart_id_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 808.560 4.000 809.160 ;
    END
  END hart_id_i[23]
  PIN hart_id_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END hart_id_i[24]
  PIN hart_id_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 832.360 1200.000 832.960 ;
    END
  END hart_id_i[25]
  PIN hart_id_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 868.400 1200.000 869.000 ;
    END
  END hart_id_i[26]
  PIN hart_id_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 0.000 904.270 4.000 ;
    END
  END hart_id_i[27]
  PIN hart_id_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END hart_id_i[28]
  PIN hart_id_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.690 0.000 970.970 4.000 ;
    END
  END hart_id_i[29]
  PIN hart_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 1196.000 119.050 1200.000 ;
    END
  END hart_id_i[2]
  PIN hart_id_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 963.600 1200.000 964.200 ;
    END
  END hart_id_i[30]
  PIN hart_id_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 999.640 1200.000 1000.240 ;
    END
  END hart_id_i[31]
  PIN hart_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END hart_id_i[3]
  PIN hart_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 1196.000 204.610 1200.000 ;
    END
  END hart_id_i[4]
  PIN hart_id_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END hart_id_i[5]
  PIN hart_id_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 308.760 1200.000 309.360 ;
    END
  END hart_id_i[6]
  PIN hart_id_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END hart_id_i[7]
  PIN hart_id_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END hart_id_i[8]
  PIN hart_id_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END hart_id_i[9]
  PIN instr_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END instr_addr_o[0]
  PIN instr_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 1196.000 309.490 1200.000 ;
    END
  END instr_addr_o[10]
  PIN instr_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 446.800 1200.000 447.400 ;
    END
  END instr_addr_o[11]
  PIN instr_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 1196.000 404.710 1200.000 ;
    END
  END instr_addr_o[12]
  PIN instr_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 0.000 587.790 4.000 ;
    END
  END instr_addr_o[13]
  PIN instr_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.800 4.000 583.400 ;
    END
  END instr_addr_o[14]
  PIN instr_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END instr_addr_o[15]
  PIN instr_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END instr_addr_o[16]
  PIN instr_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END instr_addr_o[17]
  PIN instr_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 1196.000 556.970 1200.000 ;
    END
  END instr_addr_o[18]
  PIN instr_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 665.080 1200.000 665.680 ;
    END
  END instr_addr_o[19]
  PIN instr_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END instr_addr_o[1]
  PIN instr_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END instr_addr_o[20]
  PIN instr_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 1196.000 642.990 1200.000 ;
    END
  END instr_addr_o[21]
  PIN instr_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 0.000 821.010 4.000 ;
    END
  END instr_addr_o[22]
  PIN instr_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 781.360 1200.000 781.960 ;
    END
  END instr_addr_o[23]
  PIN instr_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END instr_addr_o[24]
  PIN instr_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 0.000 854.590 4.000 ;
    END
  END instr_addr_o[25]
  PIN instr_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.120 4.000 905.720 ;
    END
  END instr_addr_o[26]
  PIN instr_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 897.640 1200.000 898.240 ;
    END
  END instr_addr_o[27]
  PIN instr_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END instr_addr_o[28]
  PIN instr_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1196.000 900.130 1200.000 ;
    END
  END instr_addr_o[29]
  PIN instr_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END instr_addr_o[2]
  PIN instr_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 0.000 1012.830 4.000 ;
    END
  END instr_addr_o[30]
  PIN instr_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.000 4.000 1018.600 ;
    END
  END instr_addr_o[31]
  PIN instr_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END instr_addr_o[3]
  PIN instr_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END instr_addr_o[4]
  PIN instr_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 250.280 1200.000 250.880 ;
    END
  END instr_addr_o[5]
  PIN instr_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END instr_addr_o[6]
  PIN instr_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END instr_addr_o[7]
  PIN instr_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END instr_addr_o[8]
  PIN instr_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END instr_addr_o[9]
  PIN instr_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 25.200 1200.000 25.800 ;
    END
  END instr_err_i
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 1196.000 42.690 1200.000 ;
    END
  END instr_gnt_i
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END instr_rdata_i[0]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 1196.000 319.150 1200.000 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 1196.000 366.530 1200.000 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 497.800 1200.000 498.400 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 519.560 1200.000 520.160 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 1196.000 471.410 1200.000 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 628.360 1200.000 628.960 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 104.760 1200.000 105.360 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 1196.000 614.470 1200.000 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 730.360 1200.000 730.960 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 1196.000 681.170 1200.000 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.720 4.000 817.320 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 1196.000 738.210 1200.000 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 1196.000 766.730 1200.000 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 1196.000 833.430 1200.000 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 919.400 1200.000 920.000 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 961.560 4.000 962.160 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 970.400 1200.000 971.000 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 1196.000 947.510 1200.000 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 1196.000 242.790 1200.000 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 359.760 1200.000 360.360 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 388.320 1200.000 388.920 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END instr_rdata_i[9]
  PIN instr_rdata_intg_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 61.240 1200.000 61.840 ;
    END
  END instr_rdata_intg_i[0]
  PIN instr_rdata_intg_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END instr_rdata_intg_i[1]
  PIN instr_rdata_intg_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END instr_rdata_intg_i[2]
  PIN instr_rdata_intg_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END instr_rdata_intg_i[3]
  PIN instr_rdata_intg_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END instr_rdata_intg_i[4]
  PIN instr_rdata_intg_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 257.760 1200.000 258.360 ;
    END
  END instr_rdata_intg_i[5]
  PIN instr_rdata_intg_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 315.560 1200.000 316.160 ;
    END
  END instr_rdata_intg_i[6]
  PIN instr_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END instr_req_o
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END instr_rvalid_i
  PIN irq_external_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END irq_external_i
  PIN irq_fast_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END irq_fast_i[0]
  PIN irq_fast_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END irq_fast_i[10]
  PIN irq_fast_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END irq_fast_i[11]
  PIN irq_fast_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END irq_fast_i[12]
  PIN irq_fast_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END irq_fast_i[13]
  PIN irq_fast_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END irq_fast_i[14]
  PIN irq_fast_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END irq_fast_i[1]
  PIN irq_fast_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END irq_fast_i[2]
  PIN irq_fast_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END irq_fast_i[3]
  PIN irq_fast_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END irq_fast_i[4]
  PIN irq_fast_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END irq_fast_i[5]
  PIN irq_fast_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END irq_fast_i[6]
  PIN irq_fast_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END irq_fast_i[7]
  PIN irq_fast_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END irq_fast_i[8]
  PIN irq_fast_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END irq_fast_i[9]
  PIN irq_nm_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END irq_nm_i
  PIN irq_software_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END irq_software_i
  PIN irq_timer_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END irq_timer_i
  PIN ram_cfg_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END ram_cfg_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END rst_ni
  PIN scan_rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 32.000 1200.000 32.600 ;
    END
  END scan_rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 39.480 1200.000 40.080 ;
    END
  END test_en_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 1188.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.040 10.640 147.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 10.640 247.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.040 10.640 297.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.040 10.640 347.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 10.640 397.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.040 10.640 447.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.040 10.640 497.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 10.640 547.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.040 10.640 597.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.040 10.640 647.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 10.640 697.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.040 10.640 747.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.040 10.640 797.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 10.640 847.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 896.040 10.640 897.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.040 10.640 947.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.040 10.640 997.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1046.040 10.640 1047.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.040 10.640 1097.640 1188.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.040 10.640 1147.640 1188.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 3.825 1195.855 1188.725 ;
      LAYER met1 ;
        RECT 0.070 3.780 1195.930 1189.620 ;
      LAYER met2 ;
        RECT 0.100 1195.720 4.410 1196.645 ;
        RECT 5.250 1195.720 13.610 1196.645 ;
        RECT 14.450 1195.720 23.270 1196.645 ;
        RECT 24.110 1195.720 32.930 1196.645 ;
        RECT 33.770 1195.720 42.130 1196.645 ;
        RECT 42.970 1195.720 51.790 1196.645 ;
        RECT 52.630 1195.720 61.450 1196.645 ;
        RECT 62.290 1195.720 70.650 1196.645 ;
        RECT 71.490 1195.720 80.310 1196.645 ;
        RECT 81.150 1195.720 89.970 1196.645 ;
        RECT 90.810 1195.720 99.630 1196.645 ;
        RECT 100.470 1195.720 108.830 1196.645 ;
        RECT 109.670 1195.720 118.490 1196.645 ;
        RECT 119.330 1195.720 128.150 1196.645 ;
        RECT 128.990 1195.720 137.350 1196.645 ;
        RECT 138.190 1195.720 147.010 1196.645 ;
        RECT 147.850 1195.720 156.670 1196.645 ;
        RECT 157.510 1195.720 166.330 1196.645 ;
        RECT 167.170 1195.720 175.530 1196.645 ;
        RECT 176.370 1195.720 185.190 1196.645 ;
        RECT 186.030 1195.720 194.850 1196.645 ;
        RECT 195.690 1195.720 204.050 1196.645 ;
        RECT 204.890 1195.720 213.710 1196.645 ;
        RECT 214.550 1195.720 223.370 1196.645 ;
        RECT 224.210 1195.720 232.570 1196.645 ;
        RECT 233.410 1195.720 242.230 1196.645 ;
        RECT 243.070 1195.720 251.890 1196.645 ;
        RECT 252.730 1195.720 261.550 1196.645 ;
        RECT 262.390 1195.720 270.750 1196.645 ;
        RECT 271.590 1195.720 280.410 1196.645 ;
        RECT 281.250 1195.720 290.070 1196.645 ;
        RECT 290.910 1195.720 299.270 1196.645 ;
        RECT 300.110 1195.720 308.930 1196.645 ;
        RECT 309.770 1195.720 318.590 1196.645 ;
        RECT 319.430 1195.720 328.250 1196.645 ;
        RECT 329.090 1195.720 337.450 1196.645 ;
        RECT 338.290 1195.720 347.110 1196.645 ;
        RECT 347.950 1195.720 356.770 1196.645 ;
        RECT 357.610 1195.720 365.970 1196.645 ;
        RECT 366.810 1195.720 375.630 1196.645 ;
        RECT 376.470 1195.720 385.290 1196.645 ;
        RECT 386.130 1195.720 394.490 1196.645 ;
        RECT 395.330 1195.720 404.150 1196.645 ;
        RECT 404.990 1195.720 413.810 1196.645 ;
        RECT 414.650 1195.720 423.470 1196.645 ;
        RECT 424.310 1195.720 432.670 1196.645 ;
        RECT 433.510 1195.720 442.330 1196.645 ;
        RECT 443.170 1195.720 451.990 1196.645 ;
        RECT 452.830 1195.720 461.190 1196.645 ;
        RECT 462.030 1195.720 470.850 1196.645 ;
        RECT 471.690 1195.720 480.510 1196.645 ;
        RECT 481.350 1195.720 490.170 1196.645 ;
        RECT 491.010 1195.720 499.370 1196.645 ;
        RECT 500.210 1195.720 509.030 1196.645 ;
        RECT 509.870 1195.720 518.690 1196.645 ;
        RECT 519.530 1195.720 527.890 1196.645 ;
        RECT 528.730 1195.720 537.550 1196.645 ;
        RECT 538.390 1195.720 547.210 1196.645 ;
        RECT 548.050 1195.720 556.410 1196.645 ;
        RECT 557.250 1195.720 566.070 1196.645 ;
        RECT 566.910 1195.720 575.730 1196.645 ;
        RECT 576.570 1195.720 585.390 1196.645 ;
        RECT 586.230 1195.720 594.590 1196.645 ;
        RECT 595.430 1195.720 604.250 1196.645 ;
        RECT 605.090 1195.720 613.910 1196.645 ;
        RECT 614.750 1195.720 623.110 1196.645 ;
        RECT 623.950 1195.720 632.770 1196.645 ;
        RECT 633.610 1195.720 642.430 1196.645 ;
        RECT 643.270 1195.720 652.090 1196.645 ;
        RECT 652.930 1195.720 661.290 1196.645 ;
        RECT 662.130 1195.720 670.950 1196.645 ;
        RECT 671.790 1195.720 680.610 1196.645 ;
        RECT 681.450 1195.720 689.810 1196.645 ;
        RECT 690.650 1195.720 699.470 1196.645 ;
        RECT 700.310 1195.720 709.130 1196.645 ;
        RECT 709.970 1195.720 718.330 1196.645 ;
        RECT 719.170 1195.720 727.990 1196.645 ;
        RECT 728.830 1195.720 737.650 1196.645 ;
        RECT 738.490 1195.720 747.310 1196.645 ;
        RECT 748.150 1195.720 756.510 1196.645 ;
        RECT 757.350 1195.720 766.170 1196.645 ;
        RECT 767.010 1195.720 775.830 1196.645 ;
        RECT 776.670 1195.720 785.030 1196.645 ;
        RECT 785.870 1195.720 794.690 1196.645 ;
        RECT 795.530 1195.720 804.350 1196.645 ;
        RECT 805.190 1195.720 814.010 1196.645 ;
        RECT 814.850 1195.720 823.210 1196.645 ;
        RECT 824.050 1195.720 832.870 1196.645 ;
        RECT 833.710 1195.720 842.530 1196.645 ;
        RECT 843.370 1195.720 851.730 1196.645 ;
        RECT 852.570 1195.720 861.390 1196.645 ;
        RECT 862.230 1195.720 871.050 1196.645 ;
        RECT 871.890 1195.720 880.250 1196.645 ;
        RECT 881.090 1195.720 889.910 1196.645 ;
        RECT 890.750 1195.720 899.570 1196.645 ;
        RECT 900.410 1195.720 909.230 1196.645 ;
        RECT 910.070 1195.720 918.430 1196.645 ;
        RECT 919.270 1195.720 928.090 1196.645 ;
        RECT 928.930 1195.720 937.750 1196.645 ;
        RECT 938.590 1195.720 946.950 1196.645 ;
        RECT 947.790 1195.720 956.610 1196.645 ;
        RECT 957.450 1195.720 966.270 1196.645 ;
        RECT 967.110 1195.720 975.930 1196.645 ;
        RECT 976.770 1195.720 985.130 1196.645 ;
        RECT 985.970 1195.720 994.790 1196.645 ;
        RECT 995.630 1195.720 1004.450 1196.645 ;
        RECT 1005.290 1195.720 1013.650 1196.645 ;
        RECT 1014.490 1195.720 1023.310 1196.645 ;
        RECT 1024.150 1195.720 1032.970 1196.645 ;
        RECT 1033.810 1195.720 1042.170 1196.645 ;
        RECT 1043.010 1195.720 1051.830 1196.645 ;
        RECT 1052.670 1195.720 1061.490 1196.645 ;
        RECT 1062.330 1195.720 1071.150 1196.645 ;
        RECT 1071.990 1195.720 1080.350 1196.645 ;
        RECT 1081.190 1195.720 1090.010 1196.645 ;
        RECT 1090.850 1195.720 1099.670 1196.645 ;
        RECT 1100.510 1195.720 1108.870 1196.645 ;
        RECT 1109.710 1195.720 1118.530 1196.645 ;
        RECT 1119.370 1195.720 1128.190 1196.645 ;
        RECT 1129.030 1195.720 1137.850 1196.645 ;
        RECT 1138.690 1195.720 1147.050 1196.645 ;
        RECT 1147.890 1195.720 1156.710 1196.645 ;
        RECT 1157.550 1195.720 1166.370 1196.645 ;
        RECT 1167.210 1195.720 1175.570 1196.645 ;
        RECT 1176.410 1195.720 1185.230 1196.645 ;
        RECT 1186.070 1195.720 1194.890 1196.645 ;
        RECT 1195.730 1195.720 1195.900 1196.645 ;
        RECT 0.100 4.280 1195.900 1195.720 ;
        RECT 0.100 3.555 3.950 4.280 ;
        RECT 4.790 3.555 12.230 4.280 ;
        RECT 13.070 3.555 20.510 4.280 ;
        RECT 21.350 3.555 28.790 4.280 ;
        RECT 29.630 3.555 37.070 4.280 ;
        RECT 37.910 3.555 45.350 4.280 ;
        RECT 46.190 3.555 53.630 4.280 ;
        RECT 54.470 3.555 61.910 4.280 ;
        RECT 62.750 3.555 70.190 4.280 ;
        RECT 71.030 3.555 78.930 4.280 ;
        RECT 79.770 3.555 87.210 4.280 ;
        RECT 88.050 3.555 95.490 4.280 ;
        RECT 96.330 3.555 103.770 4.280 ;
        RECT 104.610 3.555 112.050 4.280 ;
        RECT 112.890 3.555 120.330 4.280 ;
        RECT 121.170 3.555 128.610 4.280 ;
        RECT 129.450 3.555 136.890 4.280 ;
        RECT 137.730 3.555 145.630 4.280 ;
        RECT 146.470 3.555 153.910 4.280 ;
        RECT 154.750 3.555 162.190 4.280 ;
        RECT 163.030 3.555 170.470 4.280 ;
        RECT 171.310 3.555 178.750 4.280 ;
        RECT 179.590 3.555 187.030 4.280 ;
        RECT 187.870 3.555 195.310 4.280 ;
        RECT 196.150 3.555 203.590 4.280 ;
        RECT 204.430 3.555 211.870 4.280 ;
        RECT 212.710 3.555 220.610 4.280 ;
        RECT 221.450 3.555 228.890 4.280 ;
        RECT 229.730 3.555 237.170 4.280 ;
        RECT 238.010 3.555 245.450 4.280 ;
        RECT 246.290 3.555 253.730 4.280 ;
        RECT 254.570 3.555 262.010 4.280 ;
        RECT 262.850 3.555 270.290 4.280 ;
        RECT 271.130 3.555 278.570 4.280 ;
        RECT 279.410 3.555 287.310 4.280 ;
        RECT 288.150 3.555 295.590 4.280 ;
        RECT 296.430 3.555 303.870 4.280 ;
        RECT 304.710 3.555 312.150 4.280 ;
        RECT 312.990 3.555 320.430 4.280 ;
        RECT 321.270 3.555 328.710 4.280 ;
        RECT 329.550 3.555 336.990 4.280 ;
        RECT 337.830 3.555 345.270 4.280 ;
        RECT 346.110 3.555 353.550 4.280 ;
        RECT 354.390 3.555 362.290 4.280 ;
        RECT 363.130 3.555 370.570 4.280 ;
        RECT 371.410 3.555 378.850 4.280 ;
        RECT 379.690 3.555 387.130 4.280 ;
        RECT 387.970 3.555 395.410 4.280 ;
        RECT 396.250 3.555 403.690 4.280 ;
        RECT 404.530 3.555 411.970 4.280 ;
        RECT 412.810 3.555 420.250 4.280 ;
        RECT 421.090 3.555 428.990 4.280 ;
        RECT 429.830 3.555 437.270 4.280 ;
        RECT 438.110 3.555 445.550 4.280 ;
        RECT 446.390 3.555 453.830 4.280 ;
        RECT 454.670 3.555 462.110 4.280 ;
        RECT 462.950 3.555 470.390 4.280 ;
        RECT 471.230 3.555 478.670 4.280 ;
        RECT 479.510 3.555 486.950 4.280 ;
        RECT 487.790 3.555 495.230 4.280 ;
        RECT 496.070 3.555 503.970 4.280 ;
        RECT 504.810 3.555 512.250 4.280 ;
        RECT 513.090 3.555 520.530 4.280 ;
        RECT 521.370 3.555 528.810 4.280 ;
        RECT 529.650 3.555 537.090 4.280 ;
        RECT 537.930 3.555 545.370 4.280 ;
        RECT 546.210 3.555 553.650 4.280 ;
        RECT 554.490 3.555 561.930 4.280 ;
        RECT 562.770 3.555 570.670 4.280 ;
        RECT 571.510 3.555 578.950 4.280 ;
        RECT 579.790 3.555 587.230 4.280 ;
        RECT 588.070 3.555 595.510 4.280 ;
        RECT 596.350 3.555 603.790 4.280 ;
        RECT 604.630 3.555 612.070 4.280 ;
        RECT 612.910 3.555 620.350 4.280 ;
        RECT 621.190 3.555 628.630 4.280 ;
        RECT 629.470 3.555 636.910 4.280 ;
        RECT 637.750 3.555 645.650 4.280 ;
        RECT 646.490 3.555 653.930 4.280 ;
        RECT 654.770 3.555 662.210 4.280 ;
        RECT 663.050 3.555 670.490 4.280 ;
        RECT 671.330 3.555 678.770 4.280 ;
        RECT 679.610 3.555 687.050 4.280 ;
        RECT 687.890 3.555 695.330 4.280 ;
        RECT 696.170 3.555 703.610 4.280 ;
        RECT 704.450 3.555 712.350 4.280 ;
        RECT 713.190 3.555 720.630 4.280 ;
        RECT 721.470 3.555 728.910 4.280 ;
        RECT 729.750 3.555 737.190 4.280 ;
        RECT 738.030 3.555 745.470 4.280 ;
        RECT 746.310 3.555 753.750 4.280 ;
        RECT 754.590 3.555 762.030 4.280 ;
        RECT 762.870 3.555 770.310 4.280 ;
        RECT 771.150 3.555 778.590 4.280 ;
        RECT 779.430 3.555 787.330 4.280 ;
        RECT 788.170 3.555 795.610 4.280 ;
        RECT 796.450 3.555 803.890 4.280 ;
        RECT 804.730 3.555 812.170 4.280 ;
        RECT 813.010 3.555 820.450 4.280 ;
        RECT 821.290 3.555 828.730 4.280 ;
        RECT 829.570 3.555 837.010 4.280 ;
        RECT 837.850 3.555 845.290 4.280 ;
        RECT 846.130 3.555 854.030 4.280 ;
        RECT 854.870 3.555 862.310 4.280 ;
        RECT 863.150 3.555 870.590 4.280 ;
        RECT 871.430 3.555 878.870 4.280 ;
        RECT 879.710 3.555 887.150 4.280 ;
        RECT 887.990 3.555 895.430 4.280 ;
        RECT 896.270 3.555 903.710 4.280 ;
        RECT 904.550 3.555 911.990 4.280 ;
        RECT 912.830 3.555 920.270 4.280 ;
        RECT 921.110 3.555 929.010 4.280 ;
        RECT 929.850 3.555 937.290 4.280 ;
        RECT 938.130 3.555 945.570 4.280 ;
        RECT 946.410 3.555 953.850 4.280 ;
        RECT 954.690 3.555 962.130 4.280 ;
        RECT 962.970 3.555 970.410 4.280 ;
        RECT 971.250 3.555 978.690 4.280 ;
        RECT 979.530 3.555 986.970 4.280 ;
        RECT 987.810 3.555 995.710 4.280 ;
        RECT 996.550 3.555 1003.990 4.280 ;
        RECT 1004.830 3.555 1012.270 4.280 ;
        RECT 1013.110 3.555 1020.550 4.280 ;
        RECT 1021.390 3.555 1028.830 4.280 ;
        RECT 1029.670 3.555 1037.110 4.280 ;
        RECT 1037.950 3.555 1045.390 4.280 ;
        RECT 1046.230 3.555 1053.670 4.280 ;
        RECT 1054.510 3.555 1061.950 4.280 ;
        RECT 1062.790 3.555 1070.690 4.280 ;
        RECT 1071.530 3.555 1078.970 4.280 ;
        RECT 1079.810 3.555 1087.250 4.280 ;
        RECT 1088.090 3.555 1095.530 4.280 ;
        RECT 1096.370 3.555 1103.810 4.280 ;
        RECT 1104.650 3.555 1112.090 4.280 ;
        RECT 1112.930 3.555 1120.370 4.280 ;
        RECT 1121.210 3.555 1128.650 4.280 ;
        RECT 1129.490 3.555 1137.390 4.280 ;
        RECT 1138.230 3.555 1145.670 4.280 ;
        RECT 1146.510 3.555 1153.950 4.280 ;
        RECT 1154.790 3.555 1162.230 4.280 ;
        RECT 1163.070 3.555 1170.510 4.280 ;
        RECT 1171.350 3.555 1178.790 4.280 ;
        RECT 1179.630 3.555 1187.070 4.280 ;
        RECT 1187.910 3.555 1195.350 4.280 ;
      LAYER met3 ;
        RECT 0.525 1196.480 1195.600 1196.625 ;
        RECT 4.400 1195.760 1195.600 1196.480 ;
        RECT 4.400 1195.080 1196.610 1195.760 ;
        RECT 0.525 1189.680 1196.610 1195.080 ;
        RECT 0.525 1188.320 1195.600 1189.680 ;
        RECT 4.400 1188.280 1195.600 1188.320 ;
        RECT 4.400 1186.920 1196.610 1188.280 ;
        RECT 0.525 1182.200 1196.610 1186.920 ;
        RECT 0.525 1180.800 1195.600 1182.200 ;
        RECT 0.525 1180.160 1196.610 1180.800 ;
        RECT 4.400 1178.760 1196.610 1180.160 ;
        RECT 0.525 1175.400 1196.610 1178.760 ;
        RECT 0.525 1174.000 1195.600 1175.400 ;
        RECT 0.525 1172.000 1196.610 1174.000 ;
        RECT 4.400 1170.600 1196.610 1172.000 ;
        RECT 0.525 1167.920 1196.610 1170.600 ;
        RECT 0.525 1166.520 1195.600 1167.920 ;
        RECT 0.525 1163.840 1196.610 1166.520 ;
        RECT 4.400 1162.440 1196.610 1163.840 ;
        RECT 0.525 1160.440 1196.610 1162.440 ;
        RECT 0.525 1159.040 1195.600 1160.440 ;
        RECT 0.525 1155.680 1196.610 1159.040 ;
        RECT 4.400 1154.280 1196.610 1155.680 ;
        RECT 0.525 1153.640 1196.610 1154.280 ;
        RECT 0.525 1152.240 1195.600 1153.640 ;
        RECT 0.525 1148.200 1196.610 1152.240 ;
        RECT 4.400 1146.800 1196.610 1148.200 ;
        RECT 0.525 1146.160 1196.610 1146.800 ;
        RECT 0.525 1144.760 1195.600 1146.160 ;
        RECT 0.525 1140.040 1196.610 1144.760 ;
        RECT 4.400 1138.680 1196.610 1140.040 ;
        RECT 4.400 1138.640 1195.600 1138.680 ;
        RECT 0.525 1137.280 1195.600 1138.640 ;
        RECT 0.525 1131.880 1196.610 1137.280 ;
        RECT 4.400 1130.480 1195.600 1131.880 ;
        RECT 0.525 1124.400 1196.610 1130.480 ;
        RECT 0.525 1123.720 1195.600 1124.400 ;
        RECT 4.400 1123.000 1195.600 1123.720 ;
        RECT 4.400 1122.320 1196.610 1123.000 ;
        RECT 0.525 1116.920 1196.610 1122.320 ;
        RECT 0.525 1115.560 1195.600 1116.920 ;
        RECT 4.400 1115.520 1195.600 1115.560 ;
        RECT 4.400 1114.160 1196.610 1115.520 ;
        RECT 0.525 1109.440 1196.610 1114.160 ;
        RECT 0.525 1108.040 1195.600 1109.440 ;
        RECT 0.525 1107.400 1196.610 1108.040 ;
        RECT 4.400 1106.000 1196.610 1107.400 ;
        RECT 0.525 1102.640 1196.610 1106.000 ;
        RECT 0.525 1101.240 1195.600 1102.640 ;
        RECT 0.525 1099.920 1196.610 1101.240 ;
        RECT 4.400 1098.520 1196.610 1099.920 ;
        RECT 0.525 1095.160 1196.610 1098.520 ;
        RECT 0.525 1093.760 1195.600 1095.160 ;
        RECT 0.525 1091.760 1196.610 1093.760 ;
        RECT 4.400 1090.360 1196.610 1091.760 ;
        RECT 0.525 1087.680 1196.610 1090.360 ;
        RECT 0.525 1086.280 1195.600 1087.680 ;
        RECT 0.525 1083.600 1196.610 1086.280 ;
        RECT 4.400 1082.200 1196.610 1083.600 ;
        RECT 0.525 1080.880 1196.610 1082.200 ;
        RECT 0.525 1079.480 1195.600 1080.880 ;
        RECT 0.525 1075.440 1196.610 1079.480 ;
        RECT 4.400 1074.040 1196.610 1075.440 ;
        RECT 0.525 1073.400 1196.610 1074.040 ;
        RECT 0.525 1072.000 1195.600 1073.400 ;
        RECT 0.525 1067.280 1196.610 1072.000 ;
        RECT 4.400 1065.920 1196.610 1067.280 ;
        RECT 4.400 1065.880 1195.600 1065.920 ;
        RECT 0.525 1064.520 1195.600 1065.880 ;
        RECT 0.525 1059.120 1196.610 1064.520 ;
        RECT 4.400 1057.720 1195.600 1059.120 ;
        RECT 0.525 1051.640 1196.610 1057.720 ;
        RECT 0.525 1050.960 1195.600 1051.640 ;
        RECT 4.400 1050.240 1195.600 1050.960 ;
        RECT 4.400 1049.560 1196.610 1050.240 ;
        RECT 0.525 1044.160 1196.610 1049.560 ;
        RECT 0.525 1043.480 1195.600 1044.160 ;
        RECT 4.400 1042.760 1195.600 1043.480 ;
        RECT 4.400 1042.080 1196.610 1042.760 ;
        RECT 0.525 1036.680 1196.610 1042.080 ;
        RECT 0.525 1035.320 1195.600 1036.680 ;
        RECT 4.400 1035.280 1195.600 1035.320 ;
        RECT 4.400 1033.920 1196.610 1035.280 ;
        RECT 0.525 1029.880 1196.610 1033.920 ;
        RECT 0.525 1028.480 1195.600 1029.880 ;
        RECT 0.525 1027.160 1196.610 1028.480 ;
        RECT 4.400 1025.760 1196.610 1027.160 ;
        RECT 0.525 1022.400 1196.610 1025.760 ;
        RECT 0.525 1021.000 1195.600 1022.400 ;
        RECT 0.525 1019.000 1196.610 1021.000 ;
        RECT 4.400 1017.600 1196.610 1019.000 ;
        RECT 0.525 1014.920 1196.610 1017.600 ;
        RECT 0.525 1013.520 1195.600 1014.920 ;
        RECT 0.525 1010.840 1196.610 1013.520 ;
        RECT 4.400 1009.440 1196.610 1010.840 ;
        RECT 0.525 1008.120 1196.610 1009.440 ;
        RECT 0.525 1006.720 1195.600 1008.120 ;
        RECT 0.525 1002.680 1196.610 1006.720 ;
        RECT 4.400 1001.280 1196.610 1002.680 ;
        RECT 0.525 1000.640 1196.610 1001.280 ;
        RECT 0.525 999.240 1195.600 1000.640 ;
        RECT 0.525 995.200 1196.610 999.240 ;
        RECT 4.400 993.800 1196.610 995.200 ;
        RECT 0.525 993.160 1196.610 993.800 ;
        RECT 0.525 991.760 1195.600 993.160 ;
        RECT 0.525 987.040 1196.610 991.760 ;
        RECT 4.400 986.360 1196.610 987.040 ;
        RECT 4.400 985.640 1195.600 986.360 ;
        RECT 0.525 984.960 1195.600 985.640 ;
        RECT 0.525 978.880 1196.610 984.960 ;
        RECT 4.400 977.480 1195.600 978.880 ;
        RECT 0.525 971.400 1196.610 977.480 ;
        RECT 0.525 970.720 1195.600 971.400 ;
        RECT 4.400 970.000 1195.600 970.720 ;
        RECT 4.400 969.320 1196.610 970.000 ;
        RECT 0.525 964.600 1196.610 969.320 ;
        RECT 0.525 963.200 1195.600 964.600 ;
        RECT 0.525 962.560 1196.610 963.200 ;
        RECT 4.400 961.160 1196.610 962.560 ;
        RECT 0.525 957.120 1196.610 961.160 ;
        RECT 0.525 955.720 1195.600 957.120 ;
        RECT 0.525 954.400 1196.610 955.720 ;
        RECT 4.400 953.000 1196.610 954.400 ;
        RECT 0.525 949.640 1196.610 953.000 ;
        RECT 0.525 948.240 1195.600 949.640 ;
        RECT 0.525 946.240 1196.610 948.240 ;
        RECT 4.400 944.840 1196.610 946.240 ;
        RECT 0.525 942.160 1196.610 944.840 ;
        RECT 0.525 940.760 1195.600 942.160 ;
        RECT 0.525 938.760 1196.610 940.760 ;
        RECT 4.400 937.360 1196.610 938.760 ;
        RECT 0.525 935.360 1196.610 937.360 ;
        RECT 0.525 933.960 1195.600 935.360 ;
        RECT 0.525 930.600 1196.610 933.960 ;
        RECT 4.400 929.200 1196.610 930.600 ;
        RECT 0.525 927.880 1196.610 929.200 ;
        RECT 0.525 926.480 1195.600 927.880 ;
        RECT 0.525 922.440 1196.610 926.480 ;
        RECT 4.400 921.040 1196.610 922.440 ;
        RECT 0.525 920.400 1196.610 921.040 ;
        RECT 0.525 919.000 1195.600 920.400 ;
        RECT 0.525 914.280 1196.610 919.000 ;
        RECT 4.400 913.600 1196.610 914.280 ;
        RECT 4.400 912.880 1195.600 913.600 ;
        RECT 0.525 912.200 1195.600 912.880 ;
        RECT 0.525 906.120 1196.610 912.200 ;
        RECT 4.400 904.720 1195.600 906.120 ;
        RECT 0.525 898.640 1196.610 904.720 ;
        RECT 0.525 897.960 1195.600 898.640 ;
        RECT 4.400 897.240 1195.600 897.960 ;
        RECT 4.400 896.560 1196.610 897.240 ;
        RECT 0.525 891.840 1196.610 896.560 ;
        RECT 0.525 890.480 1195.600 891.840 ;
        RECT 4.400 890.440 1195.600 890.480 ;
        RECT 4.400 889.080 1196.610 890.440 ;
        RECT 0.525 884.360 1196.610 889.080 ;
        RECT 0.525 882.960 1195.600 884.360 ;
        RECT 0.525 882.320 1196.610 882.960 ;
        RECT 4.400 880.920 1196.610 882.320 ;
        RECT 0.525 876.880 1196.610 880.920 ;
        RECT 0.525 875.480 1195.600 876.880 ;
        RECT 0.525 874.160 1196.610 875.480 ;
        RECT 4.400 872.760 1196.610 874.160 ;
        RECT 0.525 869.400 1196.610 872.760 ;
        RECT 0.525 868.000 1195.600 869.400 ;
        RECT 0.525 866.000 1196.610 868.000 ;
        RECT 4.400 864.600 1196.610 866.000 ;
        RECT 0.525 862.600 1196.610 864.600 ;
        RECT 0.525 861.200 1195.600 862.600 ;
        RECT 0.525 857.840 1196.610 861.200 ;
        RECT 4.400 856.440 1196.610 857.840 ;
        RECT 0.525 855.120 1196.610 856.440 ;
        RECT 0.525 853.720 1195.600 855.120 ;
        RECT 0.525 849.680 1196.610 853.720 ;
        RECT 4.400 848.280 1196.610 849.680 ;
        RECT 0.525 847.640 1196.610 848.280 ;
        RECT 0.525 846.240 1195.600 847.640 ;
        RECT 0.525 841.520 1196.610 846.240 ;
        RECT 4.400 840.840 1196.610 841.520 ;
        RECT 4.400 840.120 1195.600 840.840 ;
        RECT 0.525 839.440 1195.600 840.120 ;
        RECT 0.525 834.040 1196.610 839.440 ;
        RECT 4.400 833.360 1196.610 834.040 ;
        RECT 4.400 832.640 1195.600 833.360 ;
        RECT 0.525 831.960 1195.600 832.640 ;
        RECT 0.525 825.880 1196.610 831.960 ;
        RECT 4.400 824.480 1195.600 825.880 ;
        RECT 0.525 819.080 1196.610 824.480 ;
        RECT 0.525 817.720 1195.600 819.080 ;
        RECT 4.400 817.680 1195.600 817.720 ;
        RECT 4.400 816.320 1196.610 817.680 ;
        RECT 0.525 811.600 1196.610 816.320 ;
        RECT 0.525 810.200 1195.600 811.600 ;
        RECT 0.525 809.560 1196.610 810.200 ;
        RECT 4.400 808.160 1196.610 809.560 ;
        RECT 0.525 804.120 1196.610 808.160 ;
        RECT 0.525 802.720 1195.600 804.120 ;
        RECT 0.525 801.400 1196.610 802.720 ;
        RECT 4.400 800.000 1196.610 801.400 ;
        RECT 0.525 796.640 1196.610 800.000 ;
        RECT 0.525 795.240 1195.600 796.640 ;
        RECT 0.525 793.240 1196.610 795.240 ;
        RECT 4.400 791.840 1196.610 793.240 ;
        RECT 0.525 789.840 1196.610 791.840 ;
        RECT 0.525 788.440 1195.600 789.840 ;
        RECT 0.525 785.760 1196.610 788.440 ;
        RECT 4.400 784.360 1196.610 785.760 ;
        RECT 0.525 782.360 1196.610 784.360 ;
        RECT 0.525 780.960 1195.600 782.360 ;
        RECT 0.525 777.600 1196.610 780.960 ;
        RECT 4.400 776.200 1196.610 777.600 ;
        RECT 0.525 774.880 1196.610 776.200 ;
        RECT 0.525 773.480 1195.600 774.880 ;
        RECT 0.525 769.440 1196.610 773.480 ;
        RECT 4.400 768.080 1196.610 769.440 ;
        RECT 4.400 768.040 1195.600 768.080 ;
        RECT 0.525 766.680 1195.600 768.040 ;
        RECT 0.525 761.280 1196.610 766.680 ;
        RECT 4.400 760.600 1196.610 761.280 ;
        RECT 4.400 759.880 1195.600 760.600 ;
        RECT 0.525 759.200 1195.600 759.880 ;
        RECT 0.525 753.120 1196.610 759.200 ;
        RECT 4.400 751.720 1195.600 753.120 ;
        RECT 0.525 746.320 1196.610 751.720 ;
        RECT 0.525 744.960 1195.600 746.320 ;
        RECT 4.400 744.920 1195.600 744.960 ;
        RECT 4.400 743.560 1196.610 744.920 ;
        RECT 0.525 738.840 1196.610 743.560 ;
        RECT 0.525 737.440 1195.600 738.840 ;
        RECT 0.525 736.800 1196.610 737.440 ;
        RECT 4.400 735.400 1196.610 736.800 ;
        RECT 0.525 731.360 1196.610 735.400 ;
        RECT 0.525 729.960 1195.600 731.360 ;
        RECT 0.525 729.320 1196.610 729.960 ;
        RECT 4.400 727.920 1196.610 729.320 ;
        RECT 0.525 724.560 1196.610 727.920 ;
        RECT 0.525 723.160 1195.600 724.560 ;
        RECT 0.525 721.160 1196.610 723.160 ;
        RECT 4.400 719.760 1196.610 721.160 ;
        RECT 0.525 717.080 1196.610 719.760 ;
        RECT 0.525 715.680 1195.600 717.080 ;
        RECT 0.525 713.000 1196.610 715.680 ;
        RECT 4.400 711.600 1196.610 713.000 ;
        RECT 0.525 709.600 1196.610 711.600 ;
        RECT 0.525 708.200 1195.600 709.600 ;
        RECT 0.525 704.840 1196.610 708.200 ;
        RECT 4.400 703.440 1196.610 704.840 ;
        RECT 0.525 702.120 1196.610 703.440 ;
        RECT 0.525 700.720 1195.600 702.120 ;
        RECT 0.525 696.680 1196.610 700.720 ;
        RECT 4.400 695.320 1196.610 696.680 ;
        RECT 4.400 695.280 1195.600 695.320 ;
        RECT 0.525 693.920 1195.600 695.280 ;
        RECT 0.525 688.520 1196.610 693.920 ;
        RECT 4.400 687.840 1196.610 688.520 ;
        RECT 4.400 687.120 1195.600 687.840 ;
        RECT 0.525 686.440 1195.600 687.120 ;
        RECT 0.525 681.040 1196.610 686.440 ;
        RECT 4.400 680.360 1196.610 681.040 ;
        RECT 4.400 679.640 1195.600 680.360 ;
        RECT 0.525 678.960 1195.600 679.640 ;
        RECT 0.525 673.560 1196.610 678.960 ;
        RECT 0.525 672.880 1195.600 673.560 ;
        RECT 4.400 672.160 1195.600 672.880 ;
        RECT 4.400 671.480 1196.610 672.160 ;
        RECT 0.525 666.080 1196.610 671.480 ;
        RECT 0.525 664.720 1195.600 666.080 ;
        RECT 4.400 664.680 1195.600 664.720 ;
        RECT 4.400 663.320 1196.610 664.680 ;
        RECT 0.525 658.600 1196.610 663.320 ;
        RECT 0.525 657.200 1195.600 658.600 ;
        RECT 0.525 656.560 1196.610 657.200 ;
        RECT 4.400 655.160 1196.610 656.560 ;
        RECT 0.525 651.800 1196.610 655.160 ;
        RECT 0.525 650.400 1195.600 651.800 ;
        RECT 0.525 648.400 1196.610 650.400 ;
        RECT 4.400 647.000 1196.610 648.400 ;
        RECT 0.525 644.320 1196.610 647.000 ;
        RECT 0.525 642.920 1195.600 644.320 ;
        RECT 0.525 640.240 1196.610 642.920 ;
        RECT 4.400 638.840 1196.610 640.240 ;
        RECT 0.525 636.840 1196.610 638.840 ;
        RECT 0.525 635.440 1195.600 636.840 ;
        RECT 0.525 632.080 1196.610 635.440 ;
        RECT 4.400 630.680 1196.610 632.080 ;
        RECT 0.525 629.360 1196.610 630.680 ;
        RECT 0.525 627.960 1195.600 629.360 ;
        RECT 0.525 624.600 1196.610 627.960 ;
        RECT 4.400 623.200 1196.610 624.600 ;
        RECT 0.525 622.560 1196.610 623.200 ;
        RECT 0.525 621.160 1195.600 622.560 ;
        RECT 0.525 616.440 1196.610 621.160 ;
        RECT 4.400 615.080 1196.610 616.440 ;
        RECT 4.400 615.040 1195.600 615.080 ;
        RECT 0.525 613.680 1195.600 615.040 ;
        RECT 0.525 608.280 1196.610 613.680 ;
        RECT 4.400 607.600 1196.610 608.280 ;
        RECT 4.400 606.880 1195.600 607.600 ;
        RECT 0.525 606.200 1195.600 606.880 ;
        RECT 0.525 600.800 1196.610 606.200 ;
        RECT 0.525 600.120 1195.600 600.800 ;
        RECT 4.400 599.400 1195.600 600.120 ;
        RECT 4.400 598.720 1196.610 599.400 ;
        RECT 0.525 593.320 1196.610 598.720 ;
        RECT 0.525 591.960 1195.600 593.320 ;
        RECT 4.400 591.920 1195.600 591.960 ;
        RECT 4.400 590.560 1196.610 591.920 ;
        RECT 0.525 585.840 1196.610 590.560 ;
        RECT 0.525 584.440 1195.600 585.840 ;
        RECT 0.525 583.800 1196.610 584.440 ;
        RECT 4.400 582.400 1196.610 583.800 ;
        RECT 0.525 579.040 1196.610 582.400 ;
        RECT 0.525 577.640 1195.600 579.040 ;
        RECT 0.525 576.320 1196.610 577.640 ;
        RECT 4.400 574.920 1196.610 576.320 ;
        RECT 0.525 571.560 1196.610 574.920 ;
        RECT 0.525 570.160 1195.600 571.560 ;
        RECT 0.525 568.160 1196.610 570.160 ;
        RECT 4.400 566.760 1196.610 568.160 ;
        RECT 0.525 564.080 1196.610 566.760 ;
        RECT 0.525 562.680 1195.600 564.080 ;
        RECT 0.525 560.000 1196.610 562.680 ;
        RECT 4.400 558.600 1196.610 560.000 ;
        RECT 0.525 556.600 1196.610 558.600 ;
        RECT 0.525 555.200 1195.600 556.600 ;
        RECT 0.525 551.840 1196.610 555.200 ;
        RECT 4.400 550.440 1196.610 551.840 ;
        RECT 0.525 549.800 1196.610 550.440 ;
        RECT 0.525 548.400 1195.600 549.800 ;
        RECT 0.525 543.680 1196.610 548.400 ;
        RECT 4.400 542.320 1196.610 543.680 ;
        RECT 4.400 542.280 1195.600 542.320 ;
        RECT 0.525 540.920 1195.600 542.280 ;
        RECT 0.525 535.520 1196.610 540.920 ;
        RECT 4.400 534.840 1196.610 535.520 ;
        RECT 4.400 534.120 1195.600 534.840 ;
        RECT 0.525 533.440 1195.600 534.120 ;
        RECT 0.525 528.040 1196.610 533.440 ;
        RECT 0.525 527.360 1195.600 528.040 ;
        RECT 4.400 526.640 1195.600 527.360 ;
        RECT 4.400 525.960 1196.610 526.640 ;
        RECT 0.525 520.560 1196.610 525.960 ;
        RECT 0.525 519.880 1195.600 520.560 ;
        RECT 4.400 519.160 1195.600 519.880 ;
        RECT 4.400 518.480 1196.610 519.160 ;
        RECT 0.525 513.080 1196.610 518.480 ;
        RECT 0.525 511.720 1195.600 513.080 ;
        RECT 4.400 511.680 1195.600 511.720 ;
        RECT 4.400 510.320 1196.610 511.680 ;
        RECT 0.525 506.280 1196.610 510.320 ;
        RECT 0.525 504.880 1195.600 506.280 ;
        RECT 0.525 503.560 1196.610 504.880 ;
        RECT 4.400 502.160 1196.610 503.560 ;
        RECT 0.525 498.800 1196.610 502.160 ;
        RECT 0.525 497.400 1195.600 498.800 ;
        RECT 0.525 495.400 1196.610 497.400 ;
        RECT 4.400 494.000 1196.610 495.400 ;
        RECT 0.525 491.320 1196.610 494.000 ;
        RECT 0.525 489.920 1195.600 491.320 ;
        RECT 0.525 487.240 1196.610 489.920 ;
        RECT 4.400 485.840 1196.610 487.240 ;
        RECT 0.525 484.520 1196.610 485.840 ;
        RECT 0.525 483.120 1195.600 484.520 ;
        RECT 0.525 479.080 1196.610 483.120 ;
        RECT 4.400 477.680 1196.610 479.080 ;
        RECT 0.525 477.040 1196.610 477.680 ;
        RECT 0.525 475.640 1195.600 477.040 ;
        RECT 0.525 471.600 1196.610 475.640 ;
        RECT 4.400 470.200 1196.610 471.600 ;
        RECT 0.525 469.560 1196.610 470.200 ;
        RECT 0.525 468.160 1195.600 469.560 ;
        RECT 0.525 463.440 1196.610 468.160 ;
        RECT 4.400 462.080 1196.610 463.440 ;
        RECT 4.400 462.040 1195.600 462.080 ;
        RECT 0.525 460.680 1195.600 462.040 ;
        RECT 0.525 455.280 1196.610 460.680 ;
        RECT 4.400 453.880 1195.600 455.280 ;
        RECT 0.525 447.800 1196.610 453.880 ;
        RECT 0.525 447.120 1195.600 447.800 ;
        RECT 4.400 446.400 1195.600 447.120 ;
        RECT 4.400 445.720 1196.610 446.400 ;
        RECT 0.525 440.320 1196.610 445.720 ;
        RECT 0.525 438.960 1195.600 440.320 ;
        RECT 4.400 438.920 1195.600 438.960 ;
        RECT 4.400 437.560 1196.610 438.920 ;
        RECT 0.525 433.520 1196.610 437.560 ;
        RECT 0.525 432.120 1195.600 433.520 ;
        RECT 0.525 430.800 1196.610 432.120 ;
        RECT 4.400 429.400 1196.610 430.800 ;
        RECT 0.525 426.040 1196.610 429.400 ;
        RECT 0.525 424.640 1195.600 426.040 ;
        RECT 0.525 422.640 1196.610 424.640 ;
        RECT 4.400 421.240 1196.610 422.640 ;
        RECT 0.525 418.560 1196.610 421.240 ;
        RECT 0.525 417.160 1195.600 418.560 ;
        RECT 0.525 415.160 1196.610 417.160 ;
        RECT 4.400 413.760 1196.610 415.160 ;
        RECT 0.525 411.760 1196.610 413.760 ;
        RECT 0.525 410.360 1195.600 411.760 ;
        RECT 0.525 407.000 1196.610 410.360 ;
        RECT 4.400 405.600 1196.610 407.000 ;
        RECT 0.525 404.280 1196.610 405.600 ;
        RECT 0.525 402.880 1195.600 404.280 ;
        RECT 0.525 398.840 1196.610 402.880 ;
        RECT 4.400 397.440 1196.610 398.840 ;
        RECT 0.525 396.800 1196.610 397.440 ;
        RECT 0.525 395.400 1195.600 396.800 ;
        RECT 0.525 390.680 1196.610 395.400 ;
        RECT 4.400 389.320 1196.610 390.680 ;
        RECT 4.400 389.280 1195.600 389.320 ;
        RECT 0.525 387.920 1195.600 389.280 ;
        RECT 0.525 382.520 1196.610 387.920 ;
        RECT 4.400 381.120 1195.600 382.520 ;
        RECT 0.525 375.040 1196.610 381.120 ;
        RECT 0.525 374.360 1195.600 375.040 ;
        RECT 4.400 373.640 1195.600 374.360 ;
        RECT 4.400 372.960 1196.610 373.640 ;
        RECT 0.525 367.560 1196.610 372.960 ;
        RECT 0.525 366.880 1195.600 367.560 ;
        RECT 4.400 366.160 1195.600 366.880 ;
        RECT 4.400 365.480 1196.610 366.160 ;
        RECT 0.525 360.760 1196.610 365.480 ;
        RECT 0.525 359.360 1195.600 360.760 ;
        RECT 0.525 358.720 1196.610 359.360 ;
        RECT 4.400 357.320 1196.610 358.720 ;
        RECT 0.525 353.280 1196.610 357.320 ;
        RECT 0.525 351.880 1195.600 353.280 ;
        RECT 0.525 350.560 1196.610 351.880 ;
        RECT 4.400 349.160 1196.610 350.560 ;
        RECT 0.525 345.800 1196.610 349.160 ;
        RECT 0.525 344.400 1195.600 345.800 ;
        RECT 0.525 342.400 1196.610 344.400 ;
        RECT 4.400 341.000 1196.610 342.400 ;
        RECT 0.525 339.000 1196.610 341.000 ;
        RECT 0.525 337.600 1195.600 339.000 ;
        RECT 0.525 334.240 1196.610 337.600 ;
        RECT 4.400 332.840 1196.610 334.240 ;
        RECT 0.525 331.520 1196.610 332.840 ;
        RECT 0.525 330.120 1195.600 331.520 ;
        RECT 0.525 326.080 1196.610 330.120 ;
        RECT 4.400 324.680 1196.610 326.080 ;
        RECT 0.525 324.040 1196.610 324.680 ;
        RECT 0.525 322.640 1195.600 324.040 ;
        RECT 0.525 317.920 1196.610 322.640 ;
        RECT 4.400 316.560 1196.610 317.920 ;
        RECT 4.400 316.520 1195.600 316.560 ;
        RECT 0.525 315.160 1195.600 316.520 ;
        RECT 0.525 310.440 1196.610 315.160 ;
        RECT 4.400 309.760 1196.610 310.440 ;
        RECT 4.400 309.040 1195.600 309.760 ;
        RECT 0.525 308.360 1195.600 309.040 ;
        RECT 0.525 302.280 1196.610 308.360 ;
        RECT 4.400 300.880 1195.600 302.280 ;
        RECT 0.525 294.800 1196.610 300.880 ;
        RECT 0.525 294.120 1195.600 294.800 ;
        RECT 4.400 293.400 1195.600 294.120 ;
        RECT 4.400 292.720 1196.610 293.400 ;
        RECT 0.525 288.000 1196.610 292.720 ;
        RECT 0.525 286.600 1195.600 288.000 ;
        RECT 0.525 285.960 1196.610 286.600 ;
        RECT 4.400 284.560 1196.610 285.960 ;
        RECT 0.525 280.520 1196.610 284.560 ;
        RECT 0.525 279.120 1195.600 280.520 ;
        RECT 0.525 277.800 1196.610 279.120 ;
        RECT 4.400 276.400 1196.610 277.800 ;
        RECT 0.525 273.040 1196.610 276.400 ;
        RECT 0.525 271.640 1195.600 273.040 ;
        RECT 0.525 269.640 1196.610 271.640 ;
        RECT 4.400 268.240 1196.610 269.640 ;
        RECT 0.525 266.240 1196.610 268.240 ;
        RECT 0.525 264.840 1195.600 266.240 ;
        RECT 0.525 262.160 1196.610 264.840 ;
        RECT 4.400 260.760 1196.610 262.160 ;
        RECT 0.525 258.760 1196.610 260.760 ;
        RECT 0.525 257.360 1195.600 258.760 ;
        RECT 0.525 254.000 1196.610 257.360 ;
        RECT 4.400 252.600 1196.610 254.000 ;
        RECT 0.525 251.280 1196.610 252.600 ;
        RECT 0.525 249.880 1195.600 251.280 ;
        RECT 0.525 245.840 1196.610 249.880 ;
        RECT 4.400 244.480 1196.610 245.840 ;
        RECT 4.400 244.440 1195.600 244.480 ;
        RECT 0.525 243.080 1195.600 244.440 ;
        RECT 0.525 237.680 1196.610 243.080 ;
        RECT 4.400 237.000 1196.610 237.680 ;
        RECT 4.400 236.280 1195.600 237.000 ;
        RECT 0.525 235.600 1195.600 236.280 ;
        RECT 0.525 229.520 1196.610 235.600 ;
        RECT 4.400 228.120 1195.600 229.520 ;
        RECT 0.525 222.040 1196.610 228.120 ;
        RECT 0.525 221.360 1195.600 222.040 ;
        RECT 4.400 220.640 1195.600 221.360 ;
        RECT 4.400 219.960 1196.610 220.640 ;
        RECT 0.525 215.240 1196.610 219.960 ;
        RECT 0.525 213.840 1195.600 215.240 ;
        RECT 0.525 213.200 1196.610 213.840 ;
        RECT 4.400 211.800 1196.610 213.200 ;
        RECT 0.525 207.760 1196.610 211.800 ;
        RECT 0.525 206.360 1195.600 207.760 ;
        RECT 0.525 205.720 1196.610 206.360 ;
        RECT 4.400 204.320 1196.610 205.720 ;
        RECT 0.525 200.280 1196.610 204.320 ;
        RECT 0.525 198.880 1195.600 200.280 ;
        RECT 0.525 197.560 1196.610 198.880 ;
        RECT 4.400 196.160 1196.610 197.560 ;
        RECT 0.525 193.480 1196.610 196.160 ;
        RECT 0.525 192.080 1195.600 193.480 ;
        RECT 0.525 189.400 1196.610 192.080 ;
        RECT 4.400 188.000 1196.610 189.400 ;
        RECT 0.525 186.000 1196.610 188.000 ;
        RECT 0.525 184.600 1195.600 186.000 ;
        RECT 0.525 181.240 1196.610 184.600 ;
        RECT 4.400 179.840 1196.610 181.240 ;
        RECT 0.525 178.520 1196.610 179.840 ;
        RECT 0.525 177.120 1195.600 178.520 ;
        RECT 0.525 173.080 1196.610 177.120 ;
        RECT 4.400 171.720 1196.610 173.080 ;
        RECT 4.400 171.680 1195.600 171.720 ;
        RECT 0.525 170.320 1195.600 171.680 ;
        RECT 0.525 164.920 1196.610 170.320 ;
        RECT 4.400 164.240 1196.610 164.920 ;
        RECT 4.400 163.520 1195.600 164.240 ;
        RECT 0.525 162.840 1195.600 163.520 ;
        RECT 0.525 157.440 1196.610 162.840 ;
        RECT 4.400 156.760 1196.610 157.440 ;
        RECT 4.400 156.040 1195.600 156.760 ;
        RECT 0.525 155.360 1195.600 156.040 ;
        RECT 0.525 149.280 1196.610 155.360 ;
        RECT 4.400 147.880 1195.600 149.280 ;
        RECT 0.525 142.480 1196.610 147.880 ;
        RECT 0.525 141.120 1195.600 142.480 ;
        RECT 4.400 141.080 1195.600 141.120 ;
        RECT 4.400 139.720 1196.610 141.080 ;
        RECT 0.525 135.000 1196.610 139.720 ;
        RECT 0.525 133.600 1195.600 135.000 ;
        RECT 0.525 132.960 1196.610 133.600 ;
        RECT 4.400 131.560 1196.610 132.960 ;
        RECT 0.525 127.520 1196.610 131.560 ;
        RECT 0.525 126.120 1195.600 127.520 ;
        RECT 0.525 124.800 1196.610 126.120 ;
        RECT 4.400 123.400 1196.610 124.800 ;
        RECT 0.525 120.720 1196.610 123.400 ;
        RECT 0.525 119.320 1195.600 120.720 ;
        RECT 0.525 116.640 1196.610 119.320 ;
        RECT 4.400 115.240 1196.610 116.640 ;
        RECT 0.525 113.240 1196.610 115.240 ;
        RECT 0.525 111.840 1195.600 113.240 ;
        RECT 0.525 108.480 1196.610 111.840 ;
        RECT 4.400 107.080 1196.610 108.480 ;
        RECT 0.525 105.760 1196.610 107.080 ;
        RECT 0.525 104.360 1195.600 105.760 ;
        RECT 0.525 101.000 1196.610 104.360 ;
        RECT 4.400 99.600 1196.610 101.000 ;
        RECT 0.525 98.960 1196.610 99.600 ;
        RECT 0.525 97.560 1195.600 98.960 ;
        RECT 0.525 92.840 1196.610 97.560 ;
        RECT 4.400 91.480 1196.610 92.840 ;
        RECT 4.400 91.440 1195.600 91.480 ;
        RECT 0.525 90.080 1195.600 91.440 ;
        RECT 0.525 84.680 1196.610 90.080 ;
        RECT 4.400 84.000 1196.610 84.680 ;
        RECT 4.400 83.280 1195.600 84.000 ;
        RECT 0.525 82.600 1195.600 83.280 ;
        RECT 0.525 76.520 1196.610 82.600 ;
        RECT 4.400 75.120 1195.600 76.520 ;
        RECT 0.525 69.720 1196.610 75.120 ;
        RECT 0.525 68.360 1195.600 69.720 ;
        RECT 4.400 68.320 1195.600 68.360 ;
        RECT 4.400 66.960 1196.610 68.320 ;
        RECT 0.525 62.240 1196.610 66.960 ;
        RECT 0.525 60.840 1195.600 62.240 ;
        RECT 0.525 60.200 1196.610 60.840 ;
        RECT 4.400 58.800 1196.610 60.200 ;
        RECT 0.525 54.760 1196.610 58.800 ;
        RECT 0.525 53.360 1195.600 54.760 ;
        RECT 0.525 52.720 1196.610 53.360 ;
        RECT 4.400 51.320 1196.610 52.720 ;
        RECT 0.525 47.960 1196.610 51.320 ;
        RECT 0.525 46.560 1195.600 47.960 ;
        RECT 0.525 44.560 1196.610 46.560 ;
        RECT 4.400 43.160 1196.610 44.560 ;
        RECT 0.525 40.480 1196.610 43.160 ;
        RECT 0.525 39.080 1195.600 40.480 ;
        RECT 0.525 36.400 1196.610 39.080 ;
        RECT 4.400 35.000 1196.610 36.400 ;
        RECT 0.525 33.000 1196.610 35.000 ;
        RECT 0.525 31.600 1195.600 33.000 ;
        RECT 0.525 28.240 1196.610 31.600 ;
        RECT 4.400 26.840 1196.610 28.240 ;
        RECT 0.525 26.200 1196.610 26.840 ;
        RECT 0.525 24.800 1195.600 26.200 ;
        RECT 0.525 20.080 1196.610 24.800 ;
        RECT 4.400 18.720 1196.610 20.080 ;
        RECT 4.400 18.680 1195.600 18.720 ;
        RECT 0.525 17.320 1195.600 18.680 ;
        RECT 0.525 11.920 1196.610 17.320 ;
        RECT 4.400 11.240 1196.610 11.920 ;
        RECT 4.400 10.520 1195.600 11.240 ;
        RECT 0.525 9.840 1195.600 10.520 ;
        RECT 0.525 4.440 1196.610 9.840 ;
        RECT 4.400 3.575 1195.600 4.440 ;
      LAYER met4 ;
        RECT 115.295 16.495 120.640 1176.905 ;
        RECT 123.040 16.495 145.640 1176.905 ;
        RECT 148.040 16.495 170.640 1176.905 ;
        RECT 173.040 16.495 195.640 1176.905 ;
        RECT 198.040 16.495 220.640 1176.905 ;
        RECT 223.040 16.495 245.640 1176.905 ;
        RECT 248.040 16.495 270.640 1176.905 ;
        RECT 273.040 16.495 295.640 1176.905 ;
        RECT 298.040 16.495 320.640 1176.905 ;
        RECT 323.040 16.495 345.640 1176.905 ;
        RECT 348.040 16.495 370.640 1176.905 ;
        RECT 373.040 16.495 395.640 1176.905 ;
        RECT 398.040 16.495 420.640 1176.905 ;
        RECT 423.040 16.495 445.640 1176.905 ;
        RECT 448.040 16.495 470.640 1176.905 ;
        RECT 473.040 16.495 495.640 1176.905 ;
        RECT 498.040 16.495 520.640 1176.905 ;
        RECT 523.040 16.495 545.640 1176.905 ;
        RECT 548.040 16.495 570.640 1176.905 ;
        RECT 573.040 16.495 595.640 1176.905 ;
        RECT 598.040 16.495 620.640 1176.905 ;
        RECT 623.040 16.495 645.640 1176.905 ;
        RECT 648.040 16.495 670.640 1176.905 ;
        RECT 673.040 16.495 695.640 1176.905 ;
        RECT 698.040 16.495 720.640 1176.905 ;
        RECT 723.040 16.495 745.640 1176.905 ;
        RECT 748.040 16.495 770.640 1176.905 ;
        RECT 773.040 16.495 795.640 1176.905 ;
        RECT 798.040 16.495 820.640 1176.905 ;
        RECT 823.040 16.495 845.640 1176.905 ;
        RECT 848.040 16.495 870.640 1176.905 ;
        RECT 873.040 16.495 895.640 1176.905 ;
        RECT 898.040 16.495 920.640 1176.905 ;
        RECT 923.040 16.495 945.640 1176.905 ;
        RECT 948.040 16.495 970.640 1176.905 ;
        RECT 973.040 16.495 995.640 1176.905 ;
        RECT 998.040 16.495 1019.065 1176.905 ;
  END
END ibex_top
END LIBRARY

