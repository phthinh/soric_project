VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO uart_to_mem
  CLASS BLOCK ;
  FOREIGN uart_to_mem ;
  ORIGIN 0.000 0.000 ;
  SIZE 152.725 BY 163.445 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END clk_i
  PIN data_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END data_addr_o[0]
  PIN data_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 159.445 69.830 163.445 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 52.400 152.725 53.000 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 159.445 62.930 163.445 ;
    END
  END data_addr_o[9]
  PIN data_be_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END data_be_o[0]
  PIN data_be_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 159.445 16.470 163.445 ;
    END
  END data_be_o[1]
  PIN data_be_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END data_be_o[2]
  PIN data_be_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 159.445 23.370 163.445 ;
    END
  END data_be_o[3]
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 159.445 3.590 163.445 ;
    END
  END data_gnt_i
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END data_rdata_i[0]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 80.960 152.725 81.560 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 91.160 152.725 91.760 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 159.445 83.170 163.445 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 159.445 102.950 163.445 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 110.200 152.725 110.800 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 159.445 129.630 163.445 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 129.240 152.725 129.840 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 148.280 152.725 148.880 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 157.800 152.725 158.400 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 159.445 29.810 163.445 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 42.880 152.725 43.480 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 159.445 36.710 163.445 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 159.445 50.050 163.445 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END data_rdata_i[9]
  PIN data_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END data_req_o
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 4.800 152.725 5.400 ;
    END
  END data_rvalid_i
  PIN data_wdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 14.320 152.725 14.920 ;
    END
  END data_wdata_o[0]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 61.920 152.725 62.520 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 71.440 152.725 72.040 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 159.445 76.270 163.445 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 100.680 152.725 101.280 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 159.445 89.610 163.445 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 159.445 96.510 163.445 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 159.445 109.390 163.445 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 159.445 116.290 163.445 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 159.445 122.730 163.445 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 119.720 152.725 120.320 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 159.445 136.070 163.445 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 138.760 152.725 139.360 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 159.445 142.970 163.445 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 23.840 152.725 24.440 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 159.445 149.410 163.445 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.725 33.360 152.725 33.960 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 159.445 43.150 163.445 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 159.445 56.490 163.445 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END data_wdata_o[9]
  PIN data_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 159.445 10.030 163.445 ;
    END
  END data_we_o
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END rst_i
  PIN rx_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END rx_i
  PIN tx_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END tx_o
  PIN uart_error
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END uart_error
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.335 10.640 29.935 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.560 10.640 77.160 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.785 10.640 124.385 152.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.945 10.640 53.545 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.170 10.640 100.770 152.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 147.975 152.405 ;
      LAYER met1 ;
        RECT 0.070 6.500 149.430 152.960 ;
      LAYER met2 ;
        RECT 0.100 159.165 3.030 160.325 ;
        RECT 3.870 159.165 9.470 160.325 ;
        RECT 10.310 159.165 15.910 160.325 ;
        RECT 16.750 159.165 22.810 160.325 ;
        RECT 23.650 159.165 29.250 160.325 ;
        RECT 30.090 159.165 36.150 160.325 ;
        RECT 36.990 159.165 42.590 160.325 ;
        RECT 43.430 159.165 49.490 160.325 ;
        RECT 50.330 159.165 55.930 160.325 ;
        RECT 56.770 159.165 62.370 160.325 ;
        RECT 63.210 159.165 69.270 160.325 ;
        RECT 70.110 159.165 75.710 160.325 ;
        RECT 76.550 159.165 82.610 160.325 ;
        RECT 83.450 159.165 89.050 160.325 ;
        RECT 89.890 159.165 95.950 160.325 ;
        RECT 96.790 159.165 102.390 160.325 ;
        RECT 103.230 159.165 108.830 160.325 ;
        RECT 109.670 159.165 115.730 160.325 ;
        RECT 116.570 159.165 122.170 160.325 ;
        RECT 123.010 159.165 129.070 160.325 ;
        RECT 129.910 159.165 135.510 160.325 ;
        RECT 136.350 159.165 142.410 160.325 ;
        RECT 143.250 159.165 148.850 160.325 ;
        RECT 0.100 4.280 149.400 159.165 ;
        RECT 0.100 3.555 2.570 4.280 ;
        RECT 3.410 3.555 8.550 4.280 ;
        RECT 9.390 3.555 14.530 4.280 ;
        RECT 15.370 3.555 20.510 4.280 ;
        RECT 21.350 3.555 26.950 4.280 ;
        RECT 27.790 3.555 32.930 4.280 ;
        RECT 33.770 3.555 38.910 4.280 ;
        RECT 39.750 3.555 44.890 4.280 ;
        RECT 45.730 3.555 51.330 4.280 ;
        RECT 52.170 3.555 57.310 4.280 ;
        RECT 58.150 3.555 63.290 4.280 ;
        RECT 64.130 3.555 69.730 4.280 ;
        RECT 70.570 3.555 75.710 4.280 ;
        RECT 76.550 3.555 81.690 4.280 ;
        RECT 82.530 3.555 87.670 4.280 ;
        RECT 88.510 3.555 94.110 4.280 ;
        RECT 94.950 3.555 100.090 4.280 ;
        RECT 100.930 3.555 106.070 4.280 ;
        RECT 106.910 3.555 112.510 4.280 ;
        RECT 113.350 3.555 118.490 4.280 ;
        RECT 119.330 3.555 124.470 4.280 ;
        RECT 125.310 3.555 130.450 4.280 ;
        RECT 131.290 3.555 136.890 4.280 ;
        RECT 137.730 3.555 142.870 4.280 ;
        RECT 143.710 3.555 148.850 4.280 ;
      LAYER met3 ;
        RECT 4.400 159.440 148.725 160.305 ;
        RECT 4.000 158.800 148.725 159.440 ;
        RECT 4.000 157.400 148.325 158.800 ;
        RECT 4.000 154.040 148.725 157.400 ;
        RECT 4.400 152.640 148.725 154.040 ;
        RECT 4.000 149.280 148.725 152.640 ;
        RECT 4.000 147.880 148.325 149.280 ;
        RECT 4.000 147.240 148.725 147.880 ;
        RECT 4.400 145.840 148.725 147.240 ;
        RECT 4.000 140.440 148.725 145.840 ;
        RECT 4.400 139.760 148.725 140.440 ;
        RECT 4.400 139.040 148.325 139.760 ;
        RECT 4.000 138.360 148.325 139.040 ;
        RECT 4.000 133.640 148.725 138.360 ;
        RECT 4.400 132.240 148.725 133.640 ;
        RECT 4.000 130.240 148.725 132.240 ;
        RECT 4.000 128.840 148.325 130.240 ;
        RECT 4.000 126.840 148.725 128.840 ;
        RECT 4.400 125.440 148.725 126.840 ;
        RECT 4.000 120.720 148.725 125.440 ;
        RECT 4.000 120.040 148.325 120.720 ;
        RECT 4.400 119.320 148.325 120.040 ;
        RECT 4.400 118.640 148.725 119.320 ;
        RECT 4.000 113.240 148.725 118.640 ;
        RECT 4.400 111.840 148.725 113.240 ;
        RECT 4.000 111.200 148.725 111.840 ;
        RECT 4.000 109.800 148.325 111.200 ;
        RECT 4.000 106.440 148.725 109.800 ;
        RECT 4.400 105.040 148.725 106.440 ;
        RECT 4.000 101.680 148.725 105.040 ;
        RECT 4.000 100.280 148.325 101.680 ;
        RECT 4.000 99.640 148.725 100.280 ;
        RECT 4.400 98.240 148.725 99.640 ;
        RECT 4.000 92.840 148.725 98.240 ;
        RECT 4.400 92.160 148.725 92.840 ;
        RECT 4.400 91.440 148.325 92.160 ;
        RECT 4.000 90.760 148.325 91.440 ;
        RECT 4.000 86.040 148.725 90.760 ;
        RECT 4.400 84.640 148.725 86.040 ;
        RECT 4.000 81.960 148.725 84.640 ;
        RECT 4.000 80.560 148.325 81.960 ;
        RECT 4.000 79.240 148.725 80.560 ;
        RECT 4.400 77.840 148.725 79.240 ;
        RECT 4.000 72.440 148.725 77.840 ;
        RECT 4.400 71.040 148.325 72.440 ;
        RECT 4.000 65.640 148.725 71.040 ;
        RECT 4.400 64.240 148.725 65.640 ;
        RECT 4.000 62.920 148.725 64.240 ;
        RECT 4.000 61.520 148.325 62.920 ;
        RECT 4.000 58.840 148.725 61.520 ;
        RECT 4.400 57.440 148.725 58.840 ;
        RECT 4.000 53.400 148.725 57.440 ;
        RECT 4.000 52.040 148.325 53.400 ;
        RECT 4.400 52.000 148.325 52.040 ;
        RECT 4.400 50.640 148.725 52.000 ;
        RECT 4.000 45.240 148.725 50.640 ;
        RECT 4.400 43.880 148.725 45.240 ;
        RECT 4.400 43.840 148.325 43.880 ;
        RECT 4.000 42.480 148.325 43.840 ;
        RECT 4.000 38.440 148.725 42.480 ;
        RECT 4.400 37.040 148.725 38.440 ;
        RECT 4.000 34.360 148.725 37.040 ;
        RECT 4.000 32.960 148.325 34.360 ;
        RECT 4.000 31.640 148.725 32.960 ;
        RECT 4.400 30.240 148.725 31.640 ;
        RECT 4.000 24.840 148.725 30.240 ;
        RECT 4.400 23.440 148.325 24.840 ;
        RECT 4.000 18.040 148.725 23.440 ;
        RECT 4.400 16.640 148.725 18.040 ;
        RECT 4.000 15.320 148.725 16.640 ;
        RECT 4.000 13.920 148.325 15.320 ;
        RECT 4.000 11.240 148.725 13.920 ;
        RECT 4.400 9.840 148.725 11.240 ;
        RECT 4.000 5.800 148.725 9.840 ;
        RECT 4.000 4.440 148.325 5.800 ;
        RECT 4.400 4.400 148.325 4.440 ;
        RECT 4.400 3.575 148.725 4.400 ;
      LAYER met4 ;
        RECT 30.335 10.640 51.545 152.560 ;
        RECT 53.945 10.640 75.160 152.560 ;
        RECT 77.560 10.640 98.770 152.560 ;
        RECT 101.170 10.640 101.825 152.560 ;
  END
END uart_to_mem
END LIBRARY

