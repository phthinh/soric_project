magic
tech sky130A
magscale 1 2
timestamp 1640734683
<< obsli1 >>
rect 1104 629 279375 279259
<< obsm1 >>
rect 14 620 279387 279268
<< metal2 >>
rect 1030 279200 1086 280000
rect 3146 279200 3202 280000
rect 5262 279200 5318 280000
rect 7378 279200 7434 280000
rect 9494 279200 9550 280000
rect 11610 279200 11666 280000
rect 13726 279200 13782 280000
rect 15842 279200 15898 280000
rect 17958 279200 18014 280000
rect 20074 279200 20130 280000
rect 22190 279200 22246 280000
rect 24306 279200 24362 280000
rect 26422 279200 26478 280000
rect 28538 279200 28594 280000
rect 30654 279200 30710 280000
rect 32770 279200 32826 280000
rect 34886 279200 34942 280000
rect 37002 279200 37058 280000
rect 39118 279200 39174 280000
rect 41326 279200 41382 280000
rect 43442 279200 43498 280000
rect 45558 279200 45614 280000
rect 47674 279200 47730 280000
rect 49790 279200 49846 280000
rect 51906 279200 51962 280000
rect 54022 279200 54078 280000
rect 56138 279200 56194 280000
rect 58254 279200 58310 280000
rect 60370 279200 60426 280000
rect 62486 279200 62542 280000
rect 64602 279200 64658 280000
rect 66718 279200 66774 280000
rect 68834 279200 68890 280000
rect 70950 279200 71006 280000
rect 73066 279200 73122 280000
rect 75182 279200 75238 280000
rect 77298 279200 77354 280000
rect 79414 279200 79470 280000
rect 81622 279200 81678 280000
rect 83738 279200 83794 280000
rect 85854 279200 85910 280000
rect 87970 279200 88026 280000
rect 90086 279200 90142 280000
rect 92202 279200 92258 280000
rect 94318 279200 94374 280000
rect 96434 279200 96490 280000
rect 98550 279200 98606 280000
rect 100666 279200 100722 280000
rect 102782 279200 102838 280000
rect 104898 279200 104954 280000
rect 107014 279200 107070 280000
rect 109130 279200 109186 280000
rect 111246 279200 111302 280000
rect 113362 279200 113418 280000
rect 115478 279200 115534 280000
rect 117594 279200 117650 280000
rect 119710 279200 119766 280000
rect 121918 279200 121974 280000
rect 124034 279200 124090 280000
rect 126150 279200 126206 280000
rect 128266 279200 128322 280000
rect 130382 279200 130438 280000
rect 132498 279200 132554 280000
rect 134614 279200 134670 280000
rect 136730 279200 136786 280000
rect 138846 279200 138902 280000
rect 140962 279200 141018 280000
rect 143078 279200 143134 280000
rect 145194 279200 145250 280000
rect 147310 279200 147366 280000
rect 149426 279200 149482 280000
rect 151542 279200 151598 280000
rect 153658 279200 153714 280000
rect 155774 279200 155830 280000
rect 157890 279200 157946 280000
rect 160006 279200 160062 280000
rect 162214 279200 162270 280000
rect 164330 279200 164386 280000
rect 166446 279200 166502 280000
rect 168562 279200 168618 280000
rect 170678 279200 170734 280000
rect 172794 279200 172850 280000
rect 174910 279200 174966 280000
rect 177026 279200 177082 280000
rect 179142 279200 179198 280000
rect 181258 279200 181314 280000
rect 183374 279200 183430 280000
rect 185490 279200 185546 280000
rect 187606 279200 187662 280000
rect 189722 279200 189778 280000
rect 191838 279200 191894 280000
rect 193954 279200 194010 280000
rect 196070 279200 196126 280000
rect 198186 279200 198242 280000
rect 200302 279200 200358 280000
rect 202510 279200 202566 280000
rect 204626 279200 204682 280000
rect 206742 279200 206798 280000
rect 208858 279200 208914 280000
rect 210974 279200 211030 280000
rect 213090 279200 213146 280000
rect 215206 279200 215262 280000
rect 217322 279200 217378 280000
rect 219438 279200 219494 280000
rect 221554 279200 221610 280000
rect 223670 279200 223726 280000
rect 225786 279200 225842 280000
rect 227902 279200 227958 280000
rect 230018 279200 230074 280000
rect 232134 279200 232190 280000
rect 234250 279200 234306 280000
rect 236366 279200 236422 280000
rect 238482 279200 238538 280000
rect 240598 279200 240654 280000
rect 242806 279200 242862 280000
rect 244922 279200 244978 280000
rect 247038 279200 247094 280000
rect 249154 279200 249210 280000
rect 251270 279200 251326 280000
rect 253386 279200 253442 280000
rect 255502 279200 255558 280000
rect 257618 279200 257674 280000
rect 259734 279200 259790 280000
rect 261850 279200 261906 280000
rect 263966 279200 264022 280000
rect 266082 279200 266138 280000
rect 268198 279200 268254 280000
rect 270314 279200 270370 280000
rect 272430 279200 272486 280000
rect 274546 279200 274602 280000
rect 276662 279200 276718 280000
rect 278778 279200 278834 280000
rect 1214 0 1270 800
rect 3606 0 3662 800
rect 5998 0 6054 800
rect 8390 0 8446 800
rect 10782 0 10838 800
rect 13266 0 13322 800
rect 15658 0 15714 800
rect 18050 0 18106 800
rect 20442 0 20498 800
rect 22926 0 22982 800
rect 25318 0 25374 800
rect 27710 0 27766 800
rect 30102 0 30158 800
rect 32586 0 32642 800
rect 34978 0 35034 800
rect 37370 0 37426 800
rect 39762 0 39818 800
rect 42154 0 42210 800
rect 44638 0 44694 800
rect 47030 0 47086 800
rect 49422 0 49478 800
rect 51814 0 51870 800
rect 54298 0 54354 800
rect 56690 0 56746 800
rect 59082 0 59138 800
rect 61474 0 61530 800
rect 63958 0 64014 800
rect 66350 0 66406 800
rect 68742 0 68798 800
rect 71134 0 71190 800
rect 73526 0 73582 800
rect 76010 0 76066 800
rect 78402 0 78458 800
rect 80794 0 80850 800
rect 83186 0 83242 800
rect 85670 0 85726 800
rect 88062 0 88118 800
rect 90454 0 90510 800
rect 92846 0 92902 800
rect 95330 0 95386 800
rect 97722 0 97778 800
rect 100114 0 100170 800
rect 102506 0 102562 800
rect 104990 0 105046 800
rect 107382 0 107438 800
rect 109774 0 109830 800
rect 112166 0 112222 800
rect 114558 0 114614 800
rect 117042 0 117098 800
rect 119434 0 119490 800
rect 121826 0 121882 800
rect 124218 0 124274 800
rect 126702 0 126758 800
rect 129094 0 129150 800
rect 131486 0 131542 800
rect 133878 0 133934 800
rect 136362 0 136418 800
rect 138754 0 138810 800
rect 141146 0 141202 800
rect 143538 0 143594 800
rect 145930 0 145986 800
rect 148414 0 148470 800
rect 150806 0 150862 800
rect 153198 0 153254 800
rect 155590 0 155646 800
rect 158074 0 158130 800
rect 160466 0 160522 800
rect 162858 0 162914 800
rect 165250 0 165306 800
rect 167734 0 167790 800
rect 170126 0 170182 800
rect 172518 0 172574 800
rect 174910 0 174966 800
rect 177302 0 177358 800
rect 179786 0 179842 800
rect 182178 0 182234 800
rect 184570 0 184626 800
rect 186962 0 187018 800
rect 189446 0 189502 800
rect 191838 0 191894 800
rect 194230 0 194286 800
rect 196622 0 196678 800
rect 199106 0 199162 800
rect 201498 0 201554 800
rect 203890 0 203946 800
rect 206282 0 206338 800
rect 208766 0 208822 800
rect 211158 0 211214 800
rect 213550 0 213606 800
rect 215942 0 215998 800
rect 218334 0 218390 800
rect 220818 0 220874 800
rect 223210 0 223266 800
rect 225602 0 225658 800
rect 227994 0 228050 800
rect 230478 0 230534 800
rect 232870 0 232926 800
rect 235262 0 235318 800
rect 237654 0 237710 800
rect 240138 0 240194 800
rect 242530 0 242586 800
rect 244922 0 244978 800
rect 247314 0 247370 800
rect 249706 0 249762 800
rect 252190 0 252246 800
rect 254582 0 254638 800
rect 256974 0 257030 800
rect 259366 0 259422 800
rect 261850 0 261906 800
rect 264242 0 264298 800
rect 266634 0 266690 800
rect 269026 0 269082 800
rect 271510 0 271566 800
rect 273902 0 273958 800
rect 276294 0 276350 800
rect 278686 0 278742 800
<< obsm2 >>
rect 20 279144 974 279313
rect 1142 279144 3090 279313
rect 3258 279144 5206 279313
rect 5374 279144 7322 279313
rect 7490 279144 9438 279313
rect 9606 279144 11554 279313
rect 11722 279144 13670 279313
rect 13838 279144 15786 279313
rect 15954 279144 17902 279313
rect 18070 279144 20018 279313
rect 20186 279144 22134 279313
rect 22302 279144 24250 279313
rect 24418 279144 26366 279313
rect 26534 279144 28482 279313
rect 28650 279144 30598 279313
rect 30766 279144 32714 279313
rect 32882 279144 34830 279313
rect 34998 279144 36946 279313
rect 37114 279144 39062 279313
rect 39230 279144 41270 279313
rect 41438 279144 43386 279313
rect 43554 279144 45502 279313
rect 45670 279144 47618 279313
rect 47786 279144 49734 279313
rect 49902 279144 51850 279313
rect 52018 279144 53966 279313
rect 54134 279144 56082 279313
rect 56250 279144 58198 279313
rect 58366 279144 60314 279313
rect 60482 279144 62430 279313
rect 62598 279144 64546 279313
rect 64714 279144 66662 279313
rect 66830 279144 68778 279313
rect 68946 279144 70894 279313
rect 71062 279144 73010 279313
rect 73178 279144 75126 279313
rect 75294 279144 77242 279313
rect 77410 279144 79358 279313
rect 79526 279144 81566 279313
rect 81734 279144 83682 279313
rect 83850 279144 85798 279313
rect 85966 279144 87914 279313
rect 88082 279144 90030 279313
rect 90198 279144 92146 279313
rect 92314 279144 94262 279313
rect 94430 279144 96378 279313
rect 96546 279144 98494 279313
rect 98662 279144 100610 279313
rect 100778 279144 102726 279313
rect 102894 279144 104842 279313
rect 105010 279144 106958 279313
rect 107126 279144 109074 279313
rect 109242 279144 111190 279313
rect 111358 279144 113306 279313
rect 113474 279144 115422 279313
rect 115590 279144 117538 279313
rect 117706 279144 119654 279313
rect 119822 279144 121862 279313
rect 122030 279144 123978 279313
rect 124146 279144 126094 279313
rect 126262 279144 128210 279313
rect 128378 279144 130326 279313
rect 130494 279144 132442 279313
rect 132610 279144 134558 279313
rect 134726 279144 136674 279313
rect 136842 279144 138790 279313
rect 138958 279144 140906 279313
rect 141074 279144 143022 279313
rect 143190 279144 145138 279313
rect 145306 279144 147254 279313
rect 147422 279144 149370 279313
rect 149538 279144 151486 279313
rect 151654 279144 153602 279313
rect 153770 279144 155718 279313
rect 155886 279144 157834 279313
rect 158002 279144 159950 279313
rect 160118 279144 162158 279313
rect 162326 279144 164274 279313
rect 164442 279144 166390 279313
rect 166558 279144 168506 279313
rect 168674 279144 170622 279313
rect 170790 279144 172738 279313
rect 172906 279144 174854 279313
rect 175022 279144 176970 279313
rect 177138 279144 179086 279313
rect 179254 279144 181202 279313
rect 181370 279144 183318 279313
rect 183486 279144 185434 279313
rect 185602 279144 187550 279313
rect 187718 279144 189666 279313
rect 189834 279144 191782 279313
rect 191950 279144 193898 279313
rect 194066 279144 196014 279313
rect 196182 279144 198130 279313
rect 198298 279144 200246 279313
rect 200414 279144 202454 279313
rect 202622 279144 204570 279313
rect 204738 279144 206686 279313
rect 206854 279144 208802 279313
rect 208970 279144 210918 279313
rect 211086 279144 213034 279313
rect 213202 279144 215150 279313
rect 215318 279144 217266 279313
rect 217434 279144 219382 279313
rect 219550 279144 221498 279313
rect 221666 279144 223614 279313
rect 223782 279144 225730 279313
rect 225898 279144 227846 279313
rect 228014 279144 229962 279313
rect 230130 279144 232078 279313
rect 232246 279144 234194 279313
rect 234362 279144 236310 279313
rect 236478 279144 238426 279313
rect 238594 279144 240542 279313
rect 240710 279144 242750 279313
rect 242918 279144 244866 279313
rect 245034 279144 246982 279313
rect 247150 279144 249098 279313
rect 249266 279144 251214 279313
rect 251382 279144 253330 279313
rect 253498 279144 255446 279313
rect 255614 279144 257562 279313
rect 257730 279144 259678 279313
rect 259846 279144 261794 279313
rect 261962 279144 263910 279313
rect 264078 279144 266026 279313
rect 266194 279144 268142 279313
rect 268310 279144 270258 279313
rect 270426 279144 272374 279313
rect 272542 279144 274490 279313
rect 274658 279144 276606 279313
rect 276774 279144 278722 279313
rect 278890 279144 279110 279313
rect 20 856 279110 279144
rect 20 575 1158 856
rect 1326 575 3550 856
rect 3718 575 5942 856
rect 6110 575 8334 856
rect 8502 575 10726 856
rect 10894 575 13210 856
rect 13378 575 15602 856
rect 15770 575 17994 856
rect 18162 575 20386 856
rect 20554 575 22870 856
rect 23038 575 25262 856
rect 25430 575 27654 856
rect 27822 575 30046 856
rect 30214 575 32530 856
rect 32698 575 34922 856
rect 35090 575 37314 856
rect 37482 575 39706 856
rect 39874 575 42098 856
rect 42266 575 44582 856
rect 44750 575 46974 856
rect 47142 575 49366 856
rect 49534 575 51758 856
rect 51926 575 54242 856
rect 54410 575 56634 856
rect 56802 575 59026 856
rect 59194 575 61418 856
rect 61586 575 63902 856
rect 64070 575 66294 856
rect 66462 575 68686 856
rect 68854 575 71078 856
rect 71246 575 73470 856
rect 73638 575 75954 856
rect 76122 575 78346 856
rect 78514 575 80738 856
rect 80906 575 83130 856
rect 83298 575 85614 856
rect 85782 575 88006 856
rect 88174 575 90398 856
rect 90566 575 92790 856
rect 92958 575 95274 856
rect 95442 575 97666 856
rect 97834 575 100058 856
rect 100226 575 102450 856
rect 102618 575 104934 856
rect 105102 575 107326 856
rect 107494 575 109718 856
rect 109886 575 112110 856
rect 112278 575 114502 856
rect 114670 575 116986 856
rect 117154 575 119378 856
rect 119546 575 121770 856
rect 121938 575 124162 856
rect 124330 575 126646 856
rect 126814 575 129038 856
rect 129206 575 131430 856
rect 131598 575 133822 856
rect 133990 575 136306 856
rect 136474 575 138698 856
rect 138866 575 141090 856
rect 141258 575 143482 856
rect 143650 575 145874 856
rect 146042 575 148358 856
rect 148526 575 150750 856
rect 150918 575 153142 856
rect 153310 575 155534 856
rect 155702 575 158018 856
rect 158186 575 160410 856
rect 160578 575 162802 856
rect 162970 575 165194 856
rect 165362 575 167678 856
rect 167846 575 170070 856
rect 170238 575 172462 856
rect 172630 575 174854 856
rect 175022 575 177246 856
rect 177414 575 179730 856
rect 179898 575 182122 856
rect 182290 575 184514 856
rect 184682 575 186906 856
rect 187074 575 189390 856
rect 189558 575 191782 856
rect 191950 575 194174 856
rect 194342 575 196566 856
rect 196734 575 199050 856
rect 199218 575 201442 856
rect 201610 575 203834 856
rect 204002 575 206226 856
rect 206394 575 208710 856
rect 208878 575 211102 856
rect 211270 575 213494 856
rect 213662 575 215886 856
rect 216054 575 218278 856
rect 218446 575 220762 856
rect 220930 575 223154 856
rect 223322 575 225546 856
rect 225714 575 227938 856
rect 228106 575 230422 856
rect 230590 575 232814 856
rect 232982 575 235206 856
rect 235374 575 237598 856
rect 237766 575 240082 856
rect 240250 575 242474 856
rect 242642 575 244866 856
rect 245034 575 247258 856
rect 247426 575 249650 856
rect 249818 575 252134 856
rect 252302 575 254526 856
rect 254694 575 256918 856
rect 257086 575 259310 856
rect 259478 575 261794 856
rect 261962 575 264186 856
rect 264354 575 266578 856
rect 266746 575 268970 856
rect 269138 575 271454 856
rect 271622 575 273846 856
rect 274014 575 276238 856
rect 276406 575 278630 856
rect 278798 575 279110 856
<< metal3 >>
rect 279200 279216 280000 279336
rect 0 278672 800 278792
rect 279200 277992 280000 278112
rect 279200 276632 280000 276752
rect 0 276224 800 276344
rect 279200 275408 280000 275528
rect 0 273912 800 274032
rect 279200 274048 280000 274168
rect 279200 272824 280000 272944
rect 0 271464 800 271584
rect 279200 271600 280000 271720
rect 279200 270240 280000 270360
rect 0 269152 800 269272
rect 279200 269016 280000 269136
rect 279200 267656 280000 267776
rect 0 266704 800 266824
rect 279200 266432 280000 266552
rect 279200 265208 280000 265328
rect 0 264256 800 264376
rect 279200 263848 280000 263968
rect 279200 262624 280000 262744
rect 0 261944 800 262064
rect 279200 261264 280000 261384
rect 279200 260040 280000 260160
rect 0 259496 800 259616
rect 279200 258816 280000 258936
rect 279200 257456 280000 257576
rect 0 257184 800 257304
rect 279200 256232 280000 256352
rect 0 254736 800 254856
rect 279200 254872 280000 254992
rect 279200 253648 280000 253768
rect 0 252288 800 252408
rect 279200 252424 280000 252544
rect 279200 251064 280000 251184
rect 0 249976 800 250096
rect 279200 249840 280000 249960
rect 279200 248480 280000 248600
rect 0 247528 800 247648
rect 279200 247256 280000 247376
rect 279200 246032 280000 246152
rect 0 245216 800 245336
rect 279200 244672 280000 244792
rect 279200 243448 280000 243568
rect 0 242768 800 242888
rect 279200 242088 280000 242208
rect 279200 240864 280000 240984
rect 0 240320 800 240440
rect 279200 239640 280000 239760
rect 279200 238280 280000 238400
rect 0 238008 800 238128
rect 279200 237056 280000 237176
rect 0 235560 800 235680
rect 279200 235696 280000 235816
rect 279200 234472 280000 234592
rect 0 233248 800 233368
rect 279200 233248 280000 233368
rect 279200 231888 280000 232008
rect 0 230800 800 230920
rect 279200 230664 280000 230784
rect 279200 229304 280000 229424
rect 0 228352 800 228472
rect 279200 228080 280000 228200
rect 279200 226856 280000 226976
rect 0 226040 800 226160
rect 279200 225496 280000 225616
rect 279200 224272 280000 224392
rect 0 223592 800 223712
rect 279200 222912 280000 223032
rect 279200 221688 280000 221808
rect 0 221280 800 221400
rect 279200 220464 280000 220584
rect 279200 219104 280000 219224
rect 0 218832 800 218952
rect 279200 217880 280000 218000
rect 0 216384 800 216504
rect 279200 216520 280000 216640
rect 279200 215296 280000 215416
rect 0 214072 800 214192
rect 279200 214072 280000 214192
rect 279200 212712 280000 212832
rect 0 211624 800 211744
rect 279200 211488 280000 211608
rect 279200 210128 280000 210248
rect 0 209312 800 209432
rect 279200 208904 280000 209024
rect 279200 207680 280000 207800
rect 0 206864 800 206984
rect 279200 206320 280000 206440
rect 279200 205096 280000 205216
rect 0 204416 800 204536
rect 279200 203736 280000 203856
rect 279200 202512 280000 202632
rect 0 202104 800 202224
rect 279200 201288 280000 201408
rect 279200 199928 280000 200048
rect 0 199656 800 199776
rect 279200 198704 280000 198824
rect 0 197344 800 197464
rect 279200 197344 280000 197464
rect 279200 196120 280000 196240
rect 0 194896 800 195016
rect 279200 194896 280000 195016
rect 279200 193536 280000 193656
rect 0 192448 800 192568
rect 279200 192312 280000 192432
rect 279200 190952 280000 191072
rect 0 190136 800 190256
rect 279200 189728 280000 189848
rect 279200 188504 280000 188624
rect 0 187688 800 187808
rect 279200 187144 280000 187264
rect 279200 185920 280000 186040
rect 0 185376 800 185496
rect 279200 184560 280000 184680
rect 279200 183336 280000 183456
rect 0 182928 800 183048
rect 279200 182112 280000 182232
rect 279200 180752 280000 180872
rect 0 180480 800 180600
rect 279200 179528 280000 179648
rect 0 178168 800 178288
rect 279200 178168 280000 178288
rect 279200 176944 280000 177064
rect 0 175720 800 175840
rect 279200 175720 280000 175840
rect 279200 174360 280000 174480
rect 0 173408 800 173528
rect 279200 173136 280000 173256
rect 279200 171776 280000 171896
rect 0 170960 800 171080
rect 279200 170552 280000 170672
rect 279200 169328 280000 169448
rect 0 168512 800 168632
rect 279200 167968 280000 168088
rect 279200 166744 280000 166864
rect 0 166200 800 166320
rect 279200 165384 280000 165504
rect 279200 164160 280000 164280
rect 0 163752 800 163872
rect 279200 162936 280000 163056
rect 0 161440 800 161560
rect 279200 161576 280000 161696
rect 279200 160352 280000 160472
rect 0 158992 800 159112
rect 279200 158992 280000 159112
rect 279200 157768 280000 157888
rect 0 156544 800 156664
rect 279200 156544 280000 156664
rect 279200 155184 280000 155304
rect 0 154232 800 154352
rect 279200 153960 280000 154080
rect 279200 152600 280000 152720
rect 0 151784 800 151904
rect 279200 151376 280000 151496
rect 279200 150152 280000 150272
rect 0 149472 800 149592
rect 279200 148792 280000 148912
rect 279200 147568 280000 147688
rect 0 147024 800 147144
rect 279200 146208 280000 146328
rect 279200 144984 280000 145104
rect 0 144576 800 144696
rect 279200 143760 280000 143880
rect 0 142264 800 142384
rect 279200 142400 280000 142520
rect 279200 141176 280000 141296
rect 0 139816 800 139936
rect 279200 139816 280000 139936
rect 279200 138592 280000 138712
rect 0 137504 800 137624
rect 279200 137232 280000 137352
rect 279200 136008 280000 136128
rect 0 135056 800 135176
rect 279200 134784 280000 134904
rect 279200 133424 280000 133544
rect 0 132608 800 132728
rect 279200 132200 280000 132320
rect 279200 130840 280000 130960
rect 0 130296 800 130416
rect 279200 129616 280000 129736
rect 279200 128392 280000 128512
rect 0 127848 800 127968
rect 279200 127032 280000 127152
rect 279200 125808 280000 125928
rect 0 125536 800 125656
rect 279200 124448 280000 124568
rect 0 123088 800 123208
rect 279200 123224 280000 123344
rect 279200 122000 280000 122120
rect 0 120640 800 120760
rect 279200 120640 280000 120760
rect 279200 119416 280000 119536
rect 0 118328 800 118448
rect 279200 118056 280000 118176
rect 279200 116832 280000 116952
rect 0 115880 800 116000
rect 279200 115608 280000 115728
rect 279200 114248 280000 114368
rect 0 113568 800 113688
rect 279200 113024 280000 113144
rect 279200 111664 280000 111784
rect 0 111120 800 111240
rect 279200 110440 280000 110560
rect 279200 109216 280000 109336
rect 0 108672 800 108792
rect 279200 107856 280000 107976
rect 279200 106632 280000 106752
rect 0 106360 800 106480
rect 279200 105272 280000 105392
rect 0 103912 800 104032
rect 279200 104048 280000 104168
rect 279200 102824 280000 102944
rect 0 101600 800 101720
rect 279200 101464 280000 101584
rect 279200 100240 280000 100360
rect 0 99152 800 99272
rect 279200 98880 280000 99000
rect 279200 97656 280000 97776
rect 0 96704 800 96824
rect 279200 96432 280000 96552
rect 279200 95072 280000 95192
rect 0 94392 800 94512
rect 279200 93848 280000 93968
rect 279200 92488 280000 92608
rect 0 91944 800 92064
rect 279200 91264 280000 91384
rect 279200 90040 280000 90160
rect 0 89632 800 89752
rect 279200 88680 280000 88800
rect 279200 87456 280000 87576
rect 0 87184 800 87304
rect 279200 86096 280000 86216
rect 0 84736 800 84856
rect 279200 84872 280000 84992
rect 279200 83648 280000 83768
rect 0 82424 800 82544
rect 279200 82288 280000 82408
rect 279200 81064 280000 81184
rect 0 79976 800 80096
rect 279200 79704 280000 79824
rect 279200 78480 280000 78600
rect 0 77664 800 77784
rect 279200 77256 280000 77376
rect 279200 75896 280000 76016
rect 0 75216 800 75336
rect 279200 74672 280000 74792
rect 279200 73312 280000 73432
rect 0 72768 800 72888
rect 279200 72088 280000 72208
rect 279200 70864 280000 70984
rect 0 70456 800 70576
rect 279200 69504 280000 69624
rect 279200 68280 280000 68400
rect 0 68008 800 68128
rect 279200 66920 280000 67040
rect 0 65696 800 65816
rect 279200 65696 280000 65816
rect 279200 64472 280000 64592
rect 0 63248 800 63368
rect 279200 63112 280000 63232
rect 279200 61888 280000 62008
rect 0 60800 800 60920
rect 279200 60528 280000 60648
rect 279200 59304 280000 59424
rect 0 58488 800 58608
rect 279200 58080 280000 58200
rect 279200 56720 280000 56840
rect 0 56040 800 56160
rect 279200 55496 280000 55616
rect 279200 54136 280000 54256
rect 0 53728 800 53848
rect 279200 52912 280000 53032
rect 279200 51688 280000 51808
rect 0 51280 800 51400
rect 279200 50328 280000 50448
rect 279200 49104 280000 49224
rect 0 48832 800 48952
rect 279200 47744 280000 47864
rect 0 46520 800 46640
rect 279200 46520 280000 46640
rect 279200 45296 280000 45416
rect 0 44072 800 44192
rect 279200 43936 280000 44056
rect 279200 42712 280000 42832
rect 0 41760 800 41880
rect 279200 41352 280000 41472
rect 279200 40128 280000 40248
rect 0 39312 800 39432
rect 279200 38904 280000 39024
rect 279200 37544 280000 37664
rect 0 36864 800 36984
rect 279200 36320 280000 36440
rect 279200 34960 280000 35080
rect 0 34552 800 34672
rect 279200 33736 280000 33856
rect 279200 32512 280000 32632
rect 0 32104 800 32224
rect 279200 31152 280000 31272
rect 0 29792 800 29912
rect 279200 29928 280000 30048
rect 279200 28568 280000 28688
rect 0 27344 800 27464
rect 279200 27344 280000 27464
rect 279200 26120 280000 26240
rect 0 24896 800 25016
rect 279200 24760 280000 24880
rect 279200 23536 280000 23656
rect 0 22584 800 22704
rect 279200 22176 280000 22296
rect 279200 20952 280000 21072
rect 0 20136 800 20256
rect 279200 19728 280000 19848
rect 279200 18368 280000 18488
rect 0 17824 800 17944
rect 279200 17144 280000 17264
rect 279200 15784 280000 15904
rect 0 15376 800 15496
rect 279200 14560 280000 14680
rect 279200 13336 280000 13456
rect 0 12928 800 13048
rect 279200 11976 280000 12096
rect 0 10616 800 10736
rect 279200 10752 280000 10872
rect 279200 9392 280000 9512
rect 0 8168 800 8288
rect 279200 8168 280000 8288
rect 279200 6944 280000 7064
rect 0 5856 800 5976
rect 279200 5584 280000 5704
rect 279200 4360 280000 4480
rect 0 3408 800 3528
rect 279200 3000 280000 3120
rect 279200 1776 280000 1896
rect 0 1096 800 1216
rect 279200 552 280000 672
<< obsm3 >>
rect 800 279136 279120 279309
rect 800 278872 279200 279136
rect 880 278592 279200 278872
rect 800 278192 279200 278592
rect 800 277912 279120 278192
rect 800 276832 279200 277912
rect 800 276552 279120 276832
rect 800 276424 279200 276552
rect 880 276144 279200 276424
rect 800 275608 279200 276144
rect 800 275328 279120 275608
rect 800 274248 279200 275328
rect 800 274112 279120 274248
rect 880 273968 279120 274112
rect 880 273832 279200 273968
rect 800 273024 279200 273832
rect 800 272744 279120 273024
rect 800 271800 279200 272744
rect 800 271664 279120 271800
rect 880 271520 279120 271664
rect 880 271384 279200 271520
rect 800 270440 279200 271384
rect 800 270160 279120 270440
rect 800 269352 279200 270160
rect 880 269216 279200 269352
rect 880 269072 279120 269216
rect 800 268936 279120 269072
rect 800 267856 279200 268936
rect 800 267576 279120 267856
rect 800 266904 279200 267576
rect 880 266632 279200 266904
rect 880 266624 279120 266632
rect 800 266352 279120 266624
rect 800 265408 279200 266352
rect 800 265128 279120 265408
rect 800 264456 279200 265128
rect 880 264176 279200 264456
rect 800 264048 279200 264176
rect 800 263768 279120 264048
rect 800 262824 279200 263768
rect 800 262544 279120 262824
rect 800 262144 279200 262544
rect 880 261864 279200 262144
rect 800 261464 279200 261864
rect 800 261184 279120 261464
rect 800 260240 279200 261184
rect 800 259960 279120 260240
rect 800 259696 279200 259960
rect 880 259416 279200 259696
rect 800 259016 279200 259416
rect 800 258736 279120 259016
rect 800 257656 279200 258736
rect 800 257384 279120 257656
rect 880 257376 279120 257384
rect 880 257104 279200 257376
rect 800 256432 279200 257104
rect 800 256152 279120 256432
rect 800 255072 279200 256152
rect 800 254936 279120 255072
rect 880 254792 279120 254936
rect 880 254656 279200 254792
rect 800 253848 279200 254656
rect 800 253568 279120 253848
rect 800 252624 279200 253568
rect 800 252488 279120 252624
rect 880 252344 279120 252488
rect 880 252208 279200 252344
rect 800 251264 279200 252208
rect 800 250984 279120 251264
rect 800 250176 279200 250984
rect 880 250040 279200 250176
rect 880 249896 279120 250040
rect 800 249760 279120 249896
rect 800 248680 279200 249760
rect 800 248400 279120 248680
rect 800 247728 279200 248400
rect 880 247456 279200 247728
rect 880 247448 279120 247456
rect 800 247176 279120 247448
rect 800 246232 279200 247176
rect 800 245952 279120 246232
rect 800 245416 279200 245952
rect 880 245136 279200 245416
rect 800 244872 279200 245136
rect 800 244592 279120 244872
rect 800 243648 279200 244592
rect 800 243368 279120 243648
rect 800 242968 279200 243368
rect 880 242688 279200 242968
rect 800 242288 279200 242688
rect 800 242008 279120 242288
rect 800 241064 279200 242008
rect 800 240784 279120 241064
rect 800 240520 279200 240784
rect 880 240240 279200 240520
rect 800 239840 279200 240240
rect 800 239560 279120 239840
rect 800 238480 279200 239560
rect 800 238208 279120 238480
rect 880 238200 279120 238208
rect 880 237928 279200 238200
rect 800 237256 279200 237928
rect 800 236976 279120 237256
rect 800 235896 279200 236976
rect 800 235760 279120 235896
rect 880 235616 279120 235760
rect 880 235480 279200 235616
rect 800 234672 279200 235480
rect 800 234392 279120 234672
rect 800 233448 279200 234392
rect 880 233168 279120 233448
rect 800 232088 279200 233168
rect 800 231808 279120 232088
rect 800 231000 279200 231808
rect 880 230864 279200 231000
rect 880 230720 279120 230864
rect 800 230584 279120 230720
rect 800 229504 279200 230584
rect 800 229224 279120 229504
rect 800 228552 279200 229224
rect 880 228280 279200 228552
rect 880 228272 279120 228280
rect 800 228000 279120 228272
rect 800 227056 279200 228000
rect 800 226776 279120 227056
rect 800 226240 279200 226776
rect 880 225960 279200 226240
rect 800 225696 279200 225960
rect 800 225416 279120 225696
rect 800 224472 279200 225416
rect 800 224192 279120 224472
rect 800 223792 279200 224192
rect 880 223512 279200 223792
rect 800 223112 279200 223512
rect 800 222832 279120 223112
rect 800 221888 279200 222832
rect 800 221608 279120 221888
rect 800 221480 279200 221608
rect 880 221200 279200 221480
rect 800 220664 279200 221200
rect 800 220384 279120 220664
rect 800 219304 279200 220384
rect 800 219032 279120 219304
rect 880 219024 279120 219032
rect 880 218752 279200 219024
rect 800 218080 279200 218752
rect 800 217800 279120 218080
rect 800 216720 279200 217800
rect 800 216584 279120 216720
rect 880 216440 279120 216584
rect 880 216304 279200 216440
rect 800 215496 279200 216304
rect 800 215216 279120 215496
rect 800 214272 279200 215216
rect 880 213992 279120 214272
rect 800 212912 279200 213992
rect 800 212632 279120 212912
rect 800 211824 279200 212632
rect 880 211688 279200 211824
rect 880 211544 279120 211688
rect 800 211408 279120 211544
rect 800 210328 279200 211408
rect 800 210048 279120 210328
rect 800 209512 279200 210048
rect 880 209232 279200 209512
rect 800 209104 279200 209232
rect 800 208824 279120 209104
rect 800 207880 279200 208824
rect 800 207600 279120 207880
rect 800 207064 279200 207600
rect 880 206784 279200 207064
rect 800 206520 279200 206784
rect 800 206240 279120 206520
rect 800 205296 279200 206240
rect 800 205016 279120 205296
rect 800 204616 279200 205016
rect 880 204336 279200 204616
rect 800 203936 279200 204336
rect 800 203656 279120 203936
rect 800 202712 279200 203656
rect 800 202432 279120 202712
rect 800 202304 279200 202432
rect 880 202024 279200 202304
rect 800 201488 279200 202024
rect 800 201208 279120 201488
rect 800 200128 279200 201208
rect 800 199856 279120 200128
rect 880 199848 279120 199856
rect 880 199576 279200 199848
rect 800 198904 279200 199576
rect 800 198624 279120 198904
rect 800 197544 279200 198624
rect 880 197264 279120 197544
rect 800 196320 279200 197264
rect 800 196040 279120 196320
rect 800 195096 279200 196040
rect 880 194816 279120 195096
rect 800 193736 279200 194816
rect 800 193456 279120 193736
rect 800 192648 279200 193456
rect 880 192512 279200 192648
rect 880 192368 279120 192512
rect 800 192232 279120 192368
rect 800 191152 279200 192232
rect 800 190872 279120 191152
rect 800 190336 279200 190872
rect 880 190056 279200 190336
rect 800 189928 279200 190056
rect 800 189648 279120 189928
rect 800 188704 279200 189648
rect 800 188424 279120 188704
rect 800 187888 279200 188424
rect 880 187608 279200 187888
rect 800 187344 279200 187608
rect 800 187064 279120 187344
rect 800 186120 279200 187064
rect 800 185840 279120 186120
rect 800 185576 279200 185840
rect 880 185296 279200 185576
rect 800 184760 279200 185296
rect 800 184480 279120 184760
rect 800 183536 279200 184480
rect 800 183256 279120 183536
rect 800 183128 279200 183256
rect 880 182848 279200 183128
rect 800 182312 279200 182848
rect 800 182032 279120 182312
rect 800 180952 279200 182032
rect 800 180680 279120 180952
rect 880 180672 279120 180680
rect 880 180400 279200 180672
rect 800 179728 279200 180400
rect 800 179448 279120 179728
rect 800 178368 279200 179448
rect 880 178088 279120 178368
rect 800 177144 279200 178088
rect 800 176864 279120 177144
rect 800 175920 279200 176864
rect 880 175640 279120 175920
rect 800 174560 279200 175640
rect 800 174280 279120 174560
rect 800 173608 279200 174280
rect 880 173336 279200 173608
rect 880 173328 279120 173336
rect 800 173056 279120 173328
rect 800 171976 279200 173056
rect 800 171696 279120 171976
rect 800 171160 279200 171696
rect 880 170880 279200 171160
rect 800 170752 279200 170880
rect 800 170472 279120 170752
rect 800 169528 279200 170472
rect 800 169248 279120 169528
rect 800 168712 279200 169248
rect 880 168432 279200 168712
rect 800 168168 279200 168432
rect 800 167888 279120 168168
rect 800 166944 279200 167888
rect 800 166664 279120 166944
rect 800 166400 279200 166664
rect 880 166120 279200 166400
rect 800 165584 279200 166120
rect 800 165304 279120 165584
rect 800 164360 279200 165304
rect 800 164080 279120 164360
rect 800 163952 279200 164080
rect 880 163672 279200 163952
rect 800 163136 279200 163672
rect 800 162856 279120 163136
rect 800 161776 279200 162856
rect 800 161640 279120 161776
rect 880 161496 279120 161640
rect 880 161360 279200 161496
rect 800 160552 279200 161360
rect 800 160272 279120 160552
rect 800 159192 279200 160272
rect 880 158912 279120 159192
rect 800 157968 279200 158912
rect 800 157688 279120 157968
rect 800 156744 279200 157688
rect 880 156464 279120 156744
rect 800 155384 279200 156464
rect 800 155104 279120 155384
rect 800 154432 279200 155104
rect 880 154160 279200 154432
rect 880 154152 279120 154160
rect 800 153880 279120 154152
rect 800 152800 279200 153880
rect 800 152520 279120 152800
rect 800 151984 279200 152520
rect 880 151704 279200 151984
rect 800 151576 279200 151704
rect 800 151296 279120 151576
rect 800 150352 279200 151296
rect 800 150072 279120 150352
rect 800 149672 279200 150072
rect 880 149392 279200 149672
rect 800 148992 279200 149392
rect 800 148712 279120 148992
rect 800 147768 279200 148712
rect 800 147488 279120 147768
rect 800 147224 279200 147488
rect 880 146944 279200 147224
rect 800 146408 279200 146944
rect 800 146128 279120 146408
rect 800 145184 279200 146128
rect 800 144904 279120 145184
rect 800 144776 279200 144904
rect 880 144496 279200 144776
rect 800 143960 279200 144496
rect 800 143680 279120 143960
rect 800 142600 279200 143680
rect 800 142464 279120 142600
rect 880 142320 279120 142464
rect 880 142184 279200 142320
rect 800 141376 279200 142184
rect 800 141096 279120 141376
rect 800 140016 279200 141096
rect 880 139736 279120 140016
rect 800 138792 279200 139736
rect 800 138512 279120 138792
rect 800 137704 279200 138512
rect 880 137432 279200 137704
rect 880 137424 279120 137432
rect 800 137152 279120 137424
rect 800 136208 279200 137152
rect 800 135928 279120 136208
rect 800 135256 279200 135928
rect 880 134984 279200 135256
rect 880 134976 279120 134984
rect 800 134704 279120 134976
rect 800 133624 279200 134704
rect 800 133344 279120 133624
rect 800 132808 279200 133344
rect 880 132528 279200 132808
rect 800 132400 279200 132528
rect 800 132120 279120 132400
rect 800 131040 279200 132120
rect 800 130760 279120 131040
rect 800 130496 279200 130760
rect 880 130216 279200 130496
rect 800 129816 279200 130216
rect 800 129536 279120 129816
rect 800 128592 279200 129536
rect 800 128312 279120 128592
rect 800 128048 279200 128312
rect 880 127768 279200 128048
rect 800 127232 279200 127768
rect 800 126952 279120 127232
rect 800 126008 279200 126952
rect 800 125736 279120 126008
rect 880 125728 279120 125736
rect 880 125456 279200 125728
rect 800 124648 279200 125456
rect 800 124368 279120 124648
rect 800 123424 279200 124368
rect 800 123288 279120 123424
rect 880 123144 279120 123288
rect 880 123008 279200 123144
rect 800 122200 279200 123008
rect 800 121920 279120 122200
rect 800 120840 279200 121920
rect 880 120560 279120 120840
rect 800 119616 279200 120560
rect 800 119336 279120 119616
rect 800 118528 279200 119336
rect 880 118256 279200 118528
rect 880 118248 279120 118256
rect 800 117976 279120 118248
rect 800 117032 279200 117976
rect 800 116752 279120 117032
rect 800 116080 279200 116752
rect 880 115808 279200 116080
rect 880 115800 279120 115808
rect 800 115528 279120 115800
rect 800 114448 279200 115528
rect 800 114168 279120 114448
rect 800 113768 279200 114168
rect 880 113488 279200 113768
rect 800 113224 279200 113488
rect 800 112944 279120 113224
rect 800 111864 279200 112944
rect 800 111584 279120 111864
rect 800 111320 279200 111584
rect 880 111040 279200 111320
rect 800 110640 279200 111040
rect 800 110360 279120 110640
rect 800 109416 279200 110360
rect 800 109136 279120 109416
rect 800 108872 279200 109136
rect 880 108592 279200 108872
rect 800 108056 279200 108592
rect 800 107776 279120 108056
rect 800 106832 279200 107776
rect 800 106560 279120 106832
rect 880 106552 279120 106560
rect 880 106280 279200 106552
rect 800 105472 279200 106280
rect 800 105192 279120 105472
rect 800 104248 279200 105192
rect 800 104112 279120 104248
rect 880 103968 279120 104112
rect 880 103832 279200 103968
rect 800 103024 279200 103832
rect 800 102744 279120 103024
rect 800 101800 279200 102744
rect 880 101664 279200 101800
rect 880 101520 279120 101664
rect 800 101384 279120 101520
rect 800 100440 279200 101384
rect 800 100160 279120 100440
rect 800 99352 279200 100160
rect 880 99080 279200 99352
rect 880 99072 279120 99080
rect 800 98800 279120 99072
rect 800 97856 279200 98800
rect 800 97576 279120 97856
rect 800 96904 279200 97576
rect 880 96632 279200 96904
rect 880 96624 279120 96632
rect 800 96352 279120 96624
rect 800 95272 279200 96352
rect 800 94992 279120 95272
rect 800 94592 279200 94992
rect 880 94312 279200 94592
rect 800 94048 279200 94312
rect 800 93768 279120 94048
rect 800 92688 279200 93768
rect 800 92408 279120 92688
rect 800 92144 279200 92408
rect 880 91864 279200 92144
rect 800 91464 279200 91864
rect 800 91184 279120 91464
rect 800 90240 279200 91184
rect 800 89960 279120 90240
rect 800 89832 279200 89960
rect 880 89552 279200 89832
rect 800 88880 279200 89552
rect 800 88600 279120 88880
rect 800 87656 279200 88600
rect 800 87384 279120 87656
rect 880 87376 279120 87384
rect 880 87104 279200 87376
rect 800 86296 279200 87104
rect 800 86016 279120 86296
rect 800 85072 279200 86016
rect 800 84936 279120 85072
rect 880 84792 279120 84936
rect 880 84656 279200 84792
rect 800 83848 279200 84656
rect 800 83568 279120 83848
rect 800 82624 279200 83568
rect 880 82488 279200 82624
rect 880 82344 279120 82488
rect 800 82208 279120 82344
rect 800 81264 279200 82208
rect 800 80984 279120 81264
rect 800 80176 279200 80984
rect 880 79904 279200 80176
rect 880 79896 279120 79904
rect 800 79624 279120 79896
rect 800 78680 279200 79624
rect 800 78400 279120 78680
rect 800 77864 279200 78400
rect 880 77584 279200 77864
rect 800 77456 279200 77584
rect 800 77176 279120 77456
rect 800 76096 279200 77176
rect 800 75816 279120 76096
rect 800 75416 279200 75816
rect 880 75136 279200 75416
rect 800 74872 279200 75136
rect 800 74592 279120 74872
rect 800 73512 279200 74592
rect 800 73232 279120 73512
rect 800 72968 279200 73232
rect 880 72688 279200 72968
rect 800 72288 279200 72688
rect 800 72008 279120 72288
rect 800 71064 279200 72008
rect 800 70784 279120 71064
rect 800 70656 279200 70784
rect 880 70376 279200 70656
rect 800 69704 279200 70376
rect 800 69424 279120 69704
rect 800 68480 279200 69424
rect 800 68208 279120 68480
rect 880 68200 279120 68208
rect 880 67928 279200 68200
rect 800 67120 279200 67928
rect 800 66840 279120 67120
rect 800 65896 279200 66840
rect 880 65616 279120 65896
rect 800 64672 279200 65616
rect 800 64392 279120 64672
rect 800 63448 279200 64392
rect 880 63312 279200 63448
rect 880 63168 279120 63312
rect 800 63032 279120 63168
rect 800 62088 279200 63032
rect 800 61808 279120 62088
rect 800 61000 279200 61808
rect 880 60728 279200 61000
rect 880 60720 279120 60728
rect 800 60448 279120 60720
rect 800 59504 279200 60448
rect 800 59224 279120 59504
rect 800 58688 279200 59224
rect 880 58408 279200 58688
rect 800 58280 279200 58408
rect 800 58000 279120 58280
rect 800 56920 279200 58000
rect 800 56640 279120 56920
rect 800 56240 279200 56640
rect 880 55960 279200 56240
rect 800 55696 279200 55960
rect 800 55416 279120 55696
rect 800 54336 279200 55416
rect 800 54056 279120 54336
rect 800 53928 279200 54056
rect 880 53648 279200 53928
rect 800 53112 279200 53648
rect 800 52832 279120 53112
rect 800 51888 279200 52832
rect 800 51608 279120 51888
rect 800 51480 279200 51608
rect 880 51200 279200 51480
rect 800 50528 279200 51200
rect 800 50248 279120 50528
rect 800 49304 279200 50248
rect 800 49032 279120 49304
rect 880 49024 279120 49032
rect 880 48752 279200 49024
rect 800 47944 279200 48752
rect 800 47664 279120 47944
rect 800 46720 279200 47664
rect 880 46440 279120 46720
rect 800 45496 279200 46440
rect 800 45216 279120 45496
rect 800 44272 279200 45216
rect 880 44136 279200 44272
rect 880 43992 279120 44136
rect 800 43856 279120 43992
rect 800 42912 279200 43856
rect 800 42632 279120 42912
rect 800 41960 279200 42632
rect 880 41680 279200 41960
rect 800 41552 279200 41680
rect 800 41272 279120 41552
rect 800 40328 279200 41272
rect 800 40048 279120 40328
rect 800 39512 279200 40048
rect 880 39232 279200 39512
rect 800 39104 279200 39232
rect 800 38824 279120 39104
rect 800 37744 279200 38824
rect 800 37464 279120 37744
rect 800 37064 279200 37464
rect 880 36784 279200 37064
rect 800 36520 279200 36784
rect 800 36240 279120 36520
rect 800 35160 279200 36240
rect 800 34880 279120 35160
rect 800 34752 279200 34880
rect 880 34472 279200 34752
rect 800 33936 279200 34472
rect 800 33656 279120 33936
rect 800 32712 279200 33656
rect 800 32432 279120 32712
rect 800 32304 279200 32432
rect 880 32024 279200 32304
rect 800 31352 279200 32024
rect 800 31072 279120 31352
rect 800 30128 279200 31072
rect 800 29992 279120 30128
rect 880 29848 279120 29992
rect 880 29712 279200 29848
rect 800 28768 279200 29712
rect 800 28488 279120 28768
rect 800 27544 279200 28488
rect 880 27264 279120 27544
rect 800 26320 279200 27264
rect 800 26040 279120 26320
rect 800 25096 279200 26040
rect 880 24960 279200 25096
rect 880 24816 279120 24960
rect 800 24680 279120 24816
rect 800 23736 279200 24680
rect 800 23456 279120 23736
rect 800 22784 279200 23456
rect 880 22504 279200 22784
rect 800 22376 279200 22504
rect 800 22096 279120 22376
rect 800 21152 279200 22096
rect 800 20872 279120 21152
rect 800 20336 279200 20872
rect 880 20056 279200 20336
rect 800 19928 279200 20056
rect 800 19648 279120 19928
rect 800 18568 279200 19648
rect 800 18288 279120 18568
rect 800 18024 279200 18288
rect 880 17744 279200 18024
rect 800 17344 279200 17744
rect 800 17064 279120 17344
rect 800 15984 279200 17064
rect 800 15704 279120 15984
rect 800 15576 279200 15704
rect 880 15296 279200 15576
rect 800 14760 279200 15296
rect 800 14480 279120 14760
rect 800 13536 279200 14480
rect 800 13256 279120 13536
rect 800 13128 279200 13256
rect 880 12848 279200 13128
rect 800 12176 279200 12848
rect 800 11896 279120 12176
rect 800 10952 279200 11896
rect 800 10816 279120 10952
rect 880 10672 279120 10816
rect 880 10536 279200 10672
rect 800 9592 279200 10536
rect 800 9312 279120 9592
rect 800 8368 279200 9312
rect 880 8088 279120 8368
rect 800 7144 279200 8088
rect 800 6864 279120 7144
rect 800 6056 279200 6864
rect 880 5784 279200 6056
rect 880 5776 279120 5784
rect 800 5504 279120 5776
rect 800 4560 279200 5504
rect 800 4280 279120 4560
rect 800 3608 279200 4280
rect 880 3328 279200 3608
rect 800 3200 279200 3328
rect 800 2920 279120 3200
rect 800 1976 279200 2920
rect 800 1696 279120 1976
rect 800 1296 279200 1696
rect 880 1016 279200 1296
rect 800 752 279200 1016
rect 800 579 279120 752
<< metal4 >>
rect 4208 2128 4528 277488
rect 9208 2128 9528 277488
rect 14208 2128 14528 277488
rect 19208 2128 19528 277488
rect 24208 2128 24528 277488
rect 29208 2128 29528 277488
rect 34208 2128 34528 277488
rect 39208 2128 39528 277488
rect 44208 2128 44528 277488
rect 49208 2128 49528 277488
rect 54208 2128 54528 277488
rect 59208 2128 59528 277488
rect 64208 2128 64528 277488
rect 69208 2128 69528 277488
rect 74208 2128 74528 277488
rect 79208 2128 79528 277488
rect 84208 2128 84528 277488
rect 89208 2128 89528 277488
rect 94208 2128 94528 277488
rect 99208 2128 99528 277488
rect 104208 2128 104528 277488
rect 109208 2128 109528 277488
rect 114208 2128 114528 277488
rect 119208 2128 119528 277488
rect 124208 2128 124528 277488
rect 129208 2128 129528 277488
rect 134208 2128 134528 277488
rect 139208 2128 139528 277488
rect 144208 2128 144528 277488
rect 149208 2128 149528 277488
rect 154208 2128 154528 277488
rect 159208 2128 159528 277488
rect 164208 2128 164528 277488
rect 169208 2128 169528 277488
rect 174208 2128 174528 277488
rect 179208 2128 179528 277488
rect 184208 2128 184528 277488
rect 189208 2128 189528 277488
rect 194208 2128 194528 277488
rect 199208 2128 199528 277488
rect 204208 2128 204528 277488
rect 209208 2128 209528 277488
rect 214208 2128 214528 277488
rect 219208 2128 219528 277488
rect 224208 2128 224528 277488
rect 229208 2128 229528 277488
rect 234208 2128 234528 277488
rect 239208 2128 239528 277488
rect 244208 2128 244528 277488
rect 249208 2128 249528 277488
rect 254208 2128 254528 277488
rect 259208 2128 259528 277488
rect 264208 2128 264528 277488
rect 269208 2128 269528 277488
rect 274208 2128 274528 277488
<< obsm4 >>
rect 66667 2048 69128 277133
rect 69608 2048 74128 277133
rect 74608 2048 79128 277133
rect 79608 2048 84128 277133
rect 84608 2048 89128 277133
rect 89608 2048 94128 277133
rect 94608 2048 99128 277133
rect 99608 2048 104128 277133
rect 104608 2048 109128 277133
rect 109608 2048 114128 277133
rect 114608 2048 119128 277133
rect 119608 2048 124128 277133
rect 124608 2048 129128 277133
rect 129608 2048 134128 277133
rect 134608 2048 139128 277133
rect 139608 2048 144128 277133
rect 144608 2048 149128 277133
rect 149608 2048 154128 277133
rect 154608 2048 159128 277133
rect 159608 2048 164128 277133
rect 164608 2048 169128 277133
rect 169608 2048 174128 277133
rect 174608 2048 179128 277133
rect 179608 2048 184128 277133
rect 184608 2048 189128 277133
rect 189608 2048 194128 277133
rect 194608 2048 199128 277133
rect 199608 2048 204128 277133
rect 204608 2048 209128 277133
rect 209608 2048 214128 277133
rect 214608 2048 219128 277133
rect 219608 2048 224128 277133
rect 224608 2048 229128 277133
rect 229608 2048 234128 277133
rect 234608 2048 239128 277133
rect 239608 2048 244128 277133
rect 244608 2048 249128 277133
rect 249608 2048 254128 277133
rect 254608 2048 257909 277133
rect 66667 1803 257909 2048
<< labels >>
rlabel metal2 s 1030 279200 1086 280000 6 alert_major_o
port 1 nsew signal output
rlabel metal2 s 3146 279200 3202 280000 6 alert_minor_o
port 2 nsew signal output
rlabel metal3 s 279200 102824 280000 102944 6 boot_addr_i[0]
port 3 nsew signal input
rlabel metal2 s 87970 279200 88026 280000 6 boot_addr_i[10]
port 4 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 boot_addr_i[11]
port 5 nsew signal input
rlabel metal3 s 279200 161576 280000 161696 6 boot_addr_i[12]
port 6 nsew signal input
rlabel metal3 s 0 115880 800 116000 6 boot_addr_i[13]
port 7 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 boot_addr_i[14]
port 8 nsew signal input
rlabel metal3 s 279200 175720 280000 175840 6 boot_addr_i[15]
port 9 nsew signal input
rlabel metal2 s 134614 279200 134670 280000 6 boot_addr_i[16]
port 10 nsew signal input
rlabel metal3 s 0 135056 800 135176 6 boot_addr_i[17]
port 11 nsew signal input
rlabel metal3 s 0 139816 800 139936 6 boot_addr_i[18]
port 12 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 boot_addr_i[19]
port 13 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 boot_addr_i[1]
port 14 nsew signal input
rlabel metal3 s 0 144576 800 144696 6 boot_addr_i[20]
port 15 nsew signal input
rlabel metal3 s 279200 202512 280000 202632 6 boot_addr_i[21]
port 16 nsew signal input
rlabel metal3 s 279200 206320 280000 206440 6 boot_addr_i[22]
port 17 nsew signal input
rlabel metal2 s 172794 279200 172850 280000 6 boot_addr_i[23]
port 18 nsew signal input
rlabel metal2 s 183374 279200 183430 280000 6 boot_addr_i[24]
port 19 nsew signal input
rlabel metal2 s 187606 279200 187662 280000 6 boot_addr_i[25]
port 20 nsew signal input
rlabel metal3 s 279200 225496 280000 225616 6 boot_addr_i[26]
port 21 nsew signal input
rlabel metal2 s 193954 279200 194010 280000 6 boot_addr_i[27]
port 22 nsew signal input
rlabel metal3 s 279200 230664 280000 230784 6 boot_addr_i[28]
port 23 nsew signal input
rlabel metal2 s 213550 0 213606 800 6 boot_addr_i[29]
port 24 nsew signal input
rlabel metal3 s 279200 114248 280000 114368 6 boot_addr_i[2]
port 25 nsew signal input
rlabel metal2 s 204626 279200 204682 280000 6 boot_addr_i[30]
port 26 nsew signal input
rlabel metal3 s 279200 239640 280000 239760 6 boot_addr_i[31]
port 27 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 boot_addr_i[3]
port 28 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 boot_addr_i[4]
port 29 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 boot_addr_i[5]
port 30 nsew signal input
rlabel metal3 s 279200 128392 280000 128512 6 boot_addr_i[6]
port 31 nsew signal input
rlabel metal3 s 279200 134784 280000 134904 6 boot_addr_i[7]
port 32 nsew signal input
rlabel metal3 s 279200 143760 280000 143880 6 boot_addr_i[8]
port 33 nsew signal input
rlabel metal2 s 81622 279200 81678 280000 6 boot_addr_i[9]
port 34 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 clk_i
port 35 nsew signal input
rlabel metal3 s 279200 96432 280000 96552 6 core_sleep_o
port 36 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 crash_dump_o[0]
port 37 nsew signal output
rlabel metal3 s 0 261944 800 262064 6 crash_dump_o[100]
port 38 nsew signal output
rlabel metal2 s 273902 0 273958 800 6 crash_dump_o[101]
port 39 nsew signal output
rlabel metal3 s 279200 267656 280000 267776 6 crash_dump_o[102]
port 40 nsew signal output
rlabel metal3 s 0 264256 800 264376 6 crash_dump_o[103]
port 41 nsew signal output
rlabel metal3 s 0 266704 800 266824 6 crash_dump_o[104]
port 42 nsew signal output
rlabel metal2 s 266082 279200 266138 280000 6 crash_dump_o[105]
port 43 nsew signal output
rlabel metal2 s 268198 279200 268254 280000 6 crash_dump_o[106]
port 44 nsew signal output
rlabel metal3 s 0 269152 800 269272 6 crash_dump_o[107]
port 45 nsew signal output
rlabel metal3 s 279200 269016 280000 269136 6 crash_dump_o[108]
port 46 nsew signal output
rlabel metal3 s 279200 270240 280000 270360 6 crash_dump_o[109]
port 47 nsew signal output
rlabel metal3 s 279200 153960 280000 154080 6 crash_dump_o[10]
port 48 nsew signal output
rlabel metal3 s 279200 271600 280000 271720 6 crash_dump_o[110]
port 49 nsew signal output
rlabel metal3 s 0 271464 800 271584 6 crash_dump_o[111]
port 50 nsew signal output
rlabel metal3 s 279200 272824 280000 272944 6 crash_dump_o[112]
port 51 nsew signal output
rlabel metal3 s 279200 274048 280000 274168 6 crash_dump_o[113]
port 52 nsew signal output
rlabel metal3 s 0 273912 800 274032 6 crash_dump_o[114]
port 53 nsew signal output
rlabel metal2 s 270314 279200 270370 280000 6 crash_dump_o[115]
port 54 nsew signal output
rlabel metal2 s 276294 0 276350 800 6 crash_dump_o[116]
port 55 nsew signal output
rlabel metal3 s 279200 275408 280000 275528 6 crash_dump_o[117]
port 56 nsew signal output
rlabel metal3 s 279200 276632 280000 276752 6 crash_dump_o[118]
port 57 nsew signal output
rlabel metal2 s 278686 0 278742 800 6 crash_dump_o[119]
port 58 nsew signal output
rlabel metal2 s 96434 279200 96490 280000 6 crash_dump_o[11]
port 59 nsew signal output
rlabel metal3 s 0 276224 800 276344 6 crash_dump_o[120]
port 60 nsew signal output
rlabel metal3 s 279200 277992 280000 278112 6 crash_dump_o[121]
port 61 nsew signal output
rlabel metal2 s 272430 279200 272486 280000 6 crash_dump_o[122]
port 62 nsew signal output
rlabel metal2 s 274546 279200 274602 280000 6 crash_dump_o[123]
port 63 nsew signal output
rlabel metal2 s 276662 279200 276718 280000 6 crash_dump_o[124]
port 64 nsew signal output
rlabel metal3 s 279200 279216 280000 279336 6 crash_dump_o[125]
port 65 nsew signal output
rlabel metal2 s 278778 279200 278834 280000 6 crash_dump_o[126]
port 66 nsew signal output
rlabel metal3 s 0 278672 800 278792 6 crash_dump_o[127]
port 67 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 crash_dump_o[12]
port 68 nsew signal output
rlabel metal2 s 119710 279200 119766 280000 6 crash_dump_o[13]
port 69 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 crash_dump_o[14]
port 70 nsew signal output
rlabel metal2 s 130382 279200 130438 280000 6 crash_dump_o[15]
port 71 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 crash_dump_o[16]
port 72 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 crash_dump_o[17]
port 73 nsew signal output
rlabel metal2 s 149426 279200 149482 280000 6 crash_dump_o[18]
port 74 nsew signal output
rlabel metal3 s 279200 197344 280000 197464 6 crash_dump_o[19]
port 75 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 crash_dump_o[1]
port 76 nsew signal output
rlabel metal3 s 0 147024 800 147144 6 crash_dump_o[20]
port 77 nsew signal output
rlabel metal3 s 0 158992 800 159112 6 crash_dump_o[21]
port 78 nsew signal output
rlabel metal3 s 279200 207680 280000 207800 6 crash_dump_o[22]
port 79 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 crash_dump_o[23]
port 80 nsew signal output
rlabel metal3 s 279200 211488 280000 211608 6 crash_dump_o[24]
port 81 nsew signal output
rlabel metal3 s 279200 220464 280000 220584 6 crash_dump_o[25]
port 82 nsew signal output
rlabel metal2 s 184570 0 184626 800 6 crash_dump_o[26]
port 83 nsew signal output
rlabel metal3 s 279200 228080 280000 228200 6 crash_dump_o[27]
port 84 nsew signal output
rlabel metal3 s 0 209312 800 209432 6 crash_dump_o[28]
port 85 nsew signal output
rlabel metal3 s 0 221280 800 221400 6 crash_dump_o[29]
port 86 nsew signal output
rlabel metal2 s 34886 279200 34942 280000 6 crash_dump_o[2]
port 87 nsew signal output
rlabel metal2 s 206742 279200 206798 280000 6 crash_dump_o[30]
port 88 nsew signal output
rlabel metal2 s 225602 0 225658 800 6 crash_dump_o[31]
port 89 nsew signal output
rlabel metal3 s 0 233248 800 233368 6 crash_dump_o[32]
port 90 nsew signal output
rlabel metal2 s 235262 0 235318 800 6 crash_dump_o[33]
port 91 nsew signal output
rlabel metal3 s 279200 243448 280000 243568 6 crash_dump_o[34]
port 92 nsew signal output
rlabel metal3 s 279200 244672 280000 244792 6 crash_dump_o[35]
port 93 nsew signal output
rlabel metal2 s 221554 279200 221610 280000 6 crash_dump_o[36]
port 94 nsew signal output
rlabel metal3 s 279200 246032 280000 246152 6 crash_dump_o[37]
port 95 nsew signal output
rlabel metal3 s 279200 247256 280000 247376 6 crash_dump_o[38]
port 96 nsew signal output
rlabel metal2 s 223670 279200 223726 280000 6 crash_dump_o[39]
port 97 nsew signal output
rlabel metal2 s 45558 279200 45614 280000 6 crash_dump_o[3]
port 98 nsew signal output
rlabel metal2 s 225786 279200 225842 280000 6 crash_dump_o[40]
port 99 nsew signal output
rlabel metal3 s 279200 248480 280000 248600 6 crash_dump_o[41]
port 100 nsew signal output
rlabel metal3 s 279200 249840 280000 249960 6 crash_dump_o[42]
port 101 nsew signal output
rlabel metal3 s 0 235560 800 235680 6 crash_dump_o[43]
port 102 nsew signal output
rlabel metal2 s 227902 279200 227958 280000 6 crash_dump_o[44]
port 103 nsew signal output
rlabel metal2 s 230018 279200 230074 280000 6 crash_dump_o[45]
port 104 nsew signal output
rlabel metal2 s 232134 279200 232190 280000 6 crash_dump_o[46]
port 105 nsew signal output
rlabel metal3 s 279200 251064 280000 251184 6 crash_dump_o[47]
port 106 nsew signal output
rlabel metal2 s 237654 0 237710 800 6 crash_dump_o[48]
port 107 nsew signal output
rlabel metal3 s 0 238008 800 238128 6 crash_dump_o[49]
port 108 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 crash_dump_o[4]
port 109 nsew signal output
rlabel metal2 s 234250 279200 234306 280000 6 crash_dump_o[50]
port 110 nsew signal output
rlabel metal2 s 240138 0 240194 800 6 crash_dump_o[51]
port 111 nsew signal output
rlabel metal2 s 236366 279200 236422 280000 6 crash_dump_o[52]
port 112 nsew signal output
rlabel metal3 s 279200 252424 280000 252544 6 crash_dump_o[53]
port 113 nsew signal output
rlabel metal3 s 279200 253648 280000 253768 6 crash_dump_o[54]
port 114 nsew signal output
rlabel metal3 s 279200 254872 280000 254992 6 crash_dump_o[55]
port 115 nsew signal output
rlabel metal2 s 242530 0 242586 800 6 crash_dump_o[56]
port 116 nsew signal output
rlabel metal3 s 0 240320 800 240440 6 crash_dump_o[57]
port 117 nsew signal output
rlabel metal2 s 244922 0 244978 800 6 crash_dump_o[58]
port 118 nsew signal output
rlabel metal3 s 0 242768 800 242888 6 crash_dump_o[59]
port 119 nsew signal output
rlabel metal3 s 0 65696 800 65816 6 crash_dump_o[5]
port 120 nsew signal output
rlabel metal3 s 279200 256232 280000 256352 6 crash_dump_o[60]
port 121 nsew signal output
rlabel metal2 s 238482 279200 238538 280000 6 crash_dump_o[61]
port 122 nsew signal output
rlabel metal3 s 0 245216 800 245336 6 crash_dump_o[62]
port 123 nsew signal output
rlabel metal2 s 240598 279200 240654 280000 6 crash_dump_o[63]
port 124 nsew signal output
rlabel metal3 s 279200 257456 280000 257576 6 crash_dump_o[64]
port 125 nsew signal output
rlabel metal2 s 242806 279200 242862 280000 6 crash_dump_o[65]
port 126 nsew signal output
rlabel metal2 s 247314 0 247370 800 6 crash_dump_o[66]
port 127 nsew signal output
rlabel metal3 s 279200 258816 280000 258936 6 crash_dump_o[67]
port 128 nsew signal output
rlabel metal3 s 0 247528 800 247648 6 crash_dump_o[68]
port 129 nsew signal output
rlabel metal3 s 279200 260040 280000 260160 6 crash_dump_o[69]
port 130 nsew signal output
rlabel metal3 s 279200 129616 280000 129736 6 crash_dump_o[6]
port 131 nsew signal output
rlabel metal3 s 279200 261264 280000 261384 6 crash_dump_o[70]
port 132 nsew signal output
rlabel metal2 s 249706 0 249762 800 6 crash_dump_o[71]
port 133 nsew signal output
rlabel metal3 s 279200 262624 280000 262744 6 crash_dump_o[72]
port 134 nsew signal output
rlabel metal2 s 244922 279200 244978 280000 6 crash_dump_o[73]
port 135 nsew signal output
rlabel metal2 s 252190 0 252246 800 6 crash_dump_o[74]
port 136 nsew signal output
rlabel metal2 s 247038 279200 247094 280000 6 crash_dump_o[75]
port 137 nsew signal output
rlabel metal3 s 0 249976 800 250096 6 crash_dump_o[76]
port 138 nsew signal output
rlabel metal2 s 249154 279200 249210 280000 6 crash_dump_o[77]
port 139 nsew signal output
rlabel metal2 s 254582 0 254638 800 6 crash_dump_o[78]
port 140 nsew signal output
rlabel metal2 s 256974 0 257030 800 6 crash_dump_o[79]
port 141 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 crash_dump_o[7]
port 142 nsew signal output
rlabel metal3 s 0 252288 800 252408 6 crash_dump_o[80]
port 143 nsew signal output
rlabel metal3 s 0 254736 800 254856 6 crash_dump_o[81]
port 144 nsew signal output
rlabel metal2 s 251270 279200 251326 280000 6 crash_dump_o[82]
port 145 nsew signal output
rlabel metal2 s 259366 0 259422 800 6 crash_dump_o[83]
port 146 nsew signal output
rlabel metal2 s 253386 279200 253442 280000 6 crash_dump_o[84]
port 147 nsew signal output
rlabel metal3 s 279200 263848 280000 263968 6 crash_dump_o[85]
port 148 nsew signal output
rlabel metal2 s 255502 279200 255558 280000 6 crash_dump_o[86]
port 149 nsew signal output
rlabel metal3 s 279200 265208 280000 265328 6 crash_dump_o[87]
port 150 nsew signal output
rlabel metal2 s 257618 279200 257674 280000 6 crash_dump_o[88]
port 151 nsew signal output
rlabel metal3 s 279200 266432 280000 266552 6 crash_dump_o[89]
port 152 nsew signal output
rlabel metal3 s 279200 144984 280000 145104 6 crash_dump_o[8]
port 153 nsew signal output
rlabel metal2 s 259734 279200 259790 280000 6 crash_dump_o[90]
port 154 nsew signal output
rlabel metal2 s 261850 0 261906 800 6 crash_dump_o[91]
port 155 nsew signal output
rlabel metal2 s 261850 279200 261906 280000 6 crash_dump_o[92]
port 156 nsew signal output
rlabel metal3 s 0 257184 800 257304 6 crash_dump_o[93]
port 157 nsew signal output
rlabel metal3 s 0 259496 800 259616 6 crash_dump_o[94]
port 158 nsew signal output
rlabel metal2 s 264242 0 264298 800 6 crash_dump_o[95]
port 159 nsew signal output
rlabel metal2 s 266634 0 266690 800 6 crash_dump_o[96]
port 160 nsew signal output
rlabel metal2 s 269026 0 269082 800 6 crash_dump_o[97]
port 161 nsew signal output
rlabel metal2 s 271510 0 271566 800 6 crash_dump_o[98]
port 162 nsew signal output
rlabel metal2 s 263966 279200 264022 280000 6 crash_dump_o[99]
port 163 nsew signal output
rlabel metal3 s 279200 151376 280000 151496 6 crash_dump_o[9]
port 164 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 data_addr_o[0]
port 165 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 data_addr_o[10]
port 166 nsew signal output
rlabel metal3 s 279200 158992 280000 159112 6 data_addr_o[11]
port 167 nsew signal output
rlabel metal3 s 279200 162936 280000 163056 6 data_addr_o[12]
port 168 nsew signal output
rlabel metal3 s 279200 165384 280000 165504 6 data_addr_o[13]
port 169 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 data_addr_o[14]
port 170 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 data_addr_o[15]
port 171 nsew signal output
rlabel metal3 s 279200 180752 280000 180872 6 data_addr_o[16]
port 172 nsew signal output
rlabel metal2 s 138846 279200 138902 280000 6 data_addr_o[17]
port 173 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 data_addr_o[18]
port 174 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 data_addr_o[19]
port 175 nsew signal output
rlabel metal2 s 26422 279200 26478 280000 6 data_addr_o[1]
port 176 nsew signal output
rlabel metal3 s 279200 199928 280000 200048 6 data_addr_o[20]
port 177 nsew signal output
rlabel metal2 s 157890 279200 157946 280000 6 data_addr_o[21]
port 178 nsew signal output
rlabel metal2 s 164330 279200 164386 280000 6 data_addr_o[22]
port 179 nsew signal output
rlabel metal3 s 0 175720 800 175840 6 data_addr_o[23]
port 180 nsew signal output
rlabel metal3 s 279200 212712 280000 212832 6 data_addr_o[24]
port 181 nsew signal output
rlabel metal3 s 0 180480 800 180600 6 data_addr_o[25]
port 182 nsew signal output
rlabel metal2 s 189722 279200 189778 280000 6 data_addr_o[26]
port 183 nsew signal output
rlabel metal2 s 194230 0 194286 800 6 data_addr_o[27]
port 184 nsew signal output
rlabel metal3 s 0 211624 800 211744 6 data_addr_o[28]
port 185 nsew signal output
rlabel metal3 s 0 223592 800 223712 6 data_addr_o[29]
port 186 nsew signal output
rlabel metal2 s 37002 279200 37058 280000 6 data_addr_o[2]
port 187 nsew signal output
rlabel metal3 s 279200 235696 280000 235816 6 data_addr_o[30]
port 188 nsew signal output
rlabel metal3 s 0 230800 800 230920 6 data_addr_o[31]
port 189 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 data_addr_o[3]
port 190 nsew signal output
rlabel metal2 s 54022 279200 54078 280000 6 data_addr_o[4]
port 191 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 data_addr_o[5]
port 192 nsew signal output
rlabel metal3 s 279200 130840 280000 130960 6 data_addr_o[6]
port 193 nsew signal output
rlabel metal3 s 0 84736 800 84856 6 data_addr_o[7]
port 194 nsew signal output
rlabel metal3 s 0 91944 800 92064 6 data_addr_o[8]
port 195 nsew signal output
rlabel metal3 s 0 96704 800 96824 6 data_addr_o[9]
port 196 nsew signal output
rlabel metal2 s 15842 279200 15898 280000 6 data_be_o[0]
port 197 nsew signal output
rlabel metal2 s 28538 279200 28594 280000 6 data_be_o[1]
port 198 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 data_be_o[2]
port 199 nsew signal output
rlabel metal3 s 279200 118056 280000 118176 6 data_be_o[3]
port 200 nsew signal output
rlabel metal2 s 5262 279200 5318 280000 6 data_err_i
port 201 nsew signal input
rlabel metal3 s 0 1096 800 1216 6 data_gnt_i
port 202 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 data_rdata_i[0]
port 203 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 data_rdata_i[10]
port 204 nsew signal input
rlabel metal3 s 279200 160352 280000 160472 6 data_rdata_i[11]
port 205 nsew signal input
rlabel metal2 s 109130 279200 109186 280000 6 data_rdata_i[12]
port 206 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 data_rdata_i[13]
port 207 nsew signal input
rlabel metal3 s 0 120640 800 120760 6 data_rdata_i[14]
port 208 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 data_rdata_i[15]
port 209 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 data_rdata_i[16]
port 210 nsew signal input
rlabel metal3 s 0 137504 800 137624 6 data_rdata_i[17]
port 211 nsew signal input
rlabel metal3 s 279200 188504 280000 188624 6 data_rdata_i[18]
port 212 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 data_rdata_i[19]
port 213 nsew signal input
rlabel metal3 s 279200 107856 280000 107976 6 data_rdata_i[1]
port 214 nsew signal input
rlabel metal3 s 0 149472 800 149592 6 data_rdata_i[20]
port 215 nsew signal input
rlabel metal3 s 0 161440 800 161560 6 data_rdata_i[21]
port 216 nsew signal input
rlabel metal3 s 0 168512 800 168632 6 data_rdata_i[22]
port 217 nsew signal input
rlabel metal3 s 279200 210128 280000 210248 6 data_rdata_i[23]
port 218 nsew signal input
rlabel metal3 s 279200 214072 280000 214192 6 data_rdata_i[24]
port 219 nsew signal input
rlabel metal3 s 0 182928 800 183048 6 data_rdata_i[25]
port 220 nsew signal input
rlabel metal3 s 0 194896 800 195016 6 data_rdata_i[26]
port 221 nsew signal input
rlabel metal2 s 196622 0 196678 800 6 data_rdata_i[27]
port 222 nsew signal input
rlabel metal2 s 206282 0 206338 800 6 data_rdata_i[28]
port 223 nsew signal input
rlabel metal3 s 279200 231888 280000 232008 6 data_rdata_i[29]
port 224 nsew signal input
rlabel metal3 s 279200 115608 280000 115728 6 data_rdata_i[2]
port 225 nsew signal input
rlabel metal2 s 208858 279200 208914 280000 6 data_rdata_i[30]
port 226 nsew signal input
rlabel metal2 s 227994 0 228050 800 6 data_rdata_i[31]
port 227 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 data_rdata_i[3]
port 228 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 data_rdata_i[4]
port 229 nsew signal input
rlabel metal3 s 0 70456 800 70576 6 data_rdata_i[5]
port 230 nsew signal input
rlabel metal2 s 68834 279200 68890 280000 6 data_rdata_i[6]
port 231 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 data_rdata_i[7]
port 232 nsew signal input
rlabel metal3 s 279200 146208 280000 146328 6 data_rdata_i[8]
port 233 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 data_rdata_i[9]
port 234 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 data_rdata_intg_i[0]
port 235 nsew signal input
rlabel metal2 s 30654 279200 30710 280000 6 data_rdata_intg_i[1]
port 236 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 data_rdata_intg_i[2]
port 237 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 data_rdata_intg_i[3]
port 238 nsew signal input
rlabel metal2 s 56138 279200 56194 280000 6 data_rdata_intg_i[4]
port 239 nsew signal input
rlabel metal2 s 60370 279200 60426 280000 6 data_rdata_intg_i[5]
port 240 nsew signal input
rlabel metal3 s 279200 132200 280000 132320 6 data_rdata_intg_i[6]
port 241 nsew signal input
rlabel metal2 s 7378 279200 7434 280000 6 data_req_o
port 242 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 data_rvalid_i
port 243 nsew signal input
rlabel metal2 s 17958 279200 18014 280000 6 data_wdata_intg_o[0]
port 244 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 data_wdata_intg_o[1]
port 245 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 data_wdata_intg_o[2]
port 246 nsew signal output
rlabel metal3 s 0 48832 800 48952 6 data_wdata_intg_o[3]
port 247 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 data_wdata_intg_o[4]
port 248 nsew signal output
rlabel metal3 s 279200 124448 280000 124568 6 data_wdata_intg_o[5]
port 249 nsew signal output
rlabel metal2 s 70950 279200 71006 280000 6 data_wdata_intg_o[6]
port 250 nsew signal output
rlabel metal2 s 20074 279200 20130 280000 6 data_wdata_o[0]
port 251 nsew signal output
rlabel metal3 s 279200 155184 280000 155304 6 data_wdata_o[10]
port 252 nsew signal output
rlabel metal3 s 0 108672 800 108792 6 data_wdata_o[11]
port 253 nsew signal output
rlabel metal2 s 111246 279200 111302 280000 6 data_wdata_o[12]
port 254 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 data_wdata_o[13]
port 255 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 data_wdata_o[14]
port 256 nsew signal output
rlabel metal2 s 132498 279200 132554 280000 6 data_wdata_o[15]
port 257 nsew signal output
rlabel metal3 s 279200 182112 280000 182232 6 data_wdata_o[16]
port 258 nsew signal output
rlabel metal2 s 140962 279200 141018 280000 6 data_wdata_o[17]
port 259 nsew signal output
rlabel metal3 s 279200 189728 280000 189848 6 data_wdata_o[18]
port 260 nsew signal output
rlabel metal3 s 0 142264 800 142384 6 data_wdata_o[19]
port 261 nsew signal output
rlabel metal2 s 32770 279200 32826 280000 6 data_wdata_o[1]
port 262 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 data_wdata_o[20]
port 263 nsew signal output
rlabel metal3 s 279200 203736 280000 203856 6 data_wdata_o[21]
port 264 nsew signal output
rlabel metal2 s 166446 279200 166502 280000 6 data_wdata_o[22]
port 265 nsew signal output
rlabel metal3 s 0 178168 800 178288 6 data_wdata_o[23]
port 266 nsew signal output
rlabel metal3 s 279200 215296 280000 215416 6 data_wdata_o[24]
port 267 nsew signal output
rlabel metal3 s 0 185376 800 185496 6 data_wdata_o[25]
port 268 nsew signal output
rlabel metal3 s 279200 226856 280000 226976 6 data_wdata_o[26]
port 269 nsew signal output
rlabel metal2 s 199106 0 199162 800 6 data_wdata_o[27]
port 270 nsew signal output
rlabel metal3 s 0 214072 800 214192 6 data_wdata_o[28]
port 271 nsew signal output
rlabel metal2 s 215942 0 215998 800 6 data_wdata_o[29]
port 272 nsew signal output
rlabel metal3 s 279200 116832 280000 116952 6 data_wdata_o[2]
port 273 nsew signal output
rlabel metal3 s 0 228352 800 228472 6 data_wdata_o[30]
port 274 nsew signal output
rlabel metal2 s 230478 0 230534 800 6 data_wdata_o[31]
port 275 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 data_wdata_o[3]
port 276 nsew signal output
rlabel metal3 s 0 60800 800 60920 6 data_wdata_o[4]
port 277 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 data_wdata_o[5]
port 278 nsew signal output
rlabel metal3 s 279200 133424 280000 133544 6 data_wdata_o[6]
port 279 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 data_wdata_o[7]
port 280 nsew signal output
rlabel metal2 s 79414 279200 79470 280000 6 data_wdata_o[8]
port 281 nsew signal output
rlabel metal3 s 279200 152600 280000 152720 6 data_wdata_o[9]
port 282 nsew signal output
rlabel metal3 s 279200 97656 280000 97776 6 data_we_o
port 283 nsew signal output
rlabel metal3 s 279200 98880 280000 99000 6 debug_req_i
port 284 nsew signal input
rlabel metal2 s 22190 279200 22246 280000 6 eFPGA_delay_o[0]
port 285 nsew signal output
rlabel metal3 s 279200 109216 280000 109336 6 eFPGA_delay_o[1]
port 286 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 eFPGA_delay_o[2]
port 287 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 eFPGA_delay_o[3]
port 288 nsew signal output
rlabel metal2 s 9494 279200 9550 280000 6 eFPGA_en_o
port 289 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 eFPGA_fpga_done_i
port 290 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 eFPGA_operand_a_o[0]
port 291 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 eFPGA_operand_a_o[10]
port 292 nsew signal output
rlabel metal3 s 0 111120 800 111240 6 eFPGA_operand_a_o[11]
port 293 nsew signal output
rlabel metal3 s 279200 164160 280000 164280 6 eFPGA_operand_a_o[12]
port 294 nsew signal output
rlabel metal3 s 279200 166744 280000 166864 6 eFPGA_operand_a_o[13]
port 295 nsew signal output
rlabel metal3 s 279200 171776 280000 171896 6 eFPGA_operand_a_o[14]
port 296 nsew signal output
rlabel metal3 s 279200 176944 280000 177064 6 eFPGA_operand_a_o[15]
port 297 nsew signal output
rlabel metal3 s 279200 183336 280000 183456 6 eFPGA_operand_a_o[16]
port 298 nsew signal output
rlabel metal2 s 141146 0 141202 800 6 eFPGA_operand_a_o[17]
port 299 nsew signal output
rlabel metal3 s 279200 190952 280000 191072 6 eFPGA_operand_a_o[18]
port 300 nsew signal output
rlabel metal2 s 153198 0 153254 800 6 eFPGA_operand_a_o[19]
port 301 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 eFPGA_operand_a_o[1]
port 302 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 eFPGA_operand_a_o[20]
port 303 nsew signal output
rlabel metal2 s 160006 279200 160062 280000 6 eFPGA_operand_a_o[21]
port 304 nsew signal output
rlabel metal2 s 168562 279200 168618 280000 6 eFPGA_operand_a_o[22]
port 305 nsew signal output
rlabel metal2 s 174910 279200 174966 280000 6 eFPGA_operand_a_o[23]
port 306 nsew signal output
rlabel metal2 s 179786 0 179842 800 6 eFPGA_operand_a_o[24]
port 307 nsew signal output
rlabel metal3 s 0 187688 800 187808 6 eFPGA_operand_a_o[25]
port 308 nsew signal output
rlabel metal2 s 191838 279200 191894 280000 6 eFPGA_operand_a_o[26]
port 309 nsew signal output
rlabel metal2 s 201498 0 201554 800 6 eFPGA_operand_a_o[27]
port 310 nsew signal output
rlabel metal2 s 196070 279200 196126 280000 6 eFPGA_operand_a_o[28]
port 311 nsew signal output
rlabel metal2 s 200302 279200 200358 280000 6 eFPGA_operand_a_o[29]
port 312 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 eFPGA_operand_a_o[2]
port 313 nsew signal output
rlabel metal2 s 220818 0 220874 800 6 eFPGA_operand_a_o[30]
port 314 nsew signal output
rlabel metal2 s 215206 279200 215262 280000 6 eFPGA_operand_a_o[31]
port 315 nsew signal output
rlabel metal2 s 47674 279200 47730 280000 6 eFPGA_operand_a_o[3]
port 316 nsew signal output
rlabel metal3 s 279200 123224 280000 123344 6 eFPGA_operand_a_o[4]
port 317 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 eFPGA_operand_a_o[5]
port 318 nsew signal output
rlabel metal3 s 0 75216 800 75336 6 eFPGA_operand_a_o[6]
port 319 nsew signal output
rlabel metal3 s 279200 136008 280000 136128 6 eFPGA_operand_a_o[7]
port 320 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 eFPGA_operand_a_o[8]
port 321 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 eFPGA_operand_a_o[9]
port 322 nsew signal output
rlabel metal3 s 279200 104048 280000 104168 6 eFPGA_operand_b_o[0]
port 323 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 eFPGA_operand_b_o[10]
port 324 nsew signal output
rlabel metal2 s 98550 279200 98606 280000 6 eFPGA_operand_b_o[11]
port 325 nsew signal output
rlabel metal2 s 113362 279200 113418 280000 6 eFPGA_operand_b_o[12]
port 326 nsew signal output
rlabel metal3 s 279200 167968 280000 168088 6 eFPGA_operand_b_o[13]
port 327 nsew signal output
rlabel metal2 s 124034 279200 124090 280000 6 eFPGA_operand_b_o[14]
port 328 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 eFPGA_operand_b_o[15]
port 329 nsew signal output
rlabel metal2 s 136730 279200 136786 280000 6 eFPGA_operand_b_o[16]
port 330 nsew signal output
rlabel metal2 s 143078 279200 143134 280000 6 eFPGA_operand_b_o[17]
port 331 nsew signal output
rlabel metal3 s 279200 192312 280000 192432 6 eFPGA_operand_b_o[18]
port 332 nsew signal output
rlabel metal2 s 153658 279200 153714 280000 6 eFPGA_operand_b_o[19]
port 333 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 eFPGA_operand_b_o[1]
port 334 nsew signal output
rlabel metal2 s 165250 0 165306 800 6 eFPGA_operand_b_o[20]
port 335 nsew signal output
rlabel metal3 s 0 163752 800 163872 6 eFPGA_operand_b_o[21]
port 336 nsew signal output
rlabel metal2 s 170678 279200 170734 280000 6 eFPGA_operand_b_o[22]
port 337 nsew signal output
rlabel metal2 s 177026 279200 177082 280000 6 eFPGA_operand_b_o[23]
port 338 nsew signal output
rlabel metal3 s 279200 216520 280000 216640 6 eFPGA_operand_b_o[24]
port 339 nsew signal output
rlabel metal3 s 0 190136 800 190256 6 eFPGA_operand_b_o[25]
port 340 nsew signal output
rlabel metal3 s 0 197344 800 197464 6 eFPGA_operand_b_o[26]
port 341 nsew signal output
rlabel metal2 s 203890 0 203946 800 6 eFPGA_operand_b_o[27]
port 342 nsew signal output
rlabel metal3 s 0 216384 800 216504 6 eFPGA_operand_b_o[28]
port 343 nsew signal output
rlabel metal2 s 218334 0 218390 800 6 eFPGA_operand_b_o[29]
port 344 nsew signal output
rlabel metal2 s 39118 279200 39174 280000 6 eFPGA_operand_b_o[2]
port 345 nsew signal output
rlabel metal2 s 210974 279200 211030 280000 6 eFPGA_operand_b_o[30]
port 346 nsew signal output
rlabel metal2 s 217322 279200 217378 280000 6 eFPGA_operand_b_o[31]
port 347 nsew signal output
rlabel metal3 s 279200 119416 280000 119536 6 eFPGA_operand_b_o[3]
port 348 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 eFPGA_operand_b_o[4]
port 349 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 eFPGA_operand_b_o[5]
port 350 nsew signal output
rlabel metal3 s 0 77664 800 77784 6 eFPGA_operand_b_o[6]
port 351 nsew signal output
rlabel metal3 s 279200 137232 280000 137352 6 eFPGA_operand_b_o[7]
port 352 nsew signal output
rlabel metal3 s 279200 147568 280000 147688 6 eFPGA_operand_b_o[8]
port 353 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 eFPGA_operand_b_o[9]
port 354 nsew signal output
rlabel metal2 s 24306 279200 24362 280000 6 eFPGA_operator_o[0]
port 355 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 eFPGA_operator_o[1]
port 356 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 eFPGA_result_a_i[0]
port 357 nsew signal input
rlabel metal2 s 90086 279200 90142 280000 6 eFPGA_result_a_i[10]
port 358 nsew signal input
rlabel metal2 s 100666 279200 100722 280000 6 eFPGA_result_a_i[11]
port 359 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 eFPGA_result_a_i[12]
port 360 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 eFPGA_result_a_i[13]
port 361 nsew signal input
rlabel metal3 s 279200 173136 280000 173256 6 eFPGA_result_a_i[14]
port 362 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 eFPGA_result_a_i[15]
port 363 nsew signal input
rlabel metal3 s 279200 184560 280000 184680 6 eFPGA_result_a_i[16]
port 364 nsew signal input
rlabel metal2 s 145194 279200 145250 280000 6 eFPGA_result_a_i[17]
port 365 nsew signal input
rlabel metal3 s 279200 193536 280000 193656 6 eFPGA_result_a_i[18]
port 366 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 eFPGA_result_a_i[19]
port 367 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 eFPGA_result_a_i[1]
port 368 nsew signal input
rlabel metal3 s 279200 201288 280000 201408 6 eFPGA_result_a_i[20]
port 369 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 eFPGA_result_a_i[21]
port 370 nsew signal input
rlabel metal3 s 0 170960 800 171080 6 eFPGA_result_a_i[22]
port 371 nsew signal input
rlabel metal2 s 179142 279200 179198 280000 6 eFPGA_result_a_i[23]
port 372 nsew signal input
rlabel metal2 s 185490 279200 185546 280000 6 eFPGA_result_a_i[24]
port 373 nsew signal input
rlabel metal3 s 279200 221688 280000 221808 6 eFPGA_result_a_i[25]
port 374 nsew signal input
rlabel metal3 s 0 199656 800 199776 6 eFPGA_result_a_i[26]
port 375 nsew signal input
rlabel metal3 s 0 202104 800 202224 6 eFPGA_result_a_i[27]
port 376 nsew signal input
rlabel metal3 s 0 218832 800 218952 6 eFPGA_result_a_i[28]
port 377 nsew signal input
rlabel metal3 s 279200 233248 280000 233368 6 eFPGA_result_a_i[29]
port 378 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 eFPGA_result_a_i[2]
port 379 nsew signal input
rlabel metal2 s 223210 0 223266 800 6 eFPGA_result_a_i[30]
port 380 nsew signal input
rlabel metal2 s 232870 0 232926 800 6 eFPGA_result_a_i[31]
port 381 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 eFPGA_result_a_i[3]
port 382 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 eFPGA_result_a_i[4]
port 383 nsew signal input
rlabel metal3 s 279200 125808 280000 125928 6 eFPGA_result_a_i[5]
port 384 nsew signal input
rlabel metal2 s 73066 279200 73122 280000 6 eFPGA_result_a_i[6]
port 385 nsew signal input
rlabel metal3 s 279200 138592 280000 138712 6 eFPGA_result_a_i[7]
port 386 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 eFPGA_result_a_i[8]
port 387 nsew signal input
rlabel metal3 s 0 101600 800 101720 6 eFPGA_result_a_i[9]
port 388 nsew signal input
rlabel metal3 s 279200 105272 280000 105392 6 eFPGA_result_b_i[0]
port 389 nsew signal input
rlabel metal2 s 92202 279200 92258 280000 6 eFPGA_result_b_i[10]
port 390 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 eFPGA_result_b_i[11]
port 391 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 eFPGA_result_b_i[12]
port 392 nsew signal input
rlabel metal2 s 121918 279200 121974 280000 6 eFPGA_result_b_i[13]
port 393 nsew signal input
rlabel metal2 s 126150 279200 126206 280000 6 eFPGA_result_b_i[14]
port 394 nsew signal input
rlabel metal3 s 279200 178168 280000 178288 6 eFPGA_result_b_i[15]
port 395 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 eFPGA_result_b_i[16]
port 396 nsew signal input
rlabel metal3 s 279200 185920 280000 186040 6 eFPGA_result_b_i[17]
port 397 nsew signal input
rlabel metal3 s 279200 194896 280000 195016 6 eFPGA_result_b_i[18]
port 398 nsew signal input
rlabel metal3 s 279200 198704 280000 198824 6 eFPGA_result_b_i[19]
port 399 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 eFPGA_result_b_i[1]
port 400 nsew signal input
rlabel metal3 s 0 151784 800 151904 6 eFPGA_result_b_i[20]
port 401 nsew signal input
rlabel metal2 s 162214 279200 162270 280000 6 eFPGA_result_b_i[21]
port 402 nsew signal input
rlabel metal3 s 0 173408 800 173528 6 eFPGA_result_b_i[22]
port 403 nsew signal input
rlabel metal2 s 181258 279200 181314 280000 6 eFPGA_result_b_i[23]
port 404 nsew signal input
rlabel metal3 s 279200 217880 280000 218000 6 eFPGA_result_b_i[24]
port 405 nsew signal input
rlabel metal3 s 0 192448 800 192568 6 eFPGA_result_b_i[25]
port 406 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 eFPGA_result_b_i[26]
port 407 nsew signal input
rlabel metal3 s 279200 229304 280000 229424 6 eFPGA_result_b_i[27]
port 408 nsew signal input
rlabel metal2 s 198186 279200 198242 280000 6 eFPGA_result_b_i[28]
port 409 nsew signal input
rlabel metal3 s 279200 234472 280000 234592 6 eFPGA_result_b_i[29]
port 410 nsew signal input
rlabel metal2 s 41326 279200 41382 280000 6 eFPGA_result_b_i[2]
port 411 nsew signal input
rlabel metal3 s 279200 237056 280000 237176 6 eFPGA_result_b_i[30]
port 412 nsew signal input
rlabel metal2 s 219438 279200 219494 280000 6 eFPGA_result_b_i[31]
port 413 nsew signal input
rlabel metal3 s 279200 120640 280000 120760 6 eFPGA_result_b_i[3]
port 414 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 eFPGA_result_b_i[4]
port 415 nsew signal input
rlabel metal2 s 62486 279200 62542 280000 6 eFPGA_result_b_i[5]
port 416 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 eFPGA_result_b_i[6]
port 417 nsew signal input
rlabel metal3 s 279200 139816 280000 139936 6 eFPGA_result_b_i[7]
port 418 nsew signal input
rlabel metal3 s 279200 148792 280000 148912 6 eFPGA_result_b_i[8]
port 419 nsew signal input
rlabel metal2 s 83738 279200 83794 280000 6 eFPGA_result_b_i[9]
port 420 nsew signal input
rlabel metal3 s 279200 106632 280000 106752 6 eFPGA_result_c_i[0]
port 421 nsew signal input
rlabel metal3 s 279200 156544 280000 156664 6 eFPGA_result_c_i[10]
port 422 nsew signal input
rlabel metal2 s 102782 279200 102838 280000 6 eFPGA_result_c_i[11]
port 423 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 eFPGA_result_c_i[12]
port 424 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 eFPGA_result_c_i[13]
port 425 nsew signal input
rlabel metal3 s 279200 174360 280000 174480 6 eFPGA_result_c_i[14]
port 426 nsew signal input
rlabel metal3 s 279200 179528 280000 179648 6 eFPGA_result_c_i[15]
port 427 nsew signal input
rlabel metal3 s 0 130296 800 130416 6 eFPGA_result_c_i[16]
port 428 nsew signal input
rlabel metal3 s 279200 187144 280000 187264 6 eFPGA_result_c_i[17]
port 429 nsew signal input
rlabel metal3 s 279200 196120 280000 196240 6 eFPGA_result_c_i[18]
port 430 nsew signal input
rlabel metal2 s 155774 279200 155830 280000 6 eFPGA_result_c_i[19]
port 431 nsew signal input
rlabel metal3 s 279200 110440 280000 110560 6 eFPGA_result_c_i[1]
port 432 nsew signal input
rlabel metal3 s 0 154232 800 154352 6 eFPGA_result_c_i[20]
port 433 nsew signal input
rlabel metal3 s 279200 205096 280000 205216 6 eFPGA_result_c_i[21]
port 434 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 eFPGA_result_c_i[22]
port 435 nsew signal input
rlabel metal2 s 174910 0 174966 800 6 eFPGA_result_c_i[23]
port 436 nsew signal input
rlabel metal2 s 182178 0 182234 800 6 eFPGA_result_c_i[24]
port 437 nsew signal input
rlabel metal3 s 279200 222912 280000 223032 6 eFPGA_result_c_i[25]
port 438 nsew signal input
rlabel metal2 s 189446 0 189502 800 6 eFPGA_result_c_i[26]
port 439 nsew signal input
rlabel metal3 s 0 204416 800 204536 6 eFPGA_result_c_i[27]
port 440 nsew signal input
rlabel metal2 s 208766 0 208822 800 6 eFPGA_result_c_i[28]
port 441 nsew signal input
rlabel metal3 s 0 226040 800 226160 6 eFPGA_result_c_i[29]
port 442 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 eFPGA_result_c_i[2]
port 443 nsew signal input
rlabel metal3 s 279200 238280 280000 238400 6 eFPGA_result_c_i[30]
port 444 nsew signal input
rlabel metal3 s 279200 240864 280000 240984 6 eFPGA_result_c_i[31]
port 445 nsew signal input
rlabel metal2 s 49790 279200 49846 280000 6 eFPGA_result_c_i[3]
port 446 nsew signal input
rlabel metal2 s 58254 279200 58310 280000 6 eFPGA_result_c_i[4]
port 447 nsew signal input
rlabel metal2 s 64602 279200 64658 280000 6 eFPGA_result_c_i[5]
port 448 nsew signal input
rlabel metal2 s 75182 279200 75238 280000 6 eFPGA_result_c_i[6]
port 449 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 eFPGA_result_c_i[7]
port 450 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 eFPGA_result_c_i[8]
port 451 nsew signal input
rlabel metal2 s 85854 279200 85910 280000 6 eFPGA_result_c_i[9]
port 452 nsew signal input
rlabel metal2 s 11610 279200 11666 280000 6 eFPGA_write_strobe_o
port 453 nsew signal output
rlabel metal3 s 279200 100240 280000 100360 6 fetch_enable_i
port 454 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 hart_id_i[0]
port 455 nsew signal input
rlabel metal3 s 279200 157768 280000 157888 6 hart_id_i[10]
port 456 nsew signal input
rlabel metal2 s 104898 279200 104954 280000 6 hart_id_i[11]
port 457 nsew signal input
rlabel metal2 s 115478 279200 115534 280000 6 hart_id_i[12]
port 458 nsew signal input
rlabel metal3 s 279200 169328 280000 169448 6 hart_id_i[13]
port 459 nsew signal input
rlabel metal2 s 128266 279200 128322 280000 6 hart_id_i[14]
port 460 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 hart_id_i[15]
port 461 nsew signal input
rlabel metal3 s 0 132608 800 132728 6 hart_id_i[16]
port 462 nsew signal input
rlabel metal2 s 147310 279200 147366 280000 6 hart_id_i[17]
port 463 nsew signal input
rlabel metal2 s 151542 279200 151598 280000 6 hart_id_i[18]
port 464 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 hart_id_i[19]
port 465 nsew signal input
rlabel metal3 s 279200 111664 280000 111784 6 hart_id_i[1]
port 466 nsew signal input
rlabel metal3 s 0 156544 800 156664 6 hart_id_i[20]
port 467 nsew signal input
rlabel metal3 s 0 166200 800 166320 6 hart_id_i[21]
port 468 nsew signal input
rlabel metal3 s 279200 208904 280000 209024 6 hart_id_i[22]
port 469 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 hart_id_i[23]
port 470 nsew signal input
rlabel metal3 s 279200 219104 280000 219224 6 hart_id_i[24]
port 471 nsew signal input
rlabel metal3 s 279200 224272 280000 224392 6 hart_id_i[25]
port 472 nsew signal input
rlabel metal2 s 191838 0 191894 800 6 hart_id_i[26]
port 473 nsew signal input
rlabel metal3 s 0 206864 800 206984 6 hart_id_i[27]
port 474 nsew signal input
rlabel metal2 s 211158 0 211214 800 6 hart_id_i[28]
port 475 nsew signal input
rlabel metal2 s 202510 279200 202566 280000 6 hart_id_i[29]
port 476 nsew signal input
rlabel metal2 s 43442 279200 43498 280000 6 hart_id_i[2]
port 477 nsew signal input
rlabel metal2 s 213090 279200 213146 280000 6 hart_id_i[30]
port 478 nsew signal input
rlabel metal3 s 279200 242088 280000 242208 6 hart_id_i[31]
port 479 nsew signal input
rlabel metal2 s 51906 279200 51962 280000 6 hart_id_i[3]
port 480 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 hart_id_i[4]
port 481 nsew signal input
rlabel metal3 s 279200 127032 280000 127152 6 hart_id_i[5]
port 482 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 hart_id_i[6]
port 483 nsew signal input
rlabel metal3 s 279200 141176 280000 141296 6 hart_id_i[7]
port 484 nsew signal input
rlabel metal3 s 279200 150152 280000 150272 6 hart_id_i[8]
port 485 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 hart_id_i[9]
port 486 nsew signal input
rlabel metal3 s 279200 5584 280000 5704 6 instr_addr_o[0]
port 487 nsew signal output
rlabel metal3 s 279200 40128 280000 40248 6 instr_addr_o[10]
port 488 nsew signal output
rlabel metal3 s 279200 42712 280000 42832 6 instr_addr_o[11]
port 489 nsew signal output
rlabel metal3 s 279200 45296 280000 45416 6 instr_addr_o[12]
port 490 nsew signal output
rlabel metal3 s 279200 47744 280000 47864 6 instr_addr_o[13]
port 491 nsew signal output
rlabel metal3 s 279200 50328 280000 50448 6 instr_addr_o[14]
port 492 nsew signal output
rlabel metal3 s 279200 52912 280000 53032 6 instr_addr_o[15]
port 493 nsew signal output
rlabel metal3 s 279200 55496 280000 55616 6 instr_addr_o[16]
port 494 nsew signal output
rlabel metal3 s 279200 58080 280000 58200 6 instr_addr_o[17]
port 495 nsew signal output
rlabel metal3 s 279200 60528 280000 60648 6 instr_addr_o[18]
port 496 nsew signal output
rlabel metal3 s 279200 63112 280000 63232 6 instr_addr_o[19]
port 497 nsew signal output
rlabel metal3 s 279200 9392 280000 9512 6 instr_addr_o[1]
port 498 nsew signal output
rlabel metal3 s 279200 65696 280000 65816 6 instr_addr_o[20]
port 499 nsew signal output
rlabel metal3 s 279200 68280 280000 68400 6 instr_addr_o[21]
port 500 nsew signal output
rlabel metal3 s 279200 70864 280000 70984 6 instr_addr_o[22]
port 501 nsew signal output
rlabel metal3 s 279200 73312 280000 73432 6 instr_addr_o[23]
port 502 nsew signal output
rlabel metal3 s 279200 75896 280000 76016 6 instr_addr_o[24]
port 503 nsew signal output
rlabel metal3 s 279200 78480 280000 78600 6 instr_addr_o[25]
port 504 nsew signal output
rlabel metal3 s 279200 81064 280000 81184 6 instr_addr_o[26]
port 505 nsew signal output
rlabel metal3 s 279200 83648 280000 83768 6 instr_addr_o[27]
port 506 nsew signal output
rlabel metal3 s 279200 86096 280000 86216 6 instr_addr_o[28]
port 507 nsew signal output
rlabel metal3 s 279200 88680 280000 88800 6 instr_addr_o[29]
port 508 nsew signal output
rlabel metal3 s 279200 13336 280000 13456 6 instr_addr_o[2]
port 509 nsew signal output
rlabel metal3 s 279200 91264 280000 91384 6 instr_addr_o[30]
port 510 nsew signal output
rlabel metal3 s 279200 93848 280000 93968 6 instr_addr_o[31]
port 511 nsew signal output
rlabel metal3 s 279200 17144 280000 17264 6 instr_addr_o[3]
port 512 nsew signal output
rlabel metal3 s 279200 20952 280000 21072 6 instr_addr_o[4]
port 513 nsew signal output
rlabel metal3 s 279200 24760 280000 24880 6 instr_addr_o[5]
port 514 nsew signal output
rlabel metal3 s 279200 28568 280000 28688 6 instr_addr_o[6]
port 515 nsew signal output
rlabel metal3 s 279200 32512 280000 32632 6 instr_addr_o[7]
port 516 nsew signal output
rlabel metal3 s 279200 34960 280000 35080 6 instr_addr_o[8]
port 517 nsew signal output
rlabel metal3 s 279200 37544 280000 37664 6 instr_addr_o[9]
port 518 nsew signal output
rlabel metal3 s 279200 552 280000 672 6 instr_err_i
port 519 nsew signal input
rlabel metal3 s 279200 1776 280000 1896 6 instr_gnt_i
port 520 nsew signal input
rlabel metal3 s 279200 6944 280000 7064 6 instr_rdata_i[0]
port 521 nsew signal input
rlabel metal3 s 279200 41352 280000 41472 6 instr_rdata_i[10]
port 522 nsew signal input
rlabel metal3 s 279200 43936 280000 44056 6 instr_rdata_i[11]
port 523 nsew signal input
rlabel metal3 s 279200 46520 280000 46640 6 instr_rdata_i[12]
port 524 nsew signal input
rlabel metal3 s 279200 49104 280000 49224 6 instr_rdata_i[13]
port 525 nsew signal input
rlabel metal3 s 279200 51688 280000 51808 6 instr_rdata_i[14]
port 526 nsew signal input
rlabel metal3 s 279200 54136 280000 54256 6 instr_rdata_i[15]
port 527 nsew signal input
rlabel metal3 s 279200 56720 280000 56840 6 instr_rdata_i[16]
port 528 nsew signal input
rlabel metal3 s 279200 59304 280000 59424 6 instr_rdata_i[17]
port 529 nsew signal input
rlabel metal3 s 279200 61888 280000 62008 6 instr_rdata_i[18]
port 530 nsew signal input
rlabel metal3 s 279200 64472 280000 64592 6 instr_rdata_i[19]
port 531 nsew signal input
rlabel metal3 s 279200 10752 280000 10872 6 instr_rdata_i[1]
port 532 nsew signal input
rlabel metal3 s 279200 66920 280000 67040 6 instr_rdata_i[20]
port 533 nsew signal input
rlabel metal3 s 279200 69504 280000 69624 6 instr_rdata_i[21]
port 534 nsew signal input
rlabel metal3 s 279200 72088 280000 72208 6 instr_rdata_i[22]
port 535 nsew signal input
rlabel metal3 s 279200 74672 280000 74792 6 instr_rdata_i[23]
port 536 nsew signal input
rlabel metal3 s 279200 77256 280000 77376 6 instr_rdata_i[24]
port 537 nsew signal input
rlabel metal3 s 279200 79704 280000 79824 6 instr_rdata_i[25]
port 538 nsew signal input
rlabel metal3 s 279200 82288 280000 82408 6 instr_rdata_i[26]
port 539 nsew signal input
rlabel metal3 s 279200 84872 280000 84992 6 instr_rdata_i[27]
port 540 nsew signal input
rlabel metal3 s 279200 87456 280000 87576 6 instr_rdata_i[28]
port 541 nsew signal input
rlabel metal3 s 279200 90040 280000 90160 6 instr_rdata_i[29]
port 542 nsew signal input
rlabel metal3 s 279200 14560 280000 14680 6 instr_rdata_i[2]
port 543 nsew signal input
rlabel metal3 s 279200 92488 280000 92608 6 instr_rdata_i[30]
port 544 nsew signal input
rlabel metal3 s 279200 95072 280000 95192 6 instr_rdata_i[31]
port 545 nsew signal input
rlabel metal3 s 279200 18368 280000 18488 6 instr_rdata_i[3]
port 546 nsew signal input
rlabel metal3 s 279200 22176 280000 22296 6 instr_rdata_i[4]
port 547 nsew signal input
rlabel metal3 s 279200 26120 280000 26240 6 instr_rdata_i[5]
port 548 nsew signal input
rlabel metal3 s 279200 29928 280000 30048 6 instr_rdata_i[6]
port 549 nsew signal input
rlabel metal3 s 279200 33736 280000 33856 6 instr_rdata_i[7]
port 550 nsew signal input
rlabel metal3 s 279200 36320 280000 36440 6 instr_rdata_i[8]
port 551 nsew signal input
rlabel metal3 s 279200 38904 280000 39024 6 instr_rdata_i[9]
port 552 nsew signal input
rlabel metal3 s 279200 8168 280000 8288 6 instr_rdata_intg_i[0]
port 553 nsew signal input
rlabel metal3 s 279200 11976 280000 12096 6 instr_rdata_intg_i[1]
port 554 nsew signal input
rlabel metal3 s 279200 15784 280000 15904 6 instr_rdata_intg_i[2]
port 555 nsew signal input
rlabel metal3 s 279200 19728 280000 19848 6 instr_rdata_intg_i[3]
port 556 nsew signal input
rlabel metal3 s 279200 23536 280000 23656 6 instr_rdata_intg_i[4]
port 557 nsew signal input
rlabel metal3 s 279200 27344 280000 27464 6 instr_rdata_intg_i[5]
port 558 nsew signal input
rlabel metal3 s 279200 31152 280000 31272 6 instr_rdata_intg_i[6]
port 559 nsew signal input
rlabel metal3 s 279200 3000 280000 3120 6 instr_req_o
port 560 nsew signal output
rlabel metal3 s 279200 4360 280000 4480 6 instr_rvalid_i
port 561 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 irq_external_i
port 562 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 irq_fast_i[0]
port 563 nsew signal input
rlabel metal2 s 94318 279200 94374 280000 6 irq_fast_i[10]
port 564 nsew signal input
rlabel metal2 s 107014 279200 107070 280000 6 irq_fast_i[11]
port 565 nsew signal input
rlabel metal2 s 117594 279200 117650 280000 6 irq_fast_i[12]
port 566 nsew signal input
rlabel metal3 s 279200 170552 280000 170672 6 irq_fast_i[13]
port 567 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 irq_fast_i[14]
port 568 nsew signal input
rlabel metal3 s 279200 113024 280000 113144 6 irq_fast_i[1]
port 569 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 irq_fast_i[2]
port 570 nsew signal input
rlabel metal3 s 279200 122000 280000 122120 6 irq_fast_i[3]
port 571 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 irq_fast_i[4]
port 572 nsew signal input
rlabel metal2 s 66718 279200 66774 280000 6 irq_fast_i[5]
port 573 nsew signal input
rlabel metal2 s 77298 279200 77354 280000 6 irq_fast_i[6]
port 574 nsew signal input
rlabel metal3 s 279200 142400 280000 142520 6 irq_fast_i[7]
port 575 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 irq_fast_i[8]
port 576 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 irq_fast_i[9]
port 577 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 irq_nm_i
port 578 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 irq_software_i
port 579 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 irq_timer_i
port 580 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 ram_cfg_i
port 581 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 rst_ni
port 582 nsew signal input
rlabel metal3 s 279200 101464 280000 101584 6 scan_rst_ni
port 583 nsew signal input
rlabel metal2 s 13726 279200 13782 280000 6 test_en_i
port 584 nsew signal input
rlabel metal4 s 4208 2128 4528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 14208 2128 14528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 24208 2128 24528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 34208 2128 34528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 44208 2128 44528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 54208 2128 54528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 64208 2128 64528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 74208 2128 74528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 84208 2128 84528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 94208 2128 94528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 104208 2128 104528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 114208 2128 114528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 124208 2128 124528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 134208 2128 134528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 144208 2128 144528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 154208 2128 154528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 164208 2128 164528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 174208 2128 174528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 184208 2128 184528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 194208 2128 194528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 204208 2128 204528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 214208 2128 214528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 224208 2128 224528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 234208 2128 234528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 244208 2128 244528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 254208 2128 254528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 264208 2128 264528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 274208 2128 274528 277488 6 vccd1
port 585 nsew power input
rlabel metal4 s 9208 2128 9528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 19208 2128 19528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 29208 2128 29528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 39208 2128 39528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 49208 2128 49528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 59208 2128 59528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 69208 2128 69528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 79208 2128 79528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 89208 2128 89528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 99208 2128 99528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 109208 2128 109528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 119208 2128 119528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 129208 2128 129528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 139208 2128 139528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 149208 2128 149528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 159208 2128 159528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 169208 2128 169528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 179208 2128 179528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 189208 2128 189528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 199208 2128 199528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 209208 2128 209528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 219208 2128 219528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 229208 2128 229528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 239208 2128 239528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 249208 2128 249528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 259208 2128 259528 277488 6 vssd1
port 586 nsew ground input
rlabel metal4 s 269208 2128 269528 277488 6 vssd1
port 586 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 280000 280000
string LEFview TRUE
string GDS_FILE /project/openlane/ibex_top/runs/ibex_top/results/magic/ibex_top.gds
string GDS_END 110642514
string GDS_START 1758614
<< end >>

