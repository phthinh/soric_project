VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO crypto_core
  CLASS BLOCK ;
  FOREIGN crypto_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 900.000 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END clk_i
  PIN data_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END data_addr_o[0]
  PIN data_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END data_addr_o[12]
  PIN data_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END data_addr_o[13]
  PIN data_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END data_addr_o[14]
  PIN data_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END data_addr_o[15]
  PIN data_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END data_addr_o[16]
  PIN data_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END data_addr_o[17]
  PIN data_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END data_addr_o[18]
  PIN data_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END data_addr_o[19]
  PIN data_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END data_addr_o[20]
  PIN data_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END data_addr_o[21]
  PIN data_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 0.000 665.070 4.000 ;
    END
  END data_addr_o[22]
  PIN data_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END data_addr_o[23]
  PIN data_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 0.000 712.910 4.000 ;
    END
  END data_addr_o[24]
  PIN data_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 0.000 736.830 4.000 ;
    END
  END data_addr_o[25]
  PIN data_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 4.000 ;
    END
  END data_addr_o[26]
  PIN data_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 0.000 784.670 4.000 ;
    END
  END data_addr_o[27]
  PIN data_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END data_addr_o[28]
  PIN data_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.230 0.000 832.510 4.000 ;
    END
  END data_addr_o[29]
  PIN data_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 0.000 856.430 4.000 ;
    END
  END data_addr_o[30]
  PIN data_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.070 0.000 880.350 4.000 ;
    END
  END data_addr_o[31]
  PIN data_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END data_addr_o[9]
  PIN data_be_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END data_be_o[0]
  PIN data_be_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END data_be_o[1]
  PIN data_be_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END data_be_o[2]
  PIN data_be_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END data_be_o[3]
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END data_gnt_i
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END data_rdata_i[0]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 4.000 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 0.000 696.810 4.000 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 0.000 816.410 4.000 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 0.000 840.330 4.000 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 0.000 864.250 4.000 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 0.000 888.170 4.000 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END data_rdata_i[9]
  PIN data_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END data_req_o
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END data_rvalid_i
  PIN data_wdata_intg_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END data_wdata_intg_o[0]
  PIN data_wdata_intg_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END data_wdata_intg_o[1]
  PIN data_wdata_intg_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END data_wdata_intg_o[2]
  PIN data_wdata_intg_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END data_wdata_intg_o[3]
  PIN data_wdata_intg_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END data_wdata_intg_o[4]
  PIN data_wdata_intg_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END data_wdata_intg_o[5]
  PIN data_wdata_intg_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 4.000 ;
    END
  END data_wdata_intg_o[6]
  PIN data_wdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END data_wdata_o[0]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 0.000 609.410 4.000 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 0.000 681.170 4.000 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 4.000 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 4.000 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 0.000 824.230 4.000 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.870 0.000 848.150 4.000 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END data_wdata_o[9]
  PIN data_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END data_we_o
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 879.960 900.000 880.560 ;
    END
  END debug_req_i
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 892.880 900.000 893.480 ;
    END
  END fetch_enable_i
  PIN instr_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 44.920 900.000 45.520 ;
    END
  END instr_addr_o[0]
  PIN instr_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 306.040 900.000 306.640 ;
    END
  END instr_addr_o[10]
  PIN instr_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 331.880 900.000 332.480 ;
    END
  END instr_addr_o[11]
  PIN instr_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 358.400 900.000 359.000 ;
    END
  END instr_addr_o[12]
  PIN instr_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 384.240 900.000 384.840 ;
    END
  END instr_addr_o[13]
  PIN instr_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 410.080 900.000 410.680 ;
    END
  END instr_addr_o[14]
  PIN instr_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 436.600 900.000 437.200 ;
    END
  END instr_addr_o[15]
  PIN instr_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 462.440 900.000 463.040 ;
    END
  END instr_addr_o[16]
  PIN instr_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 488.280 900.000 488.880 ;
    END
  END instr_addr_o[17]
  PIN instr_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 514.800 900.000 515.400 ;
    END
  END instr_addr_o[18]
  PIN instr_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 540.640 900.000 541.240 ;
    END
  END instr_addr_o[19]
  PIN instr_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 70.760 900.000 71.360 ;
    END
  END instr_addr_o[1]
  PIN instr_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 567.160 900.000 567.760 ;
    END
  END instr_addr_o[20]
  PIN instr_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 593.000 900.000 593.600 ;
    END
  END instr_addr_o[21]
  PIN instr_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 618.840 900.000 619.440 ;
    END
  END instr_addr_o[22]
  PIN instr_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 645.360 900.000 645.960 ;
    END
  END instr_addr_o[23]
  PIN instr_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 671.200 900.000 671.800 ;
    END
  END instr_addr_o[24]
  PIN instr_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 697.040 900.000 697.640 ;
    END
  END instr_addr_o[25]
  PIN instr_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 723.560 900.000 724.160 ;
    END
  END instr_addr_o[26]
  PIN instr_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 749.400 900.000 750.000 ;
    END
  END instr_addr_o[27]
  PIN instr_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 775.920 900.000 776.520 ;
    END
  END instr_addr_o[28]
  PIN instr_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 801.760 900.000 802.360 ;
    END
  END instr_addr_o[29]
  PIN instr_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 97.280 900.000 97.880 ;
    END
  END instr_addr_o[2]
  PIN instr_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 827.600 900.000 828.200 ;
    END
  END instr_addr_o[30]
  PIN instr_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 854.120 900.000 854.720 ;
    END
  END instr_addr_o[31]
  PIN instr_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 123.120 900.000 123.720 ;
    END
  END instr_addr_o[3]
  PIN instr_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 149.640 900.000 150.240 ;
    END
  END instr_addr_o[4]
  PIN instr_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 175.480 900.000 176.080 ;
    END
  END instr_addr_o[5]
  PIN instr_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 201.320 900.000 201.920 ;
    END
  END instr_addr_o[6]
  PIN instr_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 227.840 900.000 228.440 ;
    END
  END instr_addr_o[7]
  PIN instr_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 253.680 900.000 254.280 ;
    END
  END instr_addr_o[8]
  PIN instr_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 279.520 900.000 280.120 ;
    END
  END instr_addr_o[9]
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 6.160 900.000 6.760 ;
    END
  END instr_gnt_i
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 57.840 900.000 58.440 ;
    END
  END instr_rdata_i[0]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 318.960 900.000 319.560 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 344.800 900.000 345.400 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 371.320 900.000 371.920 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 397.160 900.000 397.760 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 423.680 900.000 424.280 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 449.520 900.000 450.120 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 475.360 900.000 475.960 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 501.880 900.000 502.480 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 527.720 900.000 528.320 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 553.560 900.000 554.160 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 84.360 900.000 84.960 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 580.080 900.000 580.680 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 605.920 900.000 606.520 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 632.440 900.000 633.040 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 658.280 900.000 658.880 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 684.120 900.000 684.720 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 710.640 900.000 711.240 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 736.480 900.000 737.080 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 762.320 900.000 762.920 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 788.840 900.000 789.440 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 814.680 900.000 815.280 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 110.200 900.000 110.800 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 841.200 900.000 841.800 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 867.040 900.000 867.640 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 136.040 900.000 136.640 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 162.560 900.000 163.160 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 188.400 900.000 189.000 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 214.920 900.000 215.520 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 240.760 900.000 241.360 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 266.600 900.000 267.200 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 293.120 900.000 293.720 ;
    END
  END instr_rdata_i[9]
  PIN instr_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 19.080 900.000 19.680 ;
    END
  END instr_req_o
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 32.000 900.000 32.600 ;
    END
  END instr_rvalid_i
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END rst_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 886.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 886.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 886.805 ;
      LAYER met1 ;
        RECT 3.750 7.860 896.470 886.960 ;
      LAYER met2 ;
        RECT 3.780 4.280 896.440 893.365 ;
        RECT 4.330 3.670 11.310 4.280 ;
        RECT 12.150 3.670 19.130 4.280 ;
        RECT 19.970 3.670 26.950 4.280 ;
        RECT 27.790 3.670 35.230 4.280 ;
        RECT 36.070 3.670 43.050 4.280 ;
        RECT 43.890 3.670 50.870 4.280 ;
        RECT 51.710 3.670 59.150 4.280 ;
        RECT 59.990 3.670 66.970 4.280 ;
        RECT 67.810 3.670 74.790 4.280 ;
        RECT 75.630 3.670 83.070 4.280 ;
        RECT 83.910 3.670 90.890 4.280 ;
        RECT 91.730 3.670 98.710 4.280 ;
        RECT 99.550 3.670 106.990 4.280 ;
        RECT 107.830 3.670 114.810 4.280 ;
        RECT 115.650 3.670 122.630 4.280 ;
        RECT 123.470 3.670 130.910 4.280 ;
        RECT 131.750 3.670 138.730 4.280 ;
        RECT 139.570 3.670 146.550 4.280 ;
        RECT 147.390 3.670 154.830 4.280 ;
        RECT 155.670 3.670 162.650 4.280 ;
        RECT 163.490 3.670 170.470 4.280 ;
        RECT 171.310 3.670 178.750 4.280 ;
        RECT 179.590 3.670 186.570 4.280 ;
        RECT 187.410 3.670 194.390 4.280 ;
        RECT 195.230 3.670 202.210 4.280 ;
        RECT 203.050 3.670 210.490 4.280 ;
        RECT 211.330 3.670 218.310 4.280 ;
        RECT 219.150 3.670 226.130 4.280 ;
        RECT 226.970 3.670 234.410 4.280 ;
        RECT 235.250 3.670 242.230 4.280 ;
        RECT 243.070 3.670 250.050 4.280 ;
        RECT 250.890 3.670 258.330 4.280 ;
        RECT 259.170 3.670 266.150 4.280 ;
        RECT 266.990 3.670 273.970 4.280 ;
        RECT 274.810 3.670 282.250 4.280 ;
        RECT 283.090 3.670 290.070 4.280 ;
        RECT 290.910 3.670 297.890 4.280 ;
        RECT 298.730 3.670 306.170 4.280 ;
        RECT 307.010 3.670 313.990 4.280 ;
        RECT 314.830 3.670 321.810 4.280 ;
        RECT 322.650 3.670 330.090 4.280 ;
        RECT 330.930 3.670 337.910 4.280 ;
        RECT 338.750 3.670 345.730 4.280 ;
        RECT 346.570 3.670 354.010 4.280 ;
        RECT 354.850 3.670 361.830 4.280 ;
        RECT 362.670 3.670 369.650 4.280 ;
        RECT 370.490 3.670 377.470 4.280 ;
        RECT 378.310 3.670 385.750 4.280 ;
        RECT 386.590 3.670 393.570 4.280 ;
        RECT 394.410 3.670 401.390 4.280 ;
        RECT 402.230 3.670 409.670 4.280 ;
        RECT 410.510 3.670 417.490 4.280 ;
        RECT 418.330 3.670 425.310 4.280 ;
        RECT 426.150 3.670 433.590 4.280 ;
        RECT 434.430 3.670 441.410 4.280 ;
        RECT 442.250 3.670 449.230 4.280 ;
        RECT 450.070 3.670 457.510 4.280 ;
        RECT 458.350 3.670 465.330 4.280 ;
        RECT 466.170 3.670 473.150 4.280 ;
        RECT 473.990 3.670 481.430 4.280 ;
        RECT 482.270 3.670 489.250 4.280 ;
        RECT 490.090 3.670 497.070 4.280 ;
        RECT 497.910 3.670 505.350 4.280 ;
        RECT 506.190 3.670 513.170 4.280 ;
        RECT 514.010 3.670 520.990 4.280 ;
        RECT 521.830 3.670 529.270 4.280 ;
        RECT 530.110 3.670 537.090 4.280 ;
        RECT 537.930 3.670 544.910 4.280 ;
        RECT 545.750 3.670 552.730 4.280 ;
        RECT 553.570 3.670 561.010 4.280 ;
        RECT 561.850 3.670 568.830 4.280 ;
        RECT 569.670 3.670 576.650 4.280 ;
        RECT 577.490 3.670 584.930 4.280 ;
        RECT 585.770 3.670 592.750 4.280 ;
        RECT 593.590 3.670 600.570 4.280 ;
        RECT 601.410 3.670 608.850 4.280 ;
        RECT 609.690 3.670 616.670 4.280 ;
        RECT 617.510 3.670 624.490 4.280 ;
        RECT 625.330 3.670 632.770 4.280 ;
        RECT 633.610 3.670 640.590 4.280 ;
        RECT 641.430 3.670 648.410 4.280 ;
        RECT 649.250 3.670 656.690 4.280 ;
        RECT 657.530 3.670 664.510 4.280 ;
        RECT 665.350 3.670 672.330 4.280 ;
        RECT 673.170 3.670 680.610 4.280 ;
        RECT 681.450 3.670 688.430 4.280 ;
        RECT 689.270 3.670 696.250 4.280 ;
        RECT 697.090 3.670 704.530 4.280 ;
        RECT 705.370 3.670 712.350 4.280 ;
        RECT 713.190 3.670 720.170 4.280 ;
        RECT 721.010 3.670 727.990 4.280 ;
        RECT 728.830 3.670 736.270 4.280 ;
        RECT 737.110 3.670 744.090 4.280 ;
        RECT 744.930 3.670 751.910 4.280 ;
        RECT 752.750 3.670 760.190 4.280 ;
        RECT 761.030 3.670 768.010 4.280 ;
        RECT 768.850 3.670 775.830 4.280 ;
        RECT 776.670 3.670 784.110 4.280 ;
        RECT 784.950 3.670 791.930 4.280 ;
        RECT 792.770 3.670 799.750 4.280 ;
        RECT 800.590 3.670 808.030 4.280 ;
        RECT 808.870 3.670 815.850 4.280 ;
        RECT 816.690 3.670 823.670 4.280 ;
        RECT 824.510 3.670 831.950 4.280 ;
        RECT 832.790 3.670 839.770 4.280 ;
        RECT 840.610 3.670 847.590 4.280 ;
        RECT 848.430 3.670 855.870 4.280 ;
        RECT 856.710 3.670 863.690 4.280 ;
        RECT 864.530 3.670 871.510 4.280 ;
        RECT 872.350 3.670 879.790 4.280 ;
        RECT 880.630 3.670 887.610 4.280 ;
        RECT 888.450 3.670 895.430 4.280 ;
        RECT 896.270 3.670 896.440 4.280 ;
      LAYER met3 ;
        RECT 21.040 892.480 895.600 893.345 ;
        RECT 21.040 880.960 896.000 892.480 ;
        RECT 21.040 879.560 895.600 880.960 ;
        RECT 21.040 868.040 896.000 879.560 ;
        RECT 21.040 866.640 895.600 868.040 ;
        RECT 21.040 855.120 896.000 866.640 ;
        RECT 21.040 853.720 895.600 855.120 ;
        RECT 21.040 842.200 896.000 853.720 ;
        RECT 21.040 840.800 895.600 842.200 ;
        RECT 21.040 828.600 896.000 840.800 ;
        RECT 21.040 827.200 895.600 828.600 ;
        RECT 21.040 815.680 896.000 827.200 ;
        RECT 21.040 814.280 895.600 815.680 ;
        RECT 21.040 802.760 896.000 814.280 ;
        RECT 21.040 801.360 895.600 802.760 ;
        RECT 21.040 789.840 896.000 801.360 ;
        RECT 21.040 788.440 895.600 789.840 ;
        RECT 21.040 776.920 896.000 788.440 ;
        RECT 21.040 775.520 895.600 776.920 ;
        RECT 21.040 763.320 896.000 775.520 ;
        RECT 21.040 761.920 895.600 763.320 ;
        RECT 21.040 750.400 896.000 761.920 ;
        RECT 21.040 749.000 895.600 750.400 ;
        RECT 21.040 737.480 896.000 749.000 ;
        RECT 21.040 736.080 895.600 737.480 ;
        RECT 21.040 724.560 896.000 736.080 ;
        RECT 21.040 723.160 895.600 724.560 ;
        RECT 21.040 711.640 896.000 723.160 ;
        RECT 21.040 710.240 895.600 711.640 ;
        RECT 21.040 698.040 896.000 710.240 ;
        RECT 21.040 696.640 895.600 698.040 ;
        RECT 21.040 685.120 896.000 696.640 ;
        RECT 21.040 683.720 895.600 685.120 ;
        RECT 21.040 672.200 896.000 683.720 ;
        RECT 21.040 670.800 895.600 672.200 ;
        RECT 21.040 659.280 896.000 670.800 ;
        RECT 21.040 657.880 895.600 659.280 ;
        RECT 21.040 646.360 896.000 657.880 ;
        RECT 21.040 644.960 895.600 646.360 ;
        RECT 21.040 633.440 896.000 644.960 ;
        RECT 21.040 632.040 895.600 633.440 ;
        RECT 21.040 619.840 896.000 632.040 ;
        RECT 21.040 618.440 895.600 619.840 ;
        RECT 21.040 606.920 896.000 618.440 ;
        RECT 21.040 605.520 895.600 606.920 ;
        RECT 21.040 594.000 896.000 605.520 ;
        RECT 21.040 592.600 895.600 594.000 ;
        RECT 21.040 581.080 896.000 592.600 ;
        RECT 21.040 579.680 895.600 581.080 ;
        RECT 21.040 568.160 896.000 579.680 ;
        RECT 21.040 566.760 895.600 568.160 ;
        RECT 21.040 554.560 896.000 566.760 ;
        RECT 21.040 553.160 895.600 554.560 ;
        RECT 21.040 541.640 896.000 553.160 ;
        RECT 21.040 540.240 895.600 541.640 ;
        RECT 21.040 528.720 896.000 540.240 ;
        RECT 21.040 527.320 895.600 528.720 ;
        RECT 21.040 515.800 896.000 527.320 ;
        RECT 21.040 514.400 895.600 515.800 ;
        RECT 21.040 502.880 896.000 514.400 ;
        RECT 21.040 501.480 895.600 502.880 ;
        RECT 21.040 489.280 896.000 501.480 ;
        RECT 21.040 487.880 895.600 489.280 ;
        RECT 21.040 476.360 896.000 487.880 ;
        RECT 21.040 474.960 895.600 476.360 ;
        RECT 21.040 463.440 896.000 474.960 ;
        RECT 21.040 462.040 895.600 463.440 ;
        RECT 21.040 450.520 896.000 462.040 ;
        RECT 21.040 449.120 895.600 450.520 ;
        RECT 21.040 437.600 896.000 449.120 ;
        RECT 21.040 436.200 895.600 437.600 ;
        RECT 21.040 424.680 896.000 436.200 ;
        RECT 21.040 423.280 895.600 424.680 ;
        RECT 21.040 411.080 896.000 423.280 ;
        RECT 21.040 409.680 895.600 411.080 ;
        RECT 21.040 398.160 896.000 409.680 ;
        RECT 21.040 396.760 895.600 398.160 ;
        RECT 21.040 385.240 896.000 396.760 ;
        RECT 21.040 383.840 895.600 385.240 ;
        RECT 21.040 372.320 896.000 383.840 ;
        RECT 21.040 370.920 895.600 372.320 ;
        RECT 21.040 359.400 896.000 370.920 ;
        RECT 21.040 358.000 895.600 359.400 ;
        RECT 21.040 345.800 896.000 358.000 ;
        RECT 21.040 344.400 895.600 345.800 ;
        RECT 21.040 332.880 896.000 344.400 ;
        RECT 21.040 331.480 895.600 332.880 ;
        RECT 21.040 319.960 896.000 331.480 ;
        RECT 21.040 318.560 895.600 319.960 ;
        RECT 21.040 307.040 896.000 318.560 ;
        RECT 21.040 305.640 895.600 307.040 ;
        RECT 21.040 294.120 896.000 305.640 ;
        RECT 21.040 292.720 895.600 294.120 ;
        RECT 21.040 280.520 896.000 292.720 ;
        RECT 21.040 279.120 895.600 280.520 ;
        RECT 21.040 267.600 896.000 279.120 ;
        RECT 21.040 266.200 895.600 267.600 ;
        RECT 21.040 254.680 896.000 266.200 ;
        RECT 21.040 253.280 895.600 254.680 ;
        RECT 21.040 241.760 896.000 253.280 ;
        RECT 21.040 240.360 895.600 241.760 ;
        RECT 21.040 228.840 896.000 240.360 ;
        RECT 21.040 227.440 895.600 228.840 ;
        RECT 21.040 215.920 896.000 227.440 ;
        RECT 21.040 214.520 895.600 215.920 ;
        RECT 21.040 202.320 896.000 214.520 ;
        RECT 21.040 200.920 895.600 202.320 ;
        RECT 21.040 189.400 896.000 200.920 ;
        RECT 21.040 188.000 895.600 189.400 ;
        RECT 21.040 176.480 896.000 188.000 ;
        RECT 21.040 175.080 895.600 176.480 ;
        RECT 21.040 163.560 896.000 175.080 ;
        RECT 21.040 162.160 895.600 163.560 ;
        RECT 21.040 150.640 896.000 162.160 ;
        RECT 21.040 149.240 895.600 150.640 ;
        RECT 21.040 137.040 896.000 149.240 ;
        RECT 21.040 135.640 895.600 137.040 ;
        RECT 21.040 124.120 896.000 135.640 ;
        RECT 21.040 122.720 895.600 124.120 ;
        RECT 21.040 111.200 896.000 122.720 ;
        RECT 21.040 109.800 895.600 111.200 ;
        RECT 21.040 98.280 896.000 109.800 ;
        RECT 21.040 96.880 895.600 98.280 ;
        RECT 21.040 85.360 896.000 96.880 ;
        RECT 21.040 83.960 895.600 85.360 ;
        RECT 21.040 71.760 896.000 83.960 ;
        RECT 21.040 70.360 895.600 71.760 ;
        RECT 21.040 58.840 896.000 70.360 ;
        RECT 21.040 57.440 895.600 58.840 ;
        RECT 21.040 45.920 896.000 57.440 ;
        RECT 21.040 44.520 895.600 45.920 ;
        RECT 21.040 33.000 896.000 44.520 ;
        RECT 21.040 31.600 895.600 33.000 ;
        RECT 21.040 20.080 896.000 31.600 ;
        RECT 21.040 18.680 895.600 20.080 ;
        RECT 21.040 7.160 896.000 18.680 ;
        RECT 21.040 6.295 895.600 7.160 ;
      LAYER met4 ;
        RECT 160.375 12.415 174.240 885.865 ;
        RECT 176.640 12.415 251.040 885.865 ;
        RECT 253.440 12.415 327.840 885.865 ;
        RECT 330.240 12.415 404.640 885.865 ;
        RECT 407.040 12.415 481.440 885.865 ;
        RECT 483.840 12.415 558.240 885.865 ;
        RECT 560.640 12.415 635.040 885.865 ;
        RECT 637.440 12.415 711.840 885.865 ;
        RECT 714.240 12.415 788.640 885.865 ;
        RECT 791.040 12.415 796.425 885.865 ;
  END
END crypto_core
END LIBRARY

