* NGSPICE file created from uart_to_mem.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

.subckt uart_to_mem clk_i data_addr_o[0] data_addr_o[10] data_addr_o[11] data_addr_o[1]
+ data_addr_o[2] data_addr_o[3] data_addr_o[4] data_addr_o[5] data_addr_o[6] data_addr_o[7]
+ data_addr_o[8] data_addr_o[9] data_be_o[0] data_be_o[1] data_be_o[2] data_be_o[3]
+ data_gnt_i data_rdata_i[0] data_rdata_i[10] data_rdata_i[11] data_rdata_i[12] data_rdata_i[13]
+ data_rdata_i[14] data_rdata_i[15] data_rdata_i[16] data_rdata_i[17] data_rdata_i[18]
+ data_rdata_i[19] data_rdata_i[1] data_rdata_i[20] data_rdata_i[21] data_rdata_i[22]
+ data_rdata_i[23] data_rdata_i[24] data_rdata_i[25] data_rdata_i[26] data_rdata_i[27]
+ data_rdata_i[28] data_rdata_i[29] data_rdata_i[2] data_rdata_i[30] data_rdata_i[31]
+ data_rdata_i[3] data_rdata_i[4] data_rdata_i[5] data_rdata_i[6] data_rdata_i[7]
+ data_rdata_i[8] data_rdata_i[9] data_req_o data_rvalid_i data_wdata_o[0] data_wdata_o[10]
+ data_wdata_o[11] data_wdata_o[12] data_wdata_o[13] data_wdata_o[14] data_wdata_o[15]
+ data_wdata_o[16] data_wdata_o[17] data_wdata_o[18] data_wdata_o[19] data_wdata_o[1]
+ data_wdata_o[20] data_wdata_o[21] data_wdata_o[22] data_wdata_o[23] data_wdata_o[24]
+ data_wdata_o[25] data_wdata_o[26] data_wdata_o[27] data_wdata_o[28] data_wdata_o[29]
+ data_wdata_o[2] data_wdata_o[30] data_wdata_o[31] data_wdata_o[3] data_wdata_o[4]
+ data_wdata_o[5] data_wdata_o[6] data_wdata_o[7] data_wdata_o[8] data_wdata_o[9]
+ data_we_o rst_i rx_i tx_o uart_error vccd1 vssd1
XANTENNA__1151__B1 data_rdata_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1206__A1 data_req_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1142__B1 data_rdata_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1270_ _1456_/A _1270_/B vssd1 vssd1 vccd1 vccd1 _1897_/D sky130_fd_sc_hd__nor2_2
XFILLER_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0985_ _0985_/A vssd1 vssd1 vccd1 vccd1 _0985_/X sky130_fd_sc_hd__buf_1
X_1606_ _1825_/Q _1606_/B vssd1 vssd1 vccd1 vccd1 _1617_/C sky130_fd_sc_hd__or2_2
X_1399_ _1399_/A vssd1 vssd1 vccd1 vccd1 _1400_/A sky130_fd_sc_hd__buf_1
X_1468_ _1476_/A vssd1 vssd1 vccd1 vccd1 _1468_/X sky130_fd_sc_hd__buf_1
X_1537_ _0987_/B _1486_/X _1500_/Y _1488_/X vssd1 vssd1 vccd1 vccd1 _1863_/D sky130_fd_sc_hd__o22ai_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1322_ _1893_/Q vssd1 vssd1 vccd1 vccd1 _1644_/B sky130_fd_sc_hd__inv_2
X_1253_ _1263_/B _1465_/B _1253_/C vssd1 vssd1 vccd1 vccd1 _1253_/X sky130_fd_sc_hd__or3_2
X_1184_ _1184_/A vssd1 vssd1 vccd1 vccd1 _1184_/X sky130_fd_sc_hd__buf_1
X_0968_ data_wdata_o[12] _0953_/X _0926_/X _0955_/X vssd1 vssd1 vccd1 vccd1 _1963_/D
+ sky130_fd_sc_hd__a22o_2
X_0899_ _1864_/Q vssd1 vssd1 vccd1 vccd1 _0906_/B sky130_fd_sc_hd__inv_2
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1871_ _1876_/CLK _1871_/D _1430_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[0] sky130_fd_sc_hd__dfrtp_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1940_ _1940_/CLK _1940_/D vssd1 vssd1 vccd1 vccd1 _1940_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1305_ _1812_/Q _1758_/S _1812_/Q _1758_/S vssd1 vssd1 vccd1 vccd1 _1306_/A sky130_fd_sc_hd__a2bb2o_2
X_1236_ _1243_/A _1740_/S _1246_/A _1235_/Y vssd1 vssd1 vccd1 vccd1 _1466_/B sky130_fd_sc_hd__o2bb2a_2
X_1167_ _1924_/Q _1163_/X data_rdata_i[17] _1164_/X _1161_/X vssd1 vssd1 vccd1 vccd1
+ _1924_/D sky130_fd_sc_hd__o221a_2
X_1098_ _1945_/Q _1096_/X _1096_/X _1097_/Y vssd1 vssd1 vccd1 vccd1 _1945_/D sky130_fd_sc_hd__o2bb2ai_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1021_ _1066_/A vssd1 vssd1 vccd1 vccd1 _1432_/B sky130_fd_sc_hd__inv_2
X_1923_ _1930_/CLK _1923_/D vssd1 vssd1 vccd1 vccd1 _1923_/Q sky130_fd_sc_hd__dfxtp_2
X_1854_ _1943_/CLK _1854_/D vssd1 vssd1 vccd1 vccd1 _1854_/Q sky130_fd_sc_hd__dfxtp_2
X_1785_ _1620_/B _1621_/X _1791_/S vssd1 vssd1 vccd1 vccd1 _1827_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1219_ _1804_/Q vssd1 vssd1 vccd1 vccd1 _1219_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1570_ _1838_/Q _1570_/B vssd1 vssd1 vccd1 vccd1 _1570_/Y sky130_fd_sc_hd__nor2_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1004_ _1004_/A vssd1 vssd1 vccd1 vccd1 _1004_/X sky130_fd_sc_hd__buf_1
X_1768_ _1911_/Q _1919_/Q _1862_/Q vssd1 vssd1 vccd1 vccd1 _1768_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0992__A1 data_wdata_o[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1906_ _1940_/CLK _1906_/D vssd1 vssd1 vccd1 vccd1 data_we_o sky130_fd_sc_hd__dfxtp_2
X_1837_ _1842_/CLK _1837_/D vssd1 vssd1 vccd1 vccd1 _1837_/Q sky130_fd_sc_hd__dfxtp_2
X_1699_ vssd1 vssd1 vccd1 vccd1 data_be_o[3] _1699_/LO sky130_fd_sc_hd__conb_1
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0983__A1 data_wdata_o[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1622_ _1828_/Q _1617_/X _1626_/B vssd1 vssd1 vccd1 vccd1 _1623_/A sky130_fd_sc_hd__a21bo_2
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1553_ _1553_/A vssd1 vssd1 vccd1 vccd1 _1553_/X sky130_fd_sc_hd__buf_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1484_ _1867_/Q _1333_/X _1483_/X _1349_/X vssd1 vssd1 vccd1 vccd1 _1867_/D sky130_fd_sc_hd__a31o_2
Xclkbuf_4_12_0_clk_i clkbuf_3_6_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1876_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__0965__A1 data_wdata_o[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0984_ _0984_/A vssd1 vssd1 vccd1 vccd1 _0985_/A sky130_fd_sc_hd__buf_1
X_1536_ _0906_/B _1488_/X _1364_/A _1535_/X vssd1 vssd1 vccd1 vccd1 _1864_/D sky130_fd_sc_hd__o22ai_2
X_1605_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1605_/X sky130_fd_sc_hd__buf_1
X_1398_ data_wdata_o[24] _1382_/X _1397_/X _1384_/X vssd1 vssd1 vccd1 vccd1 _1879_/D
+ sky130_fd_sc_hd__a22o_2
X_1467_ _1244_/A _1465_/X _1466_/B tx_o _1466_/Y vssd1 vssd1 vccd1 vccd1 _1851_/D
+ sky130_fd_sc_hd__a32o_2
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0938__A1 data_wdata_o[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1321_ _1894_/Q vssd1 vssd1 vccd1 vccd1 _1321_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1354__A1 data_addr_o[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1252_ _1901_/Q _1256_/A _1902_/Q vssd1 vssd1 vccd1 vccd1 _1253_/C sky130_fd_sc_hd__o21a_2
X_1183_ _1916_/Q _1179_/X data_rdata_i[9] _1180_/X _1177_/X vssd1 vssd1 vccd1 vccd1
+ _1916_/D sky130_fd_sc_hd__o221a_2
XFILLER_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0967_ _0967_/A vssd1 vssd1 vccd1 vccd1 _0967_/X sky130_fd_sc_hd__buf_1
X_1519_ _1519_/A vssd1 vssd1 vccd1 vccd1 _1791_/S sky130_fd_sc_hd__buf_1
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1870_ _1903_/CLK _1870_/D vssd1 vssd1 vccd1 vccd1 _1870_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1166_ _1925_/Q _1163_/X data_rdata_i[18] _1164_/X _1161_/X vssd1 vssd1 vccd1 vccd1
+ _1925_/D sky130_fd_sc_hd__o221a_2
X_1304_ _1304_/A _1304_/B vssd1 vssd1 vccd1 vccd1 _1758_/S sky130_fd_sc_hd__nor2_2
X_1235_ _1679_/A vssd1 vssd1 vccd1 vccd1 _1235_/Y sky130_fd_sc_hd__inv_2
X_1097_ _1075_/X _1773_/X _1846_/Q _1077_/X vssd1 vssd1 vccd1 vccd1 _1097_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1020_ _1811_/Q _1810_/Q vssd1 vssd1 vccd1 vccd1 _1066_/A sky130_fd_sc_hd__or2_2
X_1922_ _1930_/CLK _1922_/D vssd1 vssd1 vccd1 vccd1 _1922_/Q sky130_fd_sc_hd__dfxtp_2
X_1784_ _1624_/B _1625_/X _1791_/S vssd1 vssd1 vccd1 vccd1 _1828_/D sky130_fd_sc_hd__mux2_1
X_1853_ _1943_/CLK _1853_/D vssd1 vssd1 vccd1 vccd1 _1853_/Q sky130_fd_sc_hd__dfxtp_2
X_1149_ _1164_/A vssd1 vssd1 vccd1 vccd1 _1149_/X sky130_fd_sc_hd__buf_1
X_1218_ _1718_/X _1714_/X _1713_/X vssd1 vssd1 vccd1 vccd1 _1232_/C sky130_fd_sc_hd__or3_2
XFILLER_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1003_ _1003_/A vssd1 vssd1 vccd1 vccd1 _1004_/A sky130_fd_sc_hd__buf_1
X_1905_ _1940_/CLK _1905_/D vssd1 vssd1 vccd1 vccd1 data_req_o sky130_fd_sc_hd__dfxtp_2
XFILLER_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1698_ vssd1 vssd1 vccd1 vccd1 data_be_o[2] _1698_/LO sky130_fd_sc_hd__conb_1
X_1767_ _1766_/X _1932_/Q _1860_/Q vssd1 vssd1 vccd1 vccd1 _1767_/X sky130_fd_sc_hd__mux2_1
X_1836_ _1842_/CLK _1836_/D vssd1 vssd1 vccd1 vccd1 _1836_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1621_ _1621_/A vssd1 vssd1 vccd1 vccd1 _1621_/X sky130_fd_sc_hd__buf_1
X_1552_ _1557_/A _1552_/B vssd1 vssd1 vccd1 vccd1 _1553_/A sky130_fd_sc_hd__and2_2
XFILLER_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1483_ _1483_/A _1483_/B _1483_/C vssd1 vssd1 vccd1 vccd1 _1483_/X sky130_fd_sc_hd__or3_2
X_1819_ _1950_/CLK _1819_/D vssd1 vssd1 vccd1 vccd1 _1819_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0983_ data_wdata_o[8] _0971_/X _0946_/X _0972_/X vssd1 vssd1 vccd1 vccd1 _1959_/D
+ sky130_fd_sc_hd__a22o_2
X_1535_ _1535_/A _1535_/B vssd1 vssd1 vccd1 vccd1 _1535_/X sky130_fd_sc_hd__and2_2
X_1604_ _1609_/A _1604_/B vssd1 vssd1 vccd1 vccd1 _1605_/A sky130_fd_sc_hd__and2_2
X_1397_ _1843_/Q vssd1 vssd1 vccd1 vccd1 _1397_/X sky130_fd_sc_hd__buf_1
X_1466_ _1679_/B _1466_/B vssd1 vssd1 vccd1 vccd1 _1466_/Y sky130_fd_sc_hd__nand2_2
XFILLER_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1320_ _1313_/A _1313_/C _1476_/A _1319_/X vssd1 vssd1 vccd1 vccd1 _1895_/D sky130_fd_sc_hd__o22ai_2
X_1182_ _1917_/Q _1179_/X data_rdata_i[10] _1180_/X _1177_/X vssd1 vssd1 vccd1 vccd1
+ _1917_/D sky130_fd_sc_hd__o221a_2
X_1251_ _1251_/A vssd1 vssd1 vccd1 vccd1 _1465_/B sky130_fd_sc_hd__inv_2
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0966_ _0969_/A vssd1 vssd1 vccd1 vccd1 _0967_/A sky130_fd_sc_hd__buf_1
X_1449_ _1449_/A vssd1 vssd1 vccd1 vccd1 _1449_/X sky130_fd_sc_hd__buf_1
XFILLER_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1518_ _1514_/Y _1512_/Y _1817_/Q _1517_/Y _1515_/X vssd1 vssd1 vccd1 vccd1 _1518_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1303_ _1840_/Q _1841_/Q _1575_/B _1303_/D vssd1 vssd1 vccd1 vccd1 _1304_/B sky130_fd_sc_hd__or4_2
X_1165_ _1926_/Q _1163_/X data_rdata_i[19] _1164_/X _1161_/X vssd1 vssd1 vccd1 vccd1
+ _1926_/D sky130_fd_sc_hd__o221a_2
XFILLER_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1096_ _1096_/A vssd1 vssd1 vccd1 vccd1 _1096_/X sky130_fd_sc_hd__buf_1
X_1234_ _1903_/Q vssd1 vssd1 vccd1 vccd1 _1246_/A sky130_fd_sc_hd__buf_1
X_0949_ _0949_/A vssd1 vssd1 vccd1 vccd1 _0949_/X sky130_fd_sc_hd__buf_1
XFILLER_18_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1190__B1 data_rdata_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1921_ _1945_/CLK _1921_/D vssd1 vssd1 vccd1 vccd1 _1921_/Q sky130_fd_sc_hd__dfxtp_2
X_1852_ _1903_/CLK _1852_/D vssd1 vssd1 vccd1 vccd1 _1852_/Q sky130_fd_sc_hd__dfxtp_2
X_1783_ _1628_/Y _1629_/Y _1791_/S vssd1 vssd1 vccd1 vccd1 _1829_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1181__B1 data_rdata_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1148_ _1163_/A vssd1 vssd1 vccd1 vccd1 _1148_/X sky130_fd_sc_hd__buf_1
X_1079_ _1949_/Q _1073_/X _1073_/X _1078_/Y vssd1 vssd1 vccd1 vccd1 _1949_/D sky130_fd_sc_hd__o2bb2ai_2
XFILLER_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1217_ _1217_/A vssd1 vssd1 vccd1 vccd1 _1243_/A sky130_fd_sc_hd__inv_2
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1002_ data_wdata_o[4] _0989_/X _0926_/X _0991_/X vssd1 vssd1 vccd1 vccd1 _1955_/D
+ sky130_fd_sc_hd__a22o_2
X_1904_ _1943_/CLK _1904_/D vssd1 vssd1 vccd1 vccd1 _1904_/Q sky130_fd_sc_hd__dfxtp_2
X_1835_ _1842_/CLK _1835_/D vssd1 vssd1 vccd1 vccd1 _1835_/Q sky130_fd_sc_hd__dfxtp_2
X_1697_ vssd1 vssd1 vccd1 vccd1 data_be_o[1] _1697_/LO sky130_fd_sc_hd__conb_1
X_1766_ _1765_/X _1924_/Q _1864_/Q vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1154__B1 data_rdata_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1620_ _1632_/A _1620_/B vssd1 vssd1 vccd1 vccd1 _1621_/A sky130_fd_sc_hd__and2_2
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1551_ _1551_/A vssd1 vssd1 vccd1 vccd1 _1552_/B sky130_fd_sc_hd__buf_1
X_1482_ _1482_/A vssd1 vssd1 vccd1 vccd1 _1483_/B sky130_fd_sc_hd__buf_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1818_ _1950_/CLK _1818_/D vssd1 vssd1 vccd1 vccd1 _1818_/Q sky130_fd_sc_hd__dfxtp_2
X_1749_ _1663_/X _1664_/C _1749_/S vssd1 vssd1 vccd1 vccd1 _1749_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_4_6_0_clk_i clkbuf_4_7_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1945_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1469__A rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0982_ _0982_/A vssd1 vssd1 vccd1 vccd1 _0982_/X sky130_fd_sc_hd__buf_1
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1603_ _1603_/A vssd1 vssd1 vccd1 vccd1 _1604_/B sky130_fd_sc_hd__buf_1
X_1534_ _1022_/X _1036_/Y _1868_/Q _1533_/X vssd1 vssd1 vccd1 vccd1 _1868_/D sky130_fd_sc_hd__a22o_2
X_1465_ _1852_/Q _1465_/B vssd1 vssd1 vccd1 vccd1 _1465_/X sky130_fd_sc_hd__or2_2
X_1396_ _1396_/A vssd1 vssd1 vccd1 vccd1 _1396_/X sky130_fd_sc_hd__buf_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1181_ _1918_/Q _1179_/X data_rdata_i[11] _1180_/X _1177_/X vssd1 vssd1 vccd1 vccd1
+ _1918_/D sky130_fd_sc_hd__o221a_2
X_1250_ _1250_/A vssd1 vssd1 vccd1 vccd1 _1250_/X sky130_fd_sc_hd__buf_1
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0965_ data_wdata_o[13] _0953_/X _0922_/X _0955_/X vssd1 vssd1 vccd1 vccd1 _1964_/D
+ sky130_fd_sc_hd__a22o_2
X_1448_ _1452_/A vssd1 vssd1 vccd1 vccd1 _1449_/A sky130_fd_sc_hd__buf_1
X_1517_ _1817_/Q vssd1 vssd1 vccd1 vccd1 _1517_/Y sky130_fd_sc_hd__inv_2
X_1379_ data_wdata_o[28] _1365_/X _0926_/X _1367_/X vssd1 vssd1 vccd1 vccd1 _1883_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1302_ _1834_/Q _1835_/Q _1302_/C _1833_/Q vssd1 vssd1 vccd1 vccd1 _1303_/D sky130_fd_sc_hd__or4_2
X_1233_ _1233_/A vssd1 vssd1 vccd1 vccd1 _1740_/S sky130_fd_sc_hd__buf_1
X_1164_ _1164_/A vssd1 vssd1 vccd1 vccd1 _1164_/X sky130_fd_sc_hd__buf_1
X_1095_ _1095_/A vssd1 vssd1 vccd1 vccd1 _1095_/X sky130_fd_sc_hd__buf_1
X_0948_ _0948_/A vssd1 vssd1 vccd1 vccd1 _0949_/A sky130_fd_sc_hd__buf_1
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1920_ _1945_/CLK _1920_/D vssd1 vssd1 vccd1 vccd1 _1920_/Q sky130_fd_sc_hd__dfxtp_2
X_1851_ _1903_/CLK _1851_/D vssd1 vssd1 vccd1 vccd1 tx_o sky130_fd_sc_hd__dfxtp_2
X_1782_ _1632_/B _1633_/X _1791_/S vssd1 vssd1 vccd1 vccd1 _1830_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1216_ _1216_/A vssd1 vssd1 vccd1 vccd1 _1251_/A sky130_fd_sc_hd__buf_1
X_1147_ _1935_/Q _1139_/X data_rdata_i[28] _1141_/X _1146_/X vssd1 vssd1 vccd1 vccd1
+ _1935_/D sky130_fd_sc_hd__o221a_2
X_1078_ _1075_/X _1752_/X _1076_/X _1077_/X vssd1 vssd1 vccd1 vccd1 _1078_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _1001_/A vssd1 vssd1 vccd1 vccd1 _1001_/X sky130_fd_sc_hd__buf_1
X_1765_ _1908_/Q _1916_/Q _1862_/Q vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0977__A1 data_wdata_o[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1834_ _1842_/CLK _1834_/D vssd1 vssd1 vccd1 vccd1 _1834_/Q sky130_fd_sc_hd__dfxtp_2
X_1903_ _1903_/CLK _1903_/D vssd1 vssd1 vccd1 vccd1 _1903_/Q sky130_fd_sc_hd__dfxtp_2
X_1696_ vssd1 vssd1 vccd1 vccd1 data_be_o[0] _1696_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_clk_i clkbuf_4_3_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1940_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0924__A _0928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1481_ _1397_/X _1476_/X _1393_/X _1477_/X vssd1 vssd1 vccd1 vccd1 _1843_/D sky130_fd_sc_hd__a22o_2
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1550_ _1834_/Q _1296_/B _1297_/B vssd1 vssd1 vccd1 vccd1 _1551_/A sky130_fd_sc_hd__a21bo_2
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1748_ _1655_/B _1656_/X _1761_/S vssd1 vssd1 vccd1 vccd1 _1748_/X sky130_fd_sc_hd__mux2_1
X_1817_ _1950_/CLK _1817_/D vssd1 vssd1 vccd1 vccd1 _1817_/Q sky130_fd_sc_hd__dfxtp_2
X_1679_ _1679_/A _1679_/B vssd1 vssd1 vccd1 vccd1 _1732_/S sky130_fd_sc_hd__nor2_2
XFILLER_42_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0981_ _0984_/A vssd1 vssd1 vccd1 vccd1 _0982_/A sky130_fd_sc_hd__buf_1
X_1602_ _1824_/Q _1596_/X _1606_/B vssd1 vssd1 vccd1 vccd1 _1603_/A sky130_fd_sc_hd__a21bo_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1395_ _1399_/A vssd1 vssd1 vccd1 vccd1 _1396_/A sky130_fd_sc_hd__buf_1
X_1533_ _1533_/A _1533_/B vssd1 vssd1 vccd1 vccd1 _1533_/X sky130_fd_sc_hd__or2_2
X_1464_ _1852_/Q _1240_/A _1780_/X _1258_/X vssd1 vssd1 vccd1 vccd1 _1852_/D sky130_fd_sc_hd__a22o_2
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1180_ _1194_/A vssd1 vssd1 vccd1 vccd1 _1180_/X sky130_fd_sc_hd__buf_1
XFILLER_17_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0964_ _0964_/A vssd1 vssd1 vccd1 vccd1 _0964_/X sky130_fd_sc_hd__buf_1
X_1516_ _1514_/Y _1512_/Y _1515_/X vssd1 vssd1 vccd1 vccd1 _1516_/X sky130_fd_sc_hd__o21a_2
X_1447_ _1447_/A vssd1 vssd1 vccd1 vccd1 _1447_/X sky130_fd_sc_hd__buf_1
X_1378_ _1378_/A vssd1 vssd1 vccd1 vccd1 _1378_/X sky130_fd_sc_hd__buf_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1301_ _1832_/Q vssd1 vssd1 vccd1 vccd1 _1302_/C sky130_fd_sc_hd__inv_2
X_1232_ _1711_/X _1717_/X _1232_/C _1683_/B vssd1 vssd1 vccd1 vccd1 _1233_/A sky130_fd_sc_hd__or4_2
X_1163_ _1163_/A vssd1 vssd1 vccd1 vccd1 _1163_/X sky130_fd_sc_hd__buf_1
X_1094_ _1107_/A vssd1 vssd1 vccd1 vccd1 _1095_/A sky130_fd_sc_hd__buf_1
X_0947_ data_wdata_o[16] _0930_/X _0946_/X _0932_/X vssd1 vssd1 vccd1 vccd1 _1967_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1850_ _1938_/CLK _1850_/D vssd1 vssd1 vccd1 vccd1 _1850_/Q sky130_fd_sc_hd__dfxtp_2
X_1781_ _1230_/A _1634_/Y _1791_/S vssd1 vssd1 vccd1 vccd1 _1831_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1146_ _1694_/A vssd1 vssd1 vccd1 vccd1 _1146_/X sky130_fd_sc_hd__buf_1
X_1215_ _1901_/Q _1256_/A _1902_/Q vssd1 vssd1 vccd1 vccd1 _1216_/A sky130_fd_sc_hd__or3_2
X_1077_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1077_/X sky130_fd_sc_hd__buf_1
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1000_ _1003_/A vssd1 vssd1 vccd1 vccd1 _1001_/A sky130_fd_sc_hd__buf_1
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1902_ _1943_/CLK _1902_/D vssd1 vssd1 vccd1 vccd1 _1902_/Q sky130_fd_sc_hd__dfxtp_2
X_1764_ _1763_/X _1937_/Q _1860_/Q vssd1 vssd1 vccd1 vccd1 _1764_/X sky130_fd_sc_hd__mux2_1
X_1833_ _1842_/CLK _1833_/D vssd1 vssd1 vccd1 vccd1 _1833_/Q sky130_fd_sc_hd__dfxtp_2
X_1695_ _1695_/A vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_3_0_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1129_ _1115_/Y _1803_/S _1117_/A vssd1 vssd1 vccd1 vccd1 _1129_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1480_ _1393_/A _1476_/X _1389_/X _1477_/X vssd1 vssd1 vccd1 vccd1 _1844_/D sky130_fd_sc_hd__a22o_2
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1678_ _1716_/X _1650_/X _1754_/X _1658_/X vssd1 vssd1 vccd1 vccd1 _1678_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_7_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1816_ _1950_/CLK _1816_/D vssd1 vssd1 vccd1 vccd1 _1816_/Q sky130_fd_sc_hd__dfxtp_2
X_1747_ _1664_/B _1642_/A _1747_/S vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0980_ data_wdata_o[9] _0971_/X _0942_/X _0972_/X vssd1 vssd1 vccd1 vccd1 _1960_/D
+ sky130_fd_sc_hd__a22o_2
X_1532_ _1532_/A _1532_/B vssd1 vssd1 vccd1 vccd1 _1532_/Y sky130_fd_sc_hd__nor2_2
X_1601_ _1601_/A vssd1 vssd1 vccd1 vccd1 _1601_/X sky130_fd_sc_hd__buf_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1394_ data_wdata_o[25] _1382_/X _1393_/X _1384_/X vssd1 vssd1 vccd1 vccd1 _1880_/D
+ sky130_fd_sc_hd__a22o_2
X_1463_ _1779_/X _1250_/X _1853_/Q _1258_/X vssd1 vssd1 vccd1 vccd1 _1853_/D sky130_fd_sc_hd__o22a_2
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0963_ _0969_/A vssd1 vssd1 vccd1 vccd1 _0964_/A sky130_fd_sc_hd__buf_1
X_1515_ _1816_/Q _1515_/B vssd1 vssd1 vccd1 vccd1 _1515_/X sky130_fd_sc_hd__or2_2
X_1377_ _1380_/A vssd1 vssd1 vccd1 vccd1 _1378_/A sky130_fd_sc_hd__buf_1
X_1446_ _1452_/A vssd1 vssd1 vccd1 vccd1 _1447_/A sky130_fd_sc_hd__buf_1
XFILLER_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1162_ _1927_/Q _1155_/X data_rdata_i[20] _1156_/X _1161_/X vssd1 vssd1 vccd1 vccd1
+ _1927_/D sky130_fd_sc_hd__o221a_2
X_1300_ _1587_/B vssd1 vssd1 vccd1 vccd1 _1304_/A sky130_fd_sc_hd__inv_2
X_1231_ _1219_/Y _1718_/S _1219_/Y _1718_/S vssd1 vssd1 vccd1 vccd1 _1683_/B sky130_fd_sc_hd__a2bb2o_2
X_1093_ _1351_/A vssd1 vssd1 vccd1 vccd1 _1107_/A sky130_fd_sc_hd__buf_1
X_0946_ _1843_/Q vssd1 vssd1 vccd1 vccd1 _0946_/X sky130_fd_sc_hd__buf_1
X_1429_ _1434_/A vssd1 vssd1 vccd1 vccd1 _1430_/A sky130_fd_sc_hd__buf_1
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1175__B1 data_rdata_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1780_ _1942_/Q _1853_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _1780_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1166__B1 data_rdata_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1145_ _1445_/A vssd1 vssd1 vccd1 vccd1 _1694_/A sky130_fd_sc_hd__buf_1
X_1214_ _1900_/Q _1899_/Q vssd1 vssd1 vccd1 vccd1 _1256_/A sky130_fd_sc_hd__or2_2
X_1076_ _1850_/Q vssd1 vssd1 vccd1 vccd1 _1076_/X sky130_fd_sc_hd__buf_1
XANTENNA__1157__B1 data_rdata_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0929_ _0929_/A vssd1 vssd1 vccd1 vccd1 _0929_/X sky130_fd_sc_hd__buf_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1832_ _1842_/CLK _1832_/D vssd1 vssd1 vccd1 vccd1 _1832_/Q sky130_fd_sc_hd__dfxtp_2
X_1901_ _1903_/CLK _1901_/D vssd1 vssd1 vccd1 vccd1 _1901_/Q sky130_fd_sc_hd__dfxtp_2
X_1694_ _1694_/A vssd1 vssd1 vccd1 vccd1 _1695_/A sky130_fd_sc_hd__buf_1
X_1763_ _1762_/X _1929_/Q _1864_/Q vssd1 vssd1 vccd1 vccd1 _1763_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_4_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1128_ _1128_/A vssd1 vssd1 vccd1 vccd1 _1803_/S sky130_fd_sc_hd__buf_1
X_1059_ _1485_/A _1492_/C _1492_/B vssd1 vssd1 vccd1 vccd1 _1059_/X sky130_fd_sc_hd__or3_2
XFILLER_16_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1815_ _1940_/CLK _1815_/D vssd1 vssd1 vccd1 vccd1 _1815_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1746_ _1745_/X _1933_/Q _1860_/Q vssd1 vssd1 vccd1 vccd1 _1746_/X sky130_fd_sc_hd__mux2_1
X_1677_ _1677_/A vssd1 vssd1 vccd1 vccd1 _1677_/X sky130_fd_sc_hd__buf_1
XFILLER_26_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1112__A data_rvalid_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1462_ _1778_/X _1250_/X _1854_/Q _1458_/X vssd1 vssd1 vccd1 vccd1 _1854_/D sky130_fd_sc_hd__o22a_2
X_1600_ _1609_/A _1600_/B vssd1 vssd1 vccd1 vccd1 _1601_/A sky130_fd_sc_hd__and2_2
X_1531_ _1333_/A _1419_/A _0904_/A _0988_/B vssd1 vssd1 vccd1 vccd1 _1869_/D sky130_fd_sc_hd__o22ai_2
X_1393_ _1393_/A vssd1 vssd1 vccd1 vccd1 _1393_/X sky130_fd_sc_hd__buf_1
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1729_ _1678_/Y _1293_/B _1747_/X vssd1 vssd1 vccd1 vccd1 _1817_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0962_ data_wdata_o[14] _0953_/X _0916_/X _0955_/X vssd1 vssd1 vccd1 vccd1 _1965_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1445_ _1445_/A vssd1 vssd1 vccd1 vccd1 _1452_/A sky130_fd_sc_hd__buf_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1514_ _1816_/Q vssd1 vssd1 vccd1 vccd1 _1514_/Y sky130_fd_sc_hd__inv_2
X_1376_ data_wdata_o[29] _1365_/X _0922_/X _1367_/X vssd1 vssd1 vccd1 vccd1 _1884_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1161_ _1184_/A vssd1 vssd1 vccd1 vccd1 _1161_/X sky130_fd_sc_hd__buf_1
X_1092_ _1946_/Q _1073_/X _1073_/X _1091_/Y vssd1 vssd1 vccd1 vccd1 _1946_/D sky130_fd_sc_hd__o2bb2ai_2
X_1230_ _1230_/A _1230_/B vssd1 vssd1 vccd1 vccd1 _1718_/S sky130_fd_sc_hd__nor2_2
X_0945_ _0945_/A vssd1 vssd1 vccd1 vccd1 _0945_/X sky130_fd_sc_hd__buf_1
X_1428_ data_addr_o[1] _1419_/X _1393_/X _1420_/X vssd1 vssd1 vccd1 vccd1 _1872_/D
+ sky130_fd_sc_hd__a22o_2
X_1359_ _1359_/A vssd1 vssd1 vccd1 vccd1 _1359_/X sky130_fd_sc_hd__buf_1
XFILLER_50_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1213_ _1213_/A vssd1 vssd1 vccd1 vccd1 _1679_/A sky130_fd_sc_hd__buf_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1144_ _1936_/Q _1139_/X data_rdata_i[29] _1141_/X _0915_/X vssd1 vssd1 vccd1 vccd1
+ _1936_/D sky130_fd_sc_hd__o221a_2
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1075_ _1490_/A vssd1 vssd1 vccd1 vccd1 _1075_/X sky130_fd_sc_hd__buf_1
XFILLER_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0928_ _0928_/A vssd1 vssd1 vccd1 vccd1 _0929_/A sky130_fd_sc_hd__buf_1
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1831_ _1859_/CLK _1831_/D vssd1 vssd1 vccd1 vccd1 _1831_/Q sky130_fd_sc_hd__dfxtp_2
X_1900_ _1943_/CLK _1900_/D vssd1 vssd1 vccd1 vccd1 _1900_/Q sky130_fd_sc_hd__dfxtp_2
X_1762_ _1913_/Q _1921_/Q _1862_/Q vssd1 vssd1 vccd1 vccd1 _1762_/X sky130_fd_sc_hd__mux2_1
X_1693_ _1693_/A vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__buf_1
X_1058_ _1862_/Q _1863_/Q _1058_/C vssd1 vssd1 vccd1 vccd1 _1492_/B sky130_fd_sc_hd__or3_2
X_1127_ _1136_/A _1123_/Y _1483_/C _1123_/A _1456_/A vssd1 vssd1 vccd1 vccd1 _1941_/D
+ sky130_fd_sc_hd__a221oi_2
XFILLER_31_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1745_ _1744_/X _1925_/Q _1864_/Q vssd1 vssd1 vccd1 vccd1 _1745_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1814_ _1950_/CLK _1814_/D vssd1 vssd1 vccd1 vccd1 _1814_/Q sky130_fd_sc_hd__dfxtp_2
X_1676_ _1676_/A _1754_/X vssd1 vssd1 vccd1 vccd1 _1677_/A sky130_fd_sc_hd__or2_2
XFILLER_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1392_ _1392_/A vssd1 vssd1 vccd1 vccd1 _1392_/X sky130_fd_sc_hd__buf_1
X_1461_ _1777_/X _1250_/X _1855_/Q _1458_/X vssd1 vssd1 vccd1 vccd1 _1855_/D sky130_fd_sc_hd__o22a_2
X_1530_ _1809_/Q _1527_/A _1529_/Y _1527_/Y vssd1 vssd1 vccd1 vccd1 _1530_/X sky130_fd_sc_hd__a22o_2
X_1728_ _1675_/Y _1293_/C _1747_/X vssd1 vssd1 vccd1 vccd1 _1816_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1753__A1 rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1659_ _1748_/X _1650_/X _1655_/B _1658_/X vssd1 vssd1 vccd1 vccd1 _1659_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0961_ _0961_/A vssd1 vssd1 vccd1 vccd1 _0961_/X sky130_fd_sc_hd__buf_1
XFILLER_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1375_ _1375_/A vssd1 vssd1 vccd1 vccd1 _1375_/X sky130_fd_sc_hd__buf_1
XFILLER_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1513_ _1815_/Q _1511_/B _1512_/Y vssd1 vssd1 vccd1 vccd1 _1513_/Y sky130_fd_sc_hd__a21oi_2
X_1444_ _1444_/A vssd1 vssd1 vccd1 vccd1 _1444_/X sky130_fd_sc_hd__buf_1
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1091_ _1075_/X _1770_/X _1090_/X _1077_/X vssd1 vssd1 vccd1 vccd1 _1091_/Y sky130_fd_sc_hd__a22oi_2
X_1160_ _1369_/A vssd1 vssd1 vccd1 vccd1 _1184_/A sky130_fd_sc_hd__buf_1
X_0944_ _0948_/A vssd1 vssd1 vccd1 vccd1 _0945_/A sky130_fd_sc_hd__buf_1
XFILLER_9_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1427_ _1427_/A vssd1 vssd1 vccd1 vccd1 _1427_/X sky130_fd_sc_hd__buf_1
XFILLER_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1358_ _1361_/A vssd1 vssd1 vccd1 vccd1 _1359_/A sky130_fd_sc_hd__buf_1
X_1289_ _1757_/X vssd1 vssd1 vccd1 vccd1 _1308_/B sky130_fd_sc_hd__inv_2
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1212_ _1949_/Q _1263_/B vssd1 vssd1 vccd1 vccd1 _1212_/X sky130_fd_sc_hd__and2_2
X_1143_ _1937_/Q _1139_/X data_rdata_i[30] _1141_/X _0915_/X vssd1 vssd1 vccd1 vccd1
+ _1937_/D sky130_fd_sc_hd__o221a_2
XFILLER_1_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1074_ _1866_/Q vssd1 vssd1 vccd1 vccd1 _1490_/A sky130_fd_sc_hd__buf_1
X_0927_ data_wdata_o[20] _0907_/X _0926_/X _0910_/X vssd1 vssd1 vccd1 vccd1 _1971_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1830_ _1940_/CLK _1830_/D vssd1 vssd1 vccd1 vccd1 _1830_/Q sky130_fd_sc_hd__dfxtp_2
X_1761_ _1758_/X _1666_/Y _1761_/S vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__mux2_1
X_1692_ _1682_/X _1714_/X vssd1 vssd1 vccd1 vccd1 _1693_/A sky130_fd_sc_hd__and2b_2
X_1126_ _1432_/A vssd1 vssd1 vccd1 vccd1 _1456_/A sky130_fd_sc_hd__buf_1
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1057_ _1866_/Q vssd1 vssd1 vccd1 vccd1 _1485_/A sky130_fd_sc_hd__inv_2
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1959_ _1972_/CLK _1959_/D _0982_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[8] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1744_ _1909_/Q _1917_/Q _1862_/Q vssd1 vssd1 vccd1 vccd1 _1744_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1813_ _1950_/CLK _1813_/D vssd1 vssd1 vccd1 vccd1 _1813_/Q sky130_fd_sc_hd__dfxtp_2
X_1675_ _1739_/X _1650_/X _1756_/X _1658_/X vssd1 vssd1 vccd1 vccd1 _1675_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1109_ _1706_/X _1942_/Q _1109_/S vssd1 vssd1 vccd1 vccd1 _1110_/A sky130_fd_sc_hd__mux2_2
XFILLER_42_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1391_ _1399_/A vssd1 vssd1 vccd1 vccd1 _1392_/A sky130_fd_sc_hd__buf_1
X_1460_ _1776_/X _1240_/X _1856_/Q _1458_/X vssd1 vssd1 vccd1 vccd1 _1856_/D sky130_fd_sc_hd__o22a_2
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1727_ _1672_/Y _1308_/B _1747_/X vssd1 vssd1 vccd1 vccd1 _1815_/D sky130_fd_sc_hd__mux2_1
X_1658_ _1658_/A _1658_/B vssd1 vssd1 vccd1 vccd1 _1658_/X sky130_fd_sc_hd__and2_2
X_1589_ _1634_/A _1821_/Q vssd1 vssd1 vccd1 vccd1 _1589_/Y sky130_fd_sc_hd__nor2_2
XFILLER_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0960_ _0969_/A vssd1 vssd1 vccd1 vccd1 _0961_/A sky130_fd_sc_hd__buf_1
XFILLER_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1196__B1 data_rdata_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1512_ _1515_/B vssd1 vssd1 vccd1 vccd1 _1512_/Y sky130_fd_sc_hd__inv_2
X_1374_ _1380_/A vssd1 vssd1 vccd1 vccd1 _1375_/A sky130_fd_sc_hd__buf_1
X_1443_ _1443_/A vssd1 vssd1 vccd1 vccd1 _1444_/A sky130_fd_sc_hd__buf_1
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1178__B1 data_rdata_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1090_ _1847_/Q vssd1 vssd1 vccd1 vccd1 _1090_/X sky130_fd_sc_hd__buf_1
X_0943_ data_wdata_o[17] _0930_/X _0942_/X _0932_/X vssd1 vssd1 vccd1 vccd1 _1968_/D
+ sky130_fd_sc_hd__a22o_2
XANTENNA__1169__B1 data_rdata_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1426_ _1434_/A vssd1 vssd1 vccd1 vccd1 _1427_/A sky130_fd_sc_hd__buf_1
X_1288_ rx_i _1646_/A vssd1 vssd1 vccd1 vccd1 _1288_/Y sky130_fd_sc_hd__nor2_2
X_1357_ data_addr_o[9] _1347_/X _0942_/X _1349_/X vssd1 vssd1 vccd1 vccd1 _1888_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_11_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1142_ _1938_/Q _1139_/X data_rdata_i[31] _1141_/X _0915_/X vssd1 vssd1 vccd1 vccd1
+ _1938_/D sky130_fd_sc_hd__o221a_2
X_1211_ _1217_/A vssd1 vssd1 vccd1 vccd1 _1263_/B sky130_fd_sc_hd__buf_1
XFILLER_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1073_ _1096_/A vssd1 vssd1 vccd1 vccd1 _1073_/X sky130_fd_sc_hd__buf_1
X_0926_ _1847_/Q vssd1 vssd1 vccd1 vccd1 _0926_/X sky130_fd_sc_hd__buf_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1409_ data_addr_o[6] _1401_/X _1408_/X _1403_/X vssd1 vssd1 vccd1 vccd1 _1877_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1691_ _1691_/A vssd1 vssd1 vccd1 vccd1 _1691_/X sky130_fd_sc_hd__buf_1
X_1760_ _1647_/A rx_i _1761_/S vssd1 vssd1 vccd1 vccd1 _1760_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1125_ rst_i vssd1 vssd1 vccd1 vccd1 _1432_/A sky130_fd_sc_hd__buf_1
X_1056_ _1330_/A _1062_/A vssd1 vssd1 vccd1 vccd1 _1402_/A sky130_fd_sc_hd__or2_2
X_0909_ _0930_/A vssd1 vssd1 vccd1 vccd1 _0932_/A sky130_fd_sc_hd__inv_2
X_1958_ _1972_/CLK _1958_/D _0985_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[7] sky130_fd_sc_hd__dfrtp_2
X_1889_ _1972_/CLK _1889_/D _1353_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[10] sky130_fd_sc_hd__dfrtp_2
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1743_ _1742_/X _1936_/Q _1860_/Q vssd1 vssd1 vccd1 vccd1 _1743_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1674_ _1674_/A vssd1 vssd1 vccd1 vccd1 _1674_/X sky130_fd_sc_hd__buf_1
XFILLER_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1812_ _1950_/CLK _1812_/D vssd1 vssd1 vccd1 vccd1 _1812_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1039_ _1066_/A _1039_/B vssd1 vssd1 vccd1 vccd1 _1039_/X sky130_fd_sc_hd__or2_2
X_1108_ _1108_/A vssd1 vssd1 vccd1 vccd1 _1108_/X sky130_fd_sc_hd__buf_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1390_ data_wdata_o[26] _1382_/X _1389_/X _1384_/X vssd1 vssd1 vccd1 vccd1 _1881_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1726_ _1668_/Y _1666_/B _1747_/X vssd1 vssd1 vccd1 vccd1 _1814_/D sky130_fd_sc_hd__mux2_1
X_1657_ _1661_/A _1657_/B vssd1 vssd1 vccd1 vccd1 _1658_/B sky130_fd_sc_hd__or2_2
X_1588_ _1687_/A vssd1 vssd1 vccd1 vccd1 _1634_/A sky130_fd_sc_hd__buf_1
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0943__A1 data_wdata_o[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1511_ _1815_/Q _1511_/B vssd1 vssd1 vccd1 vccd1 _1515_/B sky130_fd_sc_hd__or2_2
X_1442_ _1442_/A vssd1 vssd1 vccd1 vccd1 _1442_/X sky130_fd_sc_hd__buf_1
X_1373_ data_wdata_o[30] _1365_/X _0916_/X _1367_/X vssd1 vssd1 vccd1 vccd1 _1885_/D
+ sky130_fd_sc_hd__a22o_2
Xclkbuf_4_15_0_clk_i clkbuf_3_7_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1974_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_23_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1709_ _1640_/X _1050_/X _1715_/S vssd1 vssd1 vccd1 vccd1 _1709_/X sky130_fd_sc_hd__mux2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1350__A1 data_addr_o[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0942_ _1393_/A vssd1 vssd1 vccd1 vccd1 _0942_/X sky130_fd_sc_hd__buf_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1425_ data_addr_o[2] _1419_/X _1389_/X _1420_/X vssd1 vssd1 vccd1 vccd1 _1873_/D
+ sky130_fd_sc_hd__a22o_2
X_1356_ _1356_/A vssd1 vssd1 vccd1 vccd1 _1356_/X sky130_fd_sc_hd__buf_1
X_1287_ _1647_/C _1287_/B vssd1 vssd1 vccd1 vccd1 _1646_/A sky130_fd_sc_hd__or2_2
XFILLER_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1141_ _1164_/A vssd1 vssd1 vccd1 vccd1 _1141_/X sky130_fd_sc_hd__buf_1
X_1072_ _1109_/S vssd1 vssd1 vccd1 vccd1 _1096_/A sky130_fd_sc_hd__buf_1
XFILLER_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1210_ _1213_/A _1738_/S vssd1 vssd1 vccd1 vccd1 _1217_/A sky130_fd_sc_hd__or2_2
X_1974_ _1974_/CLK _1974_/D _1695_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[23] sky130_fd_sc_hd__dfrtp_2
X_0925_ _0925_/A vssd1 vssd1 vccd1 vccd1 _0925_/X sky130_fd_sc_hd__buf_1
X_1408_ _1849_/Q vssd1 vssd1 vccd1 vccd1 _1408_/X sky130_fd_sc_hd__buf_1
X_1339_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1339_/X sky130_fd_sc_hd__buf_1
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1690_ _1682_/X _1713_/X vssd1 vssd1 vccd1 vccd1 _1691_/A sky130_fd_sc_hd__and2b_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1124_ _1941_/Q vssd1 vssd1 vccd1 vccd1 _1483_/C sky130_fd_sc_hd__inv_2
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1055_ _1867_/Q vssd1 vssd1 vccd1 vccd1 _1330_/A sky130_fd_sc_hd__inv_2
X_1957_ _1972_/CLK _1957_/D _0995_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[6] sky130_fd_sc_hd__dfrtp_2
X_0908_ _1850_/Q vssd1 vssd1 vccd1 vccd1 _0908_/X sky130_fd_sc_hd__buf_1
X_1888_ _1972_/CLK _1888_/D _1356_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[9] sky130_fd_sc_hd__dfrtp_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1811_ _1903_/CLK _1811_/D vssd1 vssd1 vccd1 vccd1 _1811_/Q sky130_fd_sc_hd__dfxtp_2
X_1742_ _1741_/X _1928_/Q _1864_/Q vssd1 vssd1 vccd1 vccd1 _1742_/X sky130_fd_sc_hd__mux2_1
X_1673_ _1676_/A _1756_/X vssd1 vssd1 vccd1 vccd1 _1674_/A sky130_fd_sc_hd__or2_2
X_1038_ _1950_/Q vssd1 vssd1 vccd1 vccd1 _1332_/A sky130_fd_sc_hd__buf_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1107_ _1107_/A vssd1 vssd1 vccd1 vccd1 _1108_/A sky130_fd_sc_hd__buf_1
XFILLER_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1725_ _1665_/Y _1755_/X _1747_/X vssd1 vssd1 vccd1 vccd1 _1813_/D sky130_fd_sc_hd__mux2_1
X_1587_ _1666_/A _1587_/B vssd1 vssd1 vccd1 vccd1 _1587_/Y sky130_fd_sc_hd__nor2_2
X_1656_ _1656_/A vssd1 vssd1 vccd1 vccd1 _1656_/X sky130_fd_sc_hd__buf_1
XANTENNA__1047__B data_rvalid_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_clk_i clkbuf_3_5_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1972_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1510_ _1815_/Q vssd1 vssd1 vccd1 vccd1 _1510_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1441_ _1443_/A vssd1 vssd1 vccd1 vccd1 _1442_/A sky130_fd_sc_hd__buf_1
X_1372_ _1372_/A vssd1 vssd1 vccd1 vccd1 _1372_/X sky130_fd_sc_hd__buf_1
XFILLER_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1708_ _1639_/X _1532_/B _1715_/S vssd1 vssd1 vccd1 vccd1 _1708_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1639_ _1490_/X _1743_/X _1412_/X _1636_/X vssd1 vssd1 vccd1 vccd1 _1639_/X sky130_fd_sc_hd__a22o_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0941_ _1844_/Q vssd1 vssd1 vccd1 vccd1 _1393_/A sky130_fd_sc_hd__buf_1
X_1424_ _1424_/A vssd1 vssd1 vccd1 vccd1 _1424_/X sky130_fd_sc_hd__buf_1
X_1355_ _1361_/A vssd1 vssd1 vccd1 vccd1 _1356_/A sky130_fd_sc_hd__buf_1
X_1286_ _1642_/A _1647_/B vssd1 vssd1 vccd1 vccd1 _1287_/B sky130_fd_sc_hd__or2_2
XFILLER_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1140_ _1172_/A vssd1 vssd1 vccd1 vccd1 _1164_/A sky130_fd_sc_hd__buf_1
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1071_ _1034_/A _1051_/X _1060_/X _1064_/Y _1070_/Y vssd1 vssd1 vccd1 vccd1 _1109_/S
+ sky130_fd_sc_hd__o2111ai_2
X_1973_ _1974_/CLK _1973_/D _0915_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[22] sky130_fd_sc_hd__dfrtp_2
X_0924_ _0928_/A vssd1 vssd1 vccd1 vccd1 _0925_/A sky130_fd_sc_hd__buf_1
X_1407_ _1407_/A vssd1 vssd1 vccd1 vccd1 _1407_/X sky130_fd_sc_hd__buf_1
X_1338_ _1344_/A vssd1 vssd1 vccd1 vccd1 _1339_/A sky130_fd_sc_hd__buf_1
XFILLER_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1269_ _1897_/Q _1119_/A _1202_/Y _1203_/X vssd1 vssd1 vccd1 vccd1 _1270_/B sky130_fd_sc_hd__o22a_2
XFILLER_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1123_ _1123_/A vssd1 vssd1 vccd1 vccd1 _1123_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1054_ _1866_/Q _1063_/A vssd1 vssd1 vccd1 vccd1 _1635_/A sky130_fd_sc_hd__or2_2
X_0907_ _0930_/A vssd1 vssd1 vccd1 vccd1 _0907_/X sky130_fd_sc_hd__buf_1
X_1887_ _1971_/CLK _1887_/D _1359_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[8] sky130_fd_sc_hd__dfrtp_2
X_1956_ _1972_/CLK _1956_/D _0998_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[5] sky130_fd_sc_hd__dfrtp_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1741_ _1912_/Q _1920_/Q _1862_/Q vssd1 vssd1 vccd1 vccd1 _1741_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1810_ _1903_/CLK _1810_/D vssd1 vssd1 vccd1 vccd1 _1810_/Q sky130_fd_sc_hd__dfxtp_2
X_1672_ _1757_/X _1658_/X _1287_/B _1671_/X vssd1 vssd1 vccd1 vccd1 _1672_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__1150__B1 data_rdata_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1106_ _1106_/A vssd1 vssd1 vccd1 vccd1 _1943_/D sky130_fd_sc_hd__buf_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1037_ _1532_/A vssd1 vssd1 vccd1 vccd1 _1067_/A sky130_fd_sc_hd__inv_2
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1939_ _1941_/CLK _1939_/D vssd1 vssd1 vccd1 vccd1 _1939_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1199__B1 data_rdata_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1724_ _1659_/Y _1308_/D _1747_/X vssd1 vssd1 vccd1 vccd1 _1812_/D sky130_fd_sc_hd__mux2_1
X_1655_ _1666_/A _1655_/B vssd1 vssd1 vccd1 vccd1 _1656_/A sky130_fd_sc_hd__or2_2
X_1586_ _1586_/A _1586_/B vssd1 vssd1 vccd1 vccd1 _1586_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__1047__C data_gnt_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1665__A1 _1557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1371_ _1380_/A vssd1 vssd1 vccd1 vccd1 _1372_/A sky130_fd_sc_hd__buf_1
X_1440_ _1440_/A vssd1 vssd1 vccd1 vccd1 _1440_/X sky130_fd_sc_hd__buf_1
XFILLER_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1638_ _1490_/X _1767_/X _1393_/X _1636_/X vssd1 vssd1 vccd1 vccd1 _1638_/X sky130_fd_sc_hd__a22o_2
X_1707_ _1638_/X _1067_/Y _1715_/S vssd1 vssd1 vccd1 vccd1 _1707_/X sky130_fd_sc_hd__mux2_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _1569_/A vssd1 vssd1 vccd1 vccd1 _1569_/X sky130_fd_sc_hd__buf_1
Xclkbuf_4_9_0_clk_i clkbuf_4_9_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1971_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0940_ _0940_/A vssd1 vssd1 vccd1 vccd1 _0940_/X sky130_fd_sc_hd__buf_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1423_ _1434_/A vssd1 vssd1 vccd1 vccd1 _1424_/A sky130_fd_sc_hd__buf_1
X_1285_ _1647_/A vssd1 vssd1 vccd1 vccd1 _1642_/A sky130_fd_sc_hd__inv_2
X_1354_ data_addr_o[10] _1347_/X _0937_/X _1349_/X vssd1 vssd1 vccd1 vccd1 _1889_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1070_ _1868_/Q _1331_/A _1533_/B _1495_/A vssd1 vssd1 vccd1 vccd1 _1070_/Y sky130_fd_sc_hd__a31oi_2
X_1972_ _1972_/CLK _1972_/D _0921_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[21] sky130_fd_sc_hd__dfrtp_2
X_0923_ data_wdata_o[21] _0907_/X _0922_/X _0910_/X vssd1 vssd1 vccd1 vccd1 _1972_/D
+ sky130_fd_sc_hd__a22o_2
X_1406_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1407_/A sky130_fd_sc_hd__buf_1
X_1337_ _1332_/A _1419_/A _1115_/B _1336_/X vssd1 vssd1 vccd1 vccd1 _1892_/D sky130_fd_sc_hd__o22ai_2
X_1268_ _1022_/X _1034_/X _1898_/Q _1039_/B vssd1 vssd1 vccd1 vccd1 _1898_/D sky130_fd_sc_hd__a2bb2o_2
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1199_ _1907_/Q _1193_/X data_rdata_i[0] _1194_/X _1198_/X vssd1 vssd1 vccd1 vccd1
+ _1907_/D sky130_fd_sc_hd__o221a_2
XFILLER_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_6_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1122_ _1128_/A _1122_/B vssd1 vssd1 vccd1 vccd1 _1123_/A sky130_fd_sc_hd__or2_2
XFILLER_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1053_ _1867_/Q _1868_/Q _1869_/Q vssd1 vssd1 vccd1 vccd1 _1063_/A sky130_fd_sc_hd__or3_2
X_0906_ _1860_/Q _0906_/B _1535_/B vssd1 vssd1 vccd1 vccd1 _0930_/A sky130_fd_sc_hd__or3_2
X_1886_ _1972_/CLK _1886_/D _1362_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[31] sky130_fd_sc_hd__dfrtp_2
X_1955_ _1972_/CLK _1955_/D _1001_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[4] sky130_fd_sc_hd__dfrtp_2
XANTENNA__1066__B uart_error vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0973__A1 data_wdata_o[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1671_ _1671_/A _1712_/X vssd1 vssd1 vccd1 vccd1 _1671_/X sky130_fd_sc_hd__and2_2
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1740_ _1465_/B _1738_/S _1740_/S vssd1 vssd1 vccd1 vccd1 _1740_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1105_ _1707_/X _1943_/Q _1109_/S vssd1 vssd1 vccd1 vccd1 _1106_/A sky130_fd_sc_hd__mux2_2
XFILLER_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1036_ _1039_/B vssd1 vssd1 vccd1 vccd1 _1036_/Y sky130_fd_sc_hd__inv_2
X_1938_ _1938_/CLK _1938_/D vssd1 vssd1 vccd1 vccd1 _1938_/Q sky130_fd_sc_hd__dfxtp_2
X_1869_ _1876_/CLK _1869_/D _1435_/X vssd1 vssd1 vccd1 vccd1 _1869_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1654_ _1749_/S _1647_/X _1287_/B _1652_/X _1653_/X vssd1 vssd1 vccd1 vccd1 _1654_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1723_ _1251_/A _1718_/X _1740_/S vssd1 vssd1 vccd1 vccd1 _1723_/X sky130_fd_sc_hd__mux2_1
X_1585_ _1586_/B vssd1 vssd1 vccd1 vccd1 _1585_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1019_ _1019_/A vssd1 vssd1 vccd1 vccd1 _1019_/X sky130_fd_sc_hd__buf_1
Xclkbuf_4_5_0_clk_i clkbuf_4_5_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1949_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1370_ _1422_/A vssd1 vssd1 vccd1 vccd1 _1380_/A sky130_fd_sc_hd__buf_1
XFILLER_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1637_ _1490_/X _1703_/X _1397_/X _1636_/X vssd1 vssd1 vccd1 vccd1 _1637_/X sky130_fd_sc_hd__a22o_2
X_1706_ _1637_/X _1532_/Y _1715_/S vssd1 vssd1 vccd1 vccd1 _1706_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1499_/A vssd1 vssd1 vccd1 vccd1 _1860_/D sky130_fd_sc_hd__buf_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ _1582_/A _1568_/B vssd1 vssd1 vccd1 vccd1 _1569_/A sky130_fd_sc_hd__and2_2
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1265__A _1351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1422_ _1422_/A vssd1 vssd1 vccd1 vccd1 _1434_/A sky130_fd_sc_hd__buf_1
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1284_ _1316_/A vssd1 vssd1 vccd1 vccd1 _1284_/Y sky130_fd_sc_hd__inv_2
X_1353_ _1353_/A vssd1 vssd1 vccd1 vccd1 _1353_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0_clk_i clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0999_ data_wdata_o[5] _0989_/X _0922_/X _0991_/X vssd1 vssd1 vccd1 vccd1 _1956_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_2_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0922_ _1848_/Q vssd1 vssd1 vccd1 vccd1 _0922_/X sky130_fd_sc_hd__buf_1
X_1971_ _1971_/CLK _1971_/D _0925_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[20] sky130_fd_sc_hd__dfrtp_2
X_1405_ _1422_/A vssd1 vssd1 vccd1 vccd1 _1417_/A sky130_fd_sc_hd__buf_1
X_1198_ _1198_/A vssd1 vssd1 vccd1 vccd1 _1198_/X sky130_fd_sc_hd__buf_1
X_1336_ _1330_/X _1334_/X _1335_/X vssd1 vssd1 vccd1 vccd1 _1336_/X sky130_fd_sc_hd__o21a_2
X_1267_ _1267_/A vssd1 vssd1 vccd1 vccd1 _1267_/X sky130_fd_sc_hd__buf_1
XFILLER_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1121_ _1940_/Q _1117_/B _1133_/A _1340_/B data_gnt_i vssd1 vssd1 vccd1 vccd1 _1122_/B
+ sky130_fd_sc_hd__a32o_2
XFILLER_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1052_ _1865_/Q vssd1 vssd1 vccd1 vccd1 _1498_/A sky130_fd_sc_hd__buf_1
XFILLER_33_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1954_ _1972_/CLK _1954_/D _1004_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[3] sky130_fd_sc_hd__dfrtp_2
X_1885_ _1974_/CLK _1885_/D _1372_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[30] sky130_fd_sc_hd__dfrtp_2
X_0905_ _0952_/C vssd1 vssd1 vccd1 vccd1 _1535_/B sky130_fd_sc_hd__buf_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1319_ _1895_/Q _1274_/A _1313_/A _1313_/B vssd1 vssd1 vccd1 vccd1 _1319_/X sky130_fd_sc_hd__o22a_2
XFILLER_21_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1670_ _1670_/A vssd1 vssd1 vccd1 vccd1 _1670_/X sky130_fd_sc_hd__buf_1
X_1104_ _1104_/A vssd1 vssd1 vccd1 vccd1 _1104_/X sky130_fd_sc_hd__buf_1
X_1035_ _1532_/A _1022_/X _1068_/C _1034_/X vssd1 vssd1 vccd1 vccd1 _1039_/B sky130_fd_sc_hd__a31o_2
X_1937_ _1938_/CLK _1937_/D vssd1 vssd1 vccd1 vccd1 _1937_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1799_ _1557_/B _1558_/X _1802_/S vssd1 vssd1 vccd1 vccd1 _1835_/D sky130_fd_sc_hd__mux2_1
X_1868_ _1971_/CLK _1868_/D _1438_/X vssd1 vssd1 vccd1 vccd1 _1868_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1093__A _1351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_clk_i clkbuf_4_1_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1903_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1584_ _1841_/Q _1579_/X _1298_/Y vssd1 vssd1 vccd1 vccd1 _1586_/B sky130_fd_sc_hd__a21oi_2
X_1653_ _1818_/Q _1819_/Q _1653_/C _1761_/S vssd1 vssd1 vccd1 vccd1 _1653_/X sky130_fd_sc_hd__or4_2
X_1722_ _1654_/Y _1664_/B _1722_/S vssd1 vssd1 vccd1 vccd1 _1820_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1018_ _1018_/A vssd1 vssd1 vccd1 vccd1 _1019_/A sky130_fd_sc_hd__buf_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1705_ _1647_/B _1586_/A _1761_/S vssd1 vssd1 vccd1 vccd1 _1705_/X sky130_fd_sc_hd__mux2_1
X_1636_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1636_/X sky130_fd_sc_hd__buf_1
X_1567_ _1567_/A vssd1 vssd1 vccd1 vccd1 _1568_/B sky130_fd_sc_hd__buf_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1498_/A _1498_/B _1498_/C vssd1 vssd1 vccd1 vccd1 _1499_/A sky130_fd_sc_hd__or3_2
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1281__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1421_ data_addr_o[3] _1419_/X _1383_/X _1420_/X vssd1 vssd1 vccd1 vccd1 _1874_/D
+ sky130_fd_sc_hd__a22o_2
XANTENNA__1191__A _1198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1283_ _1503_/A _1664_/B _1647_/A vssd1 vssd1 vccd1 vccd1 _1316_/A sky130_fd_sc_hd__or3_2
X_1352_ _1361_/A vssd1 vssd1 vccd1 vccd1 _1353_/A sky130_fd_sc_hd__buf_1
XANTENNA__1014__A1 data_wdata_o[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0998_ _0998_/A vssd1 vssd1 vccd1 vccd1 _0998_/X sky130_fd_sc_hd__buf_1
X_1619_ _1619_/A vssd1 vssd1 vccd1 vccd1 _1620_/B sky130_fd_sc_hd__buf_1
XFILLER_24_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1970_ _1974_/CLK _1970_/D _0929_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[19] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0921_ _0921_/A vssd1 vssd1 vccd1 vccd1 _0921_/X sky130_fd_sc_hd__buf_1
X_1404_ data_addr_o[7] _1401_/X _1076_/X _1403_/X vssd1 vssd1 vccd1 vccd1 _1878_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1335_ _1867_/Q _1498_/A vssd1 vssd1 vccd1 vccd1 _1335_/X sky130_fd_sc_hd__or2_2
X_1197_ _1908_/Q _1193_/X data_rdata_i[1] _1194_/X _1191_/X vssd1 vssd1 vccd1 vccd1
+ _1908_/D sky130_fd_sc_hd__o221a_2
X_1266_ _1344_/A vssd1 vssd1 vccd1 vccd1 _1267_/A sky130_fd_sc_hd__buf_1
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1162__B1 data_rdata_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1120_ _1203_/B vssd1 vssd1 vccd1 vccd1 _1128_/A sky130_fd_sc_hd__buf_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1051_ _1275_/B _1281_/B _1671_/A _1061_/B _1050_/X vssd1 vssd1 vccd1 vccd1 _1051_/X
+ sky130_fd_sc_hd__a41o_2
X_1884_ _1974_/CLK _1884_/D _1375_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[29] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0904_ _0904_/A _1062_/A vssd1 vssd1 vccd1 vccd1 _0952_/C sky130_fd_sc_hd__or2_2
X_1953_ _1972_/CLK _1953_/D _1010_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[2] sky130_fd_sc_hd__dfrtp_2
X_1318_ _1325_/A vssd1 vssd1 vccd1 vccd1 _1476_/A sky130_fd_sc_hd__buf_1
X_1249_ _1687_/A _1891_/Q _1198_/X _1248_/X vssd1 vssd1 vccd1 vccd1 _1903_/D sky130_fd_sc_hd__o211a_2
XFILLER_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1144__B1 data_rdata_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1103_ _1107_/A vssd1 vssd1 vccd1 vccd1 _1104_/A sky130_fd_sc_hd__buf_1
X_1034_ _1034_/A uart_error _1532_/B vssd1 vssd1 vccd1 vccd1 _1034_/X sky130_fd_sc_hd__or3_2
X_1936_ _1938_/CLK _1936_/D vssd1 vssd1 vccd1 vccd1 _1936_/Q sky130_fd_sc_hd__dfxtp_2
X_1867_ _1941_/CLK _1867_/D _1440_/X vssd1 vssd1 vccd1 vccd1 _1867_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1798_ _1563_/B _1564_/X _1802_/S vssd1 vssd1 vccd1 vccd1 _1836_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1721_ _1651_/Y _1642_/A _1722_/S vssd1 vssd1 vccd1 vccd1 _1819_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1583_ _1583_/A vssd1 vssd1 vccd1 vccd1 _1583_/X sky130_fd_sc_hd__buf_1
X_1652_ _1671_/A _1730_/X vssd1 vssd1 vccd1 vccd1 _1652_/X sky130_fd_sc_hd__and2_2
X_1017_ data_wdata_o[0] _1005_/X _0946_/X _1006_/X vssd1 vssd1 vccd1 vccd1 _1951_/D
+ sky130_fd_sc_hd__a22o_2
X_1919_ _1930_/CLK _1919_/D vssd1 vssd1 vccd1 vccd1 _1919_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1704_ _1647_/B _1645_/X _1761_/S vssd1 vssd1 vccd1 vccd1 _1704_/X sky130_fd_sc_hd__mux2_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _1330_/A _1487_/X _1364_/A vssd1 vssd1 vccd1 vccd1 _1498_/C sky130_fd_sc_hd__a21oi_2
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1566_ _1837_/Q _1565_/B _1570_/B vssd1 vssd1 vccd1 vccd1 _1567_/A sky130_fd_sc_hd__a21bo_2
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1635_ _1635_/A vssd1 vssd1 vccd1 vccd1 _1715_/S sky130_fd_sc_hd__inv_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1420_ _1498_/B vssd1 vssd1 vccd1 vccd1 _1420_/X sky130_fd_sc_hd__buf_1
X_1351_ _1351_/A vssd1 vssd1 vccd1 vccd1 _1361_/A sky130_fd_sc_hd__buf_1
XFILLER_48_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1282_ _1282_/A vssd1 vssd1 vccd1 vccd1 _1647_/A sky130_fd_sc_hd__buf_1
X_1618_ _1827_/Q _1611_/X _1617_/X vssd1 vssd1 vccd1 vccd1 _1619_/A sky130_fd_sc_hd__a21bo_2
X_0997_ _1003_/A vssd1 vssd1 vccd1 vccd1 _0998_/A sky130_fd_sc_hd__buf_1
X_1549_ _1549_/A vssd1 vssd1 vccd1 vccd1 _1549_/X sky130_fd_sc_hd__buf_1
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1557__A _1557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0920_ _0928_/A vssd1 vssd1 vccd1 vccd1 _0921_/A sky130_fd_sc_hd__buf_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1403_ _1498_/B vssd1 vssd1 vccd1 vccd1 _1403_/X sky130_fd_sc_hd__buf_1
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1334_ _1483_/A _1482_/A _1333_/X vssd1 vssd1 vccd1 vccd1 _1334_/X sky130_fd_sc_hd__o21a_2
X_1265_ _1351_/A vssd1 vssd1 vccd1 vccd1 _1344_/A sky130_fd_sc_hd__buf_1
XFILLER_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1196_ _1909_/Q _1193_/X data_rdata_i[2] _1194_/X _1191_/X vssd1 vssd1 vccd1 vccd1
+ _1909_/D sky130_fd_sc_hd__o221a_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1050_ _1050_/A vssd1 vssd1 vccd1 vccd1 _1050_/X sky130_fd_sc_hd__buf_1
X_1883_ _1965_/CLK _1883_/D _1378_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[28] sky130_fd_sc_hd__dfrtp_2
X_0903_ _1818_/Q _1281_/B _1046_/A vssd1 vssd1 vccd1 vccd1 _1062_/A sky130_fd_sc_hd__or3_2
X_1952_ _1972_/CLK _1952_/D _1013_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[1] sky130_fd_sc_hd__dfrtp_2
X_1317_ _1658_/A _1749_/S vssd1 vssd1 vccd1 vccd1 _1325_/A sky130_fd_sc_hd__or2_2
X_1248_ _1614_/A hold1/A _1859_/Q vssd1 vssd1 vccd1 vccd1 _1248_/X sky130_fd_sc_hd__or3_2
X_1179_ _1193_/A vssd1 vssd1 vccd1 vccd1 _1179_/X sky130_fd_sc_hd__buf_1
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1102_ _1944_/Q _1096_/X _1096_/X _1101_/Y vssd1 vssd1 vccd1 vccd1 _1944_/D sky130_fd_sc_hd__o2bb2ai_2
X_1033_ _1050_/A vssd1 vssd1 vccd1 vccd1 _1532_/B sky130_fd_sc_hd__inv_2
XFILLER_21_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1935_ _1938_/CLK _1935_/D vssd1 vssd1 vccd1 vccd1 _1935_/Q sky130_fd_sc_hd__dfxtp_2
X_1797_ _1568_/B _1569_/X _1802_/S vssd1 vssd1 vccd1 vccd1 _1837_/D sky130_fd_sc_hd__mux2_1
X_1866_ _1941_/CLK _1866_/D _1442_/X vssd1 vssd1 vccd1 vccd1 _1866_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1651_ _1760_/X _1650_/X _1759_/X _1647_/X _1658_/A vssd1 vssd1 vccd1 vccd1 _1651_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1720_ _1649_/Y _1747_/S _1722_/S vssd1 vssd1 vccd1 vccd1 _1818_/D sky130_fd_sc_hd__mux2_1
X_1582_ _1582_/A _1582_/B vssd1 vssd1 vccd1 vccd1 _1583_/A sky130_fd_sc_hd__and2_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1016_ _1016_/A vssd1 vssd1 vccd1 vccd1 _1016_/X sky130_fd_sc_hd__buf_1
X_1918_ _1949_/CLK _1918_/D vssd1 vssd1 vccd1 vccd1 _1918_/Q sky130_fd_sc_hd__dfxtp_2
X_1849_ _1938_/CLK _1849_/D vssd1 vssd1 vccd1 vccd1 _1849_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1703_ _1702_/X _1931_/Q _1860_/Q vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1634_ _1634_/A _1634_/B vssd1 vssd1 vccd1 vccd1 _1634_/Y sky130_fd_sc_hd__nor2_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _1837_/Q _1565_/B vssd1 vssd1 vccd1 vccd1 _1570_/B sky130_fd_sc_hd__or2_2
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _1496_/A vssd1 vssd1 vccd1 vccd1 _1865_/D sky130_fd_sc_hd__buf_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1281_ rst_i _1281_/B vssd1 vssd1 vccd1 vccd1 _1282_/A sky130_fd_sc_hd__or2_2
X_1350_ data_addr_o[11] _1347_/X _0931_/X _1349_/X vssd1 vssd1 vccd1 vccd1 _1890_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0996_ data_wdata_o[6] _0989_/X _0916_/X _0991_/X vssd1 vssd1 vccd1 vccd1 _1957_/D
+ sky130_fd_sc_hd__a22o_2
X_1617_ _1826_/Q _1827_/Q _1617_/C vssd1 vssd1 vccd1 vccd1 _1617_/X sky130_fd_sc_hd__or3_2
X_1479_ _1389_/X _1476_/X _1383_/X _1477_/X vssd1 vssd1 vccd1 vccd1 _1845_/D sky130_fd_sc_hd__a22o_2
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1548_ _1666_/A _1548_/B vssd1 vssd1 vccd1 vccd1 _1549_/A sky130_fd_sc_hd__or2_2
XANTENNA_clkbuf_3_7_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1402_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1498_/B sky130_fd_sc_hd__inv_2
XFILLER_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1264_ _1240_/A _1263_/Y _1899_/Q _1241_/X vssd1 vssd1 vccd1 vccd1 _1899_/D sky130_fd_sc_hd__o22a_2
X_1333_ _1333_/A _1533_/A vssd1 vssd1 vccd1 vccd1 _1333_/X sky130_fd_sc_hd__or2_2
X_1195_ _1910_/Q _1193_/X data_rdata_i[3] _1194_/X _1191_/X vssd1 vssd1 vccd1 vccd1
+ _1910_/D sky130_fd_sc_hd__o221a_2
X_0979_ _0979_/A vssd1 vssd1 vccd1 vccd1 _0979_/X sky130_fd_sc_hd__buf_1
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1882_ _1974_/CLK _1882_/D _1381_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[27] sky130_fd_sc_hd__dfrtp_2
X_0902_ _1820_/Q vssd1 vssd1 vccd1 vccd1 _1046_/A sky130_fd_sc_hd__inv_2
X_1951_ _1972_/CLK _1951_/D _1016_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[0] sky130_fd_sc_hd__dfrtp_2
X_1178_ _1919_/Q _1171_/X data_rdata_i[12] _1173_/X _1177_/X vssd1 vssd1 vccd1 vccd1
+ _1919_/D sky130_fd_sc_hd__o221a_2
X_1316_ _1316_/A vssd1 vssd1 vccd1 vccd1 _1658_/A sky130_fd_sc_hd__buf_1
X_1247_ _1870_/Q vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__inv_2
XFILLER_24_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1101_ _1490_/A _1746_/X _1845_/Q _1636_/A vssd1 vssd1 vccd1 vccd1 _1101_/Y sky130_fd_sc_hd__a22oi_2
X_1032_ _1898_/Q _1331_/A vssd1 vssd1 vccd1 vccd1 _1050_/A sky130_fd_sc_hd__or2_2
X_1934_ _1938_/CLK _1934_/D vssd1 vssd1 vccd1 vccd1 _1934_/Q sky130_fd_sc_hd__dfxtp_2
X_1796_ _1572_/Y _1573_/Y _1802_/S vssd1 vssd1 vccd1 vccd1 _1838_/D sky130_fd_sc_hd__mux2_1
X_1865_ _1941_/CLK _1865_/D _1444_/X vssd1 vssd1 vccd1 vccd1 _1865_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1581_ _1581_/A vssd1 vssd1 vccd1 vccd1 _1582_/B sky130_fd_sc_hd__buf_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1650_ _1650_/A vssd1 vssd1 vccd1 vccd1 _1650_/X sky130_fd_sc_hd__buf_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1015_ _1018_/A vssd1 vssd1 vccd1 vccd1 _1016_/A sky130_fd_sc_hd__buf_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1917_ _1949_/CLK _1917_/D vssd1 vssd1 vccd1 vccd1 _1917_/Q sky130_fd_sc_hd__dfxtp_2
X_1848_ _1876_/CLK _1848_/D vssd1 vssd1 vccd1 vccd1 _1848_/Q sky130_fd_sc_hd__dfxtp_2
X_1779_ _1943_/Q _1854_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _1779_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1702_ _1701_/X _1923_/Q _1864_/Q vssd1 vssd1 vccd1 vccd1 _1702_/X sky130_fd_sc_hd__mux2_1
X_1633_ _1633_/A vssd1 vssd1 vccd1 vccd1 _1633_/X sky130_fd_sc_hd__buf_1
X_1564_ _1564_/A vssd1 vssd1 vccd1 vccd1 _1564_/X sky130_fd_sc_hd__buf_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1495_/A _1495_/B vssd1 vssd1 vccd1 vccd1 _1496_/A sky130_fd_sc_hd__or2_2
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1192__B1 data_rdata_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1280_ _1653_/C vssd1 vssd1 vccd1 vccd1 _1664_/B sky130_fd_sc_hd__inv_2
XFILLER_8_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0995_ _0995_/A vssd1 vssd1 vccd1 vccd1 _0995_/X sky130_fd_sc_hd__buf_1
XANTENNA__1183__B1 data_rdata_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1616_ _1616_/A vssd1 vssd1 vccd1 vccd1 _1616_/X sky130_fd_sc_hd__buf_1
X_1547_ _1661_/A vssd1 vssd1 vccd1 vccd1 _1666_/A sky130_fd_sc_hd__buf_1
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1478_ _1383_/X _1476_/X _1090_/X _1477_/X vssd1 vssd1 vccd1 vccd1 _1846_/D sky130_fd_sc_hd__a22o_2
XANTENNA__1174__B1 data_rdata_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1165__B1 data_rdata_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1401_ _1419_/A vssd1 vssd1 vccd1 vccd1 _1401_/X sky130_fd_sc_hd__buf_1
X_1194_ _1194_/A vssd1 vssd1 vccd1 vccd1 _1194_/X sky130_fd_sc_hd__buf_1
X_1263_ _1899_/Q _1263_/B vssd1 vssd1 vccd1 vccd1 _1263_/Y sky130_fd_sc_hd__nor2_2
X_1332_ _1332_/A vssd1 vssd1 vccd1 vccd1 _1333_/A sky130_fd_sc_hd__inv_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0978_ _0984_/A vssd1 vssd1 vccd1 vccd1 _0979_/A sky130_fd_sc_hd__buf_1
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1147__B1 data_rdata_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0928__A _0928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1950_ _1950_/CLK _1950_/D _1019_/X vssd1 vssd1 vccd1 vccd1 _1950_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1881_ _1974_/CLK _1881_/D _1388_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[26] sky130_fd_sc_hd__dfrtp_2
X_0901_ _1819_/Q vssd1 vssd1 vccd1 vccd1 _1281_/B sky130_fd_sc_hd__inv_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1315_ _1271_/Y _1313_/X _1312_/A _1314_/X vssd1 vssd1 vccd1 vccd1 _1896_/D sky130_fd_sc_hd__o22ai_2
X_1177_ _1184_/A vssd1 vssd1 vccd1 vccd1 _1177_/X sky130_fd_sc_hd__buf_1
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1246_ _1246_/A vssd1 vssd1 vccd1 vccd1 _1614_/A sky130_fd_sc_hd__inv_2
XFILLER_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1100_ _1100_/A vssd1 vssd1 vccd1 vccd1 _1100_/X sky130_fd_sc_hd__buf_1
X_1031_ _1031_/A vssd1 vssd1 vccd1 vccd1 uart_error sky130_fd_sc_hd__buf_1
X_1933_ _1938_/CLK _1933_/D vssd1 vssd1 vccd1 vccd1 _1933_/Q sky130_fd_sc_hd__dfxtp_2
X_1864_ _1945_/CLK _1864_/D _1447_/X vssd1 vssd1 vccd1 vccd1 _1864_/Q sky130_fd_sc_hd__dfrtp_2
X_1795_ _1577_/B _1578_/X _1802_/S vssd1 vssd1 vccd1 vccd1 _1839_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1229_ _1229_/A _1822_/Q _1229_/C _1229_/D vssd1 vssd1 vccd1 vccd1 _1230_/B sky130_fd_sc_hd__or4_2
XFILLER_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1580_ _1840_/Q _1579_/B _1579_/X vssd1 vssd1 vccd1 vccd1 _1581_/A sky130_fd_sc_hd__a21bo_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1014_ data_wdata_o[1] _1005_/X _0942_/X _1006_/X vssd1 vssd1 vccd1 vccd1 _1952_/D
+ sky130_fd_sc_hd__a22o_2
X_1916_ _1949_/CLK _1916_/D vssd1 vssd1 vccd1 vccd1 _1916_/Q sky130_fd_sc_hd__dfxtp_2
X_1847_ _1876_/CLK _1847_/D vssd1 vssd1 vccd1 vccd1 _1847_/Q sky130_fd_sc_hd__dfxtp_2
X_1778_ _1944_/Q _1855_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _1778_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1701_ _1907_/Q _1915_/Q _1862_/Q vssd1 vssd1 vccd1 vccd1 _1701_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1632_ _1632_/A _1632_/B vssd1 vssd1 vccd1 vccd1 _1633_/A sky130_fd_sc_hd__and2_2
X_1563_ _1582_/A _1563_/B vssd1 vssd1 vccd1 vccd1 _1564_/A sky130_fd_sc_hd__and2_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _1034_/A _1050_/X _1485_/A _1492_/X _1005_/A vssd1 vssd1 vccd1 vccd1 _1495_/B
+ sky130_fd_sc_hd__o221ai_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0994_ _1003_/A vssd1 vssd1 vccd1 vccd1 _0995_/A sky130_fd_sc_hd__buf_1
X_1477_ _1477_/A vssd1 vssd1 vccd1 vccd1 _1477_/X sky130_fd_sc_hd__buf_1
X_1546_ _1546_/A vssd1 vssd1 vccd1 vccd1 _1548_/B sky130_fd_sc_hd__buf_1
X_1615_ _1632_/A _1615_/B vssd1 vssd1 vccd1 vccd1 _1616_/A sky130_fd_sc_hd__and2_2
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1400_ _1400_/A vssd1 vssd1 vccd1 vccd1 _1400_/X sky130_fd_sc_hd__buf_1
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1331_ _1331_/A vssd1 vssd1 vccd1 vccd1 _1482_/A sky130_fd_sc_hd__buf_1
X_1193_ _1193_/A vssd1 vssd1 vccd1 vccd1 _1193_/X sky130_fd_sc_hd__buf_1
X_1262_ _1244_/A _1261_/X _1258_/X _1900_/Q _1240_/A vssd1 vssd1 vccd1 vccd1 _1900_/D
+ sky130_fd_sc_hd__a32o_2
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0977_ data_wdata_o[10] _0971_/X _0937_/X _0972_/X vssd1 vssd1 vccd1 vccd1 _1961_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1529_ _1809_/Q vssd1 vssd1 vccd1 vccd1 _1529_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1965_/CLK _1880_/D _1392_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[25] sky130_fd_sc_hd__dfrtp_2
X_0900_ _1869_/Q vssd1 vssd1 vccd1 vccd1 _0904_/A sky130_fd_sc_hd__inv_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1314_ _1895_/Q _1274_/A _1896_/Q _1284_/Y vssd1 vssd1 vccd1 vccd1 _1314_/X sky130_fd_sc_hd__o31a_2
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1176_ _1920_/Q _1171_/X data_rdata_i[13] _1173_/X _1168_/X vssd1 vssd1 vccd1 vccd1
+ _1920_/D sky130_fd_sc_hd__o221a_2
X_1245_ _1246_/A vssd1 vssd1 vccd1 vccd1 _1687_/A sky130_fd_sc_hd__buf_1
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1368__A1 data_wdata_o[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1030_ _1818_/Q _1281_/B _1647_/C vssd1 vssd1 vccd1 vccd1 _1031_/A sky130_fd_sc_hd__and3_2
X_1932_ _1938_/CLK _1932_/D vssd1 vssd1 vccd1 vccd1 _1932_/Q sky130_fd_sc_hd__dfxtp_2
X_1863_ _1945_/CLK _1863_/D _1449_/X vssd1 vssd1 vccd1 vccd1 _1863_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1794_ _1582_/B _1583_/X _1802_/S vssd1 vssd1 vccd1 vccd1 _1840_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1228_ _1829_/Q _1830_/Q _1823_/Q _1824_/Q vssd1 vssd1 vccd1 vccd1 _1229_/C sky130_fd_sc_hd__or4_2
X_1159_ _1928_/Q _1155_/X data_rdata_i[21] _1156_/X _1153_/X vssd1 vssd1 vccd1 vccd1
+ _1928_/D sky130_fd_sc_hd__o221a_2
XFILLER_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1013_ _1013_/A vssd1 vssd1 vccd1 vccd1 _1013_/X sky130_fd_sc_hd__buf_1
X_1915_ _1949_/CLK _1915_/D vssd1 vssd1 vccd1 vccd1 _1915_/Q sky130_fd_sc_hd__dfxtp_2
X_1846_ _1974_/CLK _1846_/D vssd1 vssd1 vccd1 vccd1 _1846_/Q sky130_fd_sc_hd__dfxtp_2
X_1777_ _1945_/Q _1856_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _1777_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1203__A data_gnt_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1631_ _1630_/Y _1626_/Y _1224_/X vssd1 vssd1 vccd1 vccd1 _1632_/B sky130_fd_sc_hd__o21ai_2
X_1700_ tx_o vssd1 vssd1 vccd1 vccd1 _1700_/X sky130_fd_sc_hd__buf_2
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1562_ _1562_/A vssd1 vssd1 vccd1 vccd1 _1582_/A sky130_fd_sc_hd__buf_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _1330_/X _1483_/X _1490_/X _1492_/X vssd1 vssd1 vccd1 vccd1 _1866_/D sky130_fd_sc_hd__a2bb2o_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1829_ _1859_/CLK _1829_/D vssd1 vssd1 vccd1 vccd1 _1829_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0993_ _1008_/A vssd1 vssd1 vccd1 vccd1 _1003_/A sky130_fd_sc_hd__buf_1
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1614_ _1614_/A vssd1 vssd1 vccd1 vccd1 _1632_/A sky130_fd_sc_hd__buf_1
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_14_0_clk_i clkbuf_3_7_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1965_/CLK sky130_fd_sc_hd__clkbuf_2
X_1476_ _1476_/A vssd1 vssd1 vccd1 vccd1 _1476_/X sky130_fd_sc_hd__buf_1
X_1545_ _1758_/S _1545_/B vssd1 vssd1 vccd1 vccd1 _1546_/A sky130_fd_sc_hd__or2_2
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1330_ _1330_/A vssd1 vssd1 vccd1 vccd1 _1330_/X sky130_fd_sc_hd__buf_1
X_1261_ _1900_/Q _1899_/Q _1256_/Y vssd1 vssd1 vccd1 vccd1 _1261_/X sky130_fd_sc_hd__a21o_2
X_1192_ _1911_/Q _1186_/X data_rdata_i[4] _1187_/X _1191_/X vssd1 vssd1 vccd1 vccd1
+ _1911_/D sky130_fd_sc_hd__o221a_2
X_0976_ _0976_/A vssd1 vssd1 vccd1 vccd1 _0976_/X sky130_fd_sc_hd__buf_1
X_1459_ _1775_/X _1240_/X _1857_/Q _1458_/X vssd1 vssd1 vccd1 vccd1 _1857_/D sky130_fd_sc_hd__o22a_2
X_1528_ _1808_/Q _1526_/B _1527_/Y vssd1 vssd1 vccd1 vccd1 _1528_/X sky130_fd_sc_hd__a21o_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1313_ _1313_/A _1313_/B _1313_/C vssd1 vssd1 vccd1 vccd1 _1313_/X sky130_fd_sc_hd__and3_2
X_1244_ _1244_/A vssd1 vssd1 vccd1 vccd1 _1780_/S sky130_fd_sc_hd__buf_1
X_1175_ _1921_/Q _1171_/X data_rdata_i[14] _1173_/X _1168_/X vssd1 vssd1 vccd1 vccd1
+ _1921_/D sky130_fd_sc_hd__o221a_2
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0959_ _1008_/A vssd1 vssd1 vccd1 vccd1 _0969_/A sky130_fd_sc_hd__buf_1
XFILLER_11_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1931_ _1938_/CLK _1931_/D vssd1 vssd1 vccd1 vccd1 _1931_/Q sky130_fd_sc_hd__dfxtp_2
X_1862_ _1945_/CLK _1862_/D _1451_/X vssd1 vssd1 vccd1 vccd1 _1862_/Q sky130_fd_sc_hd__dfrtp_2
X_1793_ _1585_/Y _1586_/Y _1802_/S vssd1 vssd1 vccd1 vccd1 _1841_/D sky130_fd_sc_hd__mux2_1
X_1158_ _1929_/Q _1155_/X data_rdata_i[22] _1156_/X _1153_/X vssd1 vssd1 vccd1 vccd1
+ _1929_/D sky130_fd_sc_hd__o221a_2
X_1227_ _1821_/Q vssd1 vssd1 vccd1 vccd1 _1229_/A sky130_fd_sc_hd__inv_2
X_1089_ _1089_/A vssd1 vssd1 vccd1 vccd1 _1089_/X sky130_fd_sc_hd__buf_1
XFILLER_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1012_ _1018_/A vssd1 vssd1 vccd1 vccd1 _1013_/A sky130_fd_sc_hd__buf_1
X_1914_ _1930_/CLK _1914_/D vssd1 vssd1 vccd1 vccd1 _1914_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1845_ _1974_/CLK _1845_/D vssd1 vssd1 vccd1 vccd1 _1845_/Q sky130_fd_sc_hd__dfxtp_2
X_1776_ _1946_/Q _1857_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _1776_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1431__A1 data_addr_o[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1630_ _1830_/Q vssd1 vssd1 vccd1 vccd1 _1630_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1195__B1 data_rdata_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1561_ _1561_/A vssd1 vssd1 vccd1 vccd1 _1563_/B sky130_fd_sc_hd__buf_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1492_/A _1492_/B _1492_/C vssd1 vssd1 vccd1 vccd1 _1492_/X sky130_fd_sc_hd__or3_2
Xclkbuf_4_10_0_clk_i clkbuf_3_5_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1842_/CLK sky130_fd_sc_hd__clkbuf_2
X_1828_ _1859_/CLK _1828_/D vssd1 vssd1 vccd1 vccd1 _1828_/Q sky130_fd_sc_hd__dfxtp_2
X_1759_ _1647_/A _1586_/A _1761_/S vssd1 vssd1 vccd1 vccd1 _1759_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1413__A1 data_addr_o[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0992_ data_wdata_o[7] _0989_/X _0908_/X _0991_/X vssd1 vssd1 vccd1 vccd1 _1958_/D
+ sky130_fd_sc_hd__a22o_2
X_1613_ _1613_/A vssd1 vssd1 vccd1 vccd1 _1615_/B sky130_fd_sc_hd__buf_1
X_1544_ _1302_/C _1833_/Q _1832_/Q _1543_/Y vssd1 vssd1 vccd1 vccd1 _1545_/B sky130_fd_sc_hd__o22a_2
X_1475_ _1090_/X _1468_/X _1412_/X _1471_/X vssd1 vssd1 vccd1 vccd1 _1847_/D sky130_fd_sc_hd__a22o_2
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1159__B1 data_rdata_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1191_ _1198_/A vssd1 vssd1 vccd1 vccd1 _1191_/X sky130_fd_sc_hd__buf_1
X_1260_ _1260_/A vssd1 vssd1 vccd1 vccd1 _1901_/D sky130_fd_sc_hd__inv_2
X_0975_ _0984_/A vssd1 vssd1 vccd1 vccd1 _0976_/A sky130_fd_sc_hd__buf_1
X_1527_ _1527_/A vssd1 vssd1 vccd1 vccd1 _1527_/Y sky130_fd_sc_hd__inv_2
X_1389_ _1845_/Q vssd1 vssd1 vccd1 vccd1 _1389_/X sky130_fd_sc_hd__buf_1
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1458_ _1458_/A vssd1 vssd1 vccd1 vccd1 _1458_/X sky130_fd_sc_hd__buf_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1174_ _1922_/Q _1171_/X data_rdata_i[15] _1173_/X _1168_/X vssd1 vssd1 vccd1 vccd1
+ _1922_/D sky130_fd_sc_hd__o221a_2
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1312_ _1312_/A vssd1 vssd1 vccd1 vccd1 _1313_/C sky130_fd_sc_hd__inv_2
X_1243_ _1243_/A vssd1 vssd1 vccd1 vccd1 _1244_/A sky130_fd_sc_hd__buf_1
X_0958_ _1369_/A vssd1 vssd1 vccd1 vccd1 _1008_/A sky130_fd_sc_hd__buf_1
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1930_ _1930_/CLK _1930_/D vssd1 vssd1 vccd1 vccd1 _1930_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1792_ _1304_/A _1587_/Y _1802_/S vssd1 vssd1 vccd1 vccd1 _1842_/D sky130_fd_sc_hd__mux2_1
X_1861_ _1945_/CLK _1861_/D _1453_/X vssd1 vssd1 vccd1 vccd1 _1861_/Q sky130_fd_sc_hd__dfrtp_2
X_1157_ _1930_/Q _1155_/X data_rdata_i[23] _1156_/X _1153_/X vssd1 vssd1 vccd1 vccd1
+ _1930_/D sky130_fd_sc_hd__o221a_2
XANTENNA__1042__A _1351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1226_ _1634_/B vssd1 vssd1 vccd1 vccd1 _1230_/A sky130_fd_sc_hd__inv_2
X_1088_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1089_/A sky130_fd_sc_hd__buf_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1011_ data_wdata_o[2] _1005_/X _0937_/X _1006_/X vssd1 vssd1 vccd1 vccd1 _1953_/D
+ sky130_fd_sc_hd__a22o_2
X_1913_ _1930_/CLK _1913_/D vssd1 vssd1 vccd1 vccd1 _1913_/Q sky130_fd_sc_hd__dfxtp_2
X_1775_ _1947_/Q _1858_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _1775_/X sky130_fd_sc_hd__mux2_1
X_1844_ _1876_/CLK _1844_/D vssd1 vssd1 vccd1 vccd1 _1844_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1209_ _1679_/B vssd1 vssd1 vccd1 vccd1 _1738_/S sky130_fd_sc_hd__inv_2
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1560_ _1836_/Q _1575_/A _1565_/B vssd1 vssd1 vccd1 vccd1 _1561_/A sky130_fd_sc_hd__a21bo_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ _1861_/Q vssd1 vssd1 vccd1 vccd1 _1492_/A sky130_fd_sc_hd__inv_2
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1827_ _1940_/CLK _1827_/D vssd1 vssd1 vccd1 vccd1 _1827_/Q sky130_fd_sc_hd__dfxtp_2
X_1758_ _1507_/Y _1509_/X _1758_/S vssd1 vssd1 vccd1 vccd1 _1758_/X sky130_fd_sc_hd__mux2_1
X_1689_ _1609_/A _1791_/S _1717_/X _1719_/X _1244_/A vssd1 vssd1 vccd1 vccd1 _1689_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0991_ _1006_/A vssd1 vssd1 vccd1 vccd1 _0991_/X sky130_fd_sc_hd__buf_1
X_1474_ _1412_/X _1468_/X _1408_/X _1471_/X vssd1 vssd1 vccd1 vccd1 _1848_/D sky130_fd_sc_hd__a22o_2
X_1612_ _1826_/Q _1617_/C _1611_/X vssd1 vssd1 vccd1 vccd1 _1613_/A sky130_fd_sc_hd__a21bo_2
X_1543_ _1833_/Q vssd1 vssd1 vccd1 vccd1 _1543_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1034__B uart_error vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_8_0_clk_i clkbuf_4_9_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1950_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1398__A1 data_wdata_o[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1190_ _1912_/Q _1186_/X data_rdata_i[5] _1187_/X _1184_/X vssd1 vssd1 vccd1 vccd1
+ _1912_/D sky130_fd_sc_hd__o221a_2
X_0974_ _1008_/A vssd1 vssd1 vccd1 vccd1 _0984_/A sky130_fd_sc_hd__buf_1
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1457_ _1774_/X _1240_/X _1858_/Q _1241_/X vssd1 vssd1 vccd1 vccd1 _1858_/D sky130_fd_sc_hd__o22a_2
X_1526_ _1808_/Q _1526_/B vssd1 vssd1 vccd1 vccd1 _1527_/A sky130_fd_sc_hd__or2_2
XFILLER_42_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1388_ _1388_/A vssd1 vssd1 vccd1 vccd1 _1388_/X sky130_fd_sc_hd__buf_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1311_ _1284_/Y _1288_/Y _1761_/S vssd1 vssd1 vccd1 vccd1 _1312_/A sky130_fd_sc_hd__o21ai_2
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1173_ _1194_/A vssd1 vssd1 vccd1 vccd1 _1173_/X sky130_fd_sc_hd__buf_1
X_1242_ _1212_/X _1240_/X _1904_/Q _1241_/X vssd1 vssd1 vccd1 vccd1 _1904_/D sky130_fd_sc_hd__o22a_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0957_ _1207_/A vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__buf_1
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1509_ _1507_/Y _1505_/Y _1511_/B vssd1 vssd1 vccd1 vccd1 _1509_/X sky130_fd_sc_hd__o21a_2
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_5_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1860_ _1945_/CLK _1860_/D _1455_/X vssd1 vssd1 vccd1 vccd1 _1860_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1791_ _1229_/A _1589_/Y _1791_/S vssd1 vssd1 vccd1 vccd1 _1821_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1156_ _1164_/A vssd1 vssd1 vccd1 vccd1 _1156_/X sky130_fd_sc_hd__buf_1
X_1087_ _1087_/A vssd1 vssd1 vccd1 vccd1 _1947_/D sky130_fd_sc_hd__buf_1
X_1225_ _1831_/Q _1224_/X _1831_/Q _1224_/X vssd1 vssd1 vccd1 vccd1 _1634_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1010_ _1010_/A vssd1 vssd1 vccd1 vccd1 _1010_/X sky130_fd_sc_hd__buf_1
X_1912_ _1930_/CLK _1912_/D vssd1 vssd1 vccd1 vccd1 _1912_/Q sky130_fd_sc_hd__dfxtp_2
X_1843_ _1876_/CLK _1843_/D vssd1 vssd1 vccd1 vccd1 _1843_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1774_ _1948_/Q _1904_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _1774_/X sky130_fd_sc_hd__mux2_1
X_1208_ _1208_/A _1811_/Q vssd1 vssd1 vccd1 vccd1 _1679_/B sky130_fd_sc_hd__nand2_2
X_1139_ _1163_/A vssd1 vssd1 vccd1 vccd1 _1139_/X sky130_fd_sc_hd__buf_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1490_ _1490_/A vssd1 vssd1 vccd1 vccd1 _1490_/X sky130_fd_sc_hd__buf_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1826_ _1940_/CLK _1826_/D vssd1 vssd1 vccd1 vccd1 _1826_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1757_ _1510_/Y _1513_/Y _1758_/S vssd1 vssd1 vccd1 vccd1 _1757_/X sky130_fd_sc_hd__mux2_1
X_1688_ _1723_/X _1780_/S _1791_/S _1687_/X vssd1 vssd1 vccd1 vccd1 _1688_/X sky130_fd_sc_hd__a22o_2
XANTENNA__1048__A data_req_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_clk_i clkbuf_4_5_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1943_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1611_ _1826_/Q _1617_/C vssd1 vssd1 vccd1 vccd1 _1611_/X sky130_fd_sc_hd__or2_2
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0990_ _1005_/A vssd1 vssd1 vccd1 vccd1 _1006_/A sky130_fd_sc_hd__inv_2
X_1473_ _1408_/X _1468_/X _1076_/X _1471_/X vssd1 vssd1 vccd1 vccd1 _1849_/D sky130_fd_sc_hd__a22o_2
X_1542_ _1657_/B vssd1 vssd1 vccd1 vccd1 _1802_/S sky130_fd_sc_hd__inv_2
XFILLER_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1809_ _1859_/CLK _1809_/D vssd1 vssd1 vccd1 vccd1 _1809_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0973_ data_wdata_o[11] _0971_/X _0931_/X _0972_/X vssd1 vssd1 vccd1 vccd1 _1962_/D
+ sky130_fd_sc_hd__a22o_2
X_1387_ _1399_/A vssd1 vssd1 vccd1 vccd1 _1388_/A sky130_fd_sc_hd__buf_1
X_1525_ _1807_/Q _1524_/B _1526_/B vssd1 vssd1 vccd1 vccd1 _1525_/X sky130_fd_sc_hd__a21bo_2
X_1456_ _1456_/A hold1/X vssd1 vssd1 vccd1 vccd1 _1859_/D sky130_fd_sc_hd__nor2_2
XFILLER_19_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1241_ _1458_/A vssd1 vssd1 vccd1 vccd1 _1241_/X sky130_fd_sc_hd__buf_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1310_ _1749_/S vssd1 vssd1 vccd1 vccd1 _1761_/S sky130_fd_sc_hd__inv_2
X_1172_ _1172_/A vssd1 vssd1 vccd1 vccd1 _1194_/A sky130_fd_sc_hd__buf_1
X_0956_ data_wdata_o[15] _0953_/X _0908_/X _0955_/X vssd1 vssd1 vccd1 vccd1 _1966_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1508_ _1814_/Q _1508_/B vssd1 vssd1 vccd1 vccd1 _1511_/B sky130_fd_sc_hd__or2_2
X_1439_ _1443_/A vssd1 vssd1 vccd1 vccd1 _1440_/A sky130_fd_sc_hd__buf_1
XFILLER_11_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1790_ _1594_/B _1595_/X _1791_/S vssd1 vssd1 vccd1 vccd1 _1822_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1224_ _1829_/Q _1830_/Q _1626_/B vssd1 vssd1 vccd1 vccd1 _1224_/X sky130_fd_sc_hd__or3_2
X_1155_ _1163_/A vssd1 vssd1 vccd1 vccd1 _1155_/X sky130_fd_sc_hd__buf_1
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1086_ _1708_/X _1947_/Q _1096_/A vssd1 vssd1 vccd1 vccd1 _1087_/A sky130_fd_sc_hd__mux2_2
X_0939_ _0948_/A vssd1 vssd1 vccd1 vccd1 _0940_/A sky130_fd_sc_hd__buf_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1773_ _1772_/X _1934_/Q _1860_/Q vssd1 vssd1 vccd1 vccd1 _1773_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1911_ _1930_/CLK _1911_/D vssd1 vssd1 vccd1 vccd1 _1911_/Q sky130_fd_sc_hd__dfxtp_2
X_1842_ _1842_/CLK _1842_/D vssd1 vssd1 vccd1 vccd1 _1842_/Q sky130_fd_sc_hd__dfxtp_2
X_1207_ _1207_/A _1810_/Q vssd1 vssd1 vccd1 vccd1 _1213_/A sky130_fd_sc_hd__nand2_2
X_1138_ _1170_/A vssd1 vssd1 vccd1 vccd1 _1163_/A sky130_fd_sc_hd__buf_1
XFILLER_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1425__A1 data_addr_o[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1069_ _1498_/A _1050_/X _1066_/X _1067_/Y _1068_/X vssd1 vssd1 vccd1 vccd1 _1495_/A
+ sky130_fd_sc_hd__a32o_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1189__B1 data_rdata_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_0_0_clk_i clkbuf_4_1_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1859_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1756_ _1514_/Y _1516_/X _1758_/S vssd1 vssd1 vccd1 vccd1 _1756_/X sky130_fd_sc_hd__mux2_1
X_1825_ _1859_/CLK _1825_/D vssd1 vssd1 vccd1 vccd1 _1825_/Q sky130_fd_sc_hd__dfxtp_2
X_1687_ _1687_/A _1718_/X vssd1 vssd1 vccd1 vccd1 _1687_/X sky130_fd_sc_hd__or2_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1610_ _1610_/A vssd1 vssd1 vccd1 vccd1 _1610_/X sky130_fd_sc_hd__buf_1
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1472_ _1076_/X _1468_/X _1557_/A _1471_/X vssd1 vssd1 vccd1 vccd1 _1850_/D sky130_fd_sc_hd__a22o_2
XFILLER_5_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1541_ _1747_/S _1664_/B _1642_/A vssd1 vssd1 vccd1 vccd1 _1657_/B sky130_fd_sc_hd__or3_2
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1808_ _1859_/CLK _1808_/D vssd1 vssd1 vccd1 vccd1 _1808_/Q sky130_fd_sc_hd__dfxtp_2
X_1739_ _1756_/X _1674_/X _1761_/S vssd1 vssd1 vccd1 vccd1 _1739_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0972_ _0972_/A vssd1 vssd1 vccd1 vccd1 _0972_/X sky130_fd_sc_hd__buf_1
X_1524_ _1807_/Q _1524_/B vssd1 vssd1 vccd1 vccd1 _1526_/B sky130_fd_sc_hd__or2_2
X_1386_ _1422_/A vssd1 vssd1 vccd1 vccd1 _1399_/A sky130_fd_sc_hd__buf_1
X_1455_ _1455_/A vssd1 vssd1 vccd1 vccd1 _1455_/X sky130_fd_sc_hd__buf_1
XFILLER_35_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1171_ _1193_/A vssd1 vssd1 vccd1 vccd1 _1171_/X sky130_fd_sc_hd__buf_1
X_1240_ _1240_/A vssd1 vssd1 vccd1 vccd1 _1240_/X sky130_fd_sc_hd__buf_1
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0955_ _0972_/A vssd1 vssd1 vccd1 vccd1 _0955_/X sky130_fd_sc_hd__buf_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1507_ _1814_/Q vssd1 vssd1 vccd1 vccd1 _1507_/Y sky130_fd_sc_hd__inv_2
X_1369_ _1369_/A vssd1 vssd1 vccd1 vccd1 _1422_/A sky130_fd_sc_hd__buf_1
X_1438_ _1438_/A vssd1 vssd1 vccd1 vccd1 _1438_/X sky130_fd_sc_hd__buf_1
XFILLER_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1154_ _1931_/Q _1148_/X data_rdata_i[24] _1149_/X _1153_/X vssd1 vssd1 vccd1 vccd1
+ _1931_/D sky130_fd_sc_hd__o221a_2
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1223_ _1606_/B _1229_/D vssd1 vssd1 vccd1 vccd1 _1626_/B sky130_fd_sc_hd__or2_2
X_1085_ _1085_/A vssd1 vssd1 vccd1 vccd1 _1085_/X sky130_fd_sc_hd__buf_1
XFILLER_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0938_ data_wdata_o[18] _0930_/X _0937_/X _0932_/X vssd1 vssd1 vccd1 vccd1 _1969_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1910_ _1949_/CLK _1910_/D vssd1 vssd1 vccd1 vccd1 _1910_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1772_ _1771_/X _1926_/Q _1864_/Q vssd1 vssd1 vccd1 vccd1 _1772_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1841_ _1842_/CLK _1841_/D vssd1 vssd1 vccd1 vccd1 _1841_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1137_ _1172_/A vssd1 vssd1 vccd1 vccd1 _1170_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_clk_i_A clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1206_ data_req_o _1205_/A _1803_/X _1205_/Y _1198_/X vssd1 vssd1 vccd1 vccd1 _1905_/D
+ sky130_fd_sc_hd__o221a_2
X_1068_ _1066_/X _1865_/Q _1068_/C vssd1 vssd1 vccd1 vccd1 _1068_/X sky130_fd_sc_hd__and3b_2
XANTENNA_clkbuf_3_2_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0927__A1 data_wdata_o[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1755_ _1813_/Q _1506_/X _1758_/S vssd1 vssd1 vccd1 vccd1 _1755_/X sky130_fd_sc_hd__mux2_1
X_1824_ _1859_/CLK _1824_/D vssd1 vssd1 vccd1 vccd1 _1824_/Q sky130_fd_sc_hd__dfxtp_2
X_1686_ _1686_/A vssd1 vssd1 vccd1 vccd1 _1686_/X sky130_fd_sc_hd__buf_1
XFILLER_0_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1540_ _1586_/A _1832_/Q vssd1 vssd1 vccd1 vccd1 _1540_/Y sky130_fd_sc_hd__nor2_2
X_1471_ _1477_/A vssd1 vssd1 vccd1 vccd1 _1471_/X sky130_fd_sc_hd__buf_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1807_ _1903_/CLK _1807_/D vssd1 vssd1 vccd1 vccd1 _1807_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1669_ _1676_/A _1757_/X vssd1 vssd1 vccd1 vccd1 _1670_/A sky130_fd_sc_hd__or2_2
X_1738_ _1693_/X _1714_/X _1738_/S vssd1 vssd1 vccd1 vccd1 _1809_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0971_ _0971_/A vssd1 vssd1 vccd1 vccd1 _0971_/X sky130_fd_sc_hd__buf_1
X_1454_ _1694_/A vssd1 vssd1 vccd1 vccd1 _1455_/A sky130_fd_sc_hd__buf_1
X_1523_ _1806_/Q _1522_/B _1524_/B vssd1 vssd1 vccd1 vccd1 _1523_/X sky130_fd_sc_hd__a21bo_2
X_1385_ data_wdata_o[27] _1382_/X _1383_/X _1384_/X vssd1 vssd1 vccd1 vccd1 _1882_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1170_ _1170_/A vssd1 vssd1 vccd1 vccd1 _1193_/A sky130_fd_sc_hd__buf_1
XFILLER_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0954_ _0971_/A vssd1 vssd1 vccd1 vccd1 _0972_/A sky130_fd_sc_hd__inv_2
X_1506_ _1812_/Q _1813_/Q _1505_/Y vssd1 vssd1 vccd1 vccd1 _1506_/X sky130_fd_sc_hd__a21o_2
X_1437_ _1443_/A vssd1 vssd1 vccd1 vccd1 _1438_/A sky130_fd_sc_hd__buf_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1368_ data_wdata_o[31] _1365_/X _0908_/X _1367_/X vssd1 vssd1 vccd1 vccd1 _1886_/D
+ sky130_fd_sc_hd__a22o_2
X_1299_ _1842_/Q _1298_/Y _1842_/Q _1298_/Y vssd1 vssd1 vccd1 vccd1 _1587_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1153_ _1694_/A vssd1 vssd1 vccd1 vccd1 _1153_/X sky130_fd_sc_hd__buf_1
XFILLER_37_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1084_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1085_/A sky130_fd_sc_hd__buf_1
X_1222_ _1826_/Q _1827_/Q _1825_/Q _1828_/Q vssd1 vssd1 vccd1 vccd1 _1229_/D sky130_fd_sc_hd__or4_2
XFILLER_20_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0937_ _1845_/Q vssd1 vssd1 vccd1 vccd1 _0937_/X sky130_fd_sc_hd__buf_1
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1840_ _1842_/CLK _1840_/D vssd1 vssd1 vccd1 vccd1 _1840_/Q sky130_fd_sc_hd__dfxtp_2
X_1771_ _1910_/Q _1918_/Q _1862_/Q vssd1 vssd1 vccd1 vccd1 _1771_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1205_ _1205_/A vssd1 vssd1 vccd1 vccd1 _1205_/Y sky130_fd_sc_hd__inv_2
X_1136_ _1136_/A _1203_/B vssd1 vssd1 vccd1 vccd1 _1172_/A sky130_fd_sc_hd__or2_2
X_1067_ _1067_/A _1532_/B vssd1 vssd1 vccd1 vccd1 _1067_/Y sky130_fd_sc_hd__nor2_2
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1969_ _1974_/CLK _1969_/D _0936_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[18] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_6_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1823_ _1859_/CLK _1823_/D vssd1 vssd1 vccd1 vccd1 _1823_/Q sky130_fd_sc_hd__dfxtp_2
X_1754_ _1517_/Y _1518_/X _1758_/S vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__mux2_1
X_1685_ _1682_/X _1711_/X vssd1 vssd1 vccd1 vccd1 _1686_/A sky130_fd_sc_hd__and2b_2
X_1119_ _1119_/A vssd1 vssd1 vccd1 vccd1 _1203_/B sky130_fd_sc_hd__inv_2
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1470_ _1562_/A vssd1 vssd1 vccd1 vccd1 _1557_/A sky130_fd_sc_hd__buf_1
X_1806_ _1859_/CLK _1806_/D vssd1 vssd1 vccd1 vccd1 _1806_/Q sky130_fd_sc_hd__dfxtp_2
X_1737_ _1691_/X _1713_/X _1738_/S vssd1 vssd1 vccd1 vccd1 _1808_/D sky130_fd_sc_hd__mux2_1
X_1668_ _1758_/X _1658_/B _1761_/X _1650_/A _1667_/Y vssd1 vssd1 vccd1 vccd1 _1668_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1599_ _1614_/A vssd1 vssd1 vccd1 vccd1 _1609_/A sky130_fd_sc_hd__buf_1
XFILLER_5_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0970_ _0970_/A vssd1 vssd1 vccd1 vccd1 _0970_/X sky130_fd_sc_hd__buf_1
X_1522_ _1806_/Q _1522_/B vssd1 vssd1 vccd1 vccd1 _1524_/B sky130_fd_sc_hd__or2_2
X_1453_ _1453_/A vssd1 vssd1 vccd1 vccd1 _1453_/X sky130_fd_sc_hd__buf_1
X_1384_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1384_/X sky130_fd_sc_hd__buf_1
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0953_ _0971_/A vssd1 vssd1 vccd1 vccd1 _0953_/X sky130_fd_sc_hd__buf_1
X_1367_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1367_/X sky130_fd_sc_hd__buf_1
X_1505_ _1508_/B vssd1 vssd1 vccd1 vccd1 _1505_/Y sky130_fd_sc_hd__inv_2
X_1436_ _1445_/A vssd1 vssd1 vccd1 vccd1 _1443_/A sky130_fd_sc_hd__buf_1
XANTENNA__1152__B1 data_rdata_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1298_ _1840_/Q _1841_/Q _1575_/B _1554_/A vssd1 vssd1 vccd1 vccd1 _1298_/Y sky130_fd_sc_hd__nor4_2
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1143__B1 data_rdata_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1221_ _1823_/Q _1824_/Q _1596_/B vssd1 vssd1 vccd1 vccd1 _1606_/B sky130_fd_sc_hd__or3_2
X_1152_ _1932_/Q _1148_/X data_rdata_i[25] _1149_/X _1146_/X vssd1 vssd1 vccd1 vccd1
+ _1932_/D sky130_fd_sc_hd__o221a_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1083_ _1083_/A vssd1 vssd1 vccd1 vccd1 _1948_/D sky130_fd_sc_hd__buf_1
X_0936_ _0936_/A vssd1 vssd1 vccd1 vccd1 _0936_/X sky130_fd_sc_hd__buf_1
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1373__B1 _0916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1419_ _1419_/A vssd1 vssd1 vccd1 vccd1 _1419_/X sky130_fd_sc_hd__buf_1
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1428__A1 data_addr_o[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1770_ _1769_/X _1935_/Q _1860_/Q vssd1 vssd1 vccd1 vccd1 _1770_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1204_ _1202_/Y _1128_/A _1133_/Y _1203_/X vssd1 vssd1 vccd1 vccd1 _1205_/A sky130_fd_sc_hd__a211o_2
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1135_ _1456_/A _1135_/B vssd1 vssd1 vccd1 vccd1 _1939_/D sky130_fd_sc_hd__nor2_2
X_1066_ _1066_/A uart_error vssd1 vssd1 vccd1 vccd1 _1066_/X sky130_fd_sc_hd__or2_2
X_1968_ _1974_/CLK _1968_/D _0940_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[17] sky130_fd_sc_hd__dfrtp_2
X_0919_ _1445_/A vssd1 vssd1 vccd1 vccd1 _0928_/A sky130_fd_sc_hd__buf_1
X_1899_ _1943_/CLK _1899_/D vssd1 vssd1 vccd1 vccd1 _1899_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1822_ _1859_/CLK _1822_/D vssd1 vssd1 vccd1 vccd1 _1822_/Q sky130_fd_sc_hd__dfxtp_2
X_1753_ _1647_/B rx_i _1761_/S vssd1 vssd1 vccd1 vccd1 _1753_/X sky130_fd_sc_hd__mux2_1
X_1684_ _1684_/A vssd1 vssd1 vccd1 vccd1 _1684_/X sky130_fd_sc_hd__buf_1
X_1118_ _1897_/Q _1861_/Q _1950_/Q vssd1 vssd1 vccd1 vccd1 _1119_/A sky130_fd_sc_hd__o21ai_2
X_1049_ _1492_/C vssd1 vssd1 vccd1 vccd1 _1061_/B sky130_fd_sc_hd__inv_2
XANTENNA__1552__A _1557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1805_ _1859_/CLK _1805_/D vssd1 vssd1 vccd1 vccd1 _1805_/Q sky130_fd_sc_hd__dfxtp_2
X_1736_ _1689_/X _1717_/X _1738_/S vssd1 vssd1 vccd1 vccd1 _1807_/D sky130_fd_sc_hd__mux2_1
X_1598_ _1598_/A vssd1 vssd1 vccd1 vccd1 _1600_/B sky130_fd_sc_hd__buf_1
X_1667_ _1666_/B _1761_/S _1284_/Y vssd1 vssd1 vccd1 vccd1 _1667_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1383_ _1846_/Q vssd1 vssd1 vccd1 vccd1 _1383_/X sky130_fd_sc_hd__buf_1
X_1452_ _1452_/A vssd1 vssd1 vccd1 vccd1 _1453_/A sky130_fd_sc_hd__buf_1
X_1521_ _1804_/Q _1805_/Q _1522_/B vssd1 vssd1 vccd1 vccd1 _1521_/X sky130_fd_sc_hd__a21bo_2
XFILLER_35_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1719_ _1465_/B _1717_/X _1740_/S vssd1 vssd1 vccd1 vccd1 _1719_/X sky130_fd_sc_hd__mux2_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0952_ _0987_/B _1058_/C _0952_/C vssd1 vssd1 vccd1 vccd1 _0971_/A sky130_fd_sc_hd__or3_2
XFILLER_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1504_ _1812_/Q _1813_/Q vssd1 vssd1 vccd1 vccd1 _1508_/B sky130_fd_sc_hd__or2_2
X_1366_ _1382_/A vssd1 vssd1 vccd1 vccd1 _1384_/A sky130_fd_sc_hd__inv_2
X_1435_ _1435_/A vssd1 vssd1 vccd1 vccd1 _1435_/X sky130_fd_sc_hd__buf_1
X_1297_ _1835_/Q _1297_/B vssd1 vssd1 vccd1 vccd1 _1554_/A sky130_fd_sc_hd__or2_2
X_1151_ _1933_/Q _1148_/X data_rdata_i[26] _1149_/X _1146_/X vssd1 vssd1 vccd1 vccd1
+ _1933_/D sky130_fd_sc_hd__o221a_2
X_1220_ _1821_/Q _1822_/Q vssd1 vssd1 vccd1 vccd1 _1596_/B sky130_fd_sc_hd__or2_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1082_ _1709_/X _1948_/Q _1096_/A vssd1 vssd1 vccd1 vccd1 _1083_/A sky130_fd_sc_hd__mux2_2
X_0935_ _0948_/A vssd1 vssd1 vccd1 vccd1 _0936_/A sky130_fd_sc_hd__buf_1
XFILLER_9_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1418_ _1418_/A vssd1 vssd1 vccd1 vccd1 _1418_/X sky130_fd_sc_hd__buf_1
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1349_ _1349_/A vssd1 vssd1 vccd1 vccd1 _1349_/X sky130_fd_sc_hd__buf_1
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1203_ data_gnt_i _1203_/B vssd1 vssd1 vccd1 vccd1 _1203_/X sky130_fd_sc_hd__and2_2
X_1134_ _1483_/A _1115_/B _1128_/A _1132_/Y _1133_/Y vssd1 vssd1 vccd1 vccd1 _1135_/B
+ sky130_fd_sc_hd__o32a_2
X_1065_ _1850_/Q _1065_/B _1848_/Q vssd1 vssd1 vccd1 vccd1 _1533_/B sky130_fd_sc_hd__or3b_2
X_1967_ _1974_/CLK _1967_/D _0945_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[16] sky130_fd_sc_hd__dfrtp_2
X_0918_ _1207_/A vssd1 vssd1 vccd1 vccd1 _1445_/A sky130_fd_sc_hd__buf_1
X_1898_ _1971_/CLK _1898_/D _1267_/X vssd1 vssd1 vccd1 vccd1 _1898_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1752_ _1751_/X _1938_/Q _1860_/Q vssd1 vssd1 vccd1 vccd1 _1752_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1821_ _1859_/CLK _1821_/D vssd1 vssd1 vccd1 vccd1 _1821_/Q sky130_fd_sc_hd__dfxtp_2
X_1683_ _1682_/X _1683_/B vssd1 vssd1 vccd1 vccd1 _1684_/A sky130_fd_sc_hd__and2b_2
X_1117_ _1117_/A _1117_/B _1133_/A vssd1 vssd1 vccd1 vccd1 _1136_/A sky130_fd_sc_hd__or3b_2
X_1048_ data_req_o _1903_/Q _1066_/A _1048_/D vssd1 vssd1 vccd1 vccd1 _1492_/C sky130_fd_sc_hd__or4_2
XFILLER_21_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0912__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1666_ _1666_/A _1666_/B vssd1 vssd1 vccd1 vccd1 _1666_/Y sky130_fd_sc_hd__nor2_2
X_1804_ _1859_/CLK _1804_/D vssd1 vssd1 vccd1 vccd1 _1804_/Q sky130_fd_sc_hd__dfxtp_2
X_1735_ _1688_/X _1718_/X _1738_/S vssd1 vssd1 vccd1 vccd1 _1806_/D sky130_fd_sc_hd__mux2_1
X_1597_ _1823_/Q _1596_/B _1596_/X vssd1 vssd1 vccd1 vccd1 _1598_/A sky130_fd_sc_hd__a21bo_2
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1520_ _1804_/Q _1805_/Q vssd1 vssd1 vccd1 vccd1 _1522_/B sky130_fd_sc_hd__or2_2
X_1382_ _1382_/A vssd1 vssd1 vccd1 vccd1 _1382_/X sky130_fd_sc_hd__buf_1
X_1451_ _1451_/A vssd1 vssd1 vccd1 vccd1 _1451_/X sky130_fd_sc_hd__buf_1
XFILLER_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1718_ _1806_/Q _1523_/X _1718_/S vssd1 vssd1 vccd1 vccd1 _1718_/X sky130_fd_sc_hd__mux2_1
X_1649_ _1704_/X _1658_/A _1705_/X _1650_/A _1648_/X vssd1 vssd1 vccd1 vccd1 _1649_/Y
+ sky130_fd_sc_hd__o221ai_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0951_ _1860_/Q _1864_/Q vssd1 vssd1 vccd1 vccd1 _1058_/C sky130_fd_sc_hd__or2_2
X_1503_ _1503_/A vssd1 vssd1 vccd1 vccd1 _1747_/S sky130_fd_sc_hd__buf_1
X_1365_ _1382_/A vssd1 vssd1 vccd1 vccd1 _1365_/X sky130_fd_sc_hd__buf_1
X_1434_ _1434_/A vssd1 vssd1 vccd1 vccd1 _1435_/A sky130_fd_sc_hd__buf_1
X_1296_ _1834_/Q _1296_/B vssd1 vssd1 vccd1 vccd1 _1297_/B sky130_fd_sc_hd__or2_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1288__A rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0920__A _0928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1150_ _1934_/Q _1148_/X data_rdata_i[27] _1149_/X _1146_/X vssd1 vssd1 vccd1 vccd1
+ _1934_/D sky130_fd_sc_hd__o221a_2
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1081_ _1081_/A vssd1 vssd1 vccd1 vccd1 _1081_/X sky130_fd_sc_hd__buf_1
X_0934_ _1198_/A vssd1 vssd1 vccd1 vccd1 _0948_/A sky130_fd_sc_hd__buf_1
XANTENNA__1198__A _1198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1417_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1418_/A sky130_fd_sc_hd__buf_1
X_1279_ _1279_/A vssd1 vssd1 vccd1 vccd1 _1653_/C sky130_fd_sc_hd__buf_1
X_1348_ _1348_/A vssd1 vssd1 vccd1 vccd1 _1349_/A sky130_fd_sc_hd__inv_2
XANTENNA__1116__A2 data_gnt_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0915__A _1198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1202_ _1897_/Q vssd1 vssd1 vccd1 vccd1 _1202_/Y sky130_fd_sc_hd__inv_2
X_1133_ _1133_/A _1203_/B vssd1 vssd1 vccd1 vccd1 _1133_/Y sky130_fd_sc_hd__nor2_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1064_ _1866_/Q _1061_/Y _1533_/A _1636_/A vssd1 vssd1 vccd1 vccd1 _1064_/Y sky130_fd_sc_hd__a22oi_2
X_1966_ _1974_/CLK _1966_/D _0949_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[15] sky130_fd_sc_hd__dfrtp_2
X_0917_ data_wdata_o[22] _0907_/X _0916_/X _0910_/X vssd1 vssd1 vccd1 vccd1 _1973_/D
+ sky130_fd_sc_hd__a22o_2
X_1897_ _1940_/CLK _1897_/D vssd1 vssd1 vccd1 vccd1 _1897_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1820_ _1950_/CLK _1820_/D vssd1 vssd1 vccd1 vccd1 _1820_/Q sky130_fd_sc_hd__dfxtp_2
X_1751_ _1750_/X _1930_/Q _1864_/Q vssd1 vssd1 vccd1 vccd1 _1751_/X sky130_fd_sc_hd__mux2_1
X_1682_ _1246_/A _1870_/D _1217_/A vssd1 vssd1 vccd1 vccd1 _1682_/X sky130_fd_sc_hd__o21a_2
X_1047_ _1891_/Q data_rvalid_i data_gnt_i vssd1 vssd1 vccd1 vccd1 _1048_/D sky130_fd_sc_hd__or3_2
X_1116_ _1340_/B data_gnt_i _1115_/Y vssd1 vssd1 vccd1 vccd1 _1133_/A sky130_fd_sc_hd__a21oi_2
X_1949_ _1949_/CLK _1949_/D _1044_/X vssd1 vssd1 vccd1 vccd1 _1949_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1803_ _1115_/Y _1202_/Y _1803_/S vssd1 vssd1 vccd1 vccd1 _1803_/X sky130_fd_sc_hd__mux2_1
X_1596_ _1823_/Q _1596_/B vssd1 vssd1 vccd1 vccd1 _1596_/X sky130_fd_sc_hd__or2_2
X_1665_ _1557_/A _1657_/B _1749_/X _1650_/A _1664_/X vssd1 vssd1 vccd1 vccd1 _1665_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1734_ _1686_/X _1711_/X _1738_/S vssd1 vssd1 vccd1 vccd1 _1805_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1182__B1 data_rdata_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0996__B1 _0916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1450_ _1452_/A vssd1 vssd1 vccd1 vccd1 _1451_/A sky130_fd_sc_hd__buf_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1381_ _1381_/A vssd1 vssd1 vccd1 vccd1 _1381_/X sky130_fd_sc_hd__buf_1
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_13_0_clk_i clkbuf_3_6_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1938_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _1840_/Q _1579_/B vssd1 vssd1 vccd1 vccd1 _1579_/X sky130_fd_sc_hd__or2_2
X_1648_ _1753_/X _1647_/X _1562_/A _1657_/B vssd1 vssd1 vccd1 vccd1 _1648_/X sky130_fd_sc_hd__o22a_2
X_1717_ _1807_/Q _1525_/X _1718_/S vssd1 vssd1 vccd1 vccd1 _1717_/X sky130_fd_sc_hd__mux2_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0950_ _1862_/Q vssd1 vssd1 vccd1 vccd1 _0987_/B sky130_fd_sc_hd__inv_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1433_ _1519_/A vssd1 vssd1 vccd1 vccd1 _1870_/D sky130_fd_sc_hd__inv_2
X_1502_ _1500_/Y _1486_/X _1492_/A _1501_/X vssd1 vssd1 vccd1 vccd1 _1861_/D sky130_fd_sc_hd__o22ai_2
X_1364_ _1364_/A _1535_/B vssd1 vssd1 vccd1 vccd1 _1382_/A sky130_fd_sc_hd__or2_2
X_1295_ _1832_/Q _1833_/Q vssd1 vssd1 vccd1 vccd1 _1296_/B sky130_fd_sc_hd__or2_2
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1080_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1081_/A sky130_fd_sc_hd__buf_1
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0933_ data_wdata_o[19] _0930_/X _0931_/X _0932_/X vssd1 vssd1 vccd1 vccd1 _1970_/D
+ sky130_fd_sc_hd__a22o_2
X_1416_ data_addr_o[4] _1401_/X _1090_/X _1403_/X vssd1 vssd1 vccd1 vccd1 _1875_/D
+ sky130_fd_sc_hd__a22o_2
X_1347_ _1348_/A vssd1 vssd1 vccd1 vccd1 _1347_/X sky130_fd_sc_hd__buf_1
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1278_ _1432_/A _1671_/A vssd1 vssd1 vccd1 vccd1 _1279_/A sky130_fd_sc_hd__or2_2
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1201_ data_we_o _1803_/X _1200_/Y _1803_/S _1198_/X vssd1 vssd1 vccd1 vccd1 _1906_/D
+ sky130_fd_sc_hd__o221a_2
X_1132_ _1483_/A vssd1 vssd1 vccd1 vccd1 _1132_/Y sky130_fd_sc_hd__inv_2
X_1063_ _1063_/A vssd1 vssd1 vccd1 vccd1 _1636_/A sky130_fd_sc_hd__buf_1
X_0916_ _1849_/Q vssd1 vssd1 vccd1 vccd1 _0916_/X sky130_fd_sc_hd__buf_1
X_1965_ _1965_/CLK _1965_/D _0961_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[14] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1896_ _1950_/CLK _1896_/D vssd1 vssd1 vccd1 vccd1 _1896_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1750_ _1914_/Q _1922_/Q _1862_/Q vssd1 vssd1 vccd1 vccd1 _1750_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1681_ _1679_/A _1738_/S _1740_/S _1740_/X _1780_/S vssd1 vssd1 vccd1 vccd1 _1681_/X
+ sky130_fd_sc_hd__a32o_2
X_1115_ _1939_/Q _1115_/B vssd1 vssd1 vccd1 vccd1 _1115_/Y sky130_fd_sc_hd__nor2_2
X_1046_ _1046_/A vssd1 vssd1 vccd1 vccd1 _1671_/A sky130_fd_sc_hd__buf_1
X_1948_ _1949_/CLK _1948_/D _1081_/X vssd1 vssd1 vccd1 vccd1 _1948_/Q sky130_fd_sc_hd__dfrtp_2
X_1879_ _1965_/CLK _1879_/D _1396_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[24] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1802_ _1302_/C _1540_/Y _1802_/S vssd1 vssd1 vccd1 vccd1 _1832_/D sky130_fd_sc_hd__mux2_1
X_1733_ _1684_/X _1683_/B _1738_/S vssd1 vssd1 vccd1 vccd1 _1804_/D sky130_fd_sc_hd__mux2_1
X_1664_ _1747_/S _1664_/B _1664_/C vssd1 vssd1 vccd1 vccd1 _1664_/X sky130_fd_sc_hd__or3_2
X_1595_ _1595_/A vssd1 vssd1 vccd1 vccd1 _1595_/X sky130_fd_sc_hd__buf_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1029_ _1820_/Q vssd1 vssd1 vccd1 vccd1 _1647_/C sky130_fd_sc_hd__buf_1
XFILLER_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1380_ _1380_/A vssd1 vssd1 vccd1 vccd1 _1381_/A sky130_fd_sc_hd__buf_1
XFILLER_4_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1716_ _1677_/X _1754_/X _1749_/S vssd1 vssd1 vccd1 vccd1 _1716_/X sky130_fd_sc_hd__mux2_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1647_ _1647_/A _1647_/B _1647_/C vssd1 vssd1 vccd1 vccd1 _1647_/X sky130_fd_sc_hd__or3_2
X_1578_ _1578_/A vssd1 vssd1 vccd1 vccd1 _1578_/X sky130_fd_sc_hd__buf_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1394__A1 data_wdata_o[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0934__A _1198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1363_ _1860_/Q vssd1 vssd1 vccd1 vccd1 _1364_/A sky130_fd_sc_hd__inv_2
X_1432_ _1432_/A _1432_/B vssd1 vssd1 vccd1 vccd1 _1519_/A sky130_fd_sc_hd__or2_2
X_1501_ _1330_/X _1483_/B _1535_/A _0904_/A _1335_/X vssd1 vssd1 vccd1 vccd1 _1501_/X
+ sky130_fd_sc_hd__o2111a_2
X_1294_ _1836_/Q _1837_/Q _1838_/Q _1839_/Q vssd1 vssd1 vccd1 vccd1 _1575_/B sky130_fd_sc_hd__or4_2
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0932_ _0932_/A vssd1 vssd1 vccd1 vccd1 _0932_/X sky130_fd_sc_hd__buf_1
X_1415_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1415_/X sky130_fd_sc_hd__buf_1
XFILLER_3_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1346_ _1533_/A _1533_/B _1868_/Q vssd1 vssd1 vccd1 vccd1 _1348_/A sky130_fd_sc_hd__or3b_2
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1277_ _1647_/B vssd1 vssd1 vccd1 vccd1 _1503_/A sky130_fd_sc_hd__inv_2
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1200_ _1803_/X vssd1 vssd1 vccd1 vccd1 _1200_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1760__A1 rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1131_ _1340_/B vssd1 vssd1 vccd1 vccd1 _1483_/A sky130_fd_sc_hd__buf_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1062_ _1062_/A vssd1 vssd1 vccd1 vccd1 _1533_/A sky130_fd_sc_hd__buf_1
X_0915_ _1198_/A vssd1 vssd1 vccd1 vccd1 _0915_/X sky130_fd_sc_hd__buf_1
X_1964_ _1965_/CLK _1964_/D _0964_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[13] sky130_fd_sc_hd__dfrtp_2
X_1895_ _1972_/CLK _1895_/D vssd1 vssd1 vccd1 vccd1 _1895_/Q sky130_fd_sc_hd__dfxtp_2
X_1329_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1419_/A sky130_fd_sc_hd__buf_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1680_ _1710_/X _1780_/S _1634_/A _1791_/S vssd1 vssd1 vccd1 vccd1 _1680_/X sky130_fd_sc_hd__a22o_2
X_1114_ _1892_/Q vssd1 vssd1 vccd1 vccd1 _1115_/B sky130_fd_sc_hd__inv_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1045_ _1818_/Q vssd1 vssd1 vccd1 vccd1 _1275_/B sky130_fd_sc_hd__inv_2
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1878_ _1938_/CLK _1878_/D _1400_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[7] sky130_fd_sc_hd__dfrtp_2
X_1947_ _1949_/CLK _1947_/D _1085_/X vssd1 vssd1 vccd1 vccd1 _1947_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1801_ _1548_/B _1549_/X _1802_/S vssd1 vssd1 vccd1 vccd1 _1833_/D sky130_fd_sc_hd__mux2_1
X_1663_ _1663_/A vssd1 vssd1 vccd1 vccd1 _1663_/X sky130_fd_sc_hd__buf_1
X_1732_ _1681_/X _1738_/S _1732_/S vssd1 vssd1 vccd1 vccd1 _1811_/D sky130_fd_sc_hd__mux2_1
X_1594_ _1687_/A _1594_/B vssd1 vssd1 vccd1 vccd1 _1595_/A sky130_fd_sc_hd__or2_2
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1028_ _1865_/Q vssd1 vssd1 vccd1 vccd1 _1034_/A sky130_fd_sc_hd__inv_2
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1646_ _1646_/A vssd1 vssd1 vccd1 vccd1 _1650_/A sky130_fd_sc_hd__buf_1
X_1715_ _1641_/X _1051_/X _1715_/S vssd1 vssd1 vccd1 vccd1 _1715_/X sky130_fd_sc_hd__mux2_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ _1582_/A _1577_/B vssd1 vssd1 vccd1 vccd1 _1578_/A sky130_fd_sc_hd__and2_2
XFILLER_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_7_0_clk_i clkbuf_4_7_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1930_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1500_ _1863_/Q vssd1 vssd1 vccd1 vccd1 _1500_/Y sky130_fd_sc_hd__inv_2
X_1431_ data_addr_o[0] _1419_/X _1397_/X _1420_/X vssd1 vssd1 vccd1 vccd1 _1871_/D
+ sky130_fd_sc_hd__a22o_2
X_1362_ _1362_/A vssd1 vssd1 vccd1 vccd1 _1362_/X sky130_fd_sc_hd__buf_1
X_1293_ _1666_/B _1293_/B _1293_/C vssd1 vssd1 vccd1 vccd1 _1308_/C sky130_fd_sc_hd__or3_2
X_1629_ _1634_/A _1629_/B vssd1 vssd1 vccd1 vccd1 _1629_/Y sky130_fd_sc_hd__nor2_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ _1846_/Q vssd1 vssd1 vccd1 vccd1 _0931_/X sky130_fd_sc_hd__buf_1
X_1414_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1415_/A sky130_fd_sc_hd__buf_1
X_1276_ _1276_/A vssd1 vssd1 vccd1 vccd1 _1647_/B sky130_fd_sc_hd__buf_1
X_1345_ _1345_/A vssd1 vssd1 vccd1 vccd1 _1345_/X sky130_fd_sc_hd__buf_1
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_10_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1130_ _1115_/Y _1803_/S _1122_/B _0928_/A _1129_/Y vssd1 vssd1 vccd1 vccd1 _1940_/D
+ sky130_fd_sc_hd__o311a_2
XFILLER_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1061_ _1860_/Q _1061_/B vssd1 vssd1 vccd1 vccd1 _1061_/Y sky130_fd_sc_hd__nor2_2
X_1963_ _1965_/CLK _1963_/D _0967_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[12] sky130_fd_sc_hd__dfrtp_2
X_0914_ _1207_/A vssd1 vssd1 vccd1 vccd1 _1198_/A sky130_fd_sc_hd__buf_1
X_1894_ _1971_/CLK _1894_/D vssd1 vssd1 vccd1 vccd1 _1894_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1328_ _1328_/A vssd1 vssd1 vccd1 vccd1 _1328_/X sky130_fd_sc_hd__buf_1
X_1259_ _1263_/B _1257_/X _1250_/A _1255_/Y _1258_/X vssd1 vssd1 vccd1 vccd1 _1260_/A
+ sky130_fd_sc_hd__o32a_2
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1044_ _1044_/A vssd1 vssd1 vccd1 vccd1 _1044_/X sky130_fd_sc_hd__buf_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1113_ _1939_/Q vssd1 vssd1 vccd1 vccd1 _1340_/B sky130_fd_sc_hd__buf_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1877_ _1938_/CLK _1877_/D _1407_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[6] sky130_fd_sc_hd__dfrtp_2
X_1946_ _1949_/CLK _1946_/D _1089_/X vssd1 vssd1 vccd1 vccd1 _1946_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1421__A1 data_addr_o[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1185__B1 data_rdata_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1176__B1 data_rdata_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1800_ _1552_/B _1553_/X _1802_/S vssd1 vssd1 vccd1 vccd1 _1834_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1662_ _1676_/A _1664_/C vssd1 vssd1 vccd1 vccd1 _1663_/A sky130_fd_sc_hd__or2_2
X_1731_ _1680_/X _1235_/Y _1732_/S vssd1 vssd1 vccd1 vccd1 _1810_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1167__B1 data_rdata_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1593_ _1593_/A vssd1 vssd1 vccd1 vccd1 _1594_/B sky130_fd_sc_hd__buf_1
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1027_ _1027_/A _1843_/Q _1393_/A vssd1 vssd1 vccd1 vccd1 _1068_/C sky130_fd_sc_hd__or3b_2
X_1929_ _1930_/CLK _1929_/D vssd1 vssd1 vccd1 vccd1 _1929_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1158__B1 data_rdata_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_3_0_clk_i clkbuf_4_3_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1941_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1714_ _1809_/Q _1530_/X _1718_/S vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__mux2_1
X_1576_ _1574_/Y _1570_/Y _1579_/B vssd1 vssd1 vccd1 vccd1 _1577_/B sky130_fd_sc_hd__o21ai_2
X_1645_ _1645_/A vssd1 vssd1 vccd1 vccd1 _1645_/X sky130_fd_sc_hd__buf_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1430_ _1430_/A vssd1 vssd1 vccd1 vccd1 _1430_/X sky130_fd_sc_hd__buf_1
X_1361_ _1361_/A vssd1 vssd1 vccd1 vccd1 _1362_/A sky130_fd_sc_hd__buf_1
X_1292_ _1756_/X vssd1 vssd1 vccd1 vccd1 _1293_/C sky130_fd_sc_hd__inv_2
XFILLER_11_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1628_ _1629_/B vssd1 vssd1 vccd1 vccd1 _1628_/Y sky130_fd_sc_hd__inv_2
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1559_ _1836_/Q _1575_/A vssd1 vssd1 vccd1 vccd1 _1565_/B sky130_fd_sc_hd__or2_2
XFILLER_36_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_0930_ _0930_/A vssd1 vssd1 vccd1 vccd1 _0930_/X sky130_fd_sc_hd__buf_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1413_ data_addr_o[5] _1401_/X _1412_/X _1403_/X vssd1 vssd1 vccd1 vccd1 _1876_/D
+ sky130_fd_sc_hd__a22o_2
X_1275_ _1432_/A _1275_/B vssd1 vssd1 vccd1 vccd1 _1276_/A sky130_fd_sc_hd__or2_2
X_1344_ _1344_/A vssd1 vssd1 vccd1 vccd1 _1345_/A sky130_fd_sc_hd__buf_1
XFILLER_42_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1060_ _1498_/A _1635_/A _1332_/A _1402_/A _1059_/X vssd1 vssd1 vccd1 vccd1 _1060_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1962_ _1965_/CLK _1962_/D _0970_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[11] sky130_fd_sc_hd__dfrtp_2
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1893_ _1950_/CLK _1893_/D vssd1 vssd1 vccd1 vccd1 _1893_/Q sky130_fd_sc_hd__dfxtp_2
X_0913_ _1208_/A vssd1 vssd1 vccd1 vccd1 _1207_/A sky130_fd_sc_hd__buf_1
X_1189_ _1913_/Q _1186_/X data_rdata_i[6] _1187_/X _1184_/X vssd1 vssd1 vccd1 vccd1
+ _1913_/D sky130_fd_sc_hd__o221a_2
X_1327_ _1344_/A vssd1 vssd1 vccd1 vccd1 _1328_/A sky130_fd_sc_hd__buf_1
X_1258_ _1458_/A vssd1 vssd1 vccd1 vccd1 _1258_/X sky130_fd_sc_hd__buf_1
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1043_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1044_/A sky130_fd_sc_hd__buf_1
X_1112_ data_rvalid_i vssd1 vssd1 vccd1 vccd1 _1117_/B sky130_fd_sc_hd__inv_2
X_1945_ _1945_/CLK _1945_/D _1095_/X vssd1 vssd1 vccd1 vccd1 _1945_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1876_ _1876_/CLK _1876_/D _1411_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[5] sky130_fd_sc_hd__dfrtp_2
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0999__A1 data_wdata_o[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0923__A1 data_wdata_o[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1661_ _1661_/A vssd1 vssd1 vccd1 vccd1 _1676_/A sky130_fd_sc_hd__buf_1
X_1592_ _1718_/S _1592_/B vssd1 vssd1 vccd1 vccd1 _1593_/A sky130_fd_sc_hd__or2_2
X_1730_ _1653_/C _1586_/A _1761_/S vssd1 vssd1 vccd1 vccd1 _1730_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1026_ _1844_/Q _1027_/A _1843_/Q vssd1 vssd1 vccd1 vccd1 _1532_/A sky130_fd_sc_hd__or3b_2
XFILLER_14_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1928_ _1938_/CLK _1928_/D vssd1 vssd1 vccd1 vccd1 _1928_/Q sky130_fd_sc_hd__dfxtp_2
X_1859_ _1859_/CLK _1859_/D vssd1 vssd1 vccd1 vccd1 _1859_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1125__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1713_ _1808_/Q _1528_/X _1718_/S vssd1 vssd1 vccd1 vccd1 _1713_/X sky130_fd_sc_hd__mux2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1575_ _1575_/A _1575_/B vssd1 vssd1 vccd1 vccd1 _1579_/B sky130_fd_sc_hd__or2_2
X_1644_ _1894_/Q _1644_/B _1896_/Q _1895_/Q vssd1 vssd1 vccd1 vccd1 _1645_/A sky130_fd_sc_hd__or4_2
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1009_ _1018_/A vssd1 vssd1 vccd1 vccd1 _1010_/A sky130_fd_sc_hd__buf_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1379__A1 data_wdata_o[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1360_ data_addr_o[8] _1347_/X _0946_/X _1349_/A vssd1 vssd1 vccd1 vccd1 _1887_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1291_ _1754_/X vssd1 vssd1 vccd1 vccd1 _1293_/B sky130_fd_sc_hd__inv_2
XFILLER_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1489_ _0906_/B _1486_/X _0987_/B _1488_/X vssd1 vssd1 vccd1 vccd1 _1862_/D sky130_fd_sc_hd__o22ai_2
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1627_ _1829_/Q _1626_/B _1626_/Y vssd1 vssd1 vccd1 vccd1 _1629_/B sky130_fd_sc_hd__a21oi_2
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1558_ _1558_/A vssd1 vssd1 vccd1 vccd1 _1558_/X sky130_fd_sc_hd__buf_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_1_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1412_ _1848_/Q vssd1 vssd1 vccd1 vccd1 _1412_/X sky130_fd_sc_hd__buf_1
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1343_ _1343_/A vssd1 vssd1 vccd1 vccd1 _1891_/D sky130_fd_sc_hd__buf_1
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1274_ _1274_/A vssd1 vssd1 vccd1 vccd1 _1313_/B sky130_fd_sc_hd__inv_2
X_0989_ _1005_/A vssd1 vssd1 vccd1 vccd1 _0989_/X sky130_fd_sc_hd__buf_1
XFILLER_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1961_ _1965_/CLK _1961_/D _0976_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[10] sky130_fd_sc_hd__dfrtp_2
X_0912_ rst_i vssd1 vssd1 vccd1 vccd1 _1208_/A sky130_fd_sc_hd__inv_2
X_1892_ _1941_/CLK _1892_/D _1328_/X vssd1 vssd1 vccd1 vccd1 _1892_/Q sky130_fd_sc_hd__dfrtp_2
X_1326_ _1893_/Q _1477_/A _1644_/B _1312_/A vssd1 vssd1 vccd1 vccd1 _1893_/D sky130_fd_sc_hd__o22a_2
X_1188_ _1914_/Q _1186_/X data_rdata_i[7] _1187_/X _1184_/X vssd1 vssd1 vccd1 vccd1
+ _1914_/D sky130_fd_sc_hd__o221a_2
X_1257_ _1901_/Q _1256_/A _1255_/Y _1256_/Y vssd1 vssd1 vccd1 vccd1 _1257_/X sky130_fd_sc_hd__o22a_2
XFILLER_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1042_ _1351_/A vssd1 vssd1 vccd1 vccd1 _1088_/A sky130_fd_sc_hd__buf_1
X_1111_ _1940_/Q vssd1 vssd1 vccd1 vccd1 _1117_/A sky130_fd_sc_hd__inv_2
X_1875_ _1938_/CLK _1875_/D _1415_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[4] sky130_fd_sc_hd__dfrtp_2
X_1944_ _1945_/CLK _1944_/D _1100_/X vssd1 vssd1 vccd1 vccd1 _1944_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1309_ _1309_/A vssd1 vssd1 vccd1 vccd1 _1749_/S sky130_fd_sc_hd__buf_1
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1660_ _1755_/X vssd1 vssd1 vccd1 vccd1 _1664_/C sky130_fd_sc_hd__inv_2
XFILLER_7_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1591_ _1229_/A _1822_/Q _1821_/Q _1590_/Y vssd1 vssd1 vccd1 vccd1 _1592_/B sky130_fd_sc_hd__o22a_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1025_ _1850_/Q _1065_/B _1025_/C vssd1 vssd1 vccd1 vccd1 _1027_/A sky130_fd_sc_hd__or3_2
X_1927_ _1930_/CLK _1927_/D vssd1 vssd1 vccd1 vccd1 _1927_/Q sky130_fd_sc_hd__dfxtp_2
X_1858_ _1943_/CLK _1858_/D vssd1 vssd1 vccd1 vccd1 _1858_/Q sky130_fd_sc_hd__dfxtp_2
X_1789_ _1600_/B _1601_/X _1791_/S vssd1 vssd1 vccd1 vccd1 _1823_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1712_ _1670_/X _1757_/X _1749_/S vssd1 vssd1 vccd1 vccd1 _1712_/X sky130_fd_sc_hd__mux2_1
X_1643_ _1643_/A vssd1 vssd1 vccd1 vccd1 _1722_/S sky130_fd_sc_hd__buf_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1574_ _1839_/Q vssd1 vssd1 vccd1 vccd1 _1574_/Y sky130_fd_sc_hd__inv_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1008_ _1008_/A vssd1 vssd1 vccd1 vccd1 _1018_/A sky130_fd_sc_hd__buf_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1290_ _1758_/X vssd1 vssd1 vccd1 vccd1 _1666_/B sky130_fd_sc_hd__inv_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1626_ _1829_/Q _1626_/B vssd1 vssd1 vccd1 vccd1 _1626_/Y sky130_fd_sc_hd__nor2_2
X_1488_ _1485_/A _1061_/B _1330_/X _1483_/B _1487_/X vssd1 vssd1 vccd1 vccd1 _1488_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1557_ _1557_/A _1557_/B vssd1 vssd1 vccd1 vccd1 _1558_/A sky130_fd_sc_hd__and2_2
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_5_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1411_ _1411_/A vssd1 vssd1 vccd1 vccd1 _1411_/X sky130_fd_sc_hd__buf_1
XFILLER_3_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1273_ _1894_/Q _1893_/Q vssd1 vssd1 vccd1 vccd1 _1274_/A sky130_fd_sc_hd__or2_2
X_1342_ _1891_/Q _1715_/X _1342_/S vssd1 vssd1 vccd1 vccd1 _1343_/A sky130_fd_sc_hd__mux2_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0988_ _1869_/Q _0988_/B vssd1 vssd1 vccd1 vccd1 _1005_/A sky130_fd_sc_hd__nand2_2
XANTENNA__0962__B1 _0916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1609_ _1609_/A _1609_/B vssd1 vssd1 vccd1 vccd1 _1610_/A sky130_fd_sc_hd__and2_2
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1130__B1 _0928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0911_ data_wdata_o[23] _0907_/X _0908_/X _0910_/X vssd1 vssd1 vccd1 vccd1 _1974_/D
+ sky130_fd_sc_hd__a22o_2
X_1960_ _1965_/CLK _1960_/D _0979_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[9] sky130_fd_sc_hd__dfrtp_2
X_1891_ _1903_/CLK _1891_/D _1339_/X vssd1 vssd1 vccd1 vccd1 _1891_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1197__B1 data_rdata_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1325_ _1325_/A vssd1 vssd1 vccd1 vccd1 _1477_/A sky130_fd_sc_hd__inv_2
X_1256_ _1256_/A vssd1 vssd1 vccd1 vccd1 _1256_/Y sky130_fd_sc_hd__inv_2
X_1187_ _1194_/A vssd1 vssd1 vccd1 vccd1 _1187_/X sky130_fd_sc_hd__buf_1
XFILLER_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1188__B1 data_rdata_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1942_/D sky130_fd_sc_hd__buf_1
X_1041_ _1369_/A vssd1 vssd1 vccd1 vccd1 _1351_/A sky130_fd_sc_hd__buf_1
X_1874_ _1876_/CLK _1874_/D _1418_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[3] sky130_fd_sc_hd__dfrtp_2
X_1943_ _1943_/CLK _1943_/D _1104_/X vssd1 vssd1 vccd1 vccd1 _1943_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__0917__B1 _0916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1308_ _1755_/X _1308_/B _1308_/C _1308_/D vssd1 vssd1 vccd1 vccd1 _1309_/A sky130_fd_sc_hd__or4_2
X_1239_ _1250_/A vssd1 vssd1 vccd1 vccd1 _1240_/A sky130_fd_sc_hd__buf_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1590_ _1822_/Q vssd1 vssd1 vccd1 vccd1 _1590_/Y sky130_fd_sc_hd__inv_2
X_1024_ _1848_/Q _1847_/Q _1846_/Q _1845_/Q vssd1 vssd1 vccd1 vccd1 _1025_/C sky130_fd_sc_hd__or4_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1926_ _1930_/CLK _1926_/D vssd1 vssd1 vccd1 vccd1 _1926_/Q sky130_fd_sc_hd__dfxtp_2
X_1857_ _1943_/CLK _1857_/D vssd1 vssd1 vccd1 vccd1 _1857_/Q sky130_fd_sc_hd__dfxtp_2
X_1788_ _1604_/B _1605_/X _1791_/S vssd1 vssd1 vccd1 vccd1 _1824_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1711_ _1805_/Q _1521_/X _1718_/S vssd1 vssd1 vccd1 vccd1 _1711_/X sky130_fd_sc_hd__mux2_1
X_1642_ _1642_/A _1747_/S _1647_/C vssd1 vssd1 vccd1 vccd1 _1643_/A sky130_fd_sc_hd__and3_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _1586_/A _1573_/B vssd1 vssd1 vccd1 vccd1 _1573_/Y sky130_fd_sc_hd__nor2_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1007_ data_wdata_o[3] _1005_/X _0931_/X _1006_/X vssd1 vssd1 vccd1 vccd1 _1954_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1909_ _1949_/CLK _1909_/D vssd1 vssd1 vccd1 vccd1 _1909_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1625_ _1625_/A vssd1 vssd1 vccd1 vccd1 _1625_/X sky130_fd_sc_hd__buf_1
X_1556_ _1556_/A vssd1 vssd1 vccd1 vccd1 _1557_/B sky130_fd_sc_hd__buf_1
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _1490_/A _1869_/Q _1335_/X _0904_/A _1482_/A vssd1 vssd1 vccd1 vccd1 _1487_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1410_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1411_/A sky130_fd_sc_hd__buf_1
XFILLER_3_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1272_ _1895_/Q vssd1 vssd1 vccd1 vccd1 _1313_/A sky130_fd_sc_hd__inv_2
X_1341_ _1330_/A _1482_/A _1340_/Y _1060_/X _1070_/Y vssd1 vssd1 vccd1 vccd1 _1342_/S
+ sky130_fd_sc_hd__o311a_2
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0987_ _1058_/C _0987_/B _1863_/Q _1331_/A vssd1 vssd1 vccd1 vccd1 _0988_/B sky130_fd_sc_hd__and4b_2
XFILLER_22_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0962__A1 data_wdata_o[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1608_ _1608_/A vssd1 vssd1 vccd1 vccd1 _1609_/B sky130_fd_sc_hd__buf_1
X_1539_ _1661_/A vssd1 vssd1 vccd1 vccd1 _1586_/A sky130_fd_sc_hd__buf_1
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0910_ _0932_/A vssd1 vssd1 vccd1 vccd1 _0910_/X sky130_fd_sc_hd__buf_1
X_1890_ _1971_/CLK _1890_/D _1345_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[11] sky130_fd_sc_hd__dfrtp_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1186_ _1193_/A vssd1 vssd1 vccd1 vccd1 _1186_/X sky130_fd_sc_hd__buf_1
XANTENNA__1121__B2 data_gnt_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1324_ _1321_/Y _1313_/C _1476_/A _1323_/X vssd1 vssd1 vccd1 vccd1 _1894_/D sky130_fd_sc_hd__o22ai_2
X_1255_ _1901_/Q vssd1 vssd1 vccd1 vccd1 _1255_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1360__A1 data_addr_o[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1040_ _1022_/X _1036_/Y _1067_/A _1332_/A _1039_/X vssd1 vssd1 vccd1 vccd1 _1950_/D
+ sky130_fd_sc_hd__a32o_2
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1942_ _1943_/CLK _1942_/D _1108_/X vssd1 vssd1 vccd1 vccd1 _1942_/Q sky130_fd_sc_hd__dfrtp_2
X_1873_ _1876_/CLK _1873_/D _1424_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[2] sky130_fd_sc_hd__dfrtp_2
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1169_ _1923_/Q _1163_/X data_rdata_i[16] _1164_/X _1168_/X vssd1 vssd1 vccd1 vccd1
+ _1923_/D sky130_fd_sc_hd__o221a_2
X_1307_ _1655_/B vssd1 vssd1 vccd1 vccd1 _1308_/D sky130_fd_sc_hd__inv_2
X_1238_ _1458_/A vssd1 vssd1 vccd1 vccd1 _1250_/A sky130_fd_sc_hd__inv_2
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1023_ _1849_/Q vssd1 vssd1 vccd1 vccd1 _1065_/B sky130_fd_sc_hd__inv_2
X_1925_ _1949_/CLK _1925_/D vssd1 vssd1 vccd1 vccd1 _1925_/Q sky130_fd_sc_hd__dfxtp_2
X_1856_ _1943_/CLK _1856_/D vssd1 vssd1 vccd1 vccd1 _1856_/Q sky130_fd_sc_hd__dfxtp_2
X_1787_ _1609_/B _1610_/X _1791_/S vssd1 vssd1 vccd1 vccd1 _1825_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1641_ _1535_/A _1061_/Y _1483_/B _1636_/X vssd1 vssd1 vccd1 vccd1 _1641_/X sky130_fd_sc_hd__a2bb2o_2
X_1572_ _1573_/B vssd1 vssd1 vccd1 vccd1 _1572_/Y sky130_fd_sc_hd__inv_2
X_1710_ _1251_/A _1235_/Y _1740_/S vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__mux2_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1006_ _1006_/A vssd1 vssd1 vccd1 vccd1 _1006_/X sky130_fd_sc_hd__buf_1
X_1908_ _1949_/CLK _1908_/D vssd1 vssd1 vccd1 vccd1 _1908_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1839_ _1842_/CLK _1839_/D vssd1 vssd1 vccd1 vccd1 _1839_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1472__B1 _1557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1624_ _1632_/A _1624_/B vssd1 vssd1 vccd1 vccd1 _1625_/A sky130_fd_sc_hd__and2_2
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1555_ _1835_/Q _1297_/B _1575_/A vssd1 vssd1 vccd1 vccd1 _1556_/A sky130_fd_sc_hd__a21bo_2
XFILLER_39_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1486_ _1535_/A _1492_/C _1535_/B vssd1 vssd1 vccd1 vccd1 _1486_/X sky130_fd_sc_hd__o21a_2
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1340_ _1941_/Q _1340_/B vssd1 vssd1 vccd1 vccd1 _1340_/Y sky130_fd_sc_hd__nor2_2
X_1271_ _1896_/Q vssd1 vssd1 vccd1 vccd1 _1271_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0986_ _1062_/A vssd1 vssd1 vccd1 vccd1 _1331_/A sky130_fd_sc_hd__inv_2
X_1607_ _1825_/Q _1606_/B _1617_/C vssd1 vssd1 vccd1 vccd1 _1608_/A sky130_fd_sc_hd__a21bo_2
X_1538_ _1562_/A vssd1 vssd1 vccd1 vccd1 _1661_/A sky130_fd_sc_hd__inv_2
X_1469_ rx_i vssd1 vssd1 vccd1 vccd1 _1562_/A sky130_fd_sc_hd__buf_1
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1323_ _1321_/Y _1893_/Q _1894_/Q _1644_/B vssd1 vssd1 vccd1 vccd1 _1323_/X sky130_fd_sc_hd__a22o_2
X_1185_ _1915_/Q _1179_/X data_rdata_i[8] _1180_/X _1184_/X vssd1 vssd1 vccd1 vccd1
+ _1915_/D sky130_fd_sc_hd__o221a_2
X_1254_ _1902_/Q _1250_/X _1241_/X _1253_/X vssd1 vssd1 vccd1 vccd1 _1902_/D sky130_fd_sc_hd__a22o_2
XFILLER_32_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0969_ _0969_/A vssd1 vssd1 vccd1 vccd1 _0970_/A sky130_fd_sc_hd__buf_1
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1872_ _1876_/CLK _1872_/D _1427_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[1] sky130_fd_sc_hd__dfrtp_2
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1941_ _1941_/CLK _1941_/D vssd1 vssd1 vccd1 vccd1 _1941_/Q sky130_fd_sc_hd__dfxtp_2
X_1306_ _1306_/A vssd1 vssd1 vccd1 vccd1 _1655_/B sky130_fd_sc_hd__buf_1
X_1168_ _1184_/A vssd1 vssd1 vccd1 vccd1 _1168_/X sky130_fd_sc_hd__buf_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1099_ _1107_/A vssd1 vssd1 vccd1 vccd1 _1100_/A sky130_fd_sc_hd__buf_1
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1237_ _1679_/A _1251_/A _1679_/B _1466_/B vssd1 vssd1 vccd1 vccd1 _1458_/A sky130_fd_sc_hd__o211a_2
XANTENNA__1351__A _1351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1022_ _1432_/B vssd1 vssd1 vccd1 vccd1 _1022_/X sky130_fd_sc_hd__buf_1
X_1924_ _1930_/CLK _1924_/D vssd1 vssd1 vccd1 vccd1 _1924_/Q sky130_fd_sc_hd__dfxtp_2
X_1855_ _1943_/CLK _1855_/D vssd1 vssd1 vccd1 vccd1 _1855_/Q sky130_fd_sc_hd__dfxtp_2
X_1786_ _1615_/B _1616_/X _1791_/S vssd1 vssd1 vccd1 vccd1 _1826_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1640_ _1075_/X _1764_/X _1408_/X _1077_/X vssd1 vssd1 vccd1 vccd1 _1640_/X sky130_fd_sc_hd__a22o_2
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1571_ _1838_/Q _1570_/B _1570_/Y vssd1 vssd1 vccd1 vccd1 _1573_/B sky130_fd_sc_hd__a21oi_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1005_ _1005_/A vssd1 vssd1 vccd1 vccd1 _1005_/X sky130_fd_sc_hd__buf_1
X_1907_ _1949_/CLK _1907_/D vssd1 vssd1 vccd1 vccd1 _1907_/Q sky130_fd_sc_hd__dfxtp_2
X_1838_ _1842_/CLK _1838_/D vssd1 vssd1 vccd1 vccd1 _1838_/Q sky130_fd_sc_hd__dfxtp_2
X_1769_ _1768_/X _1927_/Q _1864_/Q vssd1 vssd1 vccd1 vccd1 _1769_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1485_ _1485_/A vssd1 vssd1 vccd1 vccd1 _1535_/A sky130_fd_sc_hd__buf_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1623_ _1623_/A vssd1 vssd1 vccd1 vccd1 _1624_/B sky130_fd_sc_hd__buf_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1554_ _1554_/A vssd1 vssd1 vccd1 vccd1 _1575_/A sky130_fd_sc_hd__buf_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

