magic
tech sky130A
magscale 1 2
timestamp 1640734596
<< locali >>
rect 9505 28951 9539 29257
rect 10333 28067 10367 28169
rect 10149 27319 10183 27421
rect 13921 26843 13955 27013
rect 22569 25687 22603 25857
rect 8769 24259 8803 24361
rect 24777 23579 24811 23681
rect 29653 23307 29687 28917
rect 19073 23171 19107 23273
rect 24225 20927 24259 21029
rect 19533 20315 19567 20417
rect 29653 16983 29687 17493
rect 26893 15351 26927 15589
rect 21465 15011 21499 15113
rect 19073 14331 19107 14569
rect 11345 13719 11379 14025
rect 14105 12087 14139 12189
rect 7389 10455 7423 10693
rect 20637 8959 20671 9061
rect 3341 5559 3375 5865
rect 29653 3519 29687 16949
<< viali >>
rect 10333 30277 10367 30311
rect 14289 30277 14323 30311
rect 9597 30209 9631 30243
rect 9983 30212 10017 30246
rect 10149 30209 10183 30243
rect 11713 30209 11747 30243
rect 12082 30209 12116 30243
rect 12265 30209 12299 30243
rect 14473 30209 14507 30243
rect 14638 30209 14672 30243
rect 14749 30209 14783 30243
rect 15025 30209 15059 30243
rect 16957 30209 16991 30243
rect 17140 30209 17174 30243
rect 17509 30209 17543 30243
rect 17877 30209 17911 30243
rect 9781 30141 9815 30175
rect 9873 30141 9907 30175
rect 11897 30141 11931 30175
rect 11989 30141 12023 30175
rect 14841 30141 14875 30175
rect 17233 30141 17267 30175
rect 17325 30141 17359 30175
rect 11253 30073 11287 30107
rect 9505 30005 9539 30039
rect 11621 30005 11655 30039
rect 15117 30005 15151 30039
rect 17601 30005 17635 30039
rect 17601 29733 17635 29767
rect 2973 29665 3007 29699
rect 4261 29665 4295 29699
rect 6653 29665 6687 29699
rect 13001 29665 13035 29699
rect 7113 29597 7147 29631
rect 10425 29597 10459 29631
rect 10977 29597 11011 29631
rect 12725 29597 12759 29631
rect 12909 29597 12943 29631
rect 13111 29597 13145 29631
rect 13277 29597 13311 29631
rect 13461 29597 13495 29631
rect 15577 29597 15611 29631
rect 17417 29597 17451 29631
rect 18981 29597 19015 29631
rect 7380 29529 7414 29563
rect 10158 29529 10192 29563
rect 11244 29529 11278 29563
rect 15310 29529 15344 29563
rect 17150 29529 17184 29563
rect 18714 29529 18748 29563
rect 8493 29461 8527 29495
rect 9045 29461 9079 29495
rect 12357 29461 12391 29495
rect 12633 29461 12667 29495
rect 14197 29461 14231 29495
rect 16037 29461 16071 29495
rect 8033 29257 8067 29291
rect 9505 29257 9539 29291
rect 13645 29257 13679 29291
rect 13921 29257 13955 29291
rect 14197 29257 14231 29291
rect 16773 29257 16807 29291
rect 8125 29121 8159 29155
rect 8494 29121 8528 29155
rect 8677 29121 8711 29155
rect 8309 29053 8343 29087
rect 8401 29053 8435 29087
rect 7757 28985 7791 29019
rect 12532 29189 12566 29223
rect 16138 29189 16172 29223
rect 9956 29121 9990 29155
rect 14289 29121 14323 29155
rect 14658 29121 14692 29155
rect 14841 29121 14875 29155
rect 16865 29121 16899 29155
rect 17234 29121 17268 29155
rect 17417 29147 17451 29181
rect 9689 29053 9723 29087
rect 12265 29053 12299 29087
rect 14473 29053 14507 29087
rect 14565 29053 14599 29087
rect 16405 29053 16439 29087
rect 17049 29053 17083 29087
rect 17141 29053 17175 29087
rect 15025 28985 15059 29019
rect 17601 28985 17635 29019
rect 9505 28917 9539 28951
rect 11069 28917 11103 28951
rect 29653 28917 29687 28951
rect 9873 28713 9907 28747
rect 10609 28713 10643 28747
rect 12449 28713 12483 28747
rect 14565 28713 14599 28747
rect 14841 28713 14875 28747
rect 11253 28645 11287 28679
rect 10149 28577 10183 28611
rect 16129 28577 16163 28611
rect 9965 28509 9999 28543
rect 10241 28509 10275 28543
rect 10351 28509 10385 28543
rect 10517 28509 10551 28543
rect 10793 28509 10827 28543
rect 11069 28509 11103 28543
rect 12633 28509 12667 28543
rect 14749 28509 14783 28543
rect 15025 28509 15059 28543
rect 15117 28509 15151 28543
rect 10885 28373 10919 28407
rect 15301 28373 15335 28407
rect 15577 28373 15611 28407
rect 15945 28373 15979 28407
rect 16037 28373 16071 28407
rect 17877 28373 17911 28407
rect 7757 28169 7791 28203
rect 9689 28169 9723 28203
rect 10333 28169 10367 28203
rect 12909 28169 12943 28203
rect 17877 28169 17911 28203
rect 21005 28169 21039 28203
rect 6193 28101 6227 28135
rect 6622 28101 6656 28135
rect 10425 28101 10459 28135
rect 11345 28101 11379 28135
rect 11774 28101 11808 28135
rect 5457 28033 5491 28067
rect 5640 28033 5674 28067
rect 5733 28033 5767 28067
rect 6009 28033 6043 28067
rect 6377 28033 6411 28067
rect 8208 28033 8242 28067
rect 9873 28033 9907 28067
rect 9965 28033 9999 28067
rect 10333 28033 10367 28067
rect 10609 28033 10643 28067
rect 10774 28033 10808 28067
rect 10885 28033 10919 28067
rect 11161 28033 11195 28067
rect 14298 28033 14332 28067
rect 14565 28033 14599 28067
rect 14749 28033 14783 28067
rect 16230 28033 16264 28067
rect 16957 28033 16991 28067
rect 17140 28033 17174 28067
rect 17233 28033 17267 28067
rect 17509 28033 17543 28067
rect 17693 28033 17727 28067
rect 18990 28033 19024 28067
rect 20821 28033 20855 28067
rect 21465 28033 21499 28067
rect 5825 27965 5859 27999
rect 7941 27965 7975 27999
rect 10977 27965 11011 27999
rect 11529 27965 11563 27999
rect 16497 27965 16531 27999
rect 17325 27965 17359 27999
rect 19257 27965 19291 27999
rect 9321 27829 9355 27863
rect 10149 27829 10183 27863
rect 13185 27829 13219 27863
rect 14933 27829 14967 27863
rect 15117 27829 15151 27863
rect 21649 27829 21683 27863
rect 6377 27625 6411 27659
rect 10057 27625 10091 27659
rect 8953 27557 8987 27591
rect 11253 27557 11287 27591
rect 11713 27557 11747 27591
rect 13185 27557 13219 27591
rect 13921 27557 13955 27591
rect 15853 27557 15887 27591
rect 17509 27557 17543 27591
rect 22937 27557 22971 27591
rect 7481 27489 7515 27523
rect 7665 27489 7699 27523
rect 9321 27489 9355 27523
rect 10333 27489 10367 27523
rect 10517 27489 10551 27523
rect 12725 27489 12759 27523
rect 12817 27489 12851 27523
rect 14289 27489 14323 27523
rect 14381 27489 14415 27523
rect 15485 27489 15519 27523
rect 16957 27489 16991 27523
rect 19349 27489 19383 27523
rect 9137 27421 9171 27455
rect 9413 27421 9447 27455
rect 9523 27418 9557 27452
rect 9689 27421 9723 27455
rect 9873 27421 9907 27455
rect 10149 27421 10183 27455
rect 11069 27421 11103 27455
rect 11897 27421 11931 27455
rect 12446 27421 12480 27455
rect 12632 27421 12666 27455
rect 13001 27421 13035 27455
rect 13737 27421 13771 27455
rect 15117 27421 15151 27455
rect 15300 27415 15334 27449
rect 15393 27421 15427 27455
rect 15623 27421 15657 27455
rect 16589 27421 16623 27455
rect 16772 27421 16806 27455
rect 16865 27421 16899 27455
rect 17141 27421 17175 27455
rect 18889 27421 18923 27455
rect 21097 27421 21131 27455
rect 21189 27421 21223 27455
rect 10609 27353 10643 27387
rect 17325 27353 17359 27387
rect 18622 27353 18656 27387
rect 20821 27353 20855 27387
rect 21465 27353 21499 27387
rect 7757 27285 7791 27319
rect 8125 27285 8159 27319
rect 10149 27285 10183 27319
rect 10977 27285 11011 27319
rect 13277 27285 13311 27319
rect 14473 27285 14507 27319
rect 14841 27285 14875 27319
rect 16037 27285 16071 27319
rect 6101 27081 6135 27115
rect 6745 27081 6779 27115
rect 7113 27081 7147 27115
rect 8861 27081 8895 27115
rect 12173 27081 12207 27115
rect 12633 27081 12667 27115
rect 14381 27081 14415 27115
rect 14473 27081 14507 27115
rect 15853 27081 15887 27115
rect 16865 27081 16899 27115
rect 8769 27013 8803 27047
rect 13921 27013 13955 27047
rect 15761 27013 15795 27047
rect 20453 27013 20487 27047
rect 21281 27013 21315 27047
rect 3157 26945 3191 26979
rect 3424 26945 3458 26979
rect 4721 26945 4755 26979
rect 4988 26945 5022 26979
rect 9505 26945 9539 26979
rect 9781 26945 9815 26979
rect 12265 26945 12299 26979
rect 6561 26877 6595 26911
rect 6653 26877 6687 26911
rect 8677 26877 8711 26911
rect 12081 26877 12115 26911
rect 17049 26945 17083 26979
rect 20356 26945 20390 26979
rect 20545 26945 20579 26979
rect 20729 26945 20763 26979
rect 21005 26945 21039 26979
rect 21189 26945 21223 26979
rect 21425 26945 21459 26979
rect 14657 26877 14691 26911
rect 15945 26877 15979 26911
rect 9229 26809 9263 26843
rect 13921 26809 13955 26843
rect 20177 26809 20211 26843
rect 21557 26809 21591 26843
rect 4537 26741 4571 26775
rect 9689 26741 9723 26775
rect 9873 26741 9907 26775
rect 10149 26741 10183 26775
rect 14013 26741 14047 26775
rect 15393 26741 15427 26775
rect 17509 26741 17543 26775
rect 20821 26741 20855 26775
rect 4905 26537 4939 26571
rect 6009 26537 6043 26571
rect 8401 26537 8435 26571
rect 5733 26469 5767 26503
rect 10149 26469 10183 26503
rect 13461 26469 13495 26503
rect 17509 26469 17543 26503
rect 19257 26469 19291 26503
rect 5273 26401 5307 26435
rect 6285 26401 6319 26435
rect 7021 26401 7055 26435
rect 9597 26401 9631 26435
rect 12817 26401 12851 26435
rect 13001 26401 13035 26435
rect 15485 26401 15519 26435
rect 15669 26401 15703 26435
rect 16865 26401 16899 26435
rect 16957 26401 16991 26435
rect 23489 26401 23523 26435
rect 4997 26333 5031 26367
rect 5181 26333 5215 26367
rect 5383 26333 5417 26367
rect 5549 26333 5583 26367
rect 6101 26333 6135 26367
rect 6377 26333 6411 26367
rect 6470 26333 6504 26367
rect 6653 26333 6687 26367
rect 9689 26333 9723 26367
rect 10425 26333 10459 26367
rect 15761 26333 15795 26367
rect 16589 26333 16623 26367
rect 16772 26333 16806 26367
rect 17141 26333 17175 26367
rect 18889 26333 18923 26367
rect 19441 26333 19475 26367
rect 21741 26333 21775 26367
rect 24593 26333 24627 26367
rect 7288 26265 7322 26299
rect 9781 26265 9815 26299
rect 13093 26265 13127 26299
rect 17325 26265 17359 26299
rect 18622 26265 18656 26299
rect 19533 26265 19567 26299
rect 22017 26265 22051 26299
rect 10241 26197 10275 26231
rect 16129 26197 16163 26231
rect 24409 26197 24443 26231
rect 5733 25993 5767 26027
rect 7389 25993 7423 26027
rect 8677 25993 8711 26027
rect 9137 25993 9171 26027
rect 12633 25993 12667 26027
rect 15025 25993 15059 26027
rect 19349 25993 19383 26027
rect 25145 25993 25179 26027
rect 7573 25925 7607 25959
rect 12173 25925 12207 25959
rect 14105 25925 14139 25959
rect 14933 25925 14967 25959
rect 22201 25925 22235 25959
rect 22937 25925 22971 25959
rect 4813 25857 4847 25891
rect 5182 25857 5216 25891
rect 5365 25857 5399 25891
rect 6745 25857 6779 25891
rect 6928 25857 6962 25891
rect 7297 25857 7331 25891
rect 8769 25857 8803 25891
rect 9413 25857 9447 25891
rect 10140 25857 10174 25891
rect 12265 25857 12299 25891
rect 14197 25857 14231 25891
rect 22104 25857 22138 25891
rect 22293 25857 22327 25891
rect 22477 25857 22511 25891
rect 22569 25857 22603 25891
rect 22661 25857 22695 25891
rect 22845 25857 22879 25891
rect 23034 25857 23068 25891
rect 23397 25857 23431 25891
rect 4997 25789 5031 25823
rect 5089 25789 5123 25823
rect 7021 25789 7055 25823
rect 7113 25789 7147 25823
rect 8585 25789 8619 25823
rect 9873 25789 9907 25823
rect 12081 25789 12115 25823
rect 14289 25789 14323 25823
rect 15117 25789 15151 25823
rect 20821 25789 20855 25823
rect 21097 25789 21131 25823
rect 9505 25721 9539 25755
rect 21925 25721 21959 25755
rect 23673 25789 23707 25823
rect 23213 25721 23247 25755
rect 4445 25653 4479 25687
rect 4721 25653 4755 25687
rect 9229 25653 9263 25687
rect 11253 25653 11287 25687
rect 13737 25653 13771 25687
rect 14565 25653 14599 25687
rect 17509 25653 17543 25687
rect 22569 25653 22603 25687
rect 7941 25449 7975 25483
rect 10609 25449 10643 25483
rect 11989 25449 12023 25483
rect 16957 25449 16991 25483
rect 19993 25449 20027 25483
rect 20913 25449 20947 25483
rect 23029 25449 23063 25483
rect 23213 25449 23247 25483
rect 24593 25449 24627 25483
rect 5917 25381 5951 25415
rect 10885 25381 10919 25415
rect 21833 25381 21867 25415
rect 4169 25313 4203 25347
rect 7389 25313 7423 25347
rect 11345 25313 11379 25347
rect 11529 25313 11563 25347
rect 12817 25313 12851 25347
rect 13001 25313 13035 25347
rect 14197 25313 14231 25347
rect 14381 25313 14415 25347
rect 15209 25313 15243 25347
rect 17141 25313 17175 25347
rect 4436 25245 4470 25279
rect 6101 25245 6135 25279
rect 6469 25245 6503 25279
rect 9137 25245 9171 25279
rect 9689 25245 9723 25279
rect 9965 25245 9999 25279
rect 10130 25245 10164 25279
rect 10241 25245 10275 25279
rect 10333 25245 10367 25279
rect 10517 25245 10551 25279
rect 19625 25245 19659 25279
rect 19717 25245 19751 25279
rect 20177 25245 20211 25279
rect 21092 25245 21126 25279
rect 21465 25245 21499 25279
rect 22017 25245 22051 25279
rect 22569 25245 22603 25279
rect 22845 25245 22879 25279
rect 24409 25245 24443 25279
rect 7481 25177 7515 25211
rect 14473 25177 14507 25211
rect 15485 25177 15519 25211
rect 17417 25177 17451 25211
rect 21189 25177 21223 25211
rect 21281 25177 21315 25211
rect 5549 25109 5583 25143
rect 6285 25109 6319 25143
rect 7573 25109 7607 25143
rect 8953 25109 8987 25143
rect 9873 25109 9907 25143
rect 11621 25109 11655 25143
rect 13093 25109 13127 25143
rect 13461 25109 13495 25143
rect 14841 25109 14875 25143
rect 18889 25109 18923 25143
rect 19901 25109 19935 25143
rect 22201 25109 22235 25143
rect 22753 25109 22787 25143
rect 12725 24905 12759 24939
rect 16681 24905 16715 24939
rect 22109 24905 22143 24939
rect 12357 24837 12391 24871
rect 14565 24837 14599 24871
rect 14657 24837 14691 24871
rect 3893 24769 3927 24803
rect 4537 24769 4571 24803
rect 6377 24769 6411 24803
rect 6644 24769 6678 24803
rect 8944 24769 8978 24803
rect 10333 24769 10367 24803
rect 14381 24769 14415 24803
rect 14801 24769 14835 24803
rect 15117 24769 15151 24803
rect 15301 24769 15335 24803
rect 15393 24769 15427 24803
rect 15490 24769 15524 24803
rect 16865 24769 16899 24803
rect 18236 24769 18270 24803
rect 19809 24769 19843 24803
rect 19901 24769 19935 24803
rect 20913 24769 20947 24803
rect 21005 24769 21039 24803
rect 21373 24769 21407 24803
rect 21465 24769 21499 24803
rect 21833 24769 21867 24803
rect 22293 24769 22327 24803
rect 23213 24769 23247 24803
rect 23489 24769 23523 24803
rect 24869 24769 24903 24803
rect 25145 24769 25179 24803
rect 25697 24769 25731 24803
rect 1777 24701 1811 24735
rect 2053 24701 2087 24735
rect 3709 24701 3743 24735
rect 4445 24701 4479 24735
rect 8677 24701 8711 24735
rect 12081 24701 12115 24735
rect 12265 24701 12299 24735
rect 17969 24701 18003 24735
rect 4261 24633 4295 24667
rect 10057 24633 10091 24667
rect 10517 24633 10551 24667
rect 14933 24633 14967 24667
rect 15669 24633 15703 24667
rect 19349 24633 19383 24667
rect 21649 24633 21683 24667
rect 22017 24633 22051 24667
rect 23397 24633 23431 24667
rect 25053 24633 25087 24667
rect 3525 24565 3559 24599
rect 7757 24565 7791 24599
rect 19625 24565 19659 24599
rect 20085 24565 20119 24599
rect 21189 24565 21223 24599
rect 22385 24565 22419 24599
rect 23673 24565 23707 24599
rect 25329 24565 25363 24599
rect 25881 24565 25915 24599
rect 2697 24361 2731 24395
rect 5825 24361 5859 24395
rect 6377 24361 6411 24395
rect 6561 24361 6595 24395
rect 8677 24361 8711 24395
rect 8769 24361 8803 24395
rect 9597 24361 9631 24395
rect 11437 24361 11471 24395
rect 16681 24361 16715 24395
rect 18337 24361 18371 24395
rect 24133 24361 24167 24395
rect 29101 24361 29135 24395
rect 2421 24293 2455 24327
rect 9781 24293 9815 24327
rect 13829 24293 13863 24327
rect 22201 24293 22235 24327
rect 26433 24293 26467 24327
rect 8769 24225 8803 24259
rect 9229 24225 9263 24259
rect 9321 24225 9355 24259
rect 14197 24225 14231 24259
rect 18521 24225 18555 24259
rect 19717 24225 19751 24259
rect 22385 24225 22419 24259
rect 22661 24225 22695 24259
rect 24409 24225 24443 24259
rect 2237 24157 2271 24191
rect 2513 24157 2547 24191
rect 6009 24157 6043 24191
rect 6193 24157 6227 24191
rect 6653 24157 6687 24191
rect 6837 24157 6871 24191
rect 6929 24157 6963 24191
rect 7039 24157 7073 24191
rect 7205 24157 7239 24191
rect 8502 24157 8536 24191
rect 8950 24149 8984 24183
rect 9136 24157 9170 24191
rect 9505 24157 9539 24191
rect 9965 24157 9999 24191
rect 10057 24157 10091 24191
rect 11621 24157 11655 24191
rect 13277 24157 13311 24191
rect 13461 24157 13495 24191
rect 13697 24157 13731 24191
rect 14105 24157 14139 24191
rect 14381 24157 14415 24191
rect 14565 24157 14599 24191
rect 14841 24157 14875 24191
rect 16497 24157 16531 24191
rect 17785 24157 17819 24191
rect 18158 24157 18192 24191
rect 18705 24157 18739 24191
rect 19073 24157 19107 24191
rect 19441 24157 19475 24191
rect 21465 24157 21499 24191
rect 21649 24157 21683 24191
rect 22022 24157 22056 24191
rect 26565 24157 26599 24191
rect 26709 24157 26743 24191
rect 26985 24157 27019 24191
rect 27353 24157 27387 24191
rect 10324 24089 10358 24123
rect 11888 24089 11922 24123
rect 13553 24089 13587 24123
rect 17969 24089 18003 24123
rect 18061 24089 18095 24123
rect 19962 24089 19996 24123
rect 21833 24089 21867 24123
rect 21925 24089 21959 24123
rect 24685 24089 24719 24123
rect 26801 24089 26835 24123
rect 27629 24089 27663 24123
rect 7389 24021 7423 24055
rect 8401 24021 8435 24055
rect 13001 24021 13035 24055
rect 18889 24021 18923 24055
rect 19533 24021 19567 24055
rect 21097 24021 21131 24055
rect 21281 24021 21315 24055
rect 26157 24021 26191 24055
rect 27077 24021 27111 24055
rect 6009 23817 6043 23851
rect 7205 23817 7239 23851
rect 7665 23817 7699 23851
rect 12173 23817 12207 23851
rect 14749 23817 14783 23851
rect 16865 23817 16899 23851
rect 19817 23817 19851 23851
rect 23121 23817 23155 23851
rect 24685 23817 24719 23851
rect 28549 23817 28583 23851
rect 13737 23749 13771 23783
rect 19441 23749 19475 23783
rect 25237 23749 25271 23783
rect 27261 23749 27295 23783
rect 3525 23681 3559 23715
rect 3709 23681 3743 23715
rect 4353 23681 4387 23715
rect 4629 23681 4663 23715
rect 4896 23681 4930 23715
rect 7297 23681 7331 23715
rect 9505 23681 9539 23715
rect 9597 23681 9631 23715
rect 10057 23681 10091 23715
rect 10240 23681 10274 23715
rect 10609 23681 10643 23715
rect 11529 23681 11563 23715
rect 11712 23681 11746 23715
rect 11897 23681 11931 23715
rect 12081 23681 12115 23715
rect 13461 23681 13495 23715
rect 13553 23681 13587 23715
rect 13829 23681 13863 23715
rect 14013 23681 14047 23715
rect 16497 23681 16531 23715
rect 16681 23681 16715 23715
rect 17141 23681 17175 23715
rect 17872 23681 17906 23715
rect 17969 23681 18003 23715
rect 18061 23681 18095 23715
rect 18245 23681 18279 23715
rect 18521 23681 18555 23715
rect 19303 23681 19337 23715
rect 19533 23681 19567 23715
rect 19630 23681 19664 23715
rect 20177 23681 20211 23715
rect 20545 23681 20579 23715
rect 21097 23681 21131 23715
rect 22385 23681 22419 23715
rect 23213 23681 23247 23715
rect 24501 23681 24535 23715
rect 24777 23681 24811 23715
rect 27077 23681 27111 23715
rect 27353 23681 27387 23715
rect 27450 23681 27484 23715
rect 28089 23681 28123 23715
rect 28365 23681 28399 23715
rect 1593 23613 1627 23647
rect 1869 23613 1903 23647
rect 4261 23613 4295 23647
rect 7113 23613 7147 23647
rect 10333 23613 10367 23647
rect 10425 23613 10459 23647
rect 11805 23613 11839 23647
rect 16221 23613 16255 23647
rect 24961 23613 24995 23647
rect 26709 23613 26743 23647
rect 4077 23545 4111 23579
rect 9781 23545 9815 23579
rect 10793 23545 10827 23579
rect 18337 23545 18371 23579
rect 19993 23545 20027 23579
rect 21281 23545 21315 23579
rect 22201 23545 22235 23579
rect 24777 23545 24811 23579
rect 27629 23545 27663 23579
rect 28273 23545 28307 23579
rect 3341 23477 3375 23511
rect 9321 23477 9355 23511
rect 10977 23477 11011 23511
rect 12449 23477 12483 23511
rect 16957 23477 16991 23511
rect 17693 23477 17727 23511
rect 20453 23477 20487 23511
rect 2789 23273 2823 23307
rect 3801 23273 3835 23307
rect 4905 23273 4939 23307
rect 10241 23273 10275 23307
rect 15577 23273 15611 23307
rect 18889 23273 18923 23307
rect 19073 23273 19107 23307
rect 19901 23273 19935 23307
rect 20177 23273 20211 23307
rect 29101 23273 29135 23307
rect 29653 23273 29687 23307
rect 2697 23205 2731 23239
rect 5733 23205 5767 23239
rect 22753 23205 22787 23239
rect 27169 23205 27203 23239
rect 5181 23137 5215 23171
rect 5273 23137 5307 23171
rect 6193 23137 6227 23171
rect 8309 23137 8343 23171
rect 9689 23137 9723 23171
rect 11621 23137 11655 23171
rect 14197 23137 14231 23171
rect 19073 23137 19107 23171
rect 19533 23137 19567 23171
rect 19901 23137 19935 23171
rect 20269 23137 20303 23171
rect 27353 23137 27387 23171
rect 27629 23137 27663 23171
rect 2237 23069 2271 23103
rect 2513 23069 2547 23103
rect 2973 23069 3007 23103
rect 3985 23069 4019 23103
rect 4997 23069 5031 23103
rect 5366 23069 5400 23103
rect 5549 23069 5583 23103
rect 8033 23069 8067 23103
rect 8198 23066 8232 23100
rect 8401 23069 8435 23103
rect 8585 23069 8619 23103
rect 9873 23069 9907 23103
rect 11253 23069 11287 23103
rect 11436 23069 11470 23103
rect 11529 23069 11563 23103
rect 11805 23069 11839 23103
rect 14105 23069 14139 23103
rect 14381 23069 14415 23103
rect 14565 23069 14599 23103
rect 14749 23069 14783 23103
rect 15025 23069 15059 23103
rect 15445 23069 15479 23103
rect 17509 23069 17543 23103
rect 20177 23069 20211 23103
rect 20729 23069 20763 23103
rect 21005 23069 21039 23103
rect 22569 23069 22603 23103
rect 24593 23069 24627 23103
rect 26617 23069 26651 23103
rect 27037 23069 27071 23103
rect 4721 23001 4755 23035
rect 5917 23001 5951 23035
rect 6460 23001 6494 23035
rect 9781 23001 9815 23035
rect 12081 23001 12115 23035
rect 15209 23001 15243 23035
rect 15301 23001 15335 23035
rect 17754 23001 17788 23035
rect 21250 23001 21284 23035
rect 25329 23001 25363 23035
rect 26801 23001 26835 23035
rect 26893 23001 26927 23035
rect 2421 22933 2455 22967
rect 7573 22933 7607 22967
rect 7849 22933 7883 22967
rect 8677 22933 8711 22967
rect 9413 22933 9447 22967
rect 11897 22933 11931 22967
rect 15853 22933 15887 22967
rect 19717 22933 19751 22967
rect 20545 22933 20579 22967
rect 20913 22933 20947 22967
rect 22385 22933 22419 22967
rect 24777 22933 24811 22967
rect 25513 22933 25547 22967
rect 4905 22729 4939 22763
rect 6469 22729 6503 22763
rect 9321 22729 9355 22763
rect 13737 22729 13771 22763
rect 13829 22729 13863 22763
rect 16865 22729 16899 22763
rect 20177 22729 20211 22763
rect 22661 22729 22695 22763
rect 28641 22729 28675 22763
rect 11796 22661 11830 22695
rect 15209 22661 15243 22695
rect 15301 22661 15335 22695
rect 15945 22661 15979 22695
rect 16037 22661 16071 22695
rect 23121 22661 23155 22695
rect 23213 22661 23247 22695
rect 25881 22661 25915 22695
rect 1409 22593 1443 22627
rect 4721 22593 4755 22627
rect 4997 22593 5031 22627
rect 6561 22593 6595 22627
rect 6837 22593 6871 22627
rect 6930 22593 6964 22627
rect 7113 22593 7147 22627
rect 7941 22593 7975 22627
rect 8208 22593 8242 22627
rect 9505 22593 9539 22627
rect 9688 22593 9722 22627
rect 9781 22593 9815 22627
rect 10057 22593 10091 22627
rect 11529 22593 11563 22627
rect 13553 22593 13587 22627
rect 14013 22593 14047 22627
rect 15025 22593 15059 22627
rect 15445 22593 15479 22627
rect 15761 22593 15795 22627
rect 16134 22593 16168 22627
rect 16681 22593 16715 22627
rect 17141 22593 17175 22627
rect 17417 22593 17451 22627
rect 17601 22593 17635 22627
rect 17693 22593 17727 22627
rect 17837 22593 17871 22627
rect 18153 22593 18187 22627
rect 18409 22593 18443 22627
rect 19717 22593 19751 22627
rect 19993 22593 20027 22627
rect 20545 22593 20579 22627
rect 22109 22593 22143 22627
rect 22201 22593 22235 22627
rect 22477 22593 22511 22627
rect 22937 22593 22971 22627
rect 23310 22593 23344 22627
rect 23673 22593 23707 22627
rect 25605 22593 25639 22627
rect 25789 22593 25823 22627
rect 26025 22593 26059 22627
rect 26525 22593 26559 22627
rect 28089 22593 28123 22627
rect 28457 22593 28491 22627
rect 1685 22525 1719 22559
rect 6745 22525 6779 22559
rect 9873 22525 9907 22559
rect 19809 22525 19843 22559
rect 23949 22525 23983 22559
rect 25421 22525 25455 22559
rect 6193 22457 6227 22491
rect 17969 22457 18003 22491
rect 28273 22457 28307 22491
rect 3157 22389 3191 22423
rect 5181 22389 5215 22423
rect 10149 22389 10183 22423
rect 12909 22389 12943 22423
rect 15577 22389 15611 22423
rect 16313 22389 16347 22423
rect 16957 22389 16991 22423
rect 19533 22389 19567 22423
rect 19993 22389 20027 22423
rect 20361 22389 20395 22423
rect 21925 22389 21959 22423
rect 22385 22389 22419 22423
rect 23489 22389 23523 22423
rect 26157 22389 26191 22423
rect 26341 22389 26375 22423
rect 1869 22185 1903 22219
rect 2145 22185 2179 22219
rect 20729 22185 20763 22219
rect 22569 22185 22603 22219
rect 23949 22185 23983 22219
rect 24593 22185 24627 22219
rect 26905 22185 26939 22219
rect 6377 22117 6411 22151
rect 7113 22117 7147 22151
rect 15117 22117 15151 22151
rect 17233 22117 17267 22151
rect 25421 22117 25455 22151
rect 3893 22049 3927 22083
rect 6561 22049 6595 22083
rect 7205 22049 7239 22083
rect 12633 22049 12667 22083
rect 13185 22049 13219 22083
rect 14749 22049 14783 22083
rect 21189 22049 21223 22083
rect 2053 21981 2087 22015
rect 2329 21981 2363 22015
rect 3249 21981 3283 22015
rect 6193 21981 6227 22015
rect 6653 21981 6687 22015
rect 7297 21981 7331 22015
rect 10425 21981 10459 22015
rect 10517 21981 10551 22015
rect 13093 21981 13127 22015
rect 13369 21981 13403 22015
rect 13553 21981 13587 22015
rect 13829 21981 13863 22015
rect 14473 21981 14507 22015
rect 15301 21981 15335 22015
rect 15485 21981 15519 22015
rect 19901 21981 19935 22015
rect 20177 21981 20211 22015
rect 20361 21981 20395 22015
rect 20453 21981 20487 22015
rect 20550 21981 20584 22015
rect 22845 21981 22879 22015
rect 23121 21981 23155 22015
rect 23397 21981 23431 22015
rect 23770 21981 23804 22015
rect 24409 21981 24443 22015
rect 27169 21981 27203 22015
rect 2955 21913 2989 21947
rect 3525 21913 3559 21947
rect 4169 21913 4203 21947
rect 10158 21913 10192 21947
rect 10784 21913 10818 21947
rect 12541 21913 12575 21947
rect 15761 21913 15795 21947
rect 21434 21913 21468 21947
rect 23029 21913 23063 21947
rect 23581 21913 23615 21947
rect 23673 21913 23707 21947
rect 3433 21845 3467 21879
rect 5641 21845 5675 21879
rect 9045 21845 9079 21879
rect 11897 21845 11931 21879
rect 12081 21845 12115 21879
rect 12449 21845 12483 21879
rect 14105 21845 14139 21879
rect 14565 21845 14599 21879
rect 20085 21845 20119 21879
rect 3433 21641 3467 21675
rect 4445 21641 4479 21675
rect 5733 21641 5767 21675
rect 10517 21641 10551 21675
rect 17785 21641 17819 21675
rect 19441 21641 19475 21675
rect 28825 21641 28859 21675
rect 5457 21573 5491 21607
rect 9597 21573 9631 21607
rect 15393 21573 15427 21607
rect 15485 21573 15519 21607
rect 20637 21573 20671 21607
rect 24041 21573 24075 21607
rect 26341 21573 26375 21607
rect 26433 21573 26467 21607
rect 4629 21505 4663 21539
rect 4979 21505 5013 21539
rect 5273 21505 5307 21539
rect 5917 21505 5951 21539
rect 6101 21505 6135 21539
rect 8861 21505 8895 21539
rect 9229 21505 9263 21539
rect 9413 21505 9447 21539
rect 9873 21505 9907 21539
rect 10038 21505 10072 21539
rect 10241 21505 10275 21539
rect 10425 21505 10459 21539
rect 12449 21505 12483 21539
rect 12725 21505 12759 21539
rect 13277 21505 13311 21539
rect 14105 21505 14139 21539
rect 17141 21505 17175 21539
rect 17969 21505 18003 21539
rect 18061 21505 18095 21539
rect 19625 21505 19659 21539
rect 20453 21505 20487 21539
rect 20729 21505 20763 21539
rect 20873 21505 20907 21539
rect 22845 21505 22879 21539
rect 24317 21505 24351 21539
rect 24593 21505 24627 21539
rect 25881 21505 25915 21539
rect 26157 21505 26191 21539
rect 26530 21505 26564 21539
rect 3157 21437 3191 21471
rect 3341 21437 3375 21471
rect 5549 21437 5583 21471
rect 8309 21437 8343 21471
rect 8585 21437 8619 21471
rect 9689 21437 9723 21471
rect 10149 21437 10183 21471
rect 15669 21437 15703 21471
rect 27077 21437 27111 21471
rect 27353 21437 27387 21471
rect 12633 21369 12667 21403
rect 15025 21369 15059 21403
rect 21005 21369 21039 21403
rect 24225 21369 24259 21403
rect 26065 21369 26099 21403
rect 26709 21369 26743 21403
rect 3801 21301 3835 21335
rect 6837 21301 6871 21335
rect 8677 21301 8711 21335
rect 9045 21301 9079 21335
rect 12909 21301 12943 21335
rect 13461 21301 13495 21335
rect 14289 21301 14323 21335
rect 16957 21301 16991 21335
rect 18245 21301 18279 21335
rect 22661 21301 22695 21335
rect 24501 21301 24535 21335
rect 24777 21301 24811 21335
rect 10333 21097 10367 21131
rect 11161 21097 11195 21131
rect 23857 21097 23891 21131
rect 24133 21097 24167 21131
rect 26801 21097 26835 21131
rect 27997 21097 28031 21131
rect 2789 21029 2823 21063
rect 7205 21029 7239 21063
rect 9137 21029 9171 21063
rect 9321 21029 9355 21063
rect 11253 21029 11287 21063
rect 15669 21029 15703 21063
rect 18429 21029 18463 21063
rect 20545 21029 20579 21063
rect 24225 21029 24259 21063
rect 27537 21029 27571 21063
rect 3525 20961 3559 20995
rect 6009 20961 6043 20995
rect 6745 20961 6779 20995
rect 7389 20961 7423 20995
rect 12081 20961 12115 20995
rect 15853 20961 15887 20995
rect 16129 20961 16163 20995
rect 23581 20961 23615 20995
rect 26249 20961 26283 20995
rect 1409 20893 1443 20927
rect 3249 20893 3283 20927
rect 3341 20893 3375 20927
rect 3617 20893 3651 20927
rect 3801 20893 3835 20927
rect 5825 20893 5859 20927
rect 6653 20893 6687 20927
rect 7297 20893 7331 20927
rect 8953 20893 8987 20927
rect 9781 20893 9815 20927
rect 10241 20893 10275 20927
rect 10701 20893 10735 20927
rect 10977 20893 11011 20927
rect 11437 20893 11471 20927
rect 12449 20893 12483 20927
rect 15117 20893 15151 20927
rect 15393 20893 15427 20927
rect 15537 20893 15571 20927
rect 18061 20893 18095 20927
rect 18613 20893 18647 20927
rect 18981 20893 19015 20927
rect 19441 20893 19475 20927
rect 19809 20893 19843 20927
rect 19993 20893 20027 20927
rect 20177 20893 20211 20927
rect 20366 20893 20400 20927
rect 20913 20893 20947 20927
rect 23673 20893 23707 20927
rect 23949 20893 23983 20927
rect 24225 20893 24259 20927
rect 26525 20893 26559 20927
rect 26617 20893 26651 20927
rect 27353 20893 27387 20927
rect 27813 20893 27847 20927
rect 1676 20825 1710 20859
rect 3065 20825 3099 20859
rect 4068 20825 4102 20859
rect 5917 20825 5951 20859
rect 13921 20825 13955 20859
rect 15301 20825 15335 20859
rect 20269 20825 20303 20859
rect 23305 20825 23339 20859
rect 25973 20825 26007 20859
rect 5181 20757 5215 20791
rect 5457 20757 5491 20791
rect 9597 20757 9631 20791
rect 9873 20757 9907 20791
rect 10517 20757 10551 20791
rect 17601 20757 17635 20791
rect 17877 20757 17911 20791
rect 18797 20757 18831 20791
rect 19257 20757 19291 20791
rect 19625 20757 19659 20791
rect 20729 20757 20763 20791
rect 21833 20757 21867 20791
rect 24501 20757 24535 20791
rect 26433 20757 26467 20791
rect 3065 20553 3099 20587
rect 3433 20553 3467 20587
rect 4077 20553 4111 20587
rect 7021 20553 7055 20587
rect 12817 20553 12851 20587
rect 15117 20553 15151 20587
rect 17049 20553 17083 20587
rect 19809 20553 19843 20587
rect 22017 20553 22051 20587
rect 22661 20553 22695 20587
rect 25053 20553 25087 20587
rect 26709 20553 26743 20587
rect 5365 20485 5399 20519
rect 6561 20485 6595 20519
rect 6745 20485 6779 20519
rect 14841 20485 14875 20519
rect 15945 20485 15979 20519
rect 16405 20485 16439 20519
rect 20444 20485 20478 20519
rect 23121 20485 23155 20519
rect 27169 20485 27203 20519
rect 27721 20485 27755 20519
rect 3525 20417 3559 20451
rect 3801 20417 3835 20451
rect 3893 20417 3927 20451
rect 7297 20417 7331 20451
rect 7757 20417 7791 20451
rect 8953 20417 8987 20451
rect 9229 20417 9263 20451
rect 11897 20417 11931 20451
rect 12449 20417 12483 20451
rect 13001 20417 13035 20451
rect 14105 20417 14139 20451
rect 14657 20417 14691 20451
rect 15301 20417 15335 20451
rect 15669 20417 15703 20451
rect 15853 20417 15887 20451
rect 16042 20417 16076 20451
rect 17233 20417 17267 20451
rect 19441 20417 19475 20451
rect 19533 20417 19567 20451
rect 19625 20417 19659 20451
rect 22201 20417 22235 20451
rect 22477 20417 22511 20451
rect 22845 20417 22879 20451
rect 23029 20417 23063 20451
rect 23265 20417 23299 20451
rect 23581 20417 23615 20451
rect 23765 20417 23799 20451
rect 23857 20417 23891 20451
rect 24001 20417 24035 20451
rect 24869 20417 24903 20451
rect 25973 20417 26007 20451
rect 26525 20417 26559 20451
rect 26985 20417 27019 20451
rect 27261 20417 27295 20451
rect 27358 20417 27392 20451
rect 2789 20349 2823 20383
rect 2973 20349 3007 20383
rect 11069 20349 11103 20383
rect 11345 20349 11379 20383
rect 12265 20349 12299 20383
rect 14197 20349 14231 20383
rect 15025 20349 15059 20383
rect 19165 20349 19199 20383
rect 20177 20349 20211 20383
rect 5181 20281 5215 20315
rect 7481 20281 7515 20315
rect 9137 20281 9171 20315
rect 11989 20281 12023 20315
rect 16221 20281 16255 20315
rect 19533 20281 19567 20315
rect 23397 20281 23431 20315
rect 24133 20281 24167 20315
rect 3617 20213 3651 20247
rect 7573 20213 7607 20247
rect 9413 20213 9447 20247
rect 9597 20213 9631 20247
rect 12633 20213 12667 20247
rect 14105 20213 14139 20247
rect 14473 20213 14507 20247
rect 17693 20213 17727 20247
rect 21557 20213 21591 20247
rect 22385 20213 22419 20247
rect 24317 20213 24351 20247
rect 25789 20213 25823 20247
rect 27537 20213 27571 20247
rect 6745 20009 6779 20043
rect 13737 20009 13771 20043
rect 16129 20009 16163 20043
rect 17693 20009 17727 20043
rect 18337 20009 18371 20043
rect 21281 20009 21315 20043
rect 25329 20009 25363 20043
rect 25605 20009 25639 20043
rect 26341 20009 26375 20043
rect 15117 19941 15151 19975
rect 20453 19941 20487 19975
rect 22753 19941 22787 19975
rect 8217 19873 8251 19907
rect 8493 19873 8527 19907
rect 10793 19873 10827 19907
rect 12633 19873 12667 19907
rect 14197 19873 14231 19907
rect 26617 19873 26651 19907
rect 26893 19873 26927 19907
rect 4629 19805 4663 19839
rect 8769 19805 8803 19839
rect 12357 19805 12391 19839
rect 12541 19805 12575 19839
rect 12817 19805 12851 19839
rect 13001 19805 13035 19839
rect 14105 19805 14139 19839
rect 14933 19805 14967 19839
rect 15209 19805 15243 19839
rect 15485 19805 15519 19839
rect 15582 19805 15616 19839
rect 15945 19805 15979 19839
rect 17785 19805 17819 19839
rect 18062 19805 18096 19839
rect 18158 19805 18192 19839
rect 19901 19805 19935 19839
rect 20321 19805 20355 19839
rect 21465 19805 21499 19839
rect 22569 19805 22603 19839
rect 25053 19805 25087 19839
rect 25145 19805 25179 19839
rect 25421 19805 25455 19839
rect 26157 19805 26191 19839
rect 28733 19805 28767 19839
rect 4896 19737 4930 19771
rect 10517 19737 10551 19771
rect 13461 19737 13495 19771
rect 13645 19737 13679 19771
rect 15393 19737 15427 19771
rect 17969 19737 18003 19771
rect 20085 19737 20119 19771
rect 20177 19737 20211 19771
rect 6009 19669 6043 19703
rect 8585 19669 8619 19703
rect 9045 19669 9079 19703
rect 15769 19669 15803 19703
rect 16589 19669 16623 19703
rect 24961 19669 24995 19703
rect 28365 19669 28399 19703
rect 28549 19669 28583 19703
rect 2789 19465 2823 19499
rect 4077 19465 4111 19499
rect 4997 19465 5031 19499
rect 6837 19465 6871 19499
rect 7481 19465 7515 19499
rect 7757 19465 7791 19499
rect 9505 19465 9539 19499
rect 9781 19465 9815 19499
rect 10149 19465 10183 19499
rect 12909 19465 12943 19499
rect 13461 19465 13495 19499
rect 20453 19465 20487 19499
rect 21189 19465 21223 19499
rect 21649 19465 21683 19499
rect 26065 19465 26099 19499
rect 27353 19465 27387 19499
rect 27629 19465 27663 19499
rect 6745 19397 6779 19431
rect 7941 19397 7975 19431
rect 16865 19397 16899 19431
rect 17250 19397 17284 19431
rect 18613 19397 18647 19431
rect 23765 19397 23799 19431
rect 23857 19397 23891 19431
rect 1676 19329 1710 19363
rect 3065 19329 3099 19363
rect 3249 19329 3283 19363
rect 3341 19329 3375 19363
rect 5181 19329 5215 19363
rect 5273 19329 5307 19363
rect 7297 19329 7331 19363
rect 7573 19329 7607 19363
rect 9321 19329 9355 19363
rect 9597 19329 9631 19363
rect 9873 19329 9907 19363
rect 10333 19329 10367 19363
rect 11161 19329 11195 19363
rect 11621 19329 11655 19363
rect 11805 19329 11839 19363
rect 12081 19329 12115 19363
rect 12265 19329 12299 19363
rect 13277 19329 13311 19363
rect 13369 19329 13403 19363
rect 14197 19329 14231 19363
rect 14933 19329 14967 19363
rect 16129 19329 16163 19363
rect 16405 19329 16439 19363
rect 16681 19329 16715 19363
rect 16957 19329 16991 19363
rect 17054 19329 17088 19363
rect 17693 19329 17727 19363
rect 18377 19329 18411 19363
rect 18521 19329 18555 19363
rect 18797 19329 18831 19363
rect 20269 19329 20303 19363
rect 21373 19329 21407 19363
rect 21465 19329 21499 19363
rect 21833 19329 21867 19363
rect 22425 19329 22459 19363
rect 22568 19329 22602 19363
rect 22661 19329 22695 19363
rect 22845 19329 22879 19363
rect 23305 19329 23339 19363
rect 23581 19329 23615 19363
rect 23954 19329 23988 19363
rect 24317 19329 24351 19363
rect 26525 19329 26559 19363
rect 27169 19329 27203 19363
rect 27445 19329 27479 19363
rect 28273 19329 28307 19363
rect 1409 19261 1443 19295
rect 3617 19261 3651 19295
rect 4169 19261 4203 19295
rect 4261 19261 4295 19295
rect 5549 19261 5583 19295
rect 6929 19261 6963 19295
rect 11989 19261 12023 19295
rect 13185 19261 13219 19295
rect 14289 19261 14323 19295
rect 16037 19261 16071 19295
rect 20637 19261 20671 19295
rect 24593 19261 24627 19295
rect 3709 19193 3743 19227
rect 10057 19193 10091 19227
rect 11253 19193 11287 19227
rect 14565 19193 14599 19227
rect 14749 19193 14783 19227
rect 22017 19193 22051 19227
rect 24133 19193 24167 19227
rect 3525 19125 3559 19159
rect 5457 19125 5491 19159
rect 6377 19125 6411 19159
rect 13277 19125 13311 19159
rect 14197 19125 14231 19159
rect 17509 19125 17543 19159
rect 18245 19125 18279 19159
rect 18981 19125 19015 19159
rect 20821 19125 20855 19159
rect 22293 19125 22327 19159
rect 23029 19125 23063 19159
rect 23489 19125 23523 19159
rect 26341 19125 26375 19159
rect 28457 19125 28491 19159
rect 3893 18921 3927 18955
rect 25237 18921 25271 18955
rect 13277 18853 13311 18887
rect 21557 18853 21591 18887
rect 23857 18853 23891 18887
rect 3249 18785 3283 18819
rect 3801 18785 3835 18819
rect 11161 18785 11195 18819
rect 11989 18785 12023 18819
rect 12449 18785 12483 18819
rect 12541 18785 12575 18819
rect 14105 18785 14139 18819
rect 14381 18785 14415 18819
rect 14565 18785 14599 18819
rect 15945 18785 15979 18819
rect 18061 18785 18095 18819
rect 18337 18785 18371 18819
rect 19993 18785 20027 18819
rect 22109 18785 22143 18819
rect 27353 18785 27387 18819
rect 3433 18717 3467 18751
rect 3617 18717 3651 18751
rect 4077 18717 4111 18751
rect 4169 18717 4203 18751
rect 4905 18717 4939 18751
rect 7481 18717 7515 18751
rect 9689 18717 9723 18751
rect 10793 18717 10827 18751
rect 11069 18717 11103 18751
rect 11345 18717 11379 18751
rect 11529 18717 11563 18751
rect 12173 18717 12207 18751
rect 12265 18717 12299 18751
rect 12817 18717 12851 18751
rect 13001 18717 13035 18751
rect 13093 18717 13127 18751
rect 15669 18717 15703 18751
rect 15761 18717 15795 18751
rect 18429 18717 18463 18751
rect 18797 18717 18831 18751
rect 20260 18717 20294 18751
rect 21741 18717 21775 18751
rect 24685 18717 24719 18751
rect 24777 18717 24811 18751
rect 25053 18717 25087 18751
rect 26433 18717 26467 18751
rect 5172 18649 5206 18683
rect 11805 18649 11839 18683
rect 14841 18649 14875 18683
rect 22385 18649 22419 18683
rect 27629 18649 27663 18683
rect 4353 18581 4387 18615
rect 6285 18581 6319 18615
rect 7665 18581 7699 18615
rect 9873 18581 9907 18615
rect 14473 18581 14507 18615
rect 15301 18581 15335 18615
rect 16589 18581 16623 18615
rect 18613 18581 18647 18615
rect 18981 18581 19015 18615
rect 21373 18581 21407 18615
rect 24501 18581 24535 18615
rect 24961 18581 24995 18615
rect 26249 18581 26283 18615
rect 29101 18581 29135 18615
rect 2605 18377 2639 18411
rect 4077 18377 4111 18411
rect 4537 18377 4571 18411
rect 5273 18377 5307 18411
rect 15393 18377 15427 18411
rect 15761 18377 15795 18411
rect 17601 18377 17635 18411
rect 20913 18377 20947 18411
rect 23305 18377 23339 18411
rect 23397 18377 23431 18411
rect 9229 18309 9263 18343
rect 13093 18309 13127 18343
rect 14381 18309 14415 18343
rect 18429 18309 18463 18343
rect 2421 18241 2455 18275
rect 2697 18241 2731 18275
rect 2964 18241 2998 18275
rect 4721 18241 4755 18275
rect 5457 18241 5491 18275
rect 5549 18241 5583 18275
rect 5825 18241 5859 18275
rect 10977 18241 11011 18275
rect 12173 18241 12207 18275
rect 12357 18241 12391 18275
rect 13277 18241 13311 18275
rect 14013 18241 14047 18275
rect 14197 18241 14231 18275
rect 14749 18241 14783 18275
rect 17417 18241 17451 18275
rect 17693 18241 17727 18275
rect 18153 18241 18187 18275
rect 20729 18241 20763 18275
rect 21097 18241 21131 18275
rect 23121 18241 23155 18275
rect 23581 18241 23615 18275
rect 24133 18241 24167 18275
rect 24317 18241 24351 18275
rect 24409 18241 24443 18275
rect 24506 18241 24540 18275
rect 24961 18241 24995 18275
rect 27169 18241 27203 18275
rect 27353 18241 27387 18275
rect 27445 18241 27479 18275
rect 27542 18241 27576 18275
rect 6653 18173 6687 18207
rect 6929 18173 6963 18207
rect 8953 18173 8987 18207
rect 10701 18173 10735 18207
rect 15853 18173 15887 18207
rect 16037 18173 16071 18207
rect 25237 18173 25271 18207
rect 5733 18105 5767 18139
rect 24685 18105 24719 18139
rect 27721 18105 27755 18139
rect 8401 18037 8435 18071
rect 11069 18037 11103 18071
rect 11989 18037 12023 18071
rect 12357 18037 12391 18071
rect 13001 18037 13035 18071
rect 14841 18037 14875 18071
rect 17877 18037 17911 18071
rect 19901 18037 19935 18071
rect 20637 18037 20671 18071
rect 26709 18037 26743 18071
rect 27905 18037 27939 18071
rect 4261 17833 4295 17867
rect 7205 17833 7239 17867
rect 7481 17833 7515 17867
rect 9689 17833 9723 17867
rect 12357 17833 12391 17867
rect 7849 17765 7883 17799
rect 20085 17765 20119 17799
rect 22753 17765 22787 17799
rect 27353 17765 27387 17799
rect 1409 17697 1443 17731
rect 3525 17697 3559 17731
rect 4077 17697 4111 17731
rect 6469 17697 6503 17731
rect 6561 17697 6595 17731
rect 8217 17697 8251 17731
rect 12725 17697 12759 17731
rect 14749 17697 14783 17731
rect 16221 17697 16255 17731
rect 3249 17629 3283 17663
rect 3341 17629 3375 17663
rect 3617 17629 3651 17663
rect 3801 17629 3835 17663
rect 3985 17629 4019 17663
rect 4445 17629 4479 17663
rect 7389 17629 7423 17663
rect 7665 17629 7699 17663
rect 9505 17629 9539 17663
rect 9965 17629 9999 17663
rect 12449 17629 12483 17663
rect 12587 17629 12621 17663
rect 12818 17629 12852 17663
rect 13001 17629 13035 17663
rect 13093 17629 13127 17663
rect 13599 17629 13633 17663
rect 13829 17629 13863 17663
rect 14335 17629 14369 17663
rect 14473 17629 14507 17663
rect 18337 17629 18371 17663
rect 20264 17629 20298 17663
rect 20637 17629 20671 17663
rect 22201 17629 22235 17663
rect 22621 17629 22655 17663
rect 23121 17629 23155 17663
rect 23397 17629 23431 17663
rect 24685 17629 24719 17663
rect 25329 17629 25363 17663
rect 26801 17629 26835 17663
rect 26985 17629 27019 17663
rect 27221 17629 27255 17663
rect 1676 17561 1710 17595
rect 3065 17561 3099 17595
rect 6377 17561 6411 17595
rect 8309 17561 8343 17595
rect 8401 17561 8435 17595
rect 13921 17561 13955 17595
rect 14841 17561 14875 17595
rect 16497 17561 16531 17595
rect 20361 17561 20395 17595
rect 20453 17561 20487 17595
rect 22385 17561 22419 17595
rect 22477 17561 22511 17595
rect 27077 17561 27111 17595
rect 2789 17493 2823 17527
rect 6009 17493 6043 17527
rect 9781 17493 9815 17527
rect 13277 17493 13311 17527
rect 14197 17493 14231 17527
rect 17969 17493 18003 17527
rect 18153 17493 18187 17527
rect 19809 17493 19843 17527
rect 20729 17493 20763 17527
rect 20913 17493 20947 17527
rect 22109 17493 22143 17527
rect 23305 17493 23339 17527
rect 23581 17493 23615 17527
rect 24869 17493 24903 17527
rect 25053 17493 25087 17527
rect 25145 17493 25179 17527
rect 27629 17493 27663 17527
rect 29653 17493 29687 17527
rect 7665 17289 7699 17323
rect 12909 17289 12943 17323
rect 13645 17289 13679 17323
rect 16313 17289 16347 17323
rect 16681 17289 16715 17323
rect 23949 17289 23983 17323
rect 24501 17289 24535 17323
rect 11989 17221 12023 17255
rect 14657 17221 14691 17255
rect 19717 17221 19751 17255
rect 20913 17221 20947 17255
rect 27261 17221 27295 17255
rect 4373 17153 4407 17187
rect 4629 17153 4663 17187
rect 4721 17153 4755 17187
rect 4988 17153 5022 17187
rect 7481 17153 7515 17187
rect 7849 17153 7883 17187
rect 9045 17153 9079 17187
rect 12449 17153 12483 17187
rect 13277 17153 13311 17187
rect 13553 17153 13587 17187
rect 13829 17153 13863 17187
rect 14473 17153 14507 17187
rect 14749 17153 14783 17187
rect 14841 17153 14875 17187
rect 15117 17153 15151 17187
rect 15393 17153 15427 17187
rect 15577 17153 15611 17187
rect 15761 17153 15795 17187
rect 16037 17153 16071 17187
rect 16221 17153 16255 17187
rect 16865 17153 16899 17187
rect 19993 17153 20027 17187
rect 20085 17153 20119 17187
rect 20453 17153 20487 17187
rect 20729 17153 20763 17187
rect 21005 17153 21039 17187
rect 21149 17153 21183 17187
rect 24133 17153 24167 17187
rect 9321 17085 9355 17119
rect 11897 17085 11931 17119
rect 12173 17085 12207 17119
rect 13093 17085 13127 17119
rect 13185 17085 13219 17119
rect 13369 17085 13403 17119
rect 15301 17085 15335 17119
rect 16129 17085 16163 17119
rect 23581 17085 23615 17119
rect 23857 17085 23891 17119
rect 25973 17085 26007 17119
rect 26249 17085 26283 17119
rect 26985 17085 27019 17119
rect 14289 17017 14323 17051
rect 20269 17017 20303 17051
rect 3249 16949 3283 16983
rect 6101 16949 6135 16983
rect 8033 16949 8067 16983
rect 10793 16949 10827 16983
rect 11713 16949 11747 16983
rect 12265 16949 12299 16983
rect 18245 16949 18279 16983
rect 20637 16949 20671 16983
rect 21281 16949 21315 16983
rect 22109 16949 22143 16983
rect 28733 16949 28767 16983
rect 29653 16949 29687 16983
rect 4629 16745 4663 16779
rect 5365 16745 5399 16779
rect 5825 16745 5859 16779
rect 9965 16745 9999 16779
rect 11713 16745 11747 16779
rect 12081 16745 12115 16779
rect 15485 16745 15519 16779
rect 25053 16745 25087 16779
rect 28089 16745 28123 16779
rect 4997 16677 5031 16711
rect 18613 16677 18647 16711
rect 19257 16677 19291 16711
rect 1409 16609 1443 16643
rect 5917 16609 5951 16643
rect 6469 16609 6503 16643
rect 6561 16609 6595 16643
rect 6929 16609 6963 16643
rect 10977 16609 11011 16643
rect 11621 16609 11655 16643
rect 12173 16609 12207 16643
rect 21557 16609 21591 16643
rect 21833 16609 21867 16643
rect 25237 16609 25271 16643
rect 2973 16541 3007 16575
rect 4077 16541 4111 16575
rect 4353 16541 4387 16575
rect 4497 16541 4531 16575
rect 4813 16541 4847 16575
rect 5549 16541 5583 16575
rect 5641 16541 5675 16575
rect 9781 16541 9815 16575
rect 10701 16541 10735 16575
rect 10885 16541 10919 16575
rect 11161 16541 11195 16575
rect 11345 16541 11379 16575
rect 11529 16541 11563 16575
rect 12081 16541 12115 16575
rect 12633 16541 12667 16575
rect 17141 16541 17175 16575
rect 17233 16541 17267 16575
rect 18797 16541 18831 16575
rect 19441 16541 19475 16575
rect 23673 16541 23707 16575
rect 24501 16541 24535 16575
rect 24777 16541 24811 16575
rect 24921 16541 24955 16575
rect 26709 16541 26743 16575
rect 27169 16541 27203 16575
rect 27542 16541 27576 16575
rect 27905 16541 27939 16575
rect 1676 16473 1710 16507
rect 3157 16473 3191 16507
rect 3341 16473 3375 16507
rect 4261 16473 4295 16507
rect 6377 16473 6411 16507
rect 7205 16473 7239 16507
rect 16773 16473 16807 16507
rect 24685 16473 24719 16507
rect 27353 16473 27387 16507
rect 27445 16473 27479 16507
rect 2789 16405 2823 16439
rect 6009 16405 6043 16439
rect 8677 16405 8711 16439
rect 11897 16405 11931 16439
rect 12449 16405 12483 16439
rect 12725 16405 12759 16439
rect 16865 16405 16899 16439
rect 18981 16405 19015 16439
rect 20085 16405 20119 16439
rect 23857 16405 23891 16439
rect 26893 16405 26927 16439
rect 27729 16405 27763 16439
rect 2881 16201 2915 16235
rect 5089 16201 5123 16235
rect 7481 16201 7515 16235
rect 8493 16201 8527 16235
rect 11069 16201 11103 16235
rect 14013 16201 14047 16235
rect 14565 16201 14599 16235
rect 16865 16201 16899 16235
rect 16957 16201 16991 16235
rect 20269 16201 20303 16235
rect 2329 16133 2363 16167
rect 3617 16133 3651 16167
rect 3709 16133 3743 16167
rect 9321 16133 9355 16167
rect 9413 16133 9447 16167
rect 17233 16133 17267 16167
rect 22109 16133 22143 16167
rect 27629 16133 27663 16167
rect 2513 16065 2547 16099
rect 2769 16065 2803 16099
rect 2973 16065 3007 16099
rect 3249 16065 3283 16099
rect 3433 16065 3467 16099
rect 3985 16065 4019 16099
rect 4353 16065 4387 16099
rect 4629 16065 4663 16099
rect 4905 16065 4939 16099
rect 7665 16065 7699 16099
rect 8585 16065 8619 16099
rect 10517 16065 10551 16099
rect 10977 16065 11011 16099
rect 12061 16065 12095 16099
rect 12173 16065 12207 16099
rect 12449 16065 12483 16099
rect 12633 16065 12667 16099
rect 12816 16065 12850 16099
rect 12909 16065 12943 16099
rect 13001 16065 13035 16099
rect 13185 16065 13219 16099
rect 14105 16065 14139 16099
rect 14473 16065 14507 16099
rect 14933 16065 14967 16099
rect 15301 16065 15335 16099
rect 15761 16065 15795 16099
rect 16037 16065 16071 16099
rect 16681 16065 16715 16099
rect 17049 16065 17083 16099
rect 20453 16065 20487 16099
rect 21925 16065 21959 16099
rect 22201 16065 22235 16099
rect 22298 16065 22332 16099
rect 22661 16065 22695 16099
rect 24593 16065 24627 16099
rect 24961 16065 24995 16099
rect 27353 16065 27387 16099
rect 3065 15997 3099 16031
rect 3893 15997 3927 16031
rect 8493 15997 8527 16031
rect 9229 15997 9263 16031
rect 12541 15997 12575 16031
rect 14197 15997 14231 16031
rect 15025 15997 15059 16031
rect 15209 15997 15243 16031
rect 16129 15997 16163 16031
rect 17325 15997 17359 16031
rect 17601 15997 17635 16031
rect 22937 15997 22971 16031
rect 24409 15997 24443 16031
rect 25237 15997 25271 16031
rect 8033 15929 8067 15963
rect 13645 15929 13679 15963
rect 15945 15929 15979 15963
rect 22477 15929 22511 15963
rect 4445 15861 4479 15895
rect 4813 15861 4847 15895
rect 8861 15861 8895 15895
rect 10701 15861 10735 15895
rect 11897 15861 11931 15895
rect 13277 15861 13311 15895
rect 15669 15861 15703 15895
rect 16037 15861 16071 15895
rect 16405 15861 16439 15895
rect 19073 15861 19107 15895
rect 20637 15861 20671 15895
rect 24777 15861 24811 15895
rect 26709 15861 26743 15895
rect 29101 15861 29135 15895
rect 4537 15657 4571 15691
rect 14381 15657 14415 15691
rect 17233 15657 17267 15691
rect 18429 15657 18463 15691
rect 19349 15657 19383 15691
rect 21373 15657 21407 15691
rect 23765 15657 23799 15691
rect 25145 15657 25179 15691
rect 26617 15657 26651 15691
rect 28641 15657 28675 15691
rect 5733 15589 5767 15623
rect 9229 15589 9263 15623
rect 16037 15589 16071 15623
rect 25789 15589 25823 15623
rect 26893 15589 26927 15623
rect 26985 15589 27019 15623
rect 27721 15589 27755 15623
rect 28273 15589 28307 15623
rect 2881 15521 2915 15555
rect 3065 15521 3099 15555
rect 4169 15521 4203 15555
rect 4353 15521 4387 15555
rect 9965 15521 9999 15555
rect 11437 15521 11471 15555
rect 16129 15521 16163 15555
rect 17785 15521 17819 15555
rect 17877 15521 17911 15555
rect 23121 15521 23155 15555
rect 2973 15453 3007 15487
rect 3157 15453 3191 15487
rect 3341 15453 3375 15487
rect 4445 15453 4479 15487
rect 4537 15453 4571 15487
rect 4629 15453 4663 15487
rect 5181 15453 5215 15487
rect 5365 15453 5399 15487
rect 5554 15453 5588 15487
rect 7122 15453 7156 15487
rect 7389 15453 7423 15487
rect 8125 15453 8159 15487
rect 9045 15453 9079 15487
rect 9505 15453 9539 15487
rect 9689 15453 9723 15487
rect 16313 15453 16347 15487
rect 16497 15453 16531 15487
rect 17371 15453 17405 15487
rect 17509 15453 17543 15487
rect 18245 15453 18279 15487
rect 18705 15453 18739 15487
rect 18981 15453 19015 15487
rect 21097 15453 21131 15487
rect 23397 15453 23431 15487
rect 23581 15453 23615 15487
rect 24501 15453 24535 15487
rect 25324 15453 25358 15487
rect 25697 15453 25731 15487
rect 26341 15453 26375 15487
rect 26801 15429 26835 15463
rect 5462 15385 5496 15419
rect 14105 15385 14139 15419
rect 14289 15385 14323 15419
rect 15669 15385 15703 15419
rect 15853 15385 15887 15419
rect 20821 15385 20855 15419
rect 22845 15385 22879 15419
rect 25421 15385 25455 15419
rect 25513 15385 25547 15419
rect 27169 15453 27203 15487
rect 27542 15453 27576 15487
rect 28089 15453 28123 15487
rect 28457 15453 28491 15487
rect 27353 15385 27387 15419
rect 27445 15385 27479 15419
rect 2697 15317 2731 15351
rect 3985 15317 4019 15351
rect 4905 15317 4939 15351
rect 6009 15317 6043 15351
rect 7941 15317 7975 15351
rect 9321 15317 9355 15351
rect 18521 15317 18555 15351
rect 18797 15317 18831 15351
rect 23213 15317 23247 15351
rect 24685 15317 24719 15351
rect 26525 15317 26559 15351
rect 26893 15317 26927 15351
rect 3065 15113 3099 15147
rect 4261 15113 4295 15147
rect 4721 15113 4755 15147
rect 10701 15113 10735 15147
rect 10977 15113 11011 15147
rect 12173 15113 12207 15147
rect 15485 15113 15519 15147
rect 16773 15113 16807 15147
rect 19993 15113 20027 15147
rect 21465 15113 21499 15147
rect 21557 15113 21591 15147
rect 22753 15113 22787 15147
rect 24409 15113 24443 15147
rect 26341 15113 26375 15147
rect 5457 15045 5491 15079
rect 7757 15045 7791 15079
rect 18797 15045 18831 15079
rect 19349 15045 19383 15079
rect 1409 14977 1443 15011
rect 1676 14977 1710 15011
rect 3249 14977 3283 15011
rect 3341 14977 3375 15011
rect 3617 14977 3651 15011
rect 3893 14977 3927 15011
rect 4905 14977 4939 15011
rect 5641 14977 5675 15011
rect 5733 14977 5767 15011
rect 9689 14977 9723 15011
rect 10517 14977 10551 15011
rect 10793 14977 10827 15011
rect 12357 14977 12391 15011
rect 12633 14977 12667 15011
rect 12817 14977 12851 15011
rect 13093 14977 13127 15011
rect 13369 14977 13403 15011
rect 13461 14977 13495 15011
rect 13737 14977 13771 15011
rect 13921 14977 13955 15011
rect 14289 14977 14323 15011
rect 14473 14977 14507 15011
rect 14565 14977 14599 15011
rect 14841 14977 14875 15011
rect 15025 14977 15059 15011
rect 15209 14977 15243 15011
rect 15577 14977 15611 15011
rect 16037 14977 16071 15011
rect 16865 14977 16899 15011
rect 18981 14977 19015 15011
rect 19441 14977 19475 15011
rect 19901 14977 19935 15011
rect 20269 14977 20303 15011
rect 20453 14977 20487 15011
rect 20545 14977 20579 15011
rect 20689 14977 20723 15011
rect 21097 14977 21131 15011
rect 21465 14977 21499 15011
rect 21833 14977 21867 15011
rect 21971 14977 22005 15011
rect 22106 14977 22140 15011
rect 22253 14977 22287 15011
rect 22569 14977 22603 15011
rect 24317 14977 24351 15011
rect 24593 14977 24627 15011
rect 25053 14977 25087 15011
rect 26157 14977 26191 15011
rect 26525 14977 26559 15011
rect 3985 14909 4019 14943
rect 7481 14909 7515 14943
rect 14657 14909 14691 14943
rect 15853 14909 15887 14943
rect 16313 14909 16347 14943
rect 2789 14841 2823 14875
rect 5273 14841 5307 14875
rect 12449 14841 12483 14875
rect 12541 14841 12575 14875
rect 19165 14841 19199 14875
rect 19625 14841 19659 14875
rect 20821 14841 20855 14875
rect 22385 14841 22419 14875
rect 24869 14841 24903 14875
rect 3525 14773 3559 14807
rect 4077 14773 4111 14807
rect 5825 14773 5859 14807
rect 9229 14773 9263 14807
rect 9873 14773 9907 14807
rect 12909 14773 12943 14807
rect 13185 14773 13219 14807
rect 13553 14773 13587 14807
rect 21281 14773 21315 14807
rect 24777 14773 24811 14807
rect 26709 14773 26743 14807
rect 1961 14569 1995 14603
rect 3249 14569 3283 14603
rect 3801 14569 3835 14603
rect 13001 14569 13035 14603
rect 13461 14569 13495 14603
rect 14197 14569 14231 14603
rect 14565 14569 14599 14603
rect 15577 14569 15611 14603
rect 16773 14569 16807 14603
rect 19073 14569 19107 14603
rect 19441 14569 19475 14603
rect 20361 14569 20395 14603
rect 16957 14501 16991 14535
rect 11713 14433 11747 14467
rect 12541 14433 12575 14467
rect 2053 14365 2087 14399
rect 3157 14365 3191 14399
rect 3985 14365 4019 14399
rect 5641 14365 5675 14399
rect 5917 14365 5951 14399
rect 8217 14365 8251 14399
rect 8309 14365 8343 14399
rect 8493 14365 8527 14399
rect 9965 14365 9999 14399
rect 11345 14365 11379 14399
rect 11621 14365 11655 14399
rect 11897 14365 11931 14399
rect 12081 14365 12115 14399
rect 12725 14365 12759 14399
rect 12817 14365 12851 14399
rect 13093 14365 13127 14399
rect 13553 14365 13587 14399
rect 14381 14365 14415 14399
rect 14565 14365 14599 14399
rect 15301 14365 15335 14399
rect 15485 14365 15519 14399
rect 15761 14365 15795 14399
rect 15991 14365 16025 14399
rect 16313 14365 16347 14399
rect 16405 14365 16439 14399
rect 17417 14365 17451 14399
rect 17877 14365 17911 14399
rect 24133 14501 24167 14535
rect 24685 14501 24719 14535
rect 25329 14501 25363 14535
rect 19441 14433 19475 14467
rect 25513 14433 25547 14467
rect 25789 14433 25823 14467
rect 19809 14365 19843 14399
rect 20177 14365 20211 14399
rect 21373 14365 21407 14399
rect 23213 14365 23247 14399
rect 23581 14365 23615 14399
rect 23857 14365 23891 14399
rect 23954 14365 23988 14399
rect 24777 14365 24811 14399
rect 25197 14365 25231 14399
rect 27997 14365 28031 14399
rect 28365 14365 28399 14399
rect 12357 14297 12391 14331
rect 13277 14297 13311 14331
rect 15117 14297 15151 14331
rect 16782 14297 16816 14331
rect 17233 14297 17267 14331
rect 17601 14297 17635 14331
rect 19073 14297 19107 14331
rect 23765 14297 23799 14331
rect 24501 14297 24535 14331
rect 24961 14297 24995 14331
rect 25053 14297 25087 14331
rect 5733 14229 5767 14263
rect 10149 14229 10183 14263
rect 16129 14229 16163 14263
rect 16221 14229 16255 14263
rect 17785 14229 17819 14263
rect 19625 14229 19659 14263
rect 21557 14229 21591 14263
rect 23029 14229 23063 14263
rect 23397 14229 23431 14263
rect 27261 14229 27295 14263
rect 28181 14229 28215 14263
rect 28549 14229 28583 14263
rect 3341 14025 3375 14059
rect 5089 14025 5123 14059
rect 6193 14025 6227 14059
rect 8033 14025 8067 14059
rect 11345 14025 11379 14059
rect 12541 14025 12575 14059
rect 13093 14025 13127 14059
rect 13185 14025 13219 14059
rect 15485 14025 15519 14059
rect 15853 14025 15887 14059
rect 16681 14025 16715 14059
rect 19533 14025 19567 14059
rect 21281 14025 21315 14059
rect 24225 14025 24259 14059
rect 26617 14025 26651 14059
rect 29101 14025 29135 14059
rect 3893 13957 3927 13991
rect 5825 13957 5859 13991
rect 6898 13957 6932 13991
rect 8585 13957 8619 13991
rect 8769 13957 8803 13991
rect 3157 13889 3191 13923
rect 3709 13889 3743 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 4446 13911 4480 13945
rect 4554 13889 4588 13923
rect 4813 13889 4847 13923
rect 4905 13889 4939 13923
rect 5733 13889 5767 13923
rect 8401 13889 8435 13923
rect 8861 13889 8895 13923
rect 9137 13889 9171 13923
rect 11069 13889 11103 13923
rect 4077 13821 4111 13855
rect 5641 13821 5675 13855
rect 6653 13821 6687 13855
rect 9413 13821 9447 13855
rect 10885 13821 10919 13855
rect 11161 13821 11195 13855
rect 14657 13957 14691 13991
rect 14841 13957 14875 13991
rect 15025 13957 15059 13991
rect 16313 13957 16347 13991
rect 17325 13957 17359 13991
rect 20821 13957 20855 13991
rect 27629 13957 27663 13991
rect 12081 13889 12115 13923
rect 12173 13889 12207 13923
rect 13001 13889 13035 13923
rect 13369 13889 13403 13923
rect 14105 13889 14139 13923
rect 15117 13889 15151 13923
rect 15577 13889 15611 13923
rect 15945 13889 15979 13923
rect 16129 13889 16163 13923
rect 16865 13889 16899 13923
rect 17049 13889 17083 13923
rect 17233 13889 17267 13923
rect 17469 13889 17503 13923
rect 17785 13889 17819 13923
rect 20085 13889 20119 13923
rect 20632 13889 20666 13923
rect 20729 13889 20763 13923
rect 21005 13889 21039 13923
rect 21097 13889 21131 13923
rect 24409 13889 24443 13923
rect 26433 13889 26467 13923
rect 12357 13821 12391 13855
rect 18061 13821 18095 13855
rect 20177 13821 20211 13855
rect 21373 13821 21407 13855
rect 22385 13821 22419 13855
rect 23857 13821 23891 13855
rect 24133 13821 24167 13855
rect 27353 13821 27387 13855
rect 12817 13753 12851 13787
rect 15301 13753 15335 13787
rect 17601 13753 17635 13787
rect 9045 13685 9079 13719
rect 11345 13685 11379 13719
rect 14289 13685 14323 13719
rect 20453 13685 20487 13719
rect 9045 13481 9079 13515
rect 12081 13481 12115 13515
rect 12265 13481 12299 13515
rect 18705 13481 18739 13515
rect 22293 13481 22327 13515
rect 23121 13481 23155 13515
rect 5457 13413 5491 13447
rect 8033 13413 8067 13447
rect 17325 13413 17359 13447
rect 25329 13413 25363 13447
rect 4629 13345 4663 13379
rect 6009 13345 6043 13379
rect 8677 13345 8711 13379
rect 16773 13345 16807 13379
rect 16865 13345 16899 13379
rect 20545 13345 20579 13379
rect 20821 13345 20855 13379
rect 25513 13345 25547 13379
rect 25789 13345 25823 13379
rect 2881 13277 2915 13311
rect 3157 13277 3191 13311
rect 3341 13277 3375 13311
rect 3617 13277 3651 13311
rect 4721 13277 4755 13311
rect 4813 13277 4847 13311
rect 5109 13277 5143 13311
rect 6653 13277 6687 13311
rect 8401 13277 8435 13311
rect 8585 13277 8619 13311
rect 9137 13277 9171 13311
rect 11897 13277 11931 13311
rect 11989 13277 12023 13311
rect 13645 13277 13679 13311
rect 15577 13277 15611 13311
rect 17069 13277 17103 13311
rect 17325 13277 17359 13311
rect 17601 13277 17635 13311
rect 17785 13277 17819 13311
rect 17969 13277 18003 13311
rect 18061 13277 18095 13311
rect 18521 13277 18555 13311
rect 23489 13277 23523 13311
rect 23581 13277 23615 13311
rect 23765 13277 23799 13311
rect 23954 13277 23988 13311
rect 24777 13277 24811 13311
rect 25150 13277 25184 13311
rect 2614 13209 2648 13243
rect 2973 13209 3007 13243
rect 5021 13209 5055 13243
rect 5365 13209 5399 13243
rect 6101 13209 6135 13243
rect 6898 13209 6932 13243
rect 23029 13209 23063 13243
rect 23857 13209 23891 13243
rect 24961 13209 24995 13243
rect 25053 13209 25087 13243
rect 1501 13141 1535 13175
rect 3525 13141 3559 13175
rect 4905 13141 4939 13175
rect 6193 13141 6227 13175
rect 6561 13141 6595 13175
rect 9321 13141 9355 13175
rect 13829 13141 13863 13175
rect 15393 13141 15427 13175
rect 16957 13141 16991 13175
rect 18245 13141 18279 13175
rect 22753 13141 22787 13175
rect 23305 13141 23339 13175
rect 24150 13141 24184 13175
rect 27261 13141 27295 13175
rect 2973 12937 3007 12971
rect 3525 12937 3559 12971
rect 3985 12937 4019 12971
rect 4169 12937 4203 12971
rect 4997 12937 5031 12971
rect 5457 12937 5491 12971
rect 12265 12937 12299 12971
rect 14289 12937 14323 12971
rect 16681 12937 16715 12971
rect 23029 12937 23063 12971
rect 25881 12937 25915 12971
rect 26525 12937 26559 12971
rect 2421 12869 2455 12903
rect 2605 12869 2639 12903
rect 12173 12869 12207 12903
rect 12817 12869 12851 12903
rect 16497 12869 16531 12903
rect 24409 12869 24443 12903
rect 2835 12801 2869 12835
rect 3157 12801 3191 12835
rect 3709 12801 3743 12835
rect 4167 12801 4201 12835
rect 4813 12801 4847 12835
rect 4905 12801 4939 12835
rect 5365 12801 5399 12835
rect 6561 12801 6595 12835
rect 9873 12801 9907 12835
rect 10129 12801 10163 12835
rect 11621 12801 11655 12835
rect 11805 12801 11839 12835
rect 12541 12801 12575 12835
rect 15025 12801 15059 12835
rect 16865 12801 16899 12835
rect 18521 12801 18555 12835
rect 19625 12801 19659 12835
rect 19892 12801 19926 12835
rect 22385 12801 22419 12835
rect 23213 12801 23247 12835
rect 24133 12801 24167 12835
rect 26065 12801 26099 12835
rect 26341 12801 26375 12835
rect 3065 12733 3099 12767
rect 4629 12733 4663 12767
rect 5549 12733 5583 12767
rect 14657 12733 14691 12767
rect 6377 12665 6411 12699
rect 11253 12665 11287 12699
rect 11897 12665 11931 12699
rect 26249 12665 26283 12699
rect 4537 12597 4571 12631
rect 18337 12597 18371 12631
rect 21005 12597 21039 12631
rect 22477 12597 22511 12631
rect 14289 12393 14323 12427
rect 15761 12393 15795 12427
rect 22385 12393 22419 12427
rect 25329 12393 25363 12427
rect 2973 12325 3007 12359
rect 9781 12325 9815 12359
rect 10793 12325 10827 12359
rect 13737 12325 13771 12359
rect 4445 12257 4479 12291
rect 5365 12257 5399 12291
rect 5549 12257 5583 12291
rect 9689 12257 9723 12291
rect 10241 12257 10275 12291
rect 12173 12257 12207 12291
rect 14749 12257 14783 12291
rect 17141 12257 17175 12291
rect 19625 12257 19659 12291
rect 20453 12257 20487 12291
rect 21833 12257 21867 12291
rect 23765 12257 23799 12291
rect 1593 12189 1627 12223
rect 4261 12189 4295 12223
rect 5641 12189 5675 12223
rect 7297 12189 7331 12223
rect 9597 12189 9631 12223
rect 10149 12189 10183 12223
rect 10517 12189 10551 12223
rect 10701 12189 10735 12223
rect 11805 12189 11839 12223
rect 12081 12189 12115 12223
rect 12357 12189 12391 12223
rect 13461 12189 13495 12223
rect 13921 12189 13955 12223
rect 14105 12189 14139 12223
rect 14473 12189 14507 12223
rect 14565 12189 14599 12223
rect 15577 12189 15611 12223
rect 16681 12189 16715 12223
rect 16865 12189 16899 12223
rect 19073 12189 19107 12223
rect 19257 12189 19291 12223
rect 19901 12189 19935 12223
rect 20085 12189 20119 12223
rect 20361 12189 20395 12223
rect 20637 12189 20671 12223
rect 20821 12189 20855 12223
rect 21097 12189 21131 12223
rect 21189 12189 21223 12223
rect 21373 12189 21407 12223
rect 21649 12189 21683 12223
rect 21925 12189 21959 12223
rect 22109 12189 22143 12223
rect 23498 12189 23532 12223
rect 24869 12189 24903 12223
rect 25145 12189 25179 12223
rect 1860 12121 1894 12155
rect 7564 12121 7598 12155
rect 10977 12121 11011 12155
rect 11161 12121 11195 12155
rect 12449 12121 12483 12155
rect 14841 12121 14875 12155
rect 14933 12121 14967 12155
rect 18981 12121 19015 12155
rect 19717 12121 19751 12155
rect 3801 12053 3835 12087
rect 4169 12053 4203 12087
rect 6009 12053 6043 12087
rect 8677 12053 8711 12087
rect 8953 12053 8987 12087
rect 11989 12053 12023 12087
rect 13645 12053 13679 12087
rect 14105 12053 14139 12087
rect 16589 12053 16623 12087
rect 18613 12053 18647 12087
rect 19441 12053 19475 12087
rect 25053 12053 25087 12087
rect 3801 11849 3835 11883
rect 4077 11849 4111 11883
rect 4445 11849 4479 11883
rect 7757 11849 7791 11883
rect 8401 11849 8435 11883
rect 10885 11849 10919 11883
rect 15301 11849 15335 11883
rect 15485 11849 15519 11883
rect 17049 11849 17083 11883
rect 19809 11849 19843 11883
rect 21465 11849 21499 11883
rect 22017 11849 22051 11883
rect 22845 11849 22879 11883
rect 3433 11781 3467 11815
rect 5830 11781 5864 11815
rect 8125 11781 8159 11815
rect 9781 11781 9815 11815
rect 10517 11781 10551 11815
rect 11069 11781 11103 11815
rect 13737 11781 13771 11815
rect 20545 11781 20579 11815
rect 20913 11781 20947 11815
rect 21097 11781 21131 11815
rect 22661 11781 22695 11815
rect 3249 11713 3283 11747
rect 3689 11713 3723 11747
rect 5181 11713 5215 11747
rect 5457 11713 5491 11747
rect 5549 11713 5583 11747
rect 5733 11713 5767 11747
rect 5922 11713 5956 11747
rect 6377 11713 6411 11747
rect 6633 11713 6667 11747
rect 8309 11713 8343 11747
rect 8769 11713 8803 11747
rect 8953 11713 8987 11747
rect 9137 11713 9171 11747
rect 9229 11713 9263 11747
rect 9965 11713 9999 11747
rect 10149 11713 10183 11747
rect 10333 11713 10367 11747
rect 10793 11713 10827 11747
rect 11897 11713 11931 11747
rect 11989 11713 12023 11747
rect 12173 11713 12207 11747
rect 12449 11713 12483 11747
rect 13553 11713 13587 11747
rect 15393 11713 15427 11747
rect 15669 11713 15703 11747
rect 16865 11713 16899 11747
rect 18696 11713 18730 11747
rect 20448 11713 20482 11747
rect 20637 11713 20671 11747
rect 20821 11713 20855 11747
rect 21557 11713 21591 11747
rect 22201 11713 22235 11747
rect 22293 11713 22327 11747
rect 22569 11713 22603 11747
rect 27252 11713 27286 11747
rect 3893 11645 3927 11679
rect 3985 11645 4019 11679
rect 4537 11645 4571 11679
rect 4721 11645 4755 11679
rect 18429 11645 18463 11679
rect 22477 11645 22511 11679
rect 26985 11645 27019 11679
rect 4997 11577 5031 11611
rect 5365 11577 5399 11611
rect 6101 11577 6135 11611
rect 7941 11577 7975 11611
rect 9413 11577 9447 11611
rect 10701 11577 10735 11611
rect 12265 11577 12299 11611
rect 13369 11577 13403 11611
rect 20269 11577 20303 11611
rect 8585 11509 8619 11543
rect 8953 11509 8987 11543
rect 9689 11509 9723 11543
rect 11713 11509 11747 11543
rect 12541 11509 12575 11543
rect 21189 11509 21223 11543
rect 22845 11509 22879 11543
rect 23029 11509 23063 11543
rect 28365 11509 28399 11543
rect 6929 11305 6963 11339
rect 9045 11305 9079 11339
rect 9229 11305 9263 11339
rect 11989 11305 12023 11339
rect 13921 11305 13955 11339
rect 14657 11305 14691 11339
rect 15025 11305 15059 11339
rect 15393 11305 15427 11339
rect 15577 11305 15611 11339
rect 16497 11305 16531 11339
rect 19349 11305 19383 11339
rect 19809 11305 19843 11339
rect 20913 11305 20947 11339
rect 22385 11305 22419 11339
rect 27261 11305 27295 11339
rect 1961 11237 1995 11271
rect 5733 11237 5767 11271
rect 6377 11237 6411 11271
rect 7665 11237 7699 11271
rect 27169 11237 27203 11271
rect 5089 11169 5123 11203
rect 9321 11169 9355 11203
rect 9965 11169 9999 11203
rect 10149 11169 10183 11203
rect 11713 11169 11747 11203
rect 11805 11169 11839 11203
rect 13645 11169 13679 11203
rect 19901 11169 19935 11203
rect 21097 11169 21131 11203
rect 27905 11169 27939 11203
rect 2237 11101 2271 11135
rect 5365 11101 5399 11135
rect 5825 11101 5859 11135
rect 6101 11101 6135 11135
rect 6198 11101 6232 11135
rect 7021 11101 7055 11135
rect 7389 11101 7423 11135
rect 7907 11101 7941 11135
rect 8033 11101 8067 11135
rect 8125 11101 8159 11135
rect 8309 11101 8343 11135
rect 8493 11101 8527 11135
rect 9413 11101 9447 11135
rect 9505 11101 9539 11135
rect 9781 11101 9815 11135
rect 10333 11101 10367 11135
rect 10701 11101 10735 11135
rect 11069 11101 11103 11135
rect 11253 11101 11287 11135
rect 11345 11101 11379 11135
rect 11529 11101 11563 11135
rect 11621 11101 11655 11135
rect 13378 11101 13412 11135
rect 13737 11101 13771 11135
rect 14105 11101 14139 11135
rect 14381 11101 14415 11135
rect 14657 11101 14691 11135
rect 14841 11101 14875 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 16129 11101 16163 11135
rect 16313 11101 16347 11135
rect 18153 11101 18187 11135
rect 19533 11101 19567 11135
rect 19625 11101 19659 11135
rect 20269 11101 20303 11135
rect 21189 11101 21223 11135
rect 22293 11101 22327 11135
rect 23029 11101 23063 11135
rect 23857 11101 23891 11135
rect 24041 11101 24075 11135
rect 24409 11101 24443 11135
rect 26985 11101 27019 11135
rect 27629 11101 27663 11135
rect 28089 11101 28123 11135
rect 28273 11101 28307 11135
rect 6009 11033 6043 11067
rect 8677 11033 8711 11067
rect 9597 11033 9631 11067
rect 10425 11033 10459 11067
rect 15209 11033 15243 11067
rect 17908 11033 17942 11067
rect 20177 11033 20211 11067
rect 20913 11033 20947 11067
rect 23673 11033 23707 11067
rect 24654 11033 24688 11067
rect 26065 11033 26099 11067
rect 26249 11033 26283 11067
rect 26433 11033 26467 11067
rect 1777 10965 1811 10999
rect 5273 10965 5307 10999
rect 7205 10965 7239 10999
rect 10793 10965 10827 10999
rect 12265 10965 12299 10999
rect 14565 10965 14599 10999
rect 15393 10965 15427 10999
rect 16773 10965 16807 10999
rect 21373 10965 21407 10999
rect 22937 10965 22971 10999
rect 24225 10965 24259 10999
rect 25789 10965 25823 10999
rect 27721 10965 27755 10999
rect 28457 10965 28491 10999
rect 4169 10761 4203 10795
rect 6561 10761 6595 10795
rect 7573 10761 7607 10795
rect 9045 10761 9079 10795
rect 10517 10761 10551 10795
rect 11161 10761 11195 10795
rect 12081 10761 12115 10795
rect 13093 10761 13127 10795
rect 14749 10761 14783 10795
rect 15117 10761 15151 10795
rect 17969 10761 18003 10795
rect 23673 10761 23707 10795
rect 24317 10761 24351 10795
rect 24777 10761 24811 10795
rect 25145 10761 25179 10795
rect 27721 10761 27755 10795
rect 5457 10693 5491 10727
rect 5641 10693 5675 10727
rect 7389 10693 7423 10727
rect 9965 10693 9999 10727
rect 10149 10693 10183 10727
rect 10609 10693 10643 10727
rect 19349 10693 19383 10727
rect 19533 10693 19567 10727
rect 24685 10693 24719 10727
rect 26341 10693 26375 10727
rect 26985 10693 27019 10727
rect 1501 10625 1535 10659
rect 2033 10625 2067 10659
rect 3985 10625 4019 10659
rect 5273 10625 5307 10659
rect 6377 10625 6411 10659
rect 1777 10557 1811 10591
rect 7941 10625 7975 10659
rect 8217 10625 8251 10659
rect 9413 10625 9447 10659
rect 9597 10625 9631 10659
rect 9689 10625 9723 10659
rect 9873 10625 9907 10659
rect 10405 10625 10439 10659
rect 10701 10625 10735 10659
rect 11345 10625 11379 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 11989 10625 12023 10659
rect 12173 10625 12207 10659
rect 13277 10625 13311 10659
rect 14841 10625 14875 10659
rect 14933 10625 14967 10659
rect 15209 10625 15243 10659
rect 15393 10625 15427 10659
rect 15577 10625 15611 10659
rect 15669 10625 15703 10659
rect 17601 10625 17635 10659
rect 18153 10625 18187 10659
rect 18245 10625 18279 10659
rect 18613 10625 18647 10659
rect 21097 10625 21131 10659
rect 21281 10625 21315 10659
rect 21373 10625 21407 10659
rect 22549 10625 22583 10659
rect 25329 10625 25363 10659
rect 25605 10625 25639 10659
rect 25847 10625 25881 10659
rect 26249 10625 26283 10659
rect 26525 10625 26559 10659
rect 26709 10625 26743 10659
rect 27170 10625 27204 10659
rect 27537 10625 27571 10659
rect 27905 10625 27939 10659
rect 7849 10557 7883 10591
rect 10977 10557 11011 10591
rect 17325 10557 17359 10591
rect 17509 10557 17543 10591
rect 22293 10557 22327 10591
rect 24869 10557 24903 10591
rect 26157 10557 26191 10591
rect 27629 10557 27663 10591
rect 9505 10489 9539 10523
rect 11621 10489 11655 10523
rect 21189 10489 21223 10523
rect 1685 10421 1719 10455
rect 3157 10421 3191 10455
rect 7389 10421 7423 10455
rect 7757 10421 7791 10455
rect 8125 10421 8159 10455
rect 9229 10421 9263 10455
rect 10793 10421 10827 10455
rect 15853 10421 15887 10455
rect 18429 10421 18463 10455
rect 21557 10421 21591 10455
rect 1869 10217 1903 10251
rect 3157 10217 3191 10251
rect 3617 10217 3651 10251
rect 4629 10217 4663 10251
rect 7849 10217 7883 10251
rect 10333 10217 10367 10251
rect 14197 10217 14231 10251
rect 16865 10217 16899 10251
rect 18245 10217 18279 10251
rect 24501 10217 24535 10251
rect 26709 10217 26743 10251
rect 3801 10149 3835 10183
rect 10701 10149 10735 10183
rect 12725 10149 12759 10183
rect 2329 10081 2363 10115
rect 2421 10081 2455 10115
rect 4445 10081 4479 10115
rect 5181 10081 5215 10115
rect 6009 10081 6043 10115
rect 10885 10081 10919 10115
rect 16589 10081 16623 10115
rect 18337 10081 18371 10115
rect 20085 10081 20119 10115
rect 22385 10081 22419 10115
rect 26801 10081 26835 10115
rect 27721 10081 27755 10115
rect 2237 10013 2271 10047
rect 3341 10013 3375 10047
rect 3433 10013 3467 10047
rect 5089 10013 5123 10047
rect 5825 10013 5859 10047
rect 6469 10013 6503 10047
rect 8217 10013 8251 10047
rect 8401 10013 8435 10047
rect 8953 10013 8987 10047
rect 9220 10013 9254 10047
rect 10701 10013 10735 10047
rect 11069 10013 11103 10047
rect 12725 10013 12759 10047
rect 12909 10013 12943 10047
rect 13093 10013 13127 10047
rect 15577 10013 15611 10047
rect 16773 10013 16807 10047
rect 18245 10013 18279 10047
rect 18889 10013 18923 10047
rect 19349 10013 19383 10047
rect 19809 10013 19843 10047
rect 19993 10013 20027 10047
rect 21373 10013 21407 10047
rect 22017 10013 22051 10047
rect 22293 10013 22327 10047
rect 22569 10013 22603 10047
rect 22753 10013 22787 10047
rect 24685 10013 24719 10047
rect 24869 10013 24903 10047
rect 26709 10013 26743 10047
rect 27905 10013 27939 10047
rect 28089 10013 28123 10047
rect 28273 10013 28307 10047
rect 3617 9945 3651 9979
rect 5917 9945 5951 9979
rect 6736 9945 6770 9979
rect 8033 9945 8067 9979
rect 15332 9945 15366 9979
rect 19441 9945 19475 9979
rect 20177 9945 20211 9979
rect 26985 9945 27019 9979
rect 4169 9877 4203 9911
rect 4261 9877 4295 9911
rect 4997 9877 5031 9911
rect 5457 9877 5491 9911
rect 11345 9877 11379 9911
rect 15945 9877 15979 9911
rect 16313 9877 16347 9911
rect 16405 9877 16439 9911
rect 18613 9877 18647 9911
rect 19073 9877 19107 9911
rect 21557 9877 21591 9911
rect 26525 9877 26559 9911
rect 28457 9877 28491 9911
rect 10517 9673 10551 9707
rect 14933 9673 14967 9707
rect 6745 9605 6779 9639
rect 10701 9605 10735 9639
rect 10885 9605 10919 9639
rect 12633 9605 12667 9639
rect 13921 9605 13955 9639
rect 14473 9605 14507 9639
rect 14657 9605 14691 9639
rect 17233 9605 17267 9639
rect 17417 9605 17451 9639
rect 17969 9605 18003 9639
rect 19257 9605 19291 9639
rect 19809 9605 19843 9639
rect 22293 9605 22327 9639
rect 2237 9537 2271 9571
rect 3709 9537 3743 9571
rect 4721 9537 4755 9571
rect 4988 9537 5022 9571
rect 7205 9537 7239 9571
rect 8217 9537 8251 9571
rect 10333 9537 10367 9571
rect 11161 9537 11195 9571
rect 11713 9537 11747 9571
rect 12173 9537 12207 9571
rect 12449 9537 12483 9571
rect 12725 9537 12759 9571
rect 14013 9537 14047 9571
rect 14289 9537 14323 9571
rect 15025 9537 15059 9571
rect 15577 9537 15611 9571
rect 15853 9537 15887 9571
rect 16129 9537 16163 9571
rect 17693 9537 17727 9571
rect 17785 9537 17819 9571
rect 18429 9537 18463 9571
rect 18889 9537 18923 9571
rect 19073 9537 19107 9571
rect 19533 9537 19567 9571
rect 19625 9537 19659 9571
rect 19901 9537 19935 9571
rect 20177 9537 20211 9571
rect 20637 9537 20671 9571
rect 21005 9537 21039 9571
rect 21189 9537 21223 9571
rect 22201 9537 22235 9571
rect 22753 9537 22787 9571
rect 23489 9537 23523 9571
rect 25789 9537 25823 9571
rect 25973 9537 26007 9571
rect 26249 9537 26283 9571
rect 26525 9537 26559 9571
rect 26617 9537 26651 9571
rect 27445 9537 27479 9571
rect 27988 9537 28022 9571
rect 11529 9469 11563 9503
rect 15761 9469 15795 9503
rect 15945 9469 15979 9503
rect 20729 9469 20763 9503
rect 22385 9469 22419 9503
rect 27721 9469 27755 9503
rect 1961 9401 1995 9435
rect 6561 9401 6595 9435
rect 7021 9401 7055 9435
rect 11345 9401 11379 9435
rect 12173 9401 12207 9435
rect 14197 9401 14231 9435
rect 15393 9401 15427 9435
rect 18153 9401 18187 9435
rect 20269 9401 20303 9435
rect 21833 9401 21867 9435
rect 22937 9401 22971 9435
rect 25697 9401 25731 9435
rect 26709 9401 26743 9435
rect 1777 9333 1811 9367
rect 3801 9333 3835 9367
rect 6101 9333 6135 9367
rect 8401 9333 8435 9367
rect 11897 9333 11931 9367
rect 15577 9333 15611 9367
rect 16313 9333 16347 9367
rect 17417 9333 17451 9367
rect 18245 9333 18279 9367
rect 20085 9333 20119 9367
rect 23029 9333 23063 9367
rect 23673 9333 23707 9367
rect 26157 9333 26191 9367
rect 27353 9333 27387 9367
rect 29101 9333 29135 9367
rect 3893 9129 3927 9163
rect 7757 9129 7791 9163
rect 13369 9129 13403 9163
rect 14197 9129 14231 9163
rect 16865 9129 16899 9163
rect 20085 9129 20119 9163
rect 20729 9129 20763 9163
rect 23121 9129 23155 9163
rect 27629 9129 27663 9163
rect 27905 9129 27939 9163
rect 3065 9061 3099 9095
rect 16313 9061 16347 9095
rect 18337 9061 18371 9095
rect 19257 9061 19291 9095
rect 20637 9061 20671 9095
rect 21557 9061 21591 9095
rect 26893 9061 26927 9095
rect 1685 8993 1719 9027
rect 4031 8993 4065 9027
rect 4537 8993 4571 9027
rect 10793 8993 10827 9027
rect 11989 8993 12023 9027
rect 15577 8993 15611 9027
rect 17601 8993 17635 9027
rect 18889 8993 18923 9027
rect 19901 8993 19935 9027
rect 21373 8993 21407 9027
rect 22109 8993 22143 9027
rect 22753 8993 22787 9027
rect 23765 8993 23799 9027
rect 23857 8993 23891 9027
rect 28365 8993 28399 9027
rect 28457 8993 28491 9027
rect 1409 8925 1443 8959
rect 3249 8925 3283 8959
rect 3433 8925 3467 8959
rect 4169 8925 4203 8959
rect 7205 8925 7239 8959
rect 7573 8925 7607 8959
rect 10609 8925 10643 8959
rect 11345 8925 11379 8959
rect 11437 8925 11471 8959
rect 11621 8925 11655 8959
rect 11713 8925 11747 8959
rect 12256 8925 12290 8959
rect 15669 8925 15703 8959
rect 15945 8925 15979 8959
rect 16129 8925 16163 8959
rect 16497 8925 16531 8959
rect 16589 8925 16623 8959
rect 16773 8925 16807 8959
rect 18153 8925 18187 8959
rect 18245 8925 18279 8959
rect 18613 8925 18647 8959
rect 19073 8925 19107 8959
rect 20637 8925 20671 8959
rect 22017 8925 22051 8959
rect 22385 8925 22419 8959
rect 22937 8925 22971 8959
rect 24869 8925 24903 8959
rect 26433 8925 26467 8959
rect 26617 8925 26651 8959
rect 26985 8925 27019 8959
rect 27169 8925 27203 8959
rect 27353 8925 27387 8959
rect 28273 8925 28307 8959
rect 1952 8857 1986 8891
rect 3617 8857 3651 8891
rect 4445 8857 4479 8891
rect 7021 8857 7055 8891
rect 7389 8857 7423 8891
rect 10701 8857 10735 8891
rect 15332 8857 15366 8891
rect 17417 8857 17451 8891
rect 21189 8857 21223 8891
rect 25136 8857 25170 8891
rect 27721 8857 27755 8891
rect 1593 8789 1627 8823
rect 10241 8789 10275 8823
rect 11161 8789 11195 8823
rect 17049 8789 17083 8823
rect 17509 8789 17543 8823
rect 19625 8789 19659 8823
rect 19717 8789 19751 8823
rect 21097 8789 21131 8823
rect 21925 8789 21959 8823
rect 22569 8789 22603 8823
rect 23305 8789 23339 8823
rect 23673 8789 23707 8823
rect 26249 8789 26283 8823
rect 1869 8585 1903 8619
rect 2237 8585 2271 8619
rect 2329 8585 2363 8619
rect 11805 8585 11839 8619
rect 12081 8585 12115 8619
rect 15853 8585 15887 8619
rect 16221 8585 16255 8619
rect 19073 8585 19107 8619
rect 20361 8585 20395 8619
rect 20545 8585 20579 8619
rect 23029 8585 23063 8619
rect 23213 8585 23247 8619
rect 25329 8585 25363 8619
rect 25697 8585 25731 8619
rect 4077 8517 4111 8551
rect 5365 8517 5399 8551
rect 6009 8517 6043 8551
rect 6193 8517 6227 8551
rect 9352 8517 9386 8551
rect 9689 8517 9723 8551
rect 11621 8517 11655 8551
rect 17509 8517 17543 8551
rect 17693 8517 17727 8551
rect 19533 8517 19567 8551
rect 19993 8517 20027 8551
rect 25789 8517 25823 8551
rect 3525 8449 3559 8483
rect 3835 8449 3869 8483
rect 4169 8449 4203 8483
rect 4411 8449 4445 8483
rect 5825 8449 5859 8483
rect 6377 8449 6411 8483
rect 6644 8449 6678 8483
rect 9608 8449 9642 8483
rect 9873 8449 9907 8483
rect 10242 8449 10276 8483
rect 10425 8449 10459 8483
rect 10517 8449 10551 8483
rect 10682 8449 10716 8483
rect 10793 8449 10827 8483
rect 10885 8449 10919 8483
rect 11069 8449 11103 8483
rect 11529 8449 11563 8483
rect 12265 8449 12299 8483
rect 12357 8449 12391 8483
rect 12909 8449 12943 8483
rect 17233 8449 17267 8483
rect 17325 8449 17359 8483
rect 19441 8449 19475 8483
rect 20177 8449 20211 8483
rect 20729 8449 20763 8483
rect 20821 8449 20855 8483
rect 21097 8449 21131 8483
rect 21649 8449 21683 8483
rect 22385 8449 22419 8483
rect 22661 8449 22695 8483
rect 23305 8449 23339 8483
rect 23561 8449 23595 8483
rect 27905 8449 27939 8483
rect 28089 8449 28123 8483
rect 28273 8449 28307 8483
rect 28641 8449 28675 8483
rect 2421 8381 2455 8415
rect 3433 8381 3467 8415
rect 4701 8381 4735 8415
rect 4813 8381 4847 8415
rect 5457 8381 5491 8415
rect 5641 8381 5675 8415
rect 10057 8381 10091 8415
rect 10149 8381 10183 8415
rect 12541 8381 12575 8415
rect 12633 8381 12667 8415
rect 15669 8381 15703 8415
rect 15761 8381 15795 8415
rect 17141 8381 17175 8415
rect 19625 8381 19659 8415
rect 25881 8381 25915 8415
rect 29009 8381 29043 8415
rect 8217 8313 8251 8347
rect 11253 8313 11287 8347
rect 12817 8313 12851 8347
rect 21005 8313 21039 8347
rect 22753 8313 22787 8347
rect 24685 8313 24719 8347
rect 4997 8245 5031 8279
rect 7757 8245 7791 8279
rect 16865 8245 16899 8279
rect 17233 8245 17267 8279
rect 21557 8245 21591 8279
rect 22569 8245 22603 8279
rect 28457 8245 28491 8279
rect 3801 8041 3835 8075
rect 4169 8041 4203 8075
rect 5089 8041 5123 8075
rect 6745 8041 6779 8075
rect 9413 8041 9447 8075
rect 17601 8041 17635 8075
rect 21833 8041 21867 8075
rect 22937 8041 22971 8075
rect 23949 8041 23983 8075
rect 2605 7973 2639 8007
rect 26065 7973 26099 8007
rect 28825 7973 28859 8007
rect 2237 7905 2271 7939
rect 5549 7905 5583 7939
rect 5641 7905 5675 7939
rect 7297 7905 7331 7939
rect 17693 7905 17727 7939
rect 25053 7905 25087 7939
rect 27353 7905 27387 7939
rect 28457 7905 28491 7939
rect 28549 7905 28583 7939
rect 3801 7837 3835 7871
rect 3985 7837 4019 7871
rect 4721 7837 4755 7871
rect 5239 7837 5273 7871
rect 7757 7837 7791 7871
rect 8033 7837 8067 7871
rect 9505 7837 9539 7871
rect 11354 7837 11388 7871
rect 11621 7837 11655 7871
rect 17601 7837 17635 7871
rect 19073 7837 19107 7871
rect 20913 7837 20947 7871
rect 21649 7837 21683 7871
rect 23121 7837 23155 7871
rect 23857 7837 23891 7871
rect 24133 7837 24167 7871
rect 24501 7837 24535 7871
rect 24743 7837 24777 7871
rect 25145 7837 25179 7871
rect 26249 7837 26283 7871
rect 26801 7837 26835 7871
rect 26985 7837 27019 7871
rect 27169 7837 27203 7871
rect 27721 7837 27755 7871
rect 28365 7837 28399 7871
rect 29009 7837 29043 7871
rect 4353 7769 4387 7803
rect 4537 7769 4571 7803
rect 7113 7769 7147 7803
rect 7205 7769 7239 7803
rect 21097 7769 21131 7803
rect 21281 7769 21315 7803
rect 27537 7769 27571 7803
rect 2697 7701 2731 7735
rect 7573 7701 7607 7735
rect 7849 7701 7883 7735
rect 10241 7701 10275 7735
rect 17969 7701 18003 7735
rect 18889 7701 18923 7735
rect 23305 7701 23339 7735
rect 23673 7701 23707 7735
rect 27997 7701 28031 7735
rect 2697 7497 2731 7531
rect 3157 7497 3191 7531
rect 17325 7497 17359 7531
rect 18337 7497 18371 7531
rect 22753 7497 22787 7531
rect 24593 7497 24627 7531
rect 27261 7497 27295 7531
rect 28457 7497 28491 7531
rect 1593 7429 1627 7463
rect 2789 7429 2823 7463
rect 6929 7429 6963 7463
rect 25605 7429 25639 7463
rect 25697 7429 25731 7463
rect 25881 7429 25915 7463
rect 3341 7361 3375 7395
rect 6561 7361 6595 7395
rect 6745 7361 6779 7395
rect 7205 7361 7239 7395
rect 8217 7361 8251 7395
rect 8484 7361 8518 7395
rect 14841 7361 14875 7395
rect 14933 7361 14967 7395
rect 15393 7361 15427 7395
rect 15577 7361 15611 7395
rect 15853 7361 15887 7395
rect 16037 7361 16071 7395
rect 16405 7361 16439 7395
rect 16773 7361 16807 7395
rect 17417 7361 17451 7395
rect 18797 7361 18831 7395
rect 19257 7361 19291 7395
rect 19625 7361 19659 7395
rect 19809 7361 19843 7395
rect 20085 7361 20119 7395
rect 20453 7361 20487 7395
rect 20545 7361 20579 7395
rect 21005 7361 21039 7395
rect 21373 7361 21407 7395
rect 21557 7361 21591 7395
rect 22569 7361 22603 7395
rect 22937 7361 22971 7395
rect 23193 7361 23227 7395
rect 24743 7361 24777 7395
rect 25237 7361 25271 7395
rect 25421 7361 25455 7395
rect 26065 7361 26099 7395
rect 27077 7361 27111 7395
rect 27261 7361 27295 7395
rect 27537 7361 27571 7395
rect 27721 7361 27755 7395
rect 28307 7361 28341 7395
rect 2881 7293 2915 7327
rect 15117 7293 15151 7327
rect 15669 7293 15703 7327
rect 17233 7293 17267 7327
rect 18061 7293 18095 7327
rect 18245 7293 18279 7327
rect 18981 7293 19015 7327
rect 20269 7293 20303 7327
rect 20361 7293 20395 7327
rect 21097 7293 21131 7327
rect 22385 7293 22419 7327
rect 25053 7293 25087 7327
rect 25145 7293 25179 7327
rect 27905 7293 27939 7327
rect 27997 7293 28031 7327
rect 1961 7225 1995 7259
rect 18705 7225 18739 7259
rect 19441 7225 19475 7259
rect 21189 7225 21223 7259
rect 24317 7225 24351 7259
rect 2053 7157 2087 7191
rect 2329 7157 2363 7191
rect 7113 7157 7147 7191
rect 9597 7157 9631 7191
rect 16221 7157 16255 7191
rect 16865 7157 16899 7191
rect 17785 7157 17819 7191
rect 3801 6953 3835 6987
rect 6469 6953 6503 6987
rect 6929 6953 6963 6987
rect 8769 6953 8803 6987
rect 15761 6953 15795 6987
rect 18153 6953 18187 6987
rect 18521 6953 18555 6987
rect 19901 6953 19935 6987
rect 21373 6953 21407 6987
rect 22937 6953 22971 6987
rect 25053 6953 25087 6987
rect 26617 6953 26651 6987
rect 29101 6953 29135 6987
rect 9689 6885 9723 6919
rect 19073 6885 19107 6919
rect 2053 6817 2087 6851
rect 2237 6817 2271 6851
rect 4353 6817 4387 6851
rect 7021 6817 7055 6851
rect 8217 6817 8251 6851
rect 9781 6817 9815 6851
rect 16405 6817 16439 6851
rect 16957 6817 16991 6851
rect 18245 6817 18279 6851
rect 21925 6817 21959 6851
rect 23489 6817 23523 6851
rect 24869 6817 24903 6851
rect 26525 6817 26559 6851
rect 26709 6817 26743 6851
rect 27261 6817 27295 6851
rect 27721 6817 27755 6851
rect 2605 6749 2639 6783
rect 5917 6749 5951 6783
rect 6101 6749 6135 6783
rect 6653 6749 6687 6783
rect 6745 6749 6779 6783
rect 7297 6749 7331 6783
rect 7573 6749 7607 6783
rect 7941 6749 7975 6783
rect 9319 6749 9353 6783
rect 10701 6749 10735 6783
rect 16129 6749 16163 6783
rect 18153 6749 18187 6783
rect 20821 6749 20855 6783
rect 20913 6749 20947 6783
rect 21281 6749 21315 6783
rect 21741 6749 21775 6783
rect 22293 6749 22327 6783
rect 22477 6749 22511 6783
rect 23305 6749 23339 6783
rect 25053 6749 25087 6783
rect 26341 6749 26375 6783
rect 26893 6749 26927 6783
rect 27988 6749 28022 6783
rect 1961 6681 1995 6715
rect 4261 6681 4295 6715
rect 7849 6681 7883 6715
rect 8401 6681 8435 6715
rect 16589 6681 16623 6715
rect 16773 6681 16807 6715
rect 18705 6681 18739 6715
rect 18889 6681 18923 6715
rect 21833 6681 21867 6715
rect 22201 6681 22235 6715
rect 24777 6681 24811 6715
rect 26617 6681 26651 6715
rect 1593 6613 1627 6647
rect 2421 6613 2455 6647
rect 4169 6613 4203 6647
rect 6009 6613 6043 6647
rect 7297 6613 7331 6647
rect 8309 6613 8343 6647
rect 9137 6613 9171 6647
rect 9321 6613 9355 6647
rect 10517 6613 10551 6647
rect 16221 6613 16255 6647
rect 20637 6613 20671 6647
rect 21097 6613 21131 6647
rect 23397 6613 23431 6647
rect 25237 6613 25271 6647
rect 26157 6613 26191 6647
rect 27169 6613 27203 6647
rect 3525 6409 3559 6443
rect 6101 6409 6135 6443
rect 7021 6409 7055 6443
rect 8309 6409 8343 6443
rect 19165 6409 19199 6443
rect 26709 6409 26743 6443
rect 2973 6341 3007 6375
rect 6561 6341 6595 6375
rect 6745 6341 6779 6375
rect 17601 6341 17635 6375
rect 24685 6341 24719 6375
rect 24869 6341 24903 6375
rect 3157 6273 3191 6307
rect 3341 6273 3375 6307
rect 3433 6273 3467 6307
rect 3893 6273 3927 6307
rect 4537 6273 4571 6307
rect 4988 6273 5022 6307
rect 7205 6273 7239 6307
rect 7481 6273 7515 6307
rect 8033 6273 8067 6307
rect 8309 6273 8343 6307
rect 11078 6273 11112 6307
rect 11345 6273 11379 6307
rect 15945 6273 15979 6307
rect 17785 6273 17819 6307
rect 17969 6273 18003 6307
rect 18061 6273 18095 6307
rect 19257 6273 19291 6307
rect 21833 6273 21867 6307
rect 23581 6273 23615 6307
rect 23765 6273 23799 6307
rect 24501 6273 24535 6307
rect 25596 6273 25630 6307
rect 26985 6273 27019 6307
rect 27169 6273 27203 6307
rect 3985 6205 4019 6239
rect 4077 6205 4111 6239
rect 4721 6205 4755 6239
rect 7297 6205 7331 6239
rect 25329 6205 25363 6239
rect 6377 6137 6411 6171
rect 23489 6137 23523 6171
rect 27261 6137 27295 6171
rect 4445 6069 4479 6103
rect 7205 6069 7239 6103
rect 9965 6069 9999 6103
rect 15853 6069 15887 6103
rect 18245 6069 18279 6103
rect 22017 6069 22051 6103
rect 2789 5865 2823 5899
rect 3341 5865 3375 5899
rect 4353 5865 4387 5899
rect 5365 5865 5399 5899
rect 10977 5865 11011 5899
rect 11437 5865 11471 5899
rect 19257 5865 19291 5899
rect 23857 5865 23891 5899
rect 24961 5865 24995 5899
rect 25973 5865 26007 5899
rect 1409 5661 1443 5695
rect 1676 5661 1710 5695
rect 19717 5797 19751 5831
rect 5825 5729 5859 5763
rect 6009 5729 6043 5763
rect 9689 5729 9723 5763
rect 10057 5729 10091 5763
rect 10333 5729 10367 5763
rect 10517 5729 10551 5763
rect 15393 5729 15427 5763
rect 15577 5729 15611 5763
rect 16129 5729 16163 5763
rect 17785 5729 17819 5763
rect 18981 5729 19015 5763
rect 19349 5729 19383 5763
rect 20545 5729 20579 5763
rect 21649 5729 21683 5763
rect 26433 5729 26467 5763
rect 26617 5729 26651 5763
rect 3433 5661 3467 5695
rect 3801 5661 3835 5695
rect 4077 5661 4111 5695
rect 4221 5661 4255 5695
rect 4905 5661 4939 5695
rect 6561 5661 6595 5695
rect 7849 5661 7883 5695
rect 8125 5661 8159 5695
rect 9505 5661 9539 5695
rect 9965 5661 9999 5695
rect 11161 5661 11195 5695
rect 11253 5661 11287 5695
rect 15301 5661 15335 5695
rect 15853 5661 15887 5695
rect 16037 5661 16071 5695
rect 16313 5661 16347 5695
rect 16497 5661 16531 5695
rect 16865 5661 16899 5695
rect 17049 5661 17083 5695
rect 17325 5661 17359 5695
rect 17509 5661 17543 5695
rect 17693 5661 17727 5695
rect 17969 5661 18003 5695
rect 18153 5661 18187 5695
rect 18705 5661 18739 5695
rect 19533 5661 19567 5695
rect 20085 5661 20119 5695
rect 20177 5661 20211 5695
rect 20453 5661 20487 5695
rect 20729 5661 20763 5695
rect 20913 5661 20947 5695
rect 21465 5661 21499 5695
rect 21925 5661 21959 5695
rect 22201 5661 22235 5695
rect 22477 5661 22511 5695
rect 24685 5661 24719 5695
rect 24777 5661 24811 5695
rect 25053 5661 25087 5695
rect 25145 5661 25179 5695
rect 25421 5661 25455 5695
rect 26985 5661 27019 5695
rect 3525 5593 3559 5627
rect 3985 5593 4019 5627
rect 4537 5593 4571 5627
rect 4721 5593 4755 5627
rect 5733 5593 5767 5627
rect 6469 5593 6503 5627
rect 8217 5593 8251 5627
rect 9781 5593 9815 5627
rect 9873 5593 9907 5627
rect 16681 5593 16715 5627
rect 19257 5593 19291 5627
rect 22744 5593 22778 5627
rect 25513 5593 25547 5627
rect 26341 5593 26375 5627
rect 26893 5593 26927 5627
rect 3341 5525 3375 5559
rect 10609 5525 10643 5559
rect 14933 5525 14967 5559
rect 17141 5525 17175 5559
rect 18337 5525 18371 5559
rect 18797 5525 18831 5559
rect 19901 5525 19935 5559
rect 21097 5525 21131 5559
rect 21557 5525 21591 5559
rect 22017 5525 22051 5559
rect 22385 5525 22419 5559
rect 24501 5525 24535 5559
rect 25237 5525 25271 5559
rect 3341 5321 3375 5355
rect 8401 5321 8435 5355
rect 8861 5321 8895 5355
rect 10241 5321 10275 5355
rect 11989 5321 12023 5355
rect 12357 5321 12391 5355
rect 15761 5321 15795 5355
rect 16681 5321 16715 5355
rect 17141 5321 17175 5355
rect 17969 5321 18003 5355
rect 18797 5321 18831 5355
rect 20177 5321 20211 5355
rect 21833 5321 21867 5355
rect 22293 5321 22327 5355
rect 23029 5321 23063 5355
rect 23489 5321 23523 5355
rect 2228 5253 2262 5287
rect 6377 5253 6411 5287
rect 8064 5253 8098 5287
rect 11253 5253 11287 5287
rect 15853 5253 15887 5287
rect 16313 5253 16347 5287
rect 19349 5253 19383 5287
rect 20269 5253 20303 5287
rect 20729 5253 20763 5287
rect 21649 5253 21683 5287
rect 23397 5253 23431 5287
rect 1961 5185 1995 5219
rect 4353 5185 4387 5219
rect 4997 5185 5031 5219
rect 6561 5185 6595 5219
rect 8769 5185 8803 5219
rect 9229 5185 9263 5219
rect 9597 5185 9631 5219
rect 9781 5185 9815 5219
rect 9873 5185 9907 5219
rect 10885 5185 10919 5219
rect 11069 5185 11103 5219
rect 11897 5185 11931 5219
rect 12541 5185 12575 5219
rect 16221 5185 16255 5219
rect 17049 5185 17083 5219
rect 18429 5185 18463 5219
rect 18613 5185 18647 5219
rect 20821 5185 20855 5219
rect 21281 5185 21315 5219
rect 21465 5185 21499 5219
rect 22201 5185 22235 5219
rect 25421 5185 25455 5219
rect 25697 5185 25731 5219
rect 26065 5185 26099 5219
rect 4537 5117 4571 5151
rect 8309 5117 8343 5151
rect 8953 5117 8987 5151
rect 9965 5117 9999 5151
rect 12081 5117 12115 5151
rect 16037 5117 16071 5151
rect 17325 5117 17359 5151
rect 18061 5117 18095 5151
rect 18245 5117 18279 5151
rect 19441 5117 19475 5151
rect 19625 5117 19659 5151
rect 20453 5117 20487 5151
rect 22385 5117 22419 5151
rect 23581 5117 23615 5151
rect 4813 5049 4847 5083
rect 9321 5049 9355 5083
rect 25697 5049 25731 5083
rect 4169 4981 4203 5015
rect 6653 4981 6687 5015
rect 6929 4981 6963 5015
rect 9873 4981 9907 5015
rect 11529 4981 11563 5015
rect 15393 4981 15427 5015
rect 17601 4981 17635 5015
rect 18429 4981 18463 5015
rect 18981 4981 19015 5015
rect 19809 4981 19843 5015
rect 25973 4981 26007 5015
rect 5733 4777 5767 4811
rect 6745 4777 6779 4811
rect 6929 4777 6963 4811
rect 8217 4777 8251 4811
rect 10609 4777 10643 4811
rect 11069 4777 11103 4811
rect 18061 4777 18095 4811
rect 21189 4777 21223 4811
rect 21833 4777 21867 4811
rect 28181 4777 28215 4811
rect 5457 4709 5491 4743
rect 6285 4641 6319 4675
rect 6561 4641 6595 4675
rect 9321 4641 9355 4675
rect 12909 4641 12943 4675
rect 22385 4641 22419 4675
rect 25237 4641 25271 4675
rect 25973 4641 26007 4675
rect 3801 4573 3835 4607
rect 4077 4573 4111 4607
rect 5883 4573 5917 4607
rect 6193 4573 6227 4607
rect 6745 4573 6779 4607
rect 8125 4573 8159 4607
rect 8953 4573 8987 4607
rect 9229 4573 9263 4607
rect 10425 4573 10459 4607
rect 10609 4573 10643 4607
rect 10885 4573 10919 4607
rect 12642 4573 12676 4607
rect 15945 4573 15979 4607
rect 18153 4573 18187 4607
rect 21373 4573 21407 4607
rect 23949 4573 23983 4607
rect 24409 4573 24443 4607
rect 24777 4573 24811 4607
rect 25053 4573 25087 4607
rect 25421 4573 25455 4607
rect 25513 4573 25547 4607
rect 27629 4573 27663 4607
rect 27905 4573 27939 4607
rect 28017 4573 28051 4607
rect 4344 4505 4378 4539
rect 6469 4505 6503 4539
rect 22201 4505 22235 4539
rect 23765 4505 23799 4539
rect 24133 4505 24167 4539
rect 24593 4505 24627 4539
rect 26218 4505 26252 4539
rect 27537 4505 27571 4539
rect 3985 4437 4019 4471
rect 10241 4437 10275 4471
rect 11529 4437 11563 4471
rect 16037 4437 16071 4471
rect 22293 4437 22327 4471
rect 24869 4437 24903 4471
rect 25881 4437 25915 4471
rect 27353 4437 27387 4471
rect 4445 4233 4479 4267
rect 10517 4233 10551 4267
rect 15669 4233 15703 4267
rect 16773 4233 16807 4267
rect 18613 4233 18647 4267
rect 21925 4233 21959 4267
rect 25881 4233 25915 4267
rect 8401 4165 8435 4199
rect 16405 4165 16439 4199
rect 17141 4165 17175 4199
rect 18245 4165 18279 4199
rect 19708 4165 19742 4199
rect 22477 4165 22511 4199
rect 1869 4097 1903 4131
rect 4537 4097 4571 4131
rect 6377 4097 6411 4131
rect 6561 4097 6595 4131
rect 8217 4097 8251 4131
rect 8585 4097 8619 4131
rect 9414 4097 9448 4131
rect 9873 4097 9907 4131
rect 10610 4097 10644 4131
rect 10977 4097 11011 4131
rect 14289 4097 14323 4131
rect 14556 4097 14590 4131
rect 16221 4097 16255 4131
rect 22201 4097 22235 4131
rect 22569 4097 22603 4131
rect 22937 4097 22971 4131
rect 23213 4097 23247 4131
rect 23480 4097 23514 4131
rect 25789 4097 25823 4131
rect 26065 4097 26099 4131
rect 4721 4029 4755 4063
rect 9781 4029 9815 4063
rect 11069 4029 11103 4063
rect 17233 4029 17267 4063
rect 17325 4029 17359 4063
rect 17969 4029 18003 4063
rect 18153 4029 18187 4063
rect 19441 4029 19475 4063
rect 22089 4029 22123 4063
rect 4077 3961 4111 3995
rect 20821 3961 20855 3995
rect 24593 3961 24627 3995
rect 6377 3893 6411 3927
rect 6745 3893 6779 3927
rect 9321 3893 9355 3927
rect 16129 3893 16163 3927
rect 23121 3893 23155 3927
rect 9873 3689 9907 3723
rect 10333 3689 10367 3723
rect 17785 3689 17819 3723
rect 18889 3689 18923 3723
rect 19625 3689 19659 3723
rect 22201 3689 22235 3723
rect 23489 3689 23523 3723
rect 8585 3621 8619 3655
rect 18521 3621 18555 3655
rect 4813 3553 4847 3587
rect 6101 3553 6135 3587
rect 8125 3553 8159 3587
rect 10149 3553 10183 3587
rect 11805 3553 11839 3587
rect 15945 3553 15979 3587
rect 17233 3553 17267 3587
rect 17417 3553 17451 3587
rect 18245 3553 18279 3587
rect 18337 3553 18371 3587
rect 20269 3553 20303 3587
rect 20545 3553 20579 3587
rect 22569 3553 22603 3587
rect 22845 3553 22879 3587
rect 23949 3553 23983 3587
rect 24041 3553 24075 3587
rect 4629 3485 4663 3519
rect 5699 3485 5733 3519
rect 6009 3485 6043 3519
rect 6745 3485 6779 3519
rect 6929 3485 6963 3519
rect 7205 3485 7239 3519
rect 7481 3485 7515 3519
rect 7723 3485 7757 3519
rect 8033 3485 8067 3519
rect 8217 3485 8251 3519
rect 8401 3485 8435 3519
rect 9229 3485 9263 3519
rect 9413 3485 9447 3519
rect 9689 3485 9723 3519
rect 10057 3485 10091 3519
rect 10943 3485 10977 3519
rect 11253 3485 11287 3519
rect 11345 3485 11379 3519
rect 11437 3485 11471 3519
rect 11897 3485 11931 3519
rect 16221 3485 16255 3519
rect 16681 3485 16715 3519
rect 16865 3485 16899 3519
rect 17325 3485 17359 3519
rect 18041 3485 18075 3519
rect 18428 3485 18462 3519
rect 18705 3485 18739 3519
rect 19257 3485 19291 3519
rect 20812 3485 20846 3519
rect 22385 3485 22419 3519
rect 22661 3485 22695 3519
rect 22753 3485 22787 3519
rect 23857 3485 23891 3519
rect 29653 3485 29687 3519
rect 10333 3417 10367 3451
rect 11621 3417 11655 3451
rect 16129 3417 16163 3451
rect 17785 3417 17819 3451
rect 19349 3417 19383 3451
rect 19993 3417 20027 3451
rect 4445 3349 4479 3383
rect 5549 3349 5583 3383
rect 6561 3349 6595 3383
rect 7021 3349 7055 3383
rect 9045 3349 9079 3383
rect 9505 3349 9539 3383
rect 10793 3349 10827 3383
rect 12081 3349 12115 3383
rect 16589 3349 16623 3383
rect 16865 3349 16899 3383
rect 18153 3349 18187 3383
rect 20085 3349 20119 3383
rect 21925 3349 21959 3383
rect 5733 3145 5767 3179
rect 7757 3145 7791 3179
rect 9965 3145 9999 3179
rect 11253 3145 11287 3179
rect 18613 3145 18647 3179
rect 20177 3145 20211 3179
rect 22385 3145 22419 3179
rect 20453 3077 20487 3111
rect 20821 3077 20855 3111
rect 20913 3077 20947 3111
rect 21005 3077 21039 3111
rect 21833 3077 21867 3111
rect 22017 3077 22051 3111
rect 3893 3009 3927 3043
rect 4436 3009 4470 3043
rect 5917 3009 5951 3043
rect 6009 3009 6043 3043
rect 6377 3009 6411 3043
rect 6633 3009 6667 3043
rect 8309 3009 8343 3043
rect 8585 3009 8619 3043
rect 8852 3009 8886 3043
rect 10609 3009 10643 3043
rect 11069 3009 11103 3043
rect 12734 3009 12768 3043
rect 13001 3009 13035 3043
rect 15025 3009 15059 3043
rect 15292 3009 15326 3043
rect 16681 3009 16715 3043
rect 16865 3009 16899 3043
rect 17049 3009 17083 3043
rect 17233 3009 17267 3043
rect 17500 3009 17534 3043
rect 18797 3009 18831 3043
rect 19064 3009 19098 3043
rect 20637 3009 20671 3043
rect 21189 3009 21223 3043
rect 21373 3009 21407 3043
rect 22201 3009 22235 3043
rect 22293 3009 22327 3043
rect 4169 2941 4203 2975
rect 10885 2941 10919 2975
rect 5549 2873 5583 2907
rect 10793 2873 10827 2907
rect 16405 2873 16439 2907
rect 4077 2805 4111 2839
rect 6193 2805 6227 2839
rect 8493 2805 8527 2839
rect 11621 2805 11655 2839
rect 4353 2601 4387 2635
rect 6469 2601 6503 2635
rect 8953 2601 8987 2635
rect 11529 2601 11563 2635
rect 17049 2601 17083 2635
rect 4813 2465 4847 2499
rect 4997 2465 5031 2499
rect 6929 2465 6963 2499
rect 7113 2465 7147 2499
rect 9413 2465 9447 2499
rect 9597 2465 9631 2499
rect 11989 2465 12023 2499
rect 12081 2465 12115 2499
rect 4721 2397 4755 2431
rect 6837 2397 6871 2431
rect 9321 2397 9355 2431
rect 11897 2397 11931 2431
rect 16957 2397 16991 2431
<< metal1 >>
rect 11146 30676 11152 30728
rect 11204 30716 11210 30728
rect 11606 30716 11612 30728
rect 11204 30688 11612 30716
rect 11204 30676 11210 30688
rect 11606 30676 11612 30688
rect 11664 30676 11670 30728
rect 3878 30608 3884 30660
rect 3936 30648 3942 30660
rect 13906 30648 13912 30660
rect 3936 30620 13912 30648
rect 3936 30608 3942 30620
rect 13906 30608 13912 30620
rect 13964 30608 13970 30660
rect 15286 30608 15292 30660
rect 15344 30648 15350 30660
rect 16022 30648 16028 30660
rect 15344 30620 16028 30648
rect 15344 30608 15350 30620
rect 16022 30608 16028 30620
rect 16080 30608 16086 30660
rect 10778 30540 10784 30592
rect 10836 30580 10842 30592
rect 16482 30580 16488 30592
rect 10836 30552 16488 30580
rect 10836 30540 10842 30552
rect 16482 30540 16488 30552
rect 16540 30540 16546 30592
rect 1104 30490 29532 30512
rect 1104 30438 10425 30490
rect 10477 30438 10489 30490
rect 10541 30438 10553 30490
rect 10605 30438 10617 30490
rect 10669 30438 10681 30490
rect 10733 30438 19901 30490
rect 19953 30438 19965 30490
rect 20017 30438 20029 30490
rect 20081 30438 20093 30490
rect 20145 30438 20157 30490
rect 20209 30438 29532 30490
rect 1104 30416 29532 30438
rect 4062 30336 4068 30388
rect 4120 30376 4126 30388
rect 4120 30348 14320 30376
rect 4120 30336 4126 30348
rect 10321 30311 10379 30317
rect 10321 30308 10333 30311
rect 9986 30280 10333 30308
rect 9986 30252 10014 30280
rect 10321 30277 10333 30280
rect 10367 30308 10379 30311
rect 10778 30308 10784 30320
rect 10367 30280 10784 30308
rect 10367 30277 10379 30280
rect 10321 30271 10379 30277
rect 10778 30268 10784 30280
rect 10836 30268 10842 30320
rect 14292 30317 14320 30348
rect 14277 30311 14335 30317
rect 14277 30277 14289 30311
rect 14323 30308 14335 30311
rect 14323 30280 14596 30308
rect 14323 30277 14335 30280
rect 14277 30271 14335 30277
rect 9030 30200 9036 30252
rect 9088 30240 9094 30252
rect 9585 30243 9643 30249
rect 9585 30240 9597 30243
rect 9088 30212 9597 30240
rect 9088 30200 9094 30212
rect 9585 30209 9597 30212
rect 9631 30209 9643 30243
rect 9585 30203 9643 30209
rect 9971 30246 10029 30252
rect 9971 30212 9983 30246
rect 10017 30212 10029 30246
rect 9971 30206 10029 30212
rect 10134 30200 10140 30252
rect 10192 30240 10198 30252
rect 11698 30240 11704 30252
rect 10192 30212 10237 30240
rect 11659 30212 11704 30240
rect 10192 30200 10198 30212
rect 11698 30200 11704 30212
rect 11756 30200 11762 30252
rect 12070 30243 12128 30249
rect 12070 30240 12082 30243
rect 11808 30212 12082 30240
rect 9674 30132 9680 30184
rect 9732 30172 9738 30184
rect 9769 30175 9827 30181
rect 9769 30172 9781 30175
rect 9732 30144 9781 30172
rect 9732 30132 9738 30144
rect 9769 30141 9781 30144
rect 9815 30141 9827 30175
rect 9769 30135 9827 30141
rect 9858 30132 9864 30184
rect 9916 30172 9922 30184
rect 11808 30172 11836 30212
rect 12070 30209 12082 30212
rect 12116 30209 12128 30243
rect 12070 30203 12128 30209
rect 12253 30243 12311 30249
rect 12253 30209 12265 30243
rect 12299 30240 12311 30243
rect 12526 30240 12532 30252
rect 12299 30212 12532 30240
rect 12299 30209 12311 30212
rect 12253 30203 12311 30209
rect 12526 30200 12532 30212
rect 12584 30240 12590 30252
rect 13262 30240 13268 30252
rect 12584 30212 13268 30240
rect 12584 30200 12590 30212
rect 13262 30200 13268 30212
rect 13320 30200 13326 30252
rect 14458 30240 14464 30252
rect 14419 30212 14464 30240
rect 14458 30200 14464 30212
rect 14516 30200 14522 30252
rect 14568 30240 14596 30280
rect 14752 30280 15148 30308
rect 14752 30252 14780 30280
rect 14626 30243 14684 30249
rect 14626 30240 14638 30243
rect 14568 30212 14638 30240
rect 14626 30209 14638 30212
rect 14672 30209 14684 30243
rect 14626 30203 14684 30209
rect 14734 30200 14740 30252
rect 14792 30240 14798 30252
rect 15010 30240 15016 30252
rect 14792 30212 14885 30240
rect 14971 30212 15016 30240
rect 14792 30200 14798 30212
rect 15010 30200 15016 30212
rect 15068 30200 15074 30252
rect 9916 30144 9961 30172
rect 11256 30144 11836 30172
rect 11885 30175 11943 30181
rect 9916 30132 9922 30144
rect 4062 30064 4068 30116
rect 4120 30104 4126 30116
rect 11256 30113 11284 30144
rect 11885 30141 11897 30175
rect 11931 30141 11943 30175
rect 11885 30135 11943 30141
rect 11241 30107 11299 30113
rect 11241 30104 11253 30107
rect 4120 30076 11253 30104
rect 4120 30064 4126 30076
rect 11241 30073 11253 30076
rect 11287 30073 11299 30107
rect 11900 30104 11928 30135
rect 11974 30132 11980 30184
rect 12032 30172 12038 30184
rect 14826 30172 14832 30184
rect 12032 30144 12077 30172
rect 14787 30144 14832 30172
rect 12032 30132 12038 30144
rect 14826 30132 14832 30144
rect 14884 30132 14890 30184
rect 15120 30172 15148 30280
rect 17420 30280 17908 30308
rect 16942 30240 16948 30252
rect 16903 30212 16948 30240
rect 16942 30200 16948 30212
rect 17000 30200 17006 30252
rect 17128 30243 17186 30249
rect 17128 30209 17140 30243
rect 17174 30240 17186 30243
rect 17420 30240 17448 30280
rect 17174 30212 17448 30240
rect 17497 30243 17555 30249
rect 17174 30209 17186 30212
rect 17128 30203 17186 30209
rect 17497 30209 17509 30243
rect 17543 30240 17555 30243
rect 17586 30240 17592 30252
rect 17543 30212 17592 30240
rect 17543 30209 17555 30212
rect 17497 30203 17555 30209
rect 17586 30200 17592 30212
rect 17644 30200 17650 30252
rect 17880 30249 17908 30280
rect 17865 30243 17923 30249
rect 17865 30209 17877 30243
rect 17911 30240 17923 30243
rect 27522 30240 27528 30252
rect 17911 30212 27528 30240
rect 17911 30209 17923 30212
rect 17865 30203 17923 30209
rect 27522 30200 27528 30212
rect 27580 30200 27586 30252
rect 17221 30175 17279 30181
rect 17221 30172 17233 30175
rect 15120 30144 17233 30172
rect 17221 30141 17233 30144
rect 17267 30141 17279 30175
rect 17221 30135 17279 30141
rect 17313 30175 17371 30181
rect 17313 30141 17325 30175
rect 17359 30141 17371 30175
rect 17313 30135 17371 30141
rect 12894 30104 12900 30116
rect 11900 30076 12900 30104
rect 11241 30067 11299 30073
rect 12894 30064 12900 30076
rect 12952 30064 12958 30116
rect 17126 30064 17132 30116
rect 17184 30104 17190 30116
rect 17236 30104 17264 30135
rect 17184 30076 17264 30104
rect 17184 30064 17190 30076
rect 9490 30036 9496 30048
rect 9451 30008 9496 30036
rect 9490 29996 9496 30008
rect 9548 29996 9554 30048
rect 11606 30036 11612 30048
rect 11567 30008 11612 30036
rect 11606 29996 11612 30008
rect 11664 29996 11670 30048
rect 15105 30039 15163 30045
rect 15105 30005 15117 30039
rect 15151 30036 15163 30039
rect 16114 30036 16120 30048
rect 15151 30008 16120 30036
rect 15151 30005 15163 30008
rect 15105 29999 15163 30005
rect 16114 29996 16120 30008
rect 16172 29996 16178 30048
rect 17034 29996 17040 30048
rect 17092 30036 17098 30048
rect 17328 30036 17356 30135
rect 17092 30008 17356 30036
rect 17589 30039 17647 30045
rect 17092 29996 17098 30008
rect 17589 30005 17601 30039
rect 17635 30036 17647 30039
rect 17678 30036 17684 30048
rect 17635 30008 17684 30036
rect 17635 30005 17647 30008
rect 17589 29999 17647 30005
rect 17678 29996 17684 30008
rect 17736 29996 17742 30048
rect 1104 29946 29532 29968
rect 1104 29894 5688 29946
rect 5740 29894 5752 29946
rect 5804 29894 5816 29946
rect 5868 29894 5880 29946
rect 5932 29894 5944 29946
rect 5996 29894 15163 29946
rect 15215 29894 15227 29946
rect 15279 29894 15291 29946
rect 15343 29894 15355 29946
rect 15407 29894 15419 29946
rect 15471 29894 24639 29946
rect 24691 29894 24703 29946
rect 24755 29894 24767 29946
rect 24819 29894 24831 29946
rect 24883 29894 24895 29946
rect 24947 29894 29532 29946
rect 1104 29872 29532 29894
rect 14826 29792 14832 29844
rect 14884 29832 14890 29844
rect 17034 29832 17040 29844
rect 14884 29804 17040 29832
rect 14884 29792 14890 29804
rect 17034 29792 17040 29804
rect 17092 29792 17098 29844
rect 17586 29764 17592 29776
rect 17547 29736 17592 29764
rect 17586 29724 17592 29736
rect 17644 29724 17650 29776
rect 2958 29696 2964 29708
rect 2919 29668 2964 29696
rect 2958 29656 2964 29668
rect 3016 29656 3022 29708
rect 4246 29696 4252 29708
rect 4207 29668 4252 29696
rect 4246 29656 4252 29668
rect 4304 29656 4310 29708
rect 6638 29696 6644 29708
rect 6599 29668 6644 29696
rect 6638 29656 6644 29668
rect 6696 29656 6702 29708
rect 11974 29656 11980 29708
rect 12032 29696 12038 29708
rect 12989 29699 13047 29705
rect 12989 29696 13001 29699
rect 12032 29668 13001 29696
rect 12032 29656 12038 29668
rect 12989 29665 13001 29668
rect 13035 29665 13047 29699
rect 12989 29659 13047 29665
rect 13188 29668 13492 29696
rect 6362 29588 6368 29640
rect 6420 29628 6426 29640
rect 7101 29631 7159 29637
rect 7101 29628 7113 29631
rect 6420 29600 7113 29628
rect 6420 29588 6426 29600
rect 7101 29597 7113 29600
rect 7147 29597 7159 29631
rect 7101 29591 7159 29597
rect 9582 29588 9588 29640
rect 9640 29628 9646 29640
rect 10413 29631 10471 29637
rect 10413 29628 10425 29631
rect 9640 29600 10425 29628
rect 9640 29588 9646 29600
rect 10413 29597 10425 29600
rect 10459 29628 10471 29631
rect 10965 29631 11023 29637
rect 10965 29628 10977 29631
rect 10459 29600 10977 29628
rect 10459 29597 10471 29600
rect 10413 29591 10471 29597
rect 10965 29597 10977 29600
rect 11011 29628 11023 29631
rect 11514 29628 11520 29640
rect 11011 29600 11520 29628
rect 11011 29597 11023 29600
rect 10965 29591 11023 29597
rect 11514 29588 11520 29600
rect 11572 29588 11578 29640
rect 12713 29631 12771 29637
rect 12713 29597 12725 29631
rect 12759 29597 12771 29631
rect 12894 29628 12900 29640
rect 12855 29600 12900 29628
rect 12713 29591 12771 29597
rect 7368 29563 7426 29569
rect 7368 29529 7380 29563
rect 7414 29560 7426 29563
rect 8018 29560 8024 29572
rect 7414 29532 8024 29560
rect 7414 29529 7426 29532
rect 7368 29523 7426 29529
rect 8018 29520 8024 29532
rect 8076 29520 8082 29572
rect 9490 29520 9496 29572
rect 9548 29560 9554 29572
rect 10146 29563 10204 29569
rect 10146 29560 10158 29563
rect 9548 29532 10158 29560
rect 9548 29520 9554 29532
rect 10146 29529 10158 29532
rect 10192 29529 10204 29563
rect 10146 29523 10204 29529
rect 11232 29563 11290 29569
rect 11232 29529 11244 29563
rect 11278 29560 11290 29563
rect 11606 29560 11612 29572
rect 11278 29532 11612 29560
rect 11278 29529 11290 29532
rect 11232 29523 11290 29529
rect 11606 29520 11612 29532
rect 11664 29520 11670 29572
rect 12728 29560 12756 29591
rect 12894 29588 12900 29600
rect 12952 29588 12958 29640
rect 13099 29631 13157 29637
rect 13099 29597 13111 29631
rect 13145 29628 13157 29631
rect 13188 29628 13216 29668
rect 13145 29600 13216 29628
rect 13145 29597 13157 29600
rect 13099 29591 13157 29597
rect 13262 29588 13268 29640
rect 13320 29628 13326 29640
rect 13464 29637 13492 29668
rect 13449 29631 13507 29637
rect 13320 29600 13365 29628
rect 13320 29588 13326 29600
rect 13449 29597 13461 29631
rect 13495 29628 13507 29631
rect 15565 29631 15623 29637
rect 13495 29600 15516 29628
rect 13495 29597 13507 29600
rect 13449 29591 13507 29597
rect 13630 29560 13636 29572
rect 12728 29532 13636 29560
rect 13630 29520 13636 29532
rect 13688 29520 13694 29572
rect 14274 29520 14280 29572
rect 14332 29560 14338 29572
rect 15298 29563 15356 29569
rect 15298 29560 15310 29563
rect 14332 29532 15310 29560
rect 14332 29520 14338 29532
rect 15298 29529 15310 29532
rect 15344 29529 15356 29563
rect 15488 29560 15516 29600
rect 15565 29597 15577 29631
rect 15611 29628 15623 29631
rect 17405 29631 17463 29637
rect 17405 29628 17417 29631
rect 15611 29600 17417 29628
rect 15611 29597 15623 29600
rect 15565 29591 15623 29597
rect 16500 29572 16528 29600
rect 17405 29597 17417 29600
rect 17451 29628 17463 29631
rect 18969 29631 19027 29637
rect 18969 29628 18981 29631
rect 17451 29600 18981 29628
rect 17451 29597 17463 29600
rect 17405 29591 17463 29597
rect 18969 29597 18981 29600
rect 19015 29597 19027 29631
rect 18969 29591 19027 29597
rect 15488 29532 16160 29560
rect 15298 29523 15356 29529
rect 8294 29452 8300 29504
rect 8352 29492 8358 29504
rect 8481 29495 8539 29501
rect 8481 29492 8493 29495
rect 8352 29464 8493 29492
rect 8352 29452 8358 29464
rect 8481 29461 8493 29464
rect 8527 29461 8539 29495
rect 9030 29492 9036 29504
rect 8991 29464 9036 29492
rect 8481 29455 8539 29461
rect 9030 29452 9036 29464
rect 9088 29452 9094 29504
rect 11698 29452 11704 29504
rect 11756 29492 11762 29504
rect 12158 29492 12164 29504
rect 11756 29464 12164 29492
rect 11756 29452 11762 29464
rect 12158 29452 12164 29464
rect 12216 29492 12222 29504
rect 12345 29495 12403 29501
rect 12345 29492 12357 29495
rect 12216 29464 12357 29492
rect 12216 29452 12222 29464
rect 12345 29461 12357 29464
rect 12391 29461 12403 29495
rect 12618 29492 12624 29504
rect 12579 29464 12624 29492
rect 12345 29455 12403 29461
rect 12618 29452 12624 29464
rect 12676 29452 12682 29504
rect 14185 29495 14243 29501
rect 14185 29461 14197 29495
rect 14231 29492 14243 29495
rect 14366 29492 14372 29504
rect 14231 29464 14372 29492
rect 14231 29461 14243 29464
rect 14185 29455 14243 29461
rect 14366 29452 14372 29464
rect 14424 29452 14430 29504
rect 15654 29452 15660 29504
rect 15712 29492 15718 29504
rect 16025 29495 16083 29501
rect 16025 29492 16037 29495
rect 15712 29464 16037 29492
rect 15712 29452 15718 29464
rect 16025 29461 16037 29464
rect 16071 29461 16083 29495
rect 16132 29492 16160 29532
rect 16482 29520 16488 29572
rect 16540 29520 16546 29572
rect 16758 29520 16764 29572
rect 16816 29560 16822 29572
rect 17138 29563 17196 29569
rect 17138 29560 17150 29563
rect 16816 29532 17150 29560
rect 16816 29520 16822 29532
rect 17138 29529 17150 29532
rect 17184 29529 17196 29563
rect 17138 29523 17196 29529
rect 17236 29532 17632 29560
rect 17236 29492 17264 29532
rect 16132 29464 17264 29492
rect 17604 29492 17632 29532
rect 17678 29520 17684 29572
rect 17736 29560 17742 29572
rect 18702 29563 18760 29569
rect 18702 29560 18714 29563
rect 17736 29532 18714 29560
rect 17736 29520 17742 29532
rect 18702 29529 18714 29532
rect 18748 29529 18760 29563
rect 18702 29523 18760 29529
rect 21450 29492 21456 29504
rect 17604 29464 21456 29492
rect 16025 29455 16083 29461
rect 21450 29452 21456 29464
rect 21508 29452 21514 29504
rect 1104 29402 29532 29424
rect 1104 29350 10425 29402
rect 10477 29350 10489 29402
rect 10541 29350 10553 29402
rect 10605 29350 10617 29402
rect 10669 29350 10681 29402
rect 10733 29350 19901 29402
rect 19953 29350 19965 29402
rect 20017 29350 20029 29402
rect 20081 29350 20093 29402
rect 20145 29350 20157 29402
rect 20209 29350 29532 29402
rect 1104 29328 29532 29350
rect 8018 29288 8024 29300
rect 7979 29260 8024 29288
rect 8018 29248 8024 29260
rect 8076 29248 8082 29300
rect 9493 29291 9551 29297
rect 9493 29257 9505 29291
rect 9539 29288 9551 29291
rect 13630 29288 13636 29300
rect 9539 29260 11192 29288
rect 13591 29260 13636 29288
rect 9539 29257 9551 29260
rect 9493 29251 9551 29257
rect 8294 29220 8300 29232
rect 8128 29192 8300 29220
rect 8128 29161 8156 29192
rect 8294 29180 8300 29192
rect 8352 29180 8358 29232
rect 9858 29220 9864 29232
rect 8588 29192 9864 29220
rect 8113 29155 8171 29161
rect 8113 29121 8125 29155
rect 8159 29121 8171 29155
rect 8482 29155 8540 29161
rect 8482 29152 8494 29155
rect 8113 29115 8171 29121
rect 8220 29124 8494 29152
rect 7558 28976 7564 29028
rect 7616 29016 7622 29028
rect 7745 29019 7803 29025
rect 7745 29016 7757 29019
rect 7616 28988 7757 29016
rect 7616 28976 7622 28988
rect 7745 28985 7757 28988
rect 7791 29016 7803 29019
rect 8220 29016 8248 29124
rect 8482 29121 8494 29124
rect 8528 29121 8540 29155
rect 8482 29115 8540 29121
rect 8297 29087 8355 29093
rect 8297 29053 8309 29087
rect 8343 29053 8355 29087
rect 8297 29047 8355 29053
rect 8389 29087 8447 29093
rect 8389 29053 8401 29087
rect 8435 29084 8447 29087
rect 8588 29084 8616 29192
rect 9858 29180 9864 29192
rect 9916 29220 9922 29232
rect 10226 29220 10232 29232
rect 9916 29192 10232 29220
rect 9916 29180 9922 29192
rect 10226 29180 10232 29192
rect 10284 29180 10290 29232
rect 8665 29155 8723 29161
rect 8665 29121 8677 29155
rect 8711 29152 8723 29155
rect 9766 29152 9772 29164
rect 8711 29124 9772 29152
rect 8711 29121 8723 29124
rect 8665 29115 8723 29121
rect 9766 29112 9772 29124
rect 9824 29112 9830 29164
rect 9950 29161 9956 29164
rect 9944 29115 9956 29161
rect 10008 29152 10014 29164
rect 10008 29124 10044 29152
rect 9950 29112 9956 29115
rect 10008 29112 10014 29124
rect 8435 29056 8616 29084
rect 8435 29053 8447 29056
rect 8389 29047 8447 29053
rect 7791 28988 8248 29016
rect 8312 29016 8340 29047
rect 8754 29044 8760 29096
rect 8812 29084 8818 29096
rect 9582 29084 9588 29096
rect 8812 29056 9588 29084
rect 8812 29044 8818 29056
rect 9582 29044 9588 29056
rect 9640 29084 9646 29096
rect 9677 29087 9735 29093
rect 9677 29084 9689 29087
rect 9640 29056 9689 29084
rect 9640 29044 9646 29056
rect 9677 29053 9689 29056
rect 9723 29053 9735 29087
rect 9677 29047 9735 29053
rect 8312 28988 9720 29016
rect 7791 28985 7803 28988
rect 7745 28979 7803 28985
rect 9692 28960 9720 28988
rect 566 28908 572 28960
rect 624 28948 630 28960
rect 1302 28948 1308 28960
rect 624 28920 1308 28948
rect 624 28908 630 28920
rect 1302 28908 1308 28920
rect 1360 28908 1366 28960
rect 6454 28908 6460 28960
rect 6512 28948 6518 28960
rect 9493 28951 9551 28957
rect 9493 28948 9505 28951
rect 6512 28920 9505 28948
rect 6512 28908 6518 28920
rect 9493 28917 9505 28920
rect 9539 28917 9551 28951
rect 9674 28948 9680 28960
rect 9587 28920 9680 28948
rect 9493 28911 9551 28917
rect 9674 28908 9680 28920
rect 9732 28948 9738 28960
rect 10042 28948 10048 28960
rect 9732 28920 10048 28948
rect 9732 28908 9738 28920
rect 10042 28908 10048 28920
rect 10100 28908 10106 28960
rect 11054 28948 11060 28960
rect 11015 28920 11060 28948
rect 11054 28908 11060 28920
rect 11112 28908 11118 28960
rect 11164 28948 11192 29260
rect 13630 29248 13636 29260
rect 13688 29248 13694 29300
rect 13906 29288 13912 29300
rect 13867 29260 13912 29288
rect 13906 29248 13912 29260
rect 13964 29248 13970 29300
rect 14185 29291 14243 29297
rect 14185 29257 14197 29291
rect 14231 29288 14243 29291
rect 14274 29288 14280 29300
rect 14231 29260 14280 29288
rect 14231 29257 14243 29260
rect 14185 29251 14243 29257
rect 14274 29248 14280 29260
rect 14332 29248 14338 29300
rect 16758 29288 16764 29300
rect 16719 29260 16764 29288
rect 16758 29248 16764 29260
rect 16816 29248 16822 29300
rect 17402 29288 17408 29300
rect 17328 29260 17408 29288
rect 12520 29223 12578 29229
rect 12520 29189 12532 29223
rect 12566 29220 12578 29223
rect 12618 29220 12624 29232
rect 12566 29192 12624 29220
rect 12566 29189 12578 29192
rect 12520 29183 12578 29189
rect 12618 29180 12624 29192
rect 12676 29180 12682 29232
rect 13924 29220 13952 29248
rect 13924 29192 14504 29220
rect 14277 29155 14335 29161
rect 14277 29121 14289 29155
rect 14323 29152 14335 29155
rect 14366 29152 14372 29164
rect 14323 29124 14372 29152
rect 14323 29121 14335 29124
rect 14277 29115 14335 29121
rect 14366 29112 14372 29124
rect 14424 29112 14430 29164
rect 14476 29152 14504 29192
rect 14550 29180 14556 29232
rect 14608 29220 14614 29232
rect 14608 29192 14872 29220
rect 14608 29180 14614 29192
rect 14844 29161 14872 29192
rect 16114 29180 16120 29232
rect 16172 29229 16178 29232
rect 16172 29220 16184 29229
rect 16172 29192 16217 29220
rect 16172 29183 16184 29192
rect 16172 29180 16178 29183
rect 17328 29178 17356 29260
rect 17402 29248 17408 29260
rect 17460 29248 17466 29300
rect 17405 29181 17463 29187
rect 17405 29178 17417 29181
rect 14646 29155 14704 29161
rect 14646 29152 14658 29155
rect 14476 29124 14658 29152
rect 14646 29121 14658 29124
rect 14692 29121 14704 29155
rect 14646 29115 14704 29121
rect 14829 29155 14887 29161
rect 14829 29121 14841 29155
rect 14875 29152 14887 29155
rect 14875 29124 15424 29152
rect 14875 29121 14887 29124
rect 14829 29115 14887 29121
rect 11514 29044 11520 29096
rect 11572 29084 11578 29096
rect 12253 29087 12311 29093
rect 12253 29084 12265 29087
rect 11572 29056 12265 29084
rect 11572 29044 11578 29056
rect 12253 29053 12265 29056
rect 12299 29053 12311 29087
rect 12253 29047 12311 29053
rect 14461 29087 14519 29093
rect 14461 29053 14473 29087
rect 14507 29053 14519 29087
rect 14461 29047 14519 29053
rect 14553 29087 14611 29093
rect 14553 29053 14565 29087
rect 14599 29084 14611 29087
rect 14734 29084 14740 29096
rect 14599 29056 14740 29084
rect 14599 29053 14611 29056
rect 14553 29047 14611 29053
rect 14476 29016 14504 29047
rect 14734 29044 14740 29056
rect 14792 29044 14798 29096
rect 14642 29016 14648 29028
rect 13556 28988 14044 29016
rect 14476 28988 14648 29016
rect 13556 28948 13584 28988
rect 14016 28960 14044 28988
rect 14642 28976 14648 28988
rect 14700 29016 14706 29028
rect 14826 29016 14832 29028
rect 14700 28988 14832 29016
rect 14700 28976 14706 28988
rect 14826 28976 14832 28988
rect 14884 28976 14890 29028
rect 15010 29016 15016 29028
rect 14971 28988 15016 29016
rect 15010 28976 15016 28988
rect 15068 28976 15074 29028
rect 15396 29016 15424 29124
rect 15654 29112 15660 29164
rect 15712 29152 15718 29164
rect 16853 29155 16911 29161
rect 16853 29152 16865 29155
rect 15712 29124 16865 29152
rect 15712 29112 15718 29124
rect 16853 29121 16865 29124
rect 16899 29121 16911 29155
rect 17218 29152 17224 29164
rect 17180 29124 17224 29152
rect 16853 29115 16911 29121
rect 17218 29112 17224 29124
rect 17276 29112 17282 29164
rect 17328 29150 17417 29178
rect 17405 29147 17417 29150
rect 17451 29147 17463 29181
rect 17405 29141 17463 29147
rect 16393 29087 16451 29093
rect 16393 29053 16405 29087
rect 16439 29084 16451 29087
rect 16482 29084 16488 29096
rect 16439 29056 16488 29084
rect 16439 29053 16451 29056
rect 16393 29047 16451 29053
rect 16482 29044 16488 29056
rect 16540 29044 16546 29096
rect 17034 29084 17040 29096
rect 16995 29056 17040 29084
rect 17034 29044 17040 29056
rect 17092 29044 17098 29096
rect 17126 29044 17132 29096
rect 17184 29084 17190 29096
rect 17184 29056 17229 29084
rect 17184 29044 17190 29056
rect 16574 29016 16580 29028
rect 15396 28988 15516 29016
rect 11164 28920 13584 28948
rect 13998 28908 14004 28960
rect 14056 28908 14062 28960
rect 15488 28948 15516 28988
rect 16408 28988 16580 29016
rect 16408 28948 16436 28988
rect 16574 28976 16580 28988
rect 16632 28976 16638 29028
rect 17310 28976 17316 29028
rect 17368 28976 17374 29028
rect 17589 29019 17647 29025
rect 17589 29016 17601 29019
rect 17499 28988 17601 29016
rect 17589 28985 17601 28988
rect 17635 29016 17647 29019
rect 28810 29016 28816 29028
rect 17635 28988 28816 29016
rect 17635 28985 17647 28988
rect 17589 28979 17647 28985
rect 15488 28920 16436 28948
rect 17328 28948 17356 28976
rect 17604 28948 17632 28979
rect 28810 28976 28816 28988
rect 28868 28976 28874 29028
rect 17328 28920 17632 28948
rect 29641 28951 29699 28957
rect 29641 28917 29653 28951
rect 29687 28948 29699 28951
rect 30006 28948 30012 28960
rect 29687 28920 30012 28948
rect 29687 28917 29699 28920
rect 29641 28911 29699 28917
rect 30006 28908 30012 28920
rect 30064 28908 30070 28960
rect 1104 28858 29532 28880
rect 1104 28806 5688 28858
rect 5740 28806 5752 28858
rect 5804 28806 5816 28858
rect 5868 28806 5880 28858
rect 5932 28806 5944 28858
rect 5996 28806 15163 28858
rect 15215 28806 15227 28858
rect 15279 28806 15291 28858
rect 15343 28806 15355 28858
rect 15407 28806 15419 28858
rect 15471 28806 24639 28858
rect 24691 28806 24703 28858
rect 24755 28806 24767 28858
rect 24819 28806 24831 28858
rect 24883 28806 24895 28858
rect 24947 28806 29532 28858
rect 1104 28784 29532 28806
rect 9861 28747 9919 28753
rect 9861 28713 9873 28747
rect 9907 28744 9919 28747
rect 9950 28744 9956 28756
rect 9907 28716 9956 28744
rect 9907 28713 9919 28716
rect 9861 28707 9919 28713
rect 9950 28704 9956 28716
rect 10008 28704 10014 28756
rect 10042 28704 10048 28756
rect 10100 28744 10106 28756
rect 10597 28747 10655 28753
rect 10597 28744 10609 28747
rect 10100 28716 10609 28744
rect 10100 28704 10106 28716
rect 10597 28713 10609 28716
rect 10643 28713 10655 28747
rect 10597 28707 10655 28713
rect 12434 28704 12440 28756
rect 12492 28744 12498 28756
rect 12894 28744 12900 28756
rect 12492 28716 12900 28744
rect 12492 28704 12498 28716
rect 12894 28704 12900 28716
rect 12952 28704 12958 28756
rect 14553 28747 14611 28753
rect 14553 28713 14565 28747
rect 14599 28744 14611 28747
rect 14642 28744 14648 28756
rect 14599 28716 14648 28744
rect 14599 28713 14611 28716
rect 14553 28707 14611 28713
rect 14642 28704 14648 28716
rect 14700 28704 14706 28756
rect 14734 28704 14740 28756
rect 14792 28744 14798 28756
rect 14829 28747 14887 28753
rect 14829 28744 14841 28747
rect 14792 28716 14841 28744
rect 14792 28704 14798 28716
rect 14829 28713 14841 28716
rect 14875 28713 14887 28747
rect 14829 28707 14887 28713
rect 11054 28676 11060 28688
rect 9968 28648 11060 28676
rect 7926 28500 7932 28552
rect 7984 28540 7990 28552
rect 9858 28540 9864 28552
rect 7984 28512 9864 28540
rect 7984 28500 7990 28512
rect 9858 28500 9864 28512
rect 9916 28500 9922 28552
rect 9968 28549 9996 28648
rect 11054 28636 11060 28648
rect 11112 28636 11118 28688
rect 11241 28679 11299 28685
rect 11241 28645 11253 28679
rect 11287 28676 11299 28679
rect 17770 28676 17776 28688
rect 11287 28648 17776 28676
rect 11287 28645 11299 28648
rect 11241 28639 11299 28645
rect 10042 28568 10048 28620
rect 10100 28608 10106 28620
rect 10137 28611 10195 28617
rect 10137 28608 10149 28611
rect 10100 28580 10149 28608
rect 10100 28568 10106 28580
rect 10137 28577 10149 28580
rect 10183 28577 10195 28611
rect 11256 28608 11284 28639
rect 17770 28636 17776 28648
rect 17828 28636 17834 28688
rect 10137 28571 10195 28577
rect 10428 28580 11284 28608
rect 9953 28543 10011 28549
rect 9953 28509 9965 28543
rect 9999 28509 10011 28543
rect 10226 28540 10232 28552
rect 10187 28512 10232 28540
rect 9953 28503 10011 28509
rect 10226 28500 10232 28512
rect 10284 28500 10290 28552
rect 10339 28543 10397 28549
rect 10339 28509 10351 28543
rect 10385 28540 10397 28543
rect 10428 28540 10456 28580
rect 12802 28568 12808 28620
rect 12860 28608 12866 28620
rect 16114 28608 16120 28620
rect 12860 28580 15240 28608
rect 16075 28580 16120 28608
rect 12860 28568 12866 28580
rect 10385 28512 10456 28540
rect 10505 28543 10563 28549
rect 10385 28509 10397 28512
rect 10339 28503 10397 28509
rect 10505 28509 10517 28543
rect 10551 28509 10563 28543
rect 10778 28540 10784 28552
rect 10739 28512 10784 28540
rect 10505 28503 10563 28509
rect 9766 28432 9772 28484
rect 9824 28472 9830 28484
rect 10520 28472 10548 28503
rect 10778 28500 10784 28512
rect 10836 28500 10842 28552
rect 11057 28543 11115 28549
rect 11057 28509 11069 28543
rect 11103 28509 11115 28543
rect 12618 28540 12624 28552
rect 12579 28512 12624 28540
rect 11057 28503 11115 28509
rect 9824 28444 10548 28472
rect 9824 28432 9830 28444
rect 10594 28432 10600 28484
rect 10652 28472 10658 28484
rect 11072 28472 11100 28503
rect 12618 28500 12624 28512
rect 12676 28540 12682 28552
rect 14734 28540 14740 28552
rect 12676 28512 14740 28540
rect 12676 28500 12682 28512
rect 14734 28500 14740 28512
rect 14792 28500 14798 28552
rect 15013 28543 15071 28549
rect 15013 28509 15025 28543
rect 15059 28540 15071 28543
rect 15105 28543 15163 28549
rect 15105 28540 15117 28543
rect 15059 28512 15117 28540
rect 15059 28509 15071 28512
rect 15013 28503 15071 28509
rect 15105 28509 15117 28512
rect 15151 28509 15163 28543
rect 15212 28540 15240 28580
rect 16114 28568 16120 28580
rect 16172 28568 16178 28620
rect 17770 28540 17776 28552
rect 15212 28512 17776 28540
rect 15105 28503 15163 28509
rect 11238 28472 11244 28484
rect 10652 28444 11008 28472
rect 11072 28444 11244 28472
rect 10652 28432 10658 28444
rect 9858 28364 9864 28416
rect 9916 28404 9922 28416
rect 10226 28404 10232 28416
rect 9916 28376 10232 28404
rect 9916 28364 9922 28376
rect 10226 28364 10232 28376
rect 10284 28404 10290 28416
rect 10873 28407 10931 28413
rect 10873 28404 10885 28407
rect 10284 28376 10885 28404
rect 10284 28364 10290 28376
rect 10873 28373 10885 28376
rect 10919 28373 10931 28407
rect 10980 28404 11008 28444
rect 11238 28432 11244 28444
rect 11296 28472 11302 28484
rect 15028 28472 15056 28503
rect 17770 28500 17776 28512
rect 17828 28500 17834 28552
rect 11296 28444 15056 28472
rect 11296 28432 11302 28444
rect 12250 28404 12256 28416
rect 10980 28376 12256 28404
rect 10873 28367 10931 28373
rect 12250 28364 12256 28376
rect 12308 28364 12314 28416
rect 14826 28364 14832 28416
rect 14884 28404 14890 28416
rect 15289 28407 15347 28413
rect 15289 28404 15301 28407
rect 14884 28376 15301 28404
rect 14884 28364 14890 28376
rect 15289 28373 15301 28376
rect 15335 28373 15347 28407
rect 15562 28404 15568 28416
rect 15523 28376 15568 28404
rect 15289 28367 15347 28373
rect 15562 28364 15568 28376
rect 15620 28364 15626 28416
rect 15930 28404 15936 28416
rect 15891 28376 15936 28404
rect 15930 28364 15936 28376
rect 15988 28364 15994 28416
rect 16025 28407 16083 28413
rect 16025 28373 16037 28407
rect 16071 28404 16083 28407
rect 17034 28404 17040 28416
rect 16071 28376 17040 28404
rect 16071 28373 16083 28376
rect 16025 28367 16083 28373
rect 17034 28364 17040 28376
rect 17092 28364 17098 28416
rect 17126 28364 17132 28416
rect 17184 28404 17190 28416
rect 17865 28407 17923 28413
rect 17865 28404 17877 28407
rect 17184 28376 17877 28404
rect 17184 28364 17190 28376
rect 17865 28373 17877 28376
rect 17911 28404 17923 28407
rect 26326 28404 26332 28416
rect 17911 28376 26332 28404
rect 17911 28373 17923 28376
rect 17865 28367 17923 28373
rect 26326 28364 26332 28376
rect 26384 28364 26390 28416
rect 1104 28314 29532 28336
rect 1104 28262 10425 28314
rect 10477 28262 10489 28314
rect 10541 28262 10553 28314
rect 10605 28262 10617 28314
rect 10669 28262 10681 28314
rect 10733 28262 19901 28314
rect 19953 28262 19965 28314
rect 20017 28262 20029 28314
rect 20081 28262 20093 28314
rect 20145 28262 20157 28314
rect 20209 28262 29532 28314
rect 1104 28240 29532 28262
rect 7650 28200 7656 28212
rect 6012 28172 7656 28200
rect 4062 28092 4068 28144
rect 4120 28132 4126 28144
rect 4120 28104 5948 28132
rect 4120 28092 4126 28104
rect 5445 28067 5503 28073
rect 5445 28064 5457 28067
rect 5092 28036 5457 28064
rect 5092 27860 5120 28036
rect 5445 28033 5457 28036
rect 5491 28033 5503 28067
rect 5445 28027 5503 28033
rect 5534 28024 5540 28076
rect 5592 28064 5598 28076
rect 5628 28067 5686 28073
rect 5628 28064 5640 28067
rect 5592 28036 5640 28064
rect 5592 28024 5598 28036
rect 5628 28033 5640 28036
rect 5674 28033 5686 28067
rect 5628 28027 5686 28033
rect 5718 28024 5724 28076
rect 5776 28064 5782 28076
rect 5776 28036 5821 28064
rect 5776 28024 5782 28036
rect 5166 27956 5172 28008
rect 5224 27996 5230 28008
rect 5813 27999 5871 28005
rect 5813 27996 5825 27999
rect 5224 27968 5825 27996
rect 5224 27956 5230 27968
rect 5813 27965 5825 27968
rect 5859 27965 5871 27999
rect 5920 27996 5948 28104
rect 6012 28073 6040 28172
rect 7650 28160 7656 28172
rect 7708 28200 7714 28212
rect 7745 28203 7803 28209
rect 7745 28200 7757 28203
rect 7708 28172 7757 28200
rect 7708 28160 7714 28172
rect 7745 28169 7757 28172
rect 7791 28169 7803 28203
rect 7745 28163 7803 28169
rect 9677 28203 9735 28209
rect 9677 28169 9689 28203
rect 9723 28200 9735 28203
rect 9766 28200 9772 28212
rect 9723 28172 9772 28200
rect 9723 28169 9735 28172
rect 9677 28163 9735 28169
rect 9766 28160 9772 28172
rect 9824 28200 9830 28212
rect 10321 28203 10379 28209
rect 10321 28200 10333 28203
rect 9824 28172 10333 28200
rect 9824 28160 9830 28172
rect 10321 28169 10333 28172
rect 10367 28169 10379 28203
rect 12066 28200 12072 28212
rect 10321 28163 10379 28169
rect 11164 28172 12072 28200
rect 6181 28135 6239 28141
rect 6181 28101 6193 28135
rect 6227 28132 6239 28135
rect 6610 28135 6668 28141
rect 6610 28132 6622 28135
rect 6227 28104 6622 28132
rect 6227 28101 6239 28104
rect 6181 28095 6239 28101
rect 6610 28101 6622 28104
rect 6656 28101 6668 28135
rect 10413 28135 10471 28141
rect 10413 28132 10425 28135
rect 6610 28095 6668 28101
rect 7944 28104 10425 28132
rect 5997 28067 6055 28073
rect 5997 28033 6009 28067
rect 6043 28033 6055 28067
rect 6362 28064 6368 28076
rect 6323 28036 6368 28064
rect 5997 28027 6055 28033
rect 6362 28024 6368 28036
rect 6420 28024 6426 28076
rect 7944 28064 7972 28104
rect 10413 28101 10425 28104
rect 10459 28132 10471 28135
rect 10459 28104 10732 28132
rect 10459 28101 10471 28104
rect 10413 28095 10471 28101
rect 6472 28036 7972 28064
rect 8196 28067 8254 28073
rect 6472 27996 6500 28036
rect 8196 28033 8208 28067
rect 8242 28064 8254 28067
rect 8938 28064 8944 28076
rect 8242 28036 8944 28064
rect 8242 28033 8254 28036
rect 8196 28027 8254 28033
rect 8938 28024 8944 28036
rect 8996 28024 9002 28076
rect 9398 28024 9404 28076
rect 9456 28064 9462 28076
rect 9861 28067 9919 28073
rect 9861 28064 9873 28067
rect 9456 28036 9873 28064
rect 9456 28024 9462 28036
rect 9861 28033 9873 28036
rect 9907 28064 9919 28067
rect 9953 28067 10011 28073
rect 9953 28064 9965 28067
rect 9907 28036 9965 28064
rect 9907 28033 9919 28036
rect 9861 28027 9919 28033
rect 9953 28033 9965 28036
rect 9999 28033 10011 28067
rect 9953 28027 10011 28033
rect 10321 28067 10379 28073
rect 10321 28033 10333 28067
rect 10367 28064 10379 28067
rect 10597 28067 10655 28073
rect 10597 28064 10609 28067
rect 10367 28036 10609 28064
rect 10367 28033 10379 28036
rect 10321 28027 10379 28033
rect 10597 28033 10609 28036
rect 10643 28033 10655 28067
rect 10704 28064 10732 28104
rect 11164 28073 11192 28172
rect 12066 28160 12072 28172
rect 12124 28200 12130 28212
rect 12897 28203 12955 28209
rect 12897 28200 12909 28203
rect 12124 28172 12909 28200
rect 12124 28160 12130 28172
rect 12897 28169 12909 28172
rect 12943 28169 12955 28203
rect 12897 28163 12955 28169
rect 14550 28160 14556 28212
rect 14608 28200 14614 28212
rect 17865 28203 17923 28209
rect 17865 28200 17877 28203
rect 14608 28172 17877 28200
rect 14608 28160 14614 28172
rect 11333 28135 11391 28141
rect 11333 28101 11345 28135
rect 11379 28132 11391 28135
rect 11762 28135 11820 28141
rect 11762 28132 11774 28135
rect 11379 28104 11774 28132
rect 11379 28101 11391 28104
rect 11333 28095 11391 28101
rect 11762 28101 11774 28104
rect 11808 28101 11820 28135
rect 11762 28095 11820 28101
rect 11974 28092 11980 28144
rect 12032 28092 12038 28144
rect 12250 28092 12256 28144
rect 12308 28132 12314 28144
rect 14182 28132 14188 28144
rect 12308 28104 14188 28132
rect 12308 28092 12314 28104
rect 14182 28092 14188 28104
rect 14240 28092 14246 28144
rect 16482 28132 16488 28144
rect 14568 28104 16488 28132
rect 10762 28067 10820 28073
rect 10762 28064 10774 28067
rect 10704 28036 10774 28064
rect 10597 28027 10655 28033
rect 10762 28033 10774 28036
rect 10808 28033 10820 28067
rect 10762 28027 10820 28033
rect 10873 28067 10931 28073
rect 10873 28033 10885 28067
rect 10919 28064 10931 28067
rect 11149 28067 11207 28073
rect 10919 28036 11100 28064
rect 10919 28033 10931 28036
rect 10873 28027 10931 28033
rect 5920 27968 6500 27996
rect 7929 27999 7987 28005
rect 5813 27959 5871 27965
rect 7929 27965 7941 27999
rect 7975 27965 7987 27999
rect 7929 27959 7987 27965
rect 5350 27888 5356 27940
rect 5408 27928 5414 27940
rect 5718 27928 5724 27940
rect 5408 27900 5724 27928
rect 5408 27888 5414 27900
rect 5718 27888 5724 27900
rect 5776 27888 5782 27940
rect 6270 27860 6276 27872
rect 5092 27832 6276 27860
rect 6270 27820 6276 27832
rect 6328 27820 6334 27872
rect 7944 27860 7972 27959
rect 9122 27956 9128 28008
rect 9180 27996 9186 28008
rect 10965 27999 11023 28005
rect 9180 27968 10916 27996
rect 9180 27956 9186 27968
rect 10888 27872 10916 27968
rect 10965 27965 10977 27999
rect 11011 27965 11023 27999
rect 11072 27996 11100 28036
rect 11149 28033 11161 28067
rect 11195 28033 11207 28067
rect 11992 28064 12020 28092
rect 11149 28027 11207 28033
rect 11440 28036 12020 28064
rect 11440 27996 11468 28036
rect 13814 28024 13820 28076
rect 13872 28064 13878 28076
rect 14568 28073 14596 28104
rect 16482 28092 16488 28104
rect 16540 28092 16546 28144
rect 14286 28067 14344 28073
rect 14286 28064 14298 28067
rect 13872 28036 14298 28064
rect 13872 28024 13878 28036
rect 14286 28033 14298 28036
rect 14332 28033 14344 28067
rect 14286 28027 14344 28033
rect 14553 28067 14611 28073
rect 14553 28033 14565 28067
rect 14599 28033 14611 28067
rect 14734 28064 14740 28076
rect 14695 28036 14740 28064
rect 14553 28027 14611 28033
rect 14734 28024 14740 28036
rect 14792 28024 14798 28076
rect 15838 28024 15844 28076
rect 15896 28064 15902 28076
rect 16218 28067 16276 28073
rect 16218 28064 16230 28067
rect 15896 28036 16230 28064
rect 15896 28024 15902 28036
rect 16218 28033 16230 28036
rect 16264 28033 16276 28067
rect 16218 28027 16276 28033
rect 16574 28024 16580 28076
rect 16632 28064 16638 28076
rect 16942 28064 16948 28076
rect 16632 28036 16948 28064
rect 16632 28024 16638 28036
rect 16942 28024 16948 28036
rect 17000 28024 17006 28076
rect 17126 28064 17132 28076
rect 17087 28036 17132 28064
rect 17126 28024 17132 28036
rect 17184 28024 17190 28076
rect 17218 28024 17224 28076
rect 17276 28064 17282 28076
rect 17420 28064 17448 28172
rect 17865 28169 17877 28172
rect 17911 28169 17923 28203
rect 17865 28163 17923 28169
rect 20993 28203 21051 28209
rect 20993 28169 21005 28203
rect 21039 28169 21051 28203
rect 20993 28163 21051 28169
rect 17497 28067 17555 28073
rect 17497 28064 17509 28067
rect 17276 28036 17321 28064
rect 17420 28036 17509 28064
rect 17276 28024 17282 28036
rect 17497 28033 17509 28036
rect 17543 28033 17555 28067
rect 17497 28027 17555 28033
rect 17681 28067 17739 28073
rect 17681 28033 17693 28067
rect 17727 28064 17739 28067
rect 18978 28067 19036 28073
rect 18978 28064 18990 28067
rect 17727 28036 18990 28064
rect 17727 28033 17739 28036
rect 17681 28027 17739 28033
rect 18978 28033 18990 28036
rect 19024 28033 19036 28067
rect 20806 28064 20812 28076
rect 20767 28036 20812 28064
rect 18978 28027 19036 28033
rect 20806 28024 20812 28036
rect 20864 28024 20870 28076
rect 21008 28064 21036 28163
rect 21453 28067 21511 28073
rect 21453 28064 21465 28067
rect 21008 28036 21465 28064
rect 21453 28033 21465 28036
rect 21499 28033 21511 28067
rect 21453 28027 21511 28033
rect 11072 27968 11468 27996
rect 10965 27959 11023 27965
rect 8662 27860 8668 27872
rect 7944 27832 8668 27860
rect 8662 27820 8668 27832
rect 8720 27820 8726 27872
rect 9122 27820 9128 27872
rect 9180 27860 9186 27872
rect 9309 27863 9367 27869
rect 9309 27860 9321 27863
rect 9180 27832 9321 27860
rect 9180 27820 9186 27832
rect 9309 27829 9321 27832
rect 9355 27829 9367 27863
rect 10134 27860 10140 27872
rect 10095 27832 10140 27860
rect 9309 27823 9367 27829
rect 10134 27820 10140 27832
rect 10192 27820 10198 27872
rect 10870 27820 10876 27872
rect 10928 27820 10934 27872
rect 10980 27860 11008 27959
rect 11514 27956 11520 28008
rect 11572 27996 11578 28008
rect 16482 27996 16488 28008
rect 11572 27968 11617 27996
rect 16443 27968 16488 27996
rect 11572 27956 11578 27968
rect 16482 27956 16488 27968
rect 16540 27956 16546 28008
rect 16850 27956 16856 28008
rect 16908 27996 16914 28008
rect 17313 27999 17371 28005
rect 17313 27996 17325 27999
rect 16908 27968 17325 27996
rect 16908 27956 16914 27968
rect 17313 27965 17325 27968
rect 17359 27965 17371 27999
rect 17313 27959 17371 27965
rect 19245 27999 19303 28005
rect 19245 27965 19257 27999
rect 19291 27965 19303 27999
rect 19245 27959 19303 27965
rect 12434 27860 12440 27872
rect 10980 27832 12440 27860
rect 12434 27820 12440 27832
rect 12492 27860 12498 27872
rect 12986 27860 12992 27872
rect 12492 27832 12992 27860
rect 12492 27820 12498 27832
rect 12986 27820 12992 27832
rect 13044 27820 13050 27872
rect 13170 27860 13176 27872
rect 13131 27832 13176 27860
rect 13170 27820 13176 27832
rect 13228 27820 13234 27872
rect 14918 27860 14924 27872
rect 14879 27832 14924 27860
rect 14918 27820 14924 27832
rect 14976 27820 14982 27872
rect 15105 27863 15163 27869
rect 15105 27829 15117 27863
rect 15151 27860 15163 27863
rect 15746 27860 15752 27872
rect 15151 27832 15752 27860
rect 15151 27829 15163 27832
rect 15105 27823 15163 27829
rect 15746 27820 15752 27832
rect 15804 27820 15810 27872
rect 18874 27820 18880 27872
rect 18932 27860 18938 27872
rect 19260 27860 19288 27959
rect 18932 27832 19288 27860
rect 21637 27863 21695 27869
rect 18932 27820 18938 27832
rect 21637 27829 21649 27863
rect 21683 27860 21695 27863
rect 22094 27860 22100 27872
rect 21683 27832 22100 27860
rect 21683 27829 21695 27832
rect 21637 27823 21695 27829
rect 22094 27820 22100 27832
rect 22152 27820 22158 27872
rect 1104 27770 29532 27792
rect 1104 27718 5688 27770
rect 5740 27718 5752 27770
rect 5804 27718 5816 27770
rect 5868 27718 5880 27770
rect 5932 27718 5944 27770
rect 5996 27718 15163 27770
rect 15215 27718 15227 27770
rect 15279 27718 15291 27770
rect 15343 27718 15355 27770
rect 15407 27718 15419 27770
rect 15471 27718 24639 27770
rect 24691 27718 24703 27770
rect 24755 27718 24767 27770
rect 24819 27718 24831 27770
rect 24883 27718 24895 27770
rect 24947 27718 29532 27770
rect 1104 27696 29532 27718
rect 5534 27616 5540 27668
rect 5592 27656 5598 27668
rect 6365 27659 6423 27665
rect 6365 27656 6377 27659
rect 5592 27628 6377 27656
rect 5592 27616 5598 27628
rect 6365 27625 6377 27628
rect 6411 27656 6423 27659
rect 6454 27656 6460 27668
rect 6411 27628 6460 27656
rect 6411 27625 6423 27628
rect 6365 27619 6423 27625
rect 6454 27616 6460 27628
rect 6512 27616 6518 27668
rect 9214 27616 9220 27668
rect 9272 27656 9278 27668
rect 9858 27656 9864 27668
rect 9272 27628 9864 27656
rect 9272 27616 9278 27628
rect 9858 27616 9864 27628
rect 9916 27616 9922 27668
rect 10045 27659 10103 27665
rect 10045 27625 10057 27659
rect 10091 27656 10103 27659
rect 10778 27656 10784 27668
rect 10091 27628 10784 27656
rect 10091 27625 10103 27628
rect 10045 27619 10103 27625
rect 10778 27616 10784 27628
rect 10836 27616 10842 27668
rect 10870 27616 10876 27668
rect 10928 27656 10934 27668
rect 14642 27656 14648 27668
rect 10928 27628 14648 27656
rect 10928 27616 10934 27628
rect 14642 27616 14648 27628
rect 14700 27616 14706 27668
rect 14918 27616 14924 27668
rect 14976 27656 14982 27668
rect 14976 27628 16344 27656
rect 14976 27616 14982 27628
rect 8938 27588 8944 27600
rect 8899 27560 8944 27588
rect 8938 27548 8944 27560
rect 8996 27548 9002 27600
rect 9674 27588 9680 27600
rect 9232 27560 9680 27588
rect 7466 27520 7472 27532
rect 7427 27492 7472 27520
rect 7466 27480 7472 27492
rect 7524 27480 7530 27532
rect 7650 27520 7656 27532
rect 7611 27492 7656 27520
rect 7650 27480 7656 27492
rect 7708 27480 7714 27532
rect 9232 27520 9260 27560
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 11054 27588 11060 27600
rect 10520 27560 11060 27588
rect 9309 27523 9367 27529
rect 9309 27520 9321 27523
rect 9232 27492 9321 27520
rect 9309 27489 9321 27492
rect 9355 27489 9367 27523
rect 10226 27520 10232 27532
rect 9309 27483 9367 27489
rect 9526 27492 10232 27520
rect 9122 27452 9128 27464
rect 9083 27424 9128 27452
rect 9122 27412 9128 27424
rect 9180 27412 9186 27464
rect 9214 27412 9220 27464
rect 9272 27446 9278 27464
rect 9401 27455 9459 27461
rect 9526 27458 9554 27492
rect 10226 27480 10232 27492
rect 10284 27480 10290 27532
rect 10520 27529 10548 27560
rect 11054 27548 11060 27560
rect 11112 27548 11118 27600
rect 11238 27588 11244 27600
rect 11199 27560 11244 27588
rect 11238 27548 11244 27560
rect 11296 27548 11302 27600
rect 11701 27591 11759 27597
rect 11701 27557 11713 27591
rect 11747 27588 11759 27591
rect 11974 27588 11980 27600
rect 11747 27560 11980 27588
rect 11747 27557 11759 27560
rect 11701 27551 11759 27557
rect 11974 27548 11980 27560
rect 12032 27588 12038 27600
rect 12986 27588 12992 27600
rect 12032 27560 12756 27588
rect 12032 27548 12038 27560
rect 10321 27523 10379 27529
rect 10321 27489 10333 27523
rect 10367 27489 10379 27523
rect 10321 27483 10379 27489
rect 10505 27523 10563 27529
rect 10505 27489 10517 27523
rect 10551 27489 10563 27523
rect 10505 27483 10563 27489
rect 9401 27446 9413 27455
rect 9272 27421 9413 27446
rect 9447 27421 9459 27455
rect 9272 27418 9459 27421
rect 9272 27412 9278 27418
rect 9401 27415 9459 27418
rect 9511 27452 9569 27458
rect 9511 27418 9523 27452
rect 9557 27418 9569 27452
rect 9511 27412 9569 27418
rect 9674 27412 9680 27464
rect 9732 27452 9738 27464
rect 9858 27452 9864 27464
rect 9732 27424 9777 27452
rect 9819 27424 9864 27452
rect 9732 27412 9738 27424
rect 9858 27412 9864 27424
rect 9916 27412 9922 27464
rect 10137 27455 10195 27461
rect 10137 27421 10149 27455
rect 10183 27452 10195 27455
rect 10336 27452 10364 27483
rect 10183 27424 10364 27452
rect 10183 27421 10195 27424
rect 10137 27415 10195 27421
rect 10962 27412 10968 27464
rect 11020 27452 11026 27464
rect 11057 27455 11115 27461
rect 11057 27452 11069 27455
rect 11020 27424 11069 27452
rect 11020 27412 11026 27424
rect 11057 27421 11069 27424
rect 11103 27421 11115 27455
rect 11256 27452 11284 27548
rect 12728 27529 12756 27560
rect 12820 27560 12992 27588
rect 12820 27529 12848 27560
rect 12986 27548 12992 27560
rect 13044 27548 13050 27600
rect 13173 27591 13231 27597
rect 13173 27557 13185 27591
rect 13219 27588 13231 27591
rect 13814 27588 13820 27600
rect 13219 27560 13820 27588
rect 13219 27557 13231 27560
rect 13173 27551 13231 27557
rect 13814 27548 13820 27560
rect 13872 27548 13878 27600
rect 13909 27591 13967 27597
rect 13909 27557 13921 27591
rect 13955 27557 13967 27591
rect 13909 27551 13967 27557
rect 12713 27523 12771 27529
rect 12713 27489 12725 27523
rect 12759 27489 12771 27523
rect 12713 27483 12771 27489
rect 12805 27523 12863 27529
rect 12805 27489 12817 27523
rect 12851 27489 12863 27523
rect 12805 27483 12863 27489
rect 13262 27480 13268 27532
rect 13320 27520 13326 27532
rect 13924 27520 13952 27551
rect 14826 27548 14832 27600
rect 14884 27588 14890 27600
rect 15286 27588 15292 27600
rect 14884 27560 15292 27588
rect 14884 27548 14890 27560
rect 15286 27548 15292 27560
rect 15344 27548 15350 27600
rect 14274 27520 14280 27532
rect 13320 27492 13952 27520
rect 14235 27492 14280 27520
rect 13320 27480 13326 27492
rect 11885 27455 11943 27461
rect 11885 27452 11897 27455
rect 11256 27424 11897 27452
rect 11057 27415 11115 27421
rect 11885 27421 11897 27424
rect 11931 27421 11943 27455
rect 11885 27415 11943 27421
rect 12434 27455 12492 27461
rect 12434 27421 12446 27455
rect 12480 27452 12492 27455
rect 12526 27452 12532 27464
rect 12480 27424 12532 27452
rect 12480 27421 12492 27424
rect 12434 27415 12492 27421
rect 12526 27412 12532 27424
rect 12584 27412 12590 27464
rect 12620 27455 12678 27461
rect 12620 27421 12632 27455
rect 12666 27452 12678 27455
rect 12894 27452 12900 27464
rect 12666 27424 12900 27452
rect 12666 27421 12678 27424
rect 12620 27415 12678 27421
rect 12894 27412 12900 27424
rect 12952 27412 12958 27464
rect 12989 27455 13047 27461
rect 12989 27421 13001 27455
rect 13035 27452 13047 27455
rect 13170 27452 13176 27464
rect 13035 27424 13176 27452
rect 13035 27421 13047 27424
rect 12989 27415 13047 27421
rect 13170 27412 13176 27424
rect 13228 27412 13234 27464
rect 13722 27452 13728 27464
rect 13683 27424 13728 27452
rect 13722 27412 13728 27424
rect 13780 27412 13786 27464
rect 13924 27452 13952 27492
rect 14274 27480 14280 27492
rect 14332 27480 14338 27532
rect 14369 27523 14427 27529
rect 14369 27489 14381 27523
rect 14415 27520 14427 27523
rect 14550 27520 14556 27532
rect 14415 27492 14556 27520
rect 14415 27489 14427 27492
rect 14369 27483 14427 27489
rect 14550 27480 14556 27492
rect 14608 27480 14614 27532
rect 15396 27520 15424 27628
rect 15838 27588 15844 27600
rect 15799 27560 15844 27588
rect 15838 27548 15844 27560
rect 15896 27548 15902 27600
rect 15473 27523 15531 27529
rect 15473 27520 15485 27523
rect 15396 27492 15485 27520
rect 15473 27489 15485 27492
rect 15519 27489 15531 27523
rect 15746 27520 15752 27532
rect 15473 27483 15531 27489
rect 15632 27492 15752 27520
rect 15105 27455 15163 27461
rect 15105 27452 15117 27455
rect 13924 27424 15117 27452
rect 15105 27421 15117 27424
rect 15151 27421 15163 27455
rect 15105 27415 15163 27421
rect 15288 27449 15346 27455
rect 15288 27415 15300 27449
rect 15334 27415 15346 27449
rect 15288 27409 15346 27415
rect 15378 27412 15384 27464
rect 15436 27452 15442 27464
rect 15632 27461 15660 27492
rect 15746 27480 15752 27492
rect 15804 27480 15810 27532
rect 16316 27520 16344 27628
rect 16850 27548 16856 27600
rect 16908 27548 16914 27600
rect 17497 27591 17555 27597
rect 17497 27588 17509 27591
rect 17144 27560 17509 27588
rect 16868 27520 16896 27548
rect 16945 27523 17003 27529
rect 16945 27520 16957 27523
rect 16316 27492 16957 27520
rect 16945 27489 16957 27492
rect 16991 27489 17003 27523
rect 16945 27483 17003 27489
rect 15611 27455 15669 27461
rect 15436 27424 15481 27452
rect 15436 27412 15442 27424
rect 15611 27421 15623 27455
rect 15657 27421 15669 27455
rect 16574 27452 16580 27464
rect 16535 27424 16580 27452
rect 15611 27415 15669 27421
rect 16574 27412 16580 27424
rect 16632 27412 16638 27464
rect 16666 27412 16672 27464
rect 16724 27452 16730 27464
rect 16760 27455 16818 27461
rect 16760 27452 16772 27455
rect 16724 27424 16772 27452
rect 16724 27412 16730 27424
rect 16760 27421 16772 27424
rect 16806 27421 16818 27455
rect 16760 27415 16818 27421
rect 16853 27455 16911 27461
rect 16853 27421 16865 27455
rect 16899 27421 16911 27455
rect 16853 27415 16911 27421
rect 7098 27344 7104 27396
rect 7156 27384 7162 27396
rect 10597 27387 10655 27393
rect 10597 27384 10609 27387
rect 7156 27356 10609 27384
rect 7156 27344 7162 27356
rect 10597 27353 10609 27356
rect 10643 27353 10655 27387
rect 10597 27347 10655 27353
rect 10980 27356 12434 27384
rect 4062 27276 4068 27328
rect 4120 27316 4126 27328
rect 6730 27316 6736 27328
rect 4120 27288 6736 27316
rect 4120 27276 4126 27288
rect 6730 27276 6736 27288
rect 6788 27276 6794 27328
rect 7742 27276 7748 27328
rect 7800 27316 7806 27328
rect 8113 27319 8171 27325
rect 7800 27288 7845 27316
rect 7800 27276 7806 27288
rect 8113 27285 8125 27319
rect 8159 27316 8171 27319
rect 8846 27316 8852 27328
rect 8159 27288 8852 27316
rect 8159 27285 8171 27288
rect 8113 27279 8171 27285
rect 8846 27276 8852 27288
rect 8904 27276 8910 27328
rect 9582 27276 9588 27328
rect 9640 27316 9646 27328
rect 10980 27325 11008 27356
rect 10137 27319 10195 27325
rect 10137 27316 10149 27319
rect 9640 27288 10149 27316
rect 9640 27276 9646 27288
rect 10137 27285 10149 27288
rect 10183 27285 10195 27319
rect 10137 27279 10195 27285
rect 10965 27319 11023 27325
rect 10965 27285 10977 27319
rect 11011 27285 11023 27319
rect 12406 27316 12434 27356
rect 12526 27316 12532 27328
rect 12406 27288 12532 27316
rect 10965 27279 11023 27285
rect 12526 27276 12532 27288
rect 12584 27276 12590 27328
rect 12894 27276 12900 27328
rect 12952 27316 12958 27328
rect 13262 27316 13268 27328
rect 12952 27288 13268 27316
rect 12952 27276 12958 27288
rect 13262 27276 13268 27288
rect 13320 27276 13326 27328
rect 13354 27276 13360 27328
rect 13412 27316 13418 27328
rect 14461 27319 14519 27325
rect 14461 27316 14473 27319
rect 13412 27288 14473 27316
rect 13412 27276 13418 27288
rect 14461 27285 14473 27288
rect 14507 27285 14519 27319
rect 14461 27279 14519 27285
rect 14734 27276 14740 27328
rect 14792 27316 14798 27328
rect 14829 27319 14887 27325
rect 14829 27316 14841 27319
rect 14792 27288 14841 27316
rect 14792 27276 14798 27288
rect 14829 27285 14841 27288
rect 14875 27285 14887 27319
rect 15303 27316 15331 27409
rect 16390 27344 16396 27396
rect 16448 27384 16454 27396
rect 16868 27384 16896 27415
rect 17034 27412 17040 27464
rect 17092 27452 17098 27464
rect 17144 27461 17172 27560
rect 17497 27557 17509 27560
rect 17543 27557 17555 27591
rect 17497 27551 17555 27557
rect 22646 27548 22652 27600
rect 22704 27588 22710 27600
rect 22925 27591 22983 27597
rect 22925 27588 22937 27591
rect 22704 27560 22937 27588
rect 22704 27548 22710 27560
rect 22925 27557 22937 27560
rect 22971 27557 22983 27591
rect 22925 27551 22983 27557
rect 19337 27523 19395 27529
rect 19337 27489 19349 27523
rect 19383 27520 19395 27523
rect 20254 27520 20260 27532
rect 19383 27492 20260 27520
rect 19383 27489 19395 27492
rect 19337 27483 19395 27489
rect 20254 27480 20260 27492
rect 20312 27520 20318 27532
rect 20438 27520 20444 27532
rect 20312 27492 20444 27520
rect 20312 27480 20318 27492
rect 20438 27480 20444 27492
rect 20496 27480 20502 27532
rect 17129 27455 17187 27461
rect 17129 27452 17141 27455
rect 17092 27424 17141 27452
rect 17092 27412 17098 27424
rect 17129 27421 17141 27424
rect 17175 27421 17187 27455
rect 18874 27452 18880 27464
rect 18835 27424 18880 27452
rect 17129 27415 17187 27421
rect 18874 27412 18880 27424
rect 18932 27412 18938 27464
rect 21082 27412 21088 27464
rect 21140 27452 21146 27464
rect 21177 27455 21235 27461
rect 21177 27452 21189 27455
rect 21140 27424 21189 27452
rect 21140 27412 21146 27424
rect 21177 27421 21189 27424
rect 21223 27421 21235 27455
rect 21177 27415 21235 27421
rect 17218 27384 17224 27396
rect 16448 27356 17224 27384
rect 16448 27344 16454 27356
rect 17218 27344 17224 27356
rect 17276 27344 17282 27396
rect 17313 27387 17371 27393
rect 17313 27353 17325 27387
rect 17359 27384 17371 27387
rect 18610 27387 18668 27393
rect 18610 27384 18622 27387
rect 17359 27356 18622 27384
rect 17359 27353 17371 27356
rect 17313 27347 17371 27353
rect 18610 27353 18622 27356
rect 18656 27353 18668 27387
rect 18610 27347 18668 27353
rect 18782 27344 18788 27396
rect 18840 27384 18846 27396
rect 19242 27384 19248 27396
rect 18840 27356 19248 27384
rect 18840 27344 18846 27356
rect 19242 27344 19248 27356
rect 19300 27384 19306 27396
rect 19300 27356 19642 27384
rect 19300 27344 19306 27356
rect 20714 27344 20720 27396
rect 20772 27384 20778 27396
rect 20809 27387 20867 27393
rect 20809 27384 20821 27387
rect 20772 27356 20821 27384
rect 20772 27344 20778 27356
rect 20809 27353 20821 27356
rect 20855 27353 20867 27387
rect 20809 27347 20867 27353
rect 21453 27387 21511 27393
rect 21453 27353 21465 27387
rect 21499 27384 21511 27387
rect 21542 27384 21548 27396
rect 21499 27356 21548 27384
rect 21499 27353 21511 27356
rect 21453 27347 21511 27353
rect 21542 27344 21548 27356
rect 21600 27344 21606 27396
rect 22094 27344 22100 27396
rect 22152 27344 22158 27396
rect 16025 27319 16083 27325
rect 16025 27316 16037 27319
rect 15303 27288 16037 27316
rect 14829 27279 14887 27285
rect 16025 27285 16037 27288
rect 16071 27316 16083 27319
rect 27430 27316 27436 27328
rect 16071 27288 27436 27316
rect 16071 27285 16083 27288
rect 16025 27279 16083 27285
rect 27430 27276 27436 27288
rect 27488 27276 27494 27328
rect 1104 27226 29532 27248
rect 1104 27174 10425 27226
rect 10477 27174 10489 27226
rect 10541 27174 10553 27226
rect 10605 27174 10617 27226
rect 10669 27174 10681 27226
rect 10733 27174 19901 27226
rect 19953 27174 19965 27226
rect 20017 27174 20029 27226
rect 20081 27174 20093 27226
rect 20145 27174 20157 27226
rect 20209 27174 29532 27226
rect 1104 27152 29532 27174
rect 6086 27112 6092 27124
rect 5999 27084 6092 27112
rect 6086 27072 6092 27084
rect 6144 27112 6150 27124
rect 6733 27115 6791 27121
rect 6733 27112 6745 27115
rect 6144 27084 6745 27112
rect 6144 27072 6150 27084
rect 6733 27081 6745 27084
rect 6779 27081 6791 27115
rect 7098 27112 7104 27124
rect 7059 27084 7104 27112
rect 6733 27075 6791 27081
rect 7098 27072 7104 27084
rect 7156 27072 7162 27124
rect 8846 27112 8852 27124
rect 8807 27084 8852 27112
rect 8846 27072 8852 27084
rect 8904 27072 8910 27124
rect 12066 27072 12072 27124
rect 12124 27112 12130 27124
rect 12161 27115 12219 27121
rect 12161 27112 12173 27115
rect 12124 27084 12173 27112
rect 12124 27072 12130 27084
rect 12161 27081 12173 27084
rect 12207 27081 12219 27115
rect 12161 27075 12219 27081
rect 12621 27115 12679 27121
rect 12621 27081 12633 27115
rect 12667 27112 12679 27115
rect 14369 27115 14427 27121
rect 14369 27112 14381 27115
rect 12667 27084 14381 27112
rect 12667 27081 12679 27084
rect 12621 27075 12679 27081
rect 14369 27081 14381 27084
rect 14415 27081 14427 27115
rect 14369 27075 14427 27081
rect 14458 27072 14464 27124
rect 14516 27112 14522 27124
rect 15838 27112 15844 27124
rect 14516 27084 14561 27112
rect 15799 27084 15844 27112
rect 14516 27072 14522 27084
rect 15838 27072 15844 27084
rect 15896 27072 15902 27124
rect 16853 27115 16911 27121
rect 16853 27081 16865 27115
rect 16899 27112 16911 27115
rect 16942 27112 16948 27124
rect 16899 27084 16948 27112
rect 16899 27081 16911 27084
rect 16853 27075 16911 27081
rect 16942 27072 16948 27084
rect 17000 27072 17006 27124
rect 20806 27112 20812 27124
rect 17052 27084 20812 27112
rect 4154 27044 4160 27056
rect 3160 27016 4160 27044
rect 3160 26985 3188 27016
rect 4154 27004 4160 27016
rect 4212 27044 4218 27056
rect 6362 27044 6368 27056
rect 4212 27016 6368 27044
rect 4212 27004 4218 27016
rect 3145 26979 3203 26985
rect 3145 26945 3157 26979
rect 3191 26945 3203 26979
rect 3145 26939 3203 26945
rect 3412 26979 3470 26985
rect 3412 26945 3424 26979
rect 3458 26976 3470 26979
rect 4614 26976 4620 26988
rect 3458 26948 4620 26976
rect 3458 26945 3470 26948
rect 3412 26939 3470 26945
rect 4614 26936 4620 26948
rect 4672 26936 4678 26988
rect 4724 26985 4752 27016
rect 6362 27004 6368 27016
rect 6420 27004 6426 27056
rect 7466 27044 7472 27056
rect 6564 27016 7472 27044
rect 4709 26979 4767 26985
rect 4709 26945 4721 26979
rect 4755 26945 4767 26979
rect 4709 26939 4767 26945
rect 4976 26979 5034 26985
rect 4976 26945 4988 26979
rect 5022 26976 5034 26979
rect 5534 26976 5540 26988
rect 5022 26948 5540 26976
rect 5022 26945 5034 26948
rect 4976 26939 5034 26945
rect 5534 26936 5540 26948
rect 5592 26936 5598 26988
rect 6564 26917 6592 27016
rect 7466 27004 7472 27016
rect 7524 27004 7530 27056
rect 8757 27047 8815 27053
rect 8757 27013 8769 27047
rect 8803 27044 8815 27047
rect 9122 27044 9128 27056
rect 8803 27016 9128 27044
rect 8803 27013 8815 27016
rect 8757 27007 8815 27013
rect 9122 27004 9128 27016
rect 9180 27004 9186 27056
rect 13909 27047 13967 27053
rect 13909 27044 13921 27047
rect 9324 27016 13921 27044
rect 6730 26936 6736 26988
rect 6788 26976 6794 26988
rect 9324 26976 9352 27016
rect 13909 27013 13921 27016
rect 13955 27013 13967 27047
rect 15749 27047 15807 27053
rect 15749 27044 15761 27047
rect 13909 27007 13967 27013
rect 14108 27016 15761 27044
rect 6788 26948 9352 26976
rect 6788 26936 6794 26948
rect 9398 26936 9404 26988
rect 9456 26976 9462 26988
rect 9493 26979 9551 26985
rect 9493 26976 9505 26979
rect 9456 26948 9505 26976
rect 9456 26936 9462 26948
rect 9493 26945 9505 26948
rect 9539 26945 9551 26979
rect 9493 26939 9551 26945
rect 9769 26979 9827 26985
rect 9769 26945 9781 26979
rect 9815 26976 9827 26979
rect 10042 26976 10048 26988
rect 9815 26948 10048 26976
rect 9815 26945 9827 26948
rect 9769 26939 9827 26945
rect 10042 26936 10048 26948
rect 10100 26976 10106 26988
rect 10962 26976 10968 26988
rect 10100 26948 10968 26976
rect 10100 26936 10106 26948
rect 10962 26936 10968 26948
rect 11020 26936 11026 26988
rect 12250 26976 12256 26988
rect 12211 26948 12256 26976
rect 12250 26936 12256 26948
rect 12308 26936 12314 26988
rect 12342 26936 12348 26988
rect 12400 26976 12406 26988
rect 14108 26976 14136 27016
rect 15749 27013 15761 27016
rect 15795 27013 15807 27047
rect 15749 27007 15807 27013
rect 15930 27004 15936 27056
rect 15988 27004 15994 27056
rect 15948 26976 15976 27004
rect 12400 26948 14136 26976
rect 14200 26948 15976 26976
rect 12400 26936 12406 26948
rect 6549 26911 6607 26917
rect 6549 26877 6561 26911
rect 6595 26877 6607 26911
rect 6549 26871 6607 26877
rect 6641 26911 6699 26917
rect 6641 26877 6653 26911
rect 6687 26908 6699 26911
rect 6687 26880 6776 26908
rect 6687 26877 6699 26880
rect 6641 26871 6699 26877
rect 4525 26775 4583 26781
rect 4525 26741 4537 26775
rect 4571 26772 4583 26775
rect 4982 26772 4988 26784
rect 4571 26744 4988 26772
rect 4571 26741 4583 26744
rect 4525 26735 4583 26741
rect 4982 26732 4988 26744
rect 5040 26772 5046 26784
rect 6748 26772 6776 26880
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 8665 26911 8723 26917
rect 8665 26908 8677 26911
rect 8628 26880 8677 26908
rect 8628 26868 8634 26880
rect 8665 26877 8677 26880
rect 8711 26908 8723 26911
rect 9582 26908 9588 26920
rect 8711 26880 9588 26908
rect 8711 26877 8723 26880
rect 8665 26871 8723 26877
rect 9582 26868 9588 26880
rect 9640 26868 9646 26920
rect 12066 26908 12072 26920
rect 12027 26880 12072 26908
rect 12066 26868 12072 26880
rect 12124 26868 12130 26920
rect 12526 26868 12532 26920
rect 12584 26908 12590 26920
rect 14200 26908 14228 26948
rect 16298 26936 16304 26988
rect 16356 26976 16362 26988
rect 17052 26985 17080 27084
rect 20806 27072 20812 27084
rect 20864 27072 20870 27124
rect 27522 27112 27528 27124
rect 20916 27084 27528 27112
rect 20438 27004 20444 27056
rect 20496 27044 20502 27056
rect 20496 27016 20541 27044
rect 20496 27004 20502 27016
rect 20346 26985 20352 26988
rect 17037 26979 17095 26985
rect 17037 26976 17049 26979
rect 16356 26948 17049 26976
rect 16356 26936 16362 26948
rect 17037 26945 17049 26948
rect 17083 26945 17095 26979
rect 20344 26976 20352 26985
rect 20307 26948 20352 26976
rect 17037 26939 17095 26945
rect 20344 26939 20352 26948
rect 20346 26936 20352 26939
rect 20404 26936 20410 26988
rect 20530 26976 20536 26988
rect 20491 26948 20536 26976
rect 20530 26936 20536 26948
rect 20588 26936 20594 26988
rect 20717 26979 20775 26985
rect 20717 26945 20729 26979
rect 20763 26976 20775 26979
rect 20806 26976 20812 26988
rect 20763 26948 20812 26976
rect 20763 26945 20775 26948
rect 20717 26939 20775 26945
rect 20806 26936 20812 26948
rect 20864 26936 20870 26988
rect 12584 26880 14228 26908
rect 12584 26868 12590 26880
rect 14274 26868 14280 26920
rect 14332 26908 14338 26920
rect 14645 26911 14703 26917
rect 14645 26908 14657 26911
rect 14332 26880 14657 26908
rect 14332 26868 14338 26880
rect 14645 26877 14657 26880
rect 14691 26908 14703 26911
rect 14826 26908 14832 26920
rect 14691 26880 14832 26908
rect 14691 26877 14703 26880
rect 14645 26871 14703 26877
rect 14826 26868 14832 26880
rect 14884 26908 14890 26920
rect 15933 26911 15991 26917
rect 15933 26908 15945 26911
rect 14884 26880 15945 26908
rect 14884 26868 14890 26880
rect 15933 26877 15945 26880
rect 15979 26908 15991 26911
rect 16114 26908 16120 26920
rect 15979 26880 16120 26908
rect 15979 26877 15991 26880
rect 15933 26871 15991 26877
rect 16114 26868 16120 26880
rect 16172 26868 16178 26920
rect 16850 26868 16856 26920
rect 16908 26908 16914 26920
rect 20916 26908 20944 27084
rect 27522 27072 27528 27084
rect 27580 27072 27586 27124
rect 21269 27047 21327 27053
rect 21269 27013 21281 27047
rect 21315 27044 21327 27047
rect 22646 27044 22652 27056
rect 21315 27016 22652 27044
rect 21315 27013 21327 27016
rect 21269 27007 21327 27013
rect 22646 27004 22652 27016
rect 22704 27004 22710 27056
rect 20990 26936 20996 26988
rect 21048 26976 21054 26988
rect 21174 26976 21180 26988
rect 21048 26948 21093 26976
rect 21135 26948 21180 26976
rect 21048 26936 21054 26948
rect 21174 26936 21180 26948
rect 21232 26936 21238 26988
rect 21450 26985 21456 26988
rect 21413 26979 21456 26985
rect 21413 26945 21425 26979
rect 21413 26939 21456 26945
rect 21450 26936 21456 26939
rect 21508 26936 21514 26988
rect 16908 26880 20944 26908
rect 16908 26868 16914 26880
rect 9217 26843 9275 26849
rect 9217 26809 9229 26843
rect 9263 26840 9275 26843
rect 11974 26840 11980 26852
rect 9263 26812 11980 26840
rect 9263 26809 9275 26812
rect 9217 26803 9275 26809
rect 11974 26800 11980 26812
rect 12032 26800 12038 26852
rect 13909 26843 13967 26849
rect 13909 26809 13921 26843
rect 13955 26840 13967 26843
rect 18966 26840 18972 26852
rect 13955 26812 18972 26840
rect 13955 26809 13967 26812
rect 13909 26803 13967 26809
rect 18966 26800 18972 26812
rect 19024 26800 19030 26852
rect 20165 26843 20223 26849
rect 20165 26809 20177 26843
rect 20211 26840 20223 26843
rect 20714 26840 20720 26852
rect 20211 26812 20720 26840
rect 20211 26809 20223 26812
rect 20165 26803 20223 26809
rect 20714 26800 20720 26812
rect 20772 26800 20778 26852
rect 21542 26840 21548 26852
rect 21503 26812 21548 26840
rect 21542 26800 21548 26812
rect 21600 26800 21606 26852
rect 9674 26772 9680 26784
rect 5040 26744 6776 26772
rect 9635 26744 9680 26772
rect 5040 26732 5046 26744
rect 9674 26732 9680 26744
rect 9732 26732 9738 26784
rect 9858 26772 9864 26784
rect 9819 26744 9864 26772
rect 9858 26732 9864 26744
rect 9916 26732 9922 26784
rect 10137 26775 10195 26781
rect 10137 26741 10149 26775
rect 10183 26772 10195 26775
rect 10226 26772 10232 26784
rect 10183 26744 10232 26772
rect 10183 26741 10195 26744
rect 10137 26735 10195 26741
rect 10226 26732 10232 26744
rect 10284 26732 10290 26784
rect 12526 26732 12532 26784
rect 12584 26772 12590 26784
rect 13722 26772 13728 26784
rect 12584 26744 13728 26772
rect 12584 26732 12590 26744
rect 13722 26732 13728 26744
rect 13780 26732 13786 26784
rect 13998 26772 14004 26784
rect 13959 26744 14004 26772
rect 13998 26732 14004 26744
rect 14056 26732 14062 26784
rect 15381 26775 15439 26781
rect 15381 26741 15393 26775
rect 15427 26772 15439 26775
rect 15746 26772 15752 26784
rect 15427 26744 15752 26772
rect 15427 26741 15439 26744
rect 15381 26735 15439 26741
rect 15746 26732 15752 26744
rect 15804 26732 15810 26784
rect 16666 26732 16672 26784
rect 16724 26772 16730 26784
rect 17497 26775 17555 26781
rect 17497 26772 17509 26775
rect 16724 26744 17509 26772
rect 16724 26732 16730 26744
rect 17497 26741 17509 26744
rect 17543 26772 17555 26775
rect 17586 26772 17592 26784
rect 17543 26744 17592 26772
rect 17543 26741 17555 26744
rect 17497 26735 17555 26741
rect 17586 26732 17592 26744
rect 17644 26732 17650 26784
rect 20254 26732 20260 26784
rect 20312 26772 20318 26784
rect 20530 26772 20536 26784
rect 20312 26744 20536 26772
rect 20312 26732 20318 26744
rect 20530 26732 20536 26744
rect 20588 26772 20594 26784
rect 20809 26775 20867 26781
rect 20809 26772 20821 26775
rect 20588 26744 20821 26772
rect 20588 26732 20594 26744
rect 20809 26741 20821 26744
rect 20855 26741 20867 26775
rect 20809 26735 20867 26741
rect 1104 26682 29532 26704
rect 1104 26630 5688 26682
rect 5740 26630 5752 26682
rect 5804 26630 5816 26682
rect 5868 26630 5880 26682
rect 5932 26630 5944 26682
rect 5996 26630 15163 26682
rect 15215 26630 15227 26682
rect 15279 26630 15291 26682
rect 15343 26630 15355 26682
rect 15407 26630 15419 26682
rect 15471 26630 24639 26682
rect 24691 26630 24703 26682
rect 24755 26630 24767 26682
rect 24819 26630 24831 26682
rect 24883 26630 24895 26682
rect 24947 26630 29532 26682
rect 1104 26608 29532 26630
rect 4614 26528 4620 26580
rect 4672 26568 4678 26580
rect 4893 26571 4951 26577
rect 4893 26568 4905 26571
rect 4672 26540 4905 26568
rect 4672 26528 4678 26540
rect 4893 26537 4905 26540
rect 4939 26537 4951 26571
rect 4893 26531 4951 26537
rect 5534 26528 5540 26580
rect 5592 26568 5598 26580
rect 5997 26571 6055 26577
rect 5997 26568 6009 26571
rect 5592 26540 6009 26568
rect 5592 26528 5598 26540
rect 5997 26537 6009 26540
rect 6043 26537 6055 26571
rect 5997 26531 6055 26537
rect 7282 26528 7288 26580
rect 7340 26568 7346 26580
rect 7742 26568 7748 26580
rect 7340 26540 7748 26568
rect 7340 26528 7346 26540
rect 7742 26528 7748 26540
rect 7800 26568 7806 26580
rect 8389 26571 8447 26577
rect 8389 26568 8401 26571
rect 7800 26540 8401 26568
rect 7800 26528 7806 26540
rect 8389 26537 8401 26540
rect 8435 26537 8447 26571
rect 8389 26531 8447 26537
rect 10226 26528 10232 26580
rect 10284 26568 10290 26580
rect 16850 26568 16856 26580
rect 10284 26540 16856 26568
rect 10284 26528 10290 26540
rect 16850 26528 16856 26540
rect 16908 26528 16914 26580
rect 17586 26528 17592 26580
rect 17644 26568 17650 26580
rect 23842 26568 23848 26580
rect 17644 26540 23848 26568
rect 17644 26528 17650 26540
rect 23842 26528 23848 26540
rect 23900 26528 23906 26580
rect 5350 26460 5356 26512
rect 5408 26460 5414 26512
rect 5721 26503 5779 26509
rect 5721 26469 5733 26503
rect 5767 26500 5779 26503
rect 6178 26500 6184 26512
rect 5767 26472 6184 26500
rect 5767 26469 5779 26472
rect 5721 26463 5779 26469
rect 5261 26435 5319 26441
rect 5261 26401 5273 26435
rect 5307 26432 5319 26435
rect 5368 26432 5396 26460
rect 5736 26432 5764 26463
rect 6178 26460 6184 26472
rect 6236 26460 6242 26512
rect 6362 26460 6368 26512
rect 6420 26500 6426 26512
rect 10137 26503 10195 26509
rect 6420 26472 7052 26500
rect 6420 26460 6426 26472
rect 5307 26404 5396 26432
rect 5460 26404 5764 26432
rect 6273 26435 6331 26441
rect 5307 26401 5319 26404
rect 5261 26395 5319 26401
rect 4982 26364 4988 26376
rect 4943 26336 4988 26364
rect 4982 26324 4988 26336
rect 5040 26324 5046 26376
rect 5166 26364 5172 26376
rect 5127 26336 5172 26364
rect 5166 26324 5172 26336
rect 5224 26324 5230 26376
rect 5371 26367 5429 26373
rect 5371 26333 5383 26367
rect 5417 26364 5429 26367
rect 5460 26364 5488 26404
rect 6273 26401 6285 26435
rect 6319 26432 6331 26435
rect 6914 26432 6920 26444
rect 6319 26404 6920 26432
rect 6319 26401 6331 26404
rect 6273 26395 6331 26401
rect 6914 26392 6920 26404
rect 6972 26392 6978 26444
rect 7024 26441 7052 26472
rect 10137 26469 10149 26503
rect 10183 26500 10195 26503
rect 12342 26500 12348 26512
rect 10183 26472 12348 26500
rect 10183 26469 10195 26472
rect 10137 26463 10195 26469
rect 12342 26460 12348 26472
rect 12400 26460 12406 26512
rect 13449 26503 13507 26509
rect 13449 26469 13461 26503
rect 13495 26500 13507 26503
rect 17497 26503 17555 26509
rect 13495 26472 15792 26500
rect 13495 26469 13507 26472
rect 13449 26463 13507 26469
rect 7009 26435 7067 26441
rect 7009 26401 7021 26435
rect 7055 26401 7067 26435
rect 9582 26432 9588 26444
rect 9495 26404 9588 26432
rect 7009 26395 7067 26401
rect 9582 26392 9588 26404
rect 9640 26432 9646 26444
rect 12066 26432 12072 26444
rect 9640 26404 12072 26432
rect 9640 26392 9646 26404
rect 12066 26392 12072 26404
rect 12124 26432 12130 26444
rect 12805 26435 12863 26441
rect 12805 26432 12817 26435
rect 12124 26404 12817 26432
rect 12124 26392 12130 26404
rect 12805 26401 12817 26404
rect 12851 26401 12863 26435
rect 12805 26395 12863 26401
rect 12989 26435 13047 26441
rect 12989 26401 13001 26435
rect 13035 26432 13047 26435
rect 13170 26432 13176 26444
rect 13035 26404 13176 26432
rect 13035 26401 13047 26404
rect 12989 26395 13047 26401
rect 13170 26392 13176 26404
rect 13228 26392 13234 26444
rect 14826 26392 14832 26444
rect 14884 26432 14890 26444
rect 15102 26432 15108 26444
rect 14884 26404 15108 26432
rect 14884 26392 14890 26404
rect 15102 26392 15108 26404
rect 15160 26432 15166 26444
rect 15473 26435 15531 26441
rect 15473 26432 15485 26435
rect 15160 26404 15485 26432
rect 15160 26392 15166 26404
rect 15473 26401 15485 26404
rect 15519 26401 15531 26435
rect 15654 26432 15660 26444
rect 15615 26404 15660 26432
rect 15473 26395 15531 26401
rect 15654 26392 15660 26404
rect 15712 26392 15718 26444
rect 5417 26336 5488 26364
rect 5537 26367 5595 26373
rect 5417 26333 5429 26336
rect 5371 26327 5429 26333
rect 5537 26333 5549 26367
rect 5583 26364 5595 26367
rect 5718 26364 5724 26376
rect 5583 26336 5724 26364
rect 5583 26333 5595 26336
rect 5537 26327 5595 26333
rect 5718 26324 5724 26336
rect 5776 26324 5782 26376
rect 6086 26324 6092 26376
rect 6144 26364 6150 26376
rect 6362 26364 6368 26376
rect 6144 26336 6189 26364
rect 6323 26336 6368 26364
rect 6144 26324 6150 26336
rect 6362 26324 6368 26336
rect 6420 26324 6426 26376
rect 6454 26324 6460 26376
rect 6512 26364 6518 26376
rect 6641 26367 6699 26373
rect 6512 26336 6557 26364
rect 6512 26324 6518 26336
rect 6641 26333 6653 26367
rect 6687 26364 6699 26367
rect 6730 26364 6736 26376
rect 6687 26336 6736 26364
rect 6687 26333 6699 26336
rect 6641 26327 6699 26333
rect 6730 26324 6736 26336
rect 6788 26324 6794 26376
rect 9030 26324 9036 26376
rect 9088 26364 9094 26376
rect 9677 26367 9735 26373
rect 9677 26364 9689 26367
rect 9088 26336 9689 26364
rect 9088 26324 9094 26336
rect 9677 26333 9689 26336
rect 9723 26333 9735 26367
rect 9677 26327 9735 26333
rect 9858 26324 9864 26376
rect 9916 26364 9922 26376
rect 15764 26373 15792 26472
rect 17497 26469 17509 26503
rect 17543 26469 17555 26503
rect 19242 26500 19248 26512
rect 19203 26472 19248 26500
rect 17497 26463 17555 26469
rect 16390 26392 16396 26444
rect 16448 26432 16454 26444
rect 16853 26435 16911 26441
rect 16853 26432 16865 26435
rect 16448 26404 16865 26432
rect 16448 26392 16454 26404
rect 16853 26401 16865 26404
rect 16899 26401 16911 26435
rect 16853 26395 16911 26401
rect 16942 26392 16948 26444
rect 17000 26432 17006 26444
rect 17512 26432 17540 26463
rect 19242 26460 19248 26472
rect 19300 26460 19306 26512
rect 20346 26460 20352 26512
rect 20404 26500 20410 26512
rect 21542 26500 21548 26512
rect 20404 26472 21548 26500
rect 20404 26460 20410 26472
rect 21542 26460 21548 26472
rect 21600 26460 21606 26512
rect 17000 26404 17045 26432
rect 17144 26404 17540 26432
rect 17000 26392 17006 26404
rect 10413 26367 10471 26373
rect 10413 26364 10425 26367
rect 9916 26336 10425 26364
rect 9916 26324 9922 26336
rect 10413 26333 10425 26336
rect 10459 26333 10471 26367
rect 10413 26327 10471 26333
rect 15749 26367 15807 26373
rect 15749 26333 15761 26367
rect 15795 26333 15807 26367
rect 16574 26364 16580 26376
rect 16535 26336 16580 26364
rect 15749 26327 15807 26333
rect 16574 26324 16580 26336
rect 16632 26324 16638 26376
rect 16758 26364 16764 26376
rect 16719 26336 16764 26364
rect 16758 26324 16764 26336
rect 16816 26324 16822 26376
rect 17144 26373 17172 26404
rect 18966 26392 18972 26444
rect 19024 26432 19030 26444
rect 22094 26432 22100 26444
rect 19024 26404 22100 26432
rect 19024 26392 19030 26404
rect 22094 26392 22100 26404
rect 22152 26432 22158 26444
rect 23474 26432 23480 26444
rect 22152 26404 23480 26432
rect 22152 26392 22158 26404
rect 23474 26392 23480 26404
rect 23532 26392 23538 26444
rect 17129 26367 17187 26373
rect 17129 26361 17141 26367
rect 17052 26333 17141 26361
rect 17175 26333 17187 26367
rect 18874 26364 18880 26376
rect 7276 26299 7334 26305
rect 7276 26265 7288 26299
rect 7322 26296 7334 26299
rect 7374 26296 7380 26308
rect 7322 26268 7380 26296
rect 7322 26265 7334 26268
rect 7276 26259 7334 26265
rect 7374 26256 7380 26268
rect 7432 26256 7438 26308
rect 7650 26256 7656 26308
rect 7708 26296 7714 26308
rect 9769 26299 9827 26305
rect 9769 26296 9781 26299
rect 7708 26268 9781 26296
rect 7708 26256 7714 26268
rect 9769 26265 9781 26268
rect 9815 26265 9827 26299
rect 9769 26259 9827 26265
rect 12710 26256 12716 26308
rect 12768 26296 12774 26308
rect 13081 26299 13139 26305
rect 13081 26296 13093 26299
rect 12768 26268 13093 26296
rect 12768 26256 12774 26268
rect 13081 26265 13093 26268
rect 13127 26265 13139 26299
rect 13081 26259 13139 26265
rect 13722 26256 13728 26308
rect 13780 26296 13786 26308
rect 16298 26296 16304 26308
rect 13780 26268 16304 26296
rect 13780 26256 13786 26268
rect 16298 26256 16304 26268
rect 16356 26256 16362 26308
rect 16390 26256 16396 26308
rect 16448 26296 16454 26308
rect 17052 26296 17080 26333
rect 17129 26327 17187 26333
rect 17972 26336 18880 26364
rect 17972 26308 18000 26336
rect 18874 26324 18880 26336
rect 18932 26324 18938 26376
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26364 19487 26367
rect 21729 26367 21787 26373
rect 19475 26336 19564 26364
rect 19475 26333 19487 26336
rect 19429 26327 19487 26333
rect 19536 26308 19564 26336
rect 21729 26333 21741 26367
rect 21775 26333 21787 26367
rect 21729 26327 21787 26333
rect 16448 26268 17080 26296
rect 17313 26299 17371 26305
rect 16448 26256 16454 26268
rect 17313 26265 17325 26299
rect 17359 26296 17371 26299
rect 17359 26268 17908 26296
rect 17359 26265 17371 26268
rect 17313 26259 17371 26265
rect 5718 26188 5724 26240
rect 5776 26228 5782 26240
rect 6270 26228 6276 26240
rect 5776 26200 6276 26228
rect 5776 26188 5782 26200
rect 6270 26188 6276 26200
rect 6328 26228 6334 26240
rect 9674 26228 9680 26240
rect 6328 26200 9680 26228
rect 6328 26188 6334 26200
rect 9674 26188 9680 26200
rect 9732 26188 9738 26240
rect 9858 26188 9864 26240
rect 9916 26228 9922 26240
rect 10229 26231 10287 26237
rect 10229 26228 10241 26231
rect 9916 26200 10241 26228
rect 9916 26188 9922 26200
rect 10229 26197 10241 26200
rect 10275 26197 10287 26231
rect 16114 26228 16120 26240
rect 16075 26200 16120 26228
rect 10229 26191 10287 26197
rect 16114 26188 16120 26200
rect 16172 26188 16178 26240
rect 17880 26228 17908 26268
rect 17954 26256 17960 26308
rect 18012 26256 18018 26308
rect 18610 26299 18668 26305
rect 18610 26296 18622 26299
rect 18064 26268 18622 26296
rect 18064 26228 18092 26268
rect 18610 26265 18622 26268
rect 18656 26265 18668 26299
rect 19518 26296 19524 26308
rect 19479 26268 19524 26296
rect 18610 26259 18668 26265
rect 19518 26256 19524 26268
rect 19576 26256 19582 26308
rect 17880 26200 18092 26228
rect 21082 26188 21088 26240
rect 21140 26228 21146 26240
rect 21744 26228 21772 26327
rect 24486 26324 24492 26376
rect 24544 26364 24550 26376
rect 24581 26367 24639 26373
rect 24581 26364 24593 26367
rect 24544 26336 24593 26364
rect 24544 26324 24550 26336
rect 24581 26333 24593 26336
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 21910 26256 21916 26308
rect 21968 26296 21974 26308
rect 22005 26299 22063 26305
rect 22005 26296 22017 26299
rect 21968 26268 22017 26296
rect 21968 26256 21974 26268
rect 22005 26265 22017 26268
rect 22051 26265 22063 26299
rect 22005 26259 22063 26265
rect 23014 26256 23020 26308
rect 23072 26256 23078 26308
rect 23382 26228 23388 26240
rect 21140 26200 23388 26228
rect 21140 26188 21146 26200
rect 23382 26188 23388 26200
rect 23440 26188 23446 26240
rect 24394 26228 24400 26240
rect 24355 26200 24400 26228
rect 24394 26188 24400 26200
rect 24452 26188 24458 26240
rect 1104 26138 29532 26160
rect 1104 26086 10425 26138
rect 10477 26086 10489 26138
rect 10541 26086 10553 26138
rect 10605 26086 10617 26138
rect 10669 26086 10681 26138
rect 10733 26086 19901 26138
rect 19953 26086 19965 26138
rect 20017 26086 20029 26138
rect 20081 26086 20093 26138
rect 20145 26086 20157 26138
rect 20209 26086 29532 26138
rect 1104 26064 29532 26086
rect 5350 25984 5356 26036
rect 5408 25984 5414 26036
rect 5442 25984 5448 26036
rect 5500 26024 5506 26036
rect 5721 26027 5779 26033
rect 5721 26024 5733 26027
rect 5500 25996 5733 26024
rect 5500 25984 5506 25996
rect 5721 25993 5733 25996
rect 5767 26024 5779 26027
rect 6454 26024 6460 26036
rect 5767 25996 6460 26024
rect 5767 25993 5779 25996
rect 5721 25987 5779 25993
rect 6454 25984 6460 25996
rect 6512 25984 6518 26036
rect 7374 26024 7380 26036
rect 7335 25996 7380 26024
rect 7374 25984 7380 25996
rect 7432 25984 7438 26036
rect 8294 25984 8300 26036
rect 8352 26024 8358 26036
rect 8665 26027 8723 26033
rect 8665 26024 8677 26027
rect 8352 25996 8677 26024
rect 8352 25984 8358 25996
rect 8665 25993 8677 25996
rect 8711 25993 8723 26027
rect 8665 25987 8723 25993
rect 9125 26027 9183 26033
rect 9125 25993 9137 26027
rect 9171 26024 9183 26027
rect 12621 26027 12679 26033
rect 9171 25996 12434 26024
rect 9171 25993 9183 25996
rect 9125 25987 9183 25993
rect 5368 25956 5396 25984
rect 5276 25928 5396 25956
rect 4798 25888 4804 25900
rect 4759 25860 4804 25888
rect 4798 25848 4804 25860
rect 4856 25848 4862 25900
rect 5170 25891 5228 25897
rect 5170 25888 5182 25891
rect 4908 25860 5182 25888
rect 4908 25820 4936 25860
rect 5170 25857 5182 25860
rect 5216 25857 5228 25891
rect 5170 25851 5228 25857
rect 4448 25792 4936 25820
rect 4985 25823 5043 25829
rect 4246 25644 4252 25696
rect 4304 25684 4310 25696
rect 4448 25693 4476 25792
rect 4985 25789 4997 25823
rect 5031 25789 5043 25823
rect 4985 25783 5043 25789
rect 5077 25823 5135 25829
rect 5077 25789 5089 25823
rect 5123 25820 5135 25823
rect 5276 25820 5304 25928
rect 7098 25916 7104 25968
rect 7156 25956 7162 25968
rect 7561 25959 7619 25965
rect 7561 25956 7573 25959
rect 7156 25928 7573 25956
rect 7156 25916 7162 25928
rect 7561 25925 7573 25928
rect 7607 25925 7619 25959
rect 12158 25956 12164 25968
rect 7561 25919 7619 25925
rect 9416 25928 10916 25956
rect 12119 25928 12164 25956
rect 5353 25891 5411 25897
rect 5353 25857 5365 25891
rect 5399 25888 5411 25891
rect 5718 25888 5724 25900
rect 5399 25860 5724 25888
rect 5399 25857 5411 25860
rect 5353 25851 5411 25857
rect 5718 25848 5724 25860
rect 5776 25848 5782 25900
rect 6730 25888 6736 25900
rect 6691 25860 6736 25888
rect 6730 25848 6736 25860
rect 6788 25848 6794 25900
rect 6916 25891 6974 25897
rect 6916 25857 6928 25891
rect 6962 25888 6974 25891
rect 7116 25888 7144 25916
rect 7282 25888 7288 25900
rect 6962 25860 7144 25888
rect 7243 25860 7288 25888
rect 6962 25857 6974 25860
rect 6916 25851 6974 25857
rect 7282 25848 7288 25860
rect 7340 25848 7346 25900
rect 7926 25848 7932 25900
rect 7984 25888 7990 25900
rect 9416 25897 9444 25928
rect 8757 25891 8815 25897
rect 8757 25888 8769 25891
rect 7984 25860 8769 25888
rect 7984 25848 7990 25860
rect 8757 25857 8769 25860
rect 8803 25857 8815 25891
rect 8757 25851 8815 25857
rect 9401 25891 9459 25897
rect 9401 25857 9413 25891
rect 9447 25857 9459 25891
rect 9401 25851 9459 25857
rect 10128 25891 10186 25897
rect 10128 25857 10140 25891
rect 10174 25888 10186 25891
rect 10594 25888 10600 25900
rect 10174 25860 10600 25888
rect 10174 25857 10186 25860
rect 10128 25851 10186 25857
rect 6086 25820 6092 25832
rect 5123 25792 6092 25820
rect 5123 25789 5135 25792
rect 5077 25783 5135 25789
rect 5000 25752 5028 25783
rect 6086 25780 6092 25792
rect 6144 25780 6150 25832
rect 6362 25780 6368 25832
rect 6420 25820 6426 25832
rect 7009 25823 7067 25829
rect 7009 25820 7021 25823
rect 6420 25792 7021 25820
rect 6420 25780 6426 25792
rect 7009 25789 7021 25792
rect 7055 25789 7067 25823
rect 7009 25783 7067 25789
rect 7101 25823 7159 25829
rect 7101 25789 7113 25823
rect 7147 25789 7159 25823
rect 8570 25820 8576 25832
rect 8531 25792 8576 25820
rect 7101 25783 7159 25789
rect 5166 25752 5172 25764
rect 5000 25724 5172 25752
rect 5166 25712 5172 25724
rect 5224 25712 5230 25764
rect 6914 25712 6920 25764
rect 6972 25752 6978 25764
rect 7116 25752 7144 25783
rect 8570 25780 8576 25792
rect 8628 25780 8634 25832
rect 6972 25724 7144 25752
rect 6972 25712 6978 25724
rect 9122 25712 9128 25764
rect 9180 25752 9186 25764
rect 9416 25752 9444 25851
rect 10594 25848 10600 25860
rect 10652 25848 10658 25900
rect 9766 25780 9772 25832
rect 9824 25820 9830 25832
rect 9861 25823 9919 25829
rect 9861 25820 9873 25823
rect 9824 25792 9873 25820
rect 9824 25780 9830 25792
rect 9861 25789 9873 25792
rect 9907 25789 9919 25823
rect 9861 25783 9919 25789
rect 9493 25755 9551 25761
rect 9493 25752 9505 25755
rect 9180 25724 9505 25752
rect 9180 25712 9186 25724
rect 9493 25721 9505 25724
rect 9539 25721 9551 25755
rect 10888 25752 10916 25928
rect 12158 25916 12164 25928
rect 12216 25916 12222 25968
rect 12406 25956 12434 25996
rect 12621 25993 12633 26027
rect 12667 26024 12679 26027
rect 15010 26024 15016 26036
rect 12667 25996 14228 26024
rect 14971 25996 15016 26024
rect 12667 25993 12679 25996
rect 12621 25987 12679 25993
rect 14093 25959 14151 25965
rect 14093 25956 14105 25959
rect 12406 25928 14105 25956
rect 14093 25925 14105 25928
rect 14139 25925 14151 25959
rect 14200 25956 14228 25996
rect 15010 25984 15016 25996
rect 15068 25984 15074 26036
rect 19334 26024 19340 26036
rect 19295 25996 19340 26024
rect 19334 25984 19340 25996
rect 19392 25984 19398 26036
rect 22094 25984 22100 26036
rect 22152 26024 22158 26036
rect 25133 26027 25191 26033
rect 25133 26024 25145 26027
rect 22152 25996 22232 26024
rect 22152 25984 22158 25996
rect 14921 25959 14979 25965
rect 14921 25956 14933 25959
rect 14200 25928 14933 25956
rect 14093 25919 14151 25925
rect 14921 25925 14933 25928
rect 14967 25925 14979 25959
rect 14921 25919 14979 25925
rect 20070 25916 20076 25968
rect 20128 25916 20134 25968
rect 22204 25965 22232 25996
rect 22940 25996 25145 26024
rect 22940 25965 22968 25996
rect 25133 25993 25145 25996
rect 25179 26024 25191 26027
rect 27522 26024 27528 26036
rect 25179 25996 27528 26024
rect 25179 25993 25191 25996
rect 25133 25987 25191 25993
rect 27522 25984 27528 25996
rect 27580 25984 27586 26036
rect 22189 25959 22247 25965
rect 22189 25925 22201 25959
rect 22235 25925 22247 25959
rect 22189 25919 22247 25925
rect 22925 25959 22983 25965
rect 22925 25925 22937 25959
rect 22971 25925 22983 25959
rect 22925 25919 22983 25925
rect 24394 25916 24400 25968
rect 24452 25916 24458 25968
rect 12253 25891 12311 25897
rect 12253 25857 12265 25891
rect 12299 25888 12311 25891
rect 12342 25888 12348 25900
rect 12299 25860 12348 25888
rect 12299 25857 12311 25860
rect 12253 25851 12311 25857
rect 12342 25848 12348 25860
rect 12400 25848 12406 25900
rect 14185 25891 14243 25897
rect 14185 25857 14197 25891
rect 14231 25888 14243 25891
rect 16390 25888 16396 25900
rect 14231 25860 16396 25888
rect 14231 25857 14243 25860
rect 14185 25851 14243 25857
rect 16390 25848 16396 25860
rect 16448 25848 16454 25900
rect 21634 25848 21640 25900
rect 21692 25888 21698 25900
rect 22092 25891 22150 25897
rect 22092 25888 22104 25891
rect 21692 25860 22104 25888
rect 21692 25848 21698 25860
rect 22092 25857 22104 25860
rect 22138 25857 22150 25891
rect 22278 25888 22284 25900
rect 22239 25860 22284 25888
rect 22092 25851 22150 25857
rect 12066 25820 12072 25832
rect 11979 25792 12072 25820
rect 12066 25780 12072 25792
rect 12124 25820 12130 25832
rect 12802 25820 12808 25832
rect 12124 25792 12808 25820
rect 12124 25780 12130 25792
rect 12802 25780 12808 25792
rect 12860 25780 12866 25832
rect 14274 25820 14280 25832
rect 14235 25792 14280 25820
rect 14274 25780 14280 25792
rect 14332 25820 14338 25832
rect 15102 25820 15108 25832
rect 14332 25792 15108 25820
rect 14332 25780 14338 25792
rect 15102 25780 15108 25792
rect 15160 25780 15166 25832
rect 20806 25820 20812 25832
rect 20767 25792 20812 25820
rect 20806 25780 20812 25792
rect 20864 25780 20870 25832
rect 21082 25820 21088 25832
rect 21043 25792 21088 25820
rect 21082 25780 21088 25792
rect 21140 25780 21146 25832
rect 19518 25752 19524 25764
rect 10888 25724 12020 25752
rect 9493 25715 9551 25721
rect 4433 25687 4491 25693
rect 4433 25684 4445 25687
rect 4304 25656 4445 25684
rect 4304 25644 4310 25656
rect 4433 25653 4445 25656
rect 4479 25653 4491 25687
rect 4706 25684 4712 25696
rect 4667 25656 4712 25684
rect 4433 25647 4491 25653
rect 4706 25644 4712 25656
rect 4764 25644 4770 25696
rect 6730 25644 6736 25696
rect 6788 25684 6794 25696
rect 8938 25684 8944 25696
rect 6788 25656 8944 25684
rect 6788 25644 6794 25656
rect 8938 25644 8944 25656
rect 8996 25684 9002 25696
rect 9217 25687 9275 25693
rect 9217 25684 9229 25687
rect 8996 25656 9229 25684
rect 8996 25644 9002 25656
rect 9217 25653 9229 25656
rect 9263 25653 9275 25687
rect 9217 25647 9275 25653
rect 11241 25687 11299 25693
rect 11241 25653 11253 25687
rect 11287 25684 11299 25687
rect 11514 25684 11520 25696
rect 11287 25656 11520 25684
rect 11287 25653 11299 25656
rect 11241 25647 11299 25653
rect 11514 25644 11520 25656
rect 11572 25644 11578 25696
rect 11992 25684 12020 25724
rect 12406 25724 19524 25752
rect 12406 25684 12434 25724
rect 19518 25712 19524 25724
rect 19576 25712 19582 25764
rect 21910 25752 21916 25764
rect 21871 25724 21916 25752
rect 21910 25712 21916 25724
rect 21968 25712 21974 25764
rect 22112 25752 22140 25851
rect 22278 25848 22284 25860
rect 22336 25848 22342 25900
rect 22465 25891 22523 25897
rect 22465 25857 22477 25891
rect 22511 25888 22523 25891
rect 22557 25891 22615 25897
rect 22557 25888 22569 25891
rect 22511 25860 22569 25888
rect 22511 25857 22523 25860
rect 22465 25851 22523 25857
rect 22557 25857 22569 25860
rect 22603 25888 22615 25891
rect 22649 25891 22707 25897
rect 22649 25888 22661 25891
rect 22603 25860 22661 25888
rect 22603 25857 22615 25860
rect 22557 25851 22615 25857
rect 22649 25857 22661 25860
rect 22695 25857 22707 25891
rect 22649 25851 22707 25857
rect 22738 25848 22744 25900
rect 22796 25888 22802 25900
rect 22833 25891 22891 25897
rect 22833 25888 22845 25891
rect 22796 25860 22845 25888
rect 22796 25848 22802 25860
rect 22833 25857 22845 25860
rect 22879 25857 22891 25891
rect 23022 25891 23080 25897
rect 23022 25888 23034 25891
rect 22833 25851 22891 25857
rect 22940 25860 23034 25888
rect 22940 25752 22968 25860
rect 23022 25857 23034 25860
rect 23068 25857 23080 25891
rect 23382 25888 23388 25900
rect 23343 25860 23388 25888
rect 23022 25851 23080 25857
rect 23382 25848 23388 25860
rect 23440 25848 23446 25900
rect 23661 25823 23719 25829
rect 23661 25820 23673 25823
rect 23492 25792 23673 25820
rect 22112 25724 22968 25752
rect 23201 25755 23259 25761
rect 23201 25721 23213 25755
rect 23247 25752 23259 25755
rect 23492 25752 23520 25792
rect 23661 25789 23673 25792
rect 23707 25789 23719 25823
rect 23661 25783 23719 25789
rect 23247 25724 23520 25752
rect 23247 25721 23259 25724
rect 23201 25715 23259 25721
rect 11992 25656 12434 25684
rect 13725 25687 13783 25693
rect 13725 25653 13737 25687
rect 13771 25684 13783 25687
rect 13814 25684 13820 25696
rect 13771 25656 13820 25684
rect 13771 25653 13783 25656
rect 13725 25647 13783 25653
rect 13814 25644 13820 25656
rect 13872 25644 13878 25696
rect 13906 25644 13912 25696
rect 13964 25684 13970 25696
rect 14553 25687 14611 25693
rect 14553 25684 14565 25687
rect 13964 25656 14565 25684
rect 13964 25644 13970 25656
rect 14553 25653 14565 25656
rect 14599 25653 14611 25687
rect 14553 25647 14611 25653
rect 14826 25644 14832 25696
rect 14884 25684 14890 25696
rect 16022 25684 16028 25696
rect 14884 25656 16028 25684
rect 14884 25644 14890 25656
rect 16022 25644 16028 25656
rect 16080 25644 16086 25696
rect 16758 25644 16764 25696
rect 16816 25684 16822 25696
rect 17497 25687 17555 25693
rect 17497 25684 17509 25687
rect 16816 25656 17509 25684
rect 16816 25644 16822 25656
rect 17497 25653 17509 25656
rect 17543 25684 17555 25687
rect 17586 25684 17592 25696
rect 17543 25656 17592 25684
rect 17543 25653 17555 25656
rect 17497 25647 17555 25653
rect 17586 25644 17592 25656
rect 17644 25644 17650 25696
rect 22002 25644 22008 25696
rect 22060 25684 22066 25696
rect 22557 25687 22615 25693
rect 22557 25684 22569 25687
rect 22060 25656 22569 25684
rect 22060 25644 22066 25656
rect 22557 25653 22569 25656
rect 22603 25653 22615 25687
rect 22557 25647 22615 25653
rect 1104 25594 29532 25616
rect 1104 25542 5688 25594
rect 5740 25542 5752 25594
rect 5804 25542 5816 25594
rect 5868 25542 5880 25594
rect 5932 25542 5944 25594
rect 5996 25542 15163 25594
rect 15215 25542 15227 25594
rect 15279 25542 15291 25594
rect 15343 25542 15355 25594
rect 15407 25542 15419 25594
rect 15471 25542 24639 25594
rect 24691 25542 24703 25594
rect 24755 25542 24767 25594
rect 24819 25542 24831 25594
rect 24883 25542 24895 25594
rect 24947 25542 29532 25594
rect 1104 25520 29532 25542
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 7558 25480 7564 25492
rect 4120 25452 7564 25480
rect 4120 25440 4126 25452
rect 7558 25440 7564 25452
rect 7616 25440 7622 25492
rect 7926 25480 7932 25492
rect 7887 25452 7932 25480
rect 7926 25440 7932 25452
rect 7984 25440 7990 25492
rect 10594 25480 10600 25492
rect 10555 25452 10600 25480
rect 10594 25440 10600 25452
rect 10652 25440 10658 25492
rect 11977 25483 12035 25489
rect 11977 25449 11989 25483
rect 12023 25480 12035 25483
rect 12250 25480 12256 25492
rect 12023 25452 12256 25480
rect 12023 25449 12035 25452
rect 11977 25443 12035 25449
rect 12250 25440 12256 25452
rect 12308 25440 12314 25492
rect 12406 25452 13860 25480
rect 5166 25372 5172 25424
rect 5224 25412 5230 25424
rect 5905 25415 5963 25421
rect 5905 25412 5917 25415
rect 5224 25384 5917 25412
rect 5224 25372 5230 25384
rect 5905 25381 5917 25384
rect 5951 25381 5963 25415
rect 5905 25375 5963 25381
rect 9674 25372 9680 25424
rect 9732 25412 9738 25424
rect 10873 25415 10931 25421
rect 9732 25384 9996 25412
rect 9732 25372 9738 25384
rect 4154 25344 4160 25356
rect 4115 25316 4160 25344
rect 4154 25304 4160 25316
rect 4212 25304 4218 25356
rect 7377 25347 7435 25353
rect 7377 25313 7389 25347
rect 7423 25344 7435 25347
rect 7466 25344 7472 25356
rect 7423 25316 7472 25344
rect 7423 25313 7435 25316
rect 7377 25307 7435 25313
rect 7466 25304 7472 25316
rect 7524 25304 7530 25356
rect 4424 25279 4482 25285
rect 4424 25245 4436 25279
rect 4470 25276 4482 25279
rect 4706 25276 4712 25288
rect 4470 25248 4712 25276
rect 4470 25245 4482 25248
rect 4424 25239 4482 25245
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 6089 25279 6147 25285
rect 6089 25245 6101 25279
rect 6135 25276 6147 25279
rect 6457 25279 6515 25285
rect 6457 25276 6469 25279
rect 6135 25248 6469 25276
rect 6135 25245 6147 25248
rect 6089 25239 6147 25245
rect 6457 25245 6469 25248
rect 6503 25276 6515 25279
rect 9125 25279 9183 25285
rect 9125 25276 9137 25279
rect 6503 25248 9137 25276
rect 6503 25245 6515 25248
rect 6457 25239 6515 25245
rect 9125 25245 9137 25248
rect 9171 25276 9183 25279
rect 9677 25279 9735 25285
rect 9677 25276 9689 25279
rect 9171 25248 9689 25276
rect 9171 25245 9183 25248
rect 9125 25239 9183 25245
rect 9677 25245 9689 25248
rect 9723 25276 9735 25279
rect 9858 25276 9864 25288
rect 9723 25248 9864 25276
rect 9723 25245 9735 25248
rect 9677 25239 9735 25245
rect 9858 25236 9864 25248
rect 9916 25236 9922 25288
rect 9968 25285 9996 25384
rect 10873 25381 10885 25415
rect 10919 25412 10931 25415
rect 12406 25412 12434 25452
rect 10919 25384 12434 25412
rect 13832 25412 13860 25452
rect 14642 25440 14648 25492
rect 14700 25480 14706 25492
rect 16945 25483 17003 25489
rect 16945 25480 16957 25483
rect 14700 25452 16957 25480
rect 14700 25440 14706 25452
rect 16945 25449 16957 25452
rect 16991 25449 17003 25483
rect 16945 25443 17003 25449
rect 19981 25483 20039 25489
rect 19981 25449 19993 25483
rect 20027 25480 20039 25483
rect 20070 25480 20076 25492
rect 20027 25452 20076 25480
rect 20027 25449 20039 25452
rect 19981 25443 20039 25449
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 20806 25440 20812 25492
rect 20864 25480 20870 25492
rect 20901 25483 20959 25489
rect 20901 25480 20913 25483
rect 20864 25452 20913 25480
rect 20864 25440 20870 25452
rect 20901 25449 20913 25452
rect 20947 25449 20959 25483
rect 23014 25480 23020 25492
rect 22975 25452 23020 25480
rect 20901 25443 20959 25449
rect 23014 25440 23020 25452
rect 23072 25440 23078 25492
rect 23201 25483 23259 25489
rect 23201 25449 23213 25483
rect 23247 25480 23259 25483
rect 23474 25480 23480 25492
rect 23247 25452 23480 25480
rect 23247 25449 23259 25452
rect 23201 25443 23259 25449
rect 23474 25440 23480 25452
rect 23532 25440 23538 25492
rect 24486 25440 24492 25492
rect 24544 25480 24550 25492
rect 24581 25483 24639 25489
rect 24581 25480 24593 25483
rect 24544 25452 24593 25480
rect 24544 25440 24550 25452
rect 24581 25449 24593 25452
rect 24627 25449 24639 25483
rect 24581 25443 24639 25449
rect 14826 25412 14832 25424
rect 13832 25384 14832 25412
rect 10919 25381 10931 25384
rect 10873 25375 10931 25381
rect 10888 25344 10916 25375
rect 14826 25372 14832 25384
rect 14884 25372 14890 25424
rect 19518 25372 19524 25424
rect 19576 25412 19582 25424
rect 21821 25415 21879 25421
rect 21821 25412 21833 25415
rect 19576 25384 21833 25412
rect 19576 25372 19582 25384
rect 21821 25381 21833 25384
rect 21867 25381 21879 25415
rect 21821 25375 21879 25381
rect 11330 25344 11336 25356
rect 10060 25316 10916 25344
rect 11291 25316 11336 25344
rect 9953 25279 10011 25285
rect 9953 25245 9965 25279
rect 9999 25245 10011 25279
rect 10060 25276 10088 25316
rect 11330 25304 11336 25316
rect 11388 25304 11394 25356
rect 11514 25344 11520 25356
rect 11475 25316 11520 25344
rect 11514 25304 11520 25316
rect 11572 25304 11578 25356
rect 12802 25344 12808 25356
rect 12763 25316 12808 25344
rect 12802 25304 12808 25316
rect 12860 25304 12866 25356
rect 12989 25347 13047 25353
rect 12989 25313 13001 25347
rect 13035 25344 13047 25347
rect 13630 25344 13636 25356
rect 13035 25316 13636 25344
rect 13035 25313 13047 25316
rect 12989 25307 13047 25313
rect 13630 25304 13636 25316
rect 13688 25304 13694 25356
rect 14185 25347 14243 25353
rect 14185 25313 14197 25347
rect 14231 25313 14243 25347
rect 14366 25344 14372 25356
rect 14327 25316 14372 25344
rect 14185 25307 14243 25313
rect 10118 25279 10176 25285
rect 10118 25276 10130 25279
rect 10060 25248 10130 25276
rect 9953 25239 10011 25245
rect 10118 25245 10130 25248
rect 10164 25245 10176 25279
rect 10118 25239 10176 25245
rect 10229 25279 10287 25285
rect 10229 25245 10241 25279
rect 10275 25245 10287 25279
rect 10229 25239 10287 25245
rect 4798 25168 4804 25220
rect 4856 25208 4862 25220
rect 7469 25211 7527 25217
rect 7469 25208 7481 25211
rect 4856 25180 7481 25208
rect 4856 25168 4862 25180
rect 5552 25149 5580 25180
rect 7469 25177 7481 25180
rect 7515 25177 7527 25211
rect 7469 25171 7527 25177
rect 8662 25168 8668 25220
rect 8720 25208 8726 25220
rect 9582 25208 9588 25220
rect 8720 25180 9588 25208
rect 8720 25168 8726 25180
rect 9582 25168 9588 25180
rect 9640 25168 9646 25220
rect 10244 25208 10272 25239
rect 10318 25236 10324 25288
rect 10376 25276 10382 25288
rect 10505 25279 10563 25285
rect 10376 25248 10421 25276
rect 10376 25236 10382 25248
rect 10505 25245 10517 25279
rect 10551 25276 10563 25279
rect 11532 25276 11560 25304
rect 10551 25248 11560 25276
rect 14200 25276 14228 25307
rect 14366 25304 14372 25316
rect 14424 25304 14430 25356
rect 15197 25347 15255 25353
rect 15197 25313 15209 25347
rect 15243 25344 15255 25347
rect 16482 25344 16488 25356
rect 15243 25316 16488 25344
rect 15243 25313 15255 25316
rect 15197 25307 15255 25313
rect 16482 25304 16488 25316
rect 16540 25344 16546 25356
rect 17129 25347 17187 25353
rect 17129 25344 17141 25347
rect 16540 25316 17141 25344
rect 16540 25304 16546 25316
rect 17129 25313 17141 25316
rect 17175 25344 17187 25347
rect 17954 25344 17960 25356
rect 17175 25316 17960 25344
rect 17175 25313 17187 25316
rect 17129 25307 17187 25313
rect 17954 25304 17960 25316
rect 18012 25304 18018 25356
rect 19334 25304 19340 25356
rect 19392 25344 19398 25356
rect 21634 25344 21640 25356
rect 19392 25316 20300 25344
rect 19392 25304 19398 25316
rect 14274 25276 14280 25288
rect 14200 25248 14280 25276
rect 10551 25245 10563 25248
rect 10505 25239 10563 25245
rect 14274 25236 14280 25248
rect 14332 25236 14338 25288
rect 16574 25236 16580 25288
rect 16632 25236 16638 25288
rect 19610 25276 19616 25288
rect 19571 25248 19616 25276
rect 19610 25236 19616 25248
rect 19668 25276 19674 25288
rect 19705 25279 19763 25285
rect 19705 25276 19717 25279
rect 19668 25248 19717 25276
rect 19668 25236 19674 25248
rect 19705 25245 19717 25248
rect 19751 25245 19763 25279
rect 20165 25279 20223 25285
rect 20165 25276 20177 25279
rect 19705 25239 19763 25245
rect 19904 25248 20177 25276
rect 14461 25211 14519 25217
rect 14461 25208 14473 25211
rect 9968 25180 10272 25208
rect 13464 25180 14473 25208
rect 9968 25152 9996 25180
rect 5537 25143 5595 25149
rect 5537 25109 5549 25143
rect 5583 25109 5595 25143
rect 5537 25103 5595 25109
rect 6273 25143 6331 25149
rect 6273 25109 6285 25143
rect 6319 25140 6331 25143
rect 6822 25140 6828 25152
rect 6319 25112 6828 25140
rect 6319 25109 6331 25112
rect 6273 25103 6331 25109
rect 6822 25100 6828 25112
rect 6880 25100 6886 25152
rect 7561 25143 7619 25149
rect 7561 25109 7573 25143
rect 7607 25140 7619 25143
rect 7742 25140 7748 25152
rect 7607 25112 7748 25140
rect 7607 25109 7619 25112
rect 7561 25103 7619 25109
rect 7742 25100 7748 25112
rect 7800 25100 7806 25152
rect 8941 25143 8999 25149
rect 8941 25109 8953 25143
rect 8987 25140 8999 25143
rect 9306 25140 9312 25152
rect 8987 25112 9312 25140
rect 8987 25109 8999 25112
rect 8941 25103 8999 25109
rect 9306 25100 9312 25112
rect 9364 25100 9370 25152
rect 9858 25140 9864 25152
rect 9819 25112 9864 25140
rect 9858 25100 9864 25112
rect 9916 25100 9922 25152
rect 9950 25100 9956 25152
rect 10008 25100 10014 25152
rect 10226 25100 10232 25152
rect 10284 25140 10290 25152
rect 11609 25143 11667 25149
rect 11609 25140 11621 25143
rect 10284 25112 11621 25140
rect 10284 25100 10290 25112
rect 11609 25109 11621 25112
rect 11655 25109 11667 25143
rect 11609 25103 11667 25109
rect 13078 25100 13084 25152
rect 13136 25140 13142 25152
rect 13464 25149 13492 25180
rect 14461 25177 14473 25180
rect 14507 25177 14519 25211
rect 15470 25208 15476 25220
rect 15431 25180 15476 25208
rect 14461 25171 14519 25177
rect 15470 25168 15476 25180
rect 15528 25168 15534 25220
rect 17402 25208 17408 25220
rect 17363 25180 17408 25208
rect 17402 25168 17408 25180
rect 17460 25168 17466 25220
rect 19794 25208 19800 25220
rect 18630 25180 19800 25208
rect 19794 25168 19800 25180
rect 19852 25168 19858 25220
rect 13449 25143 13507 25149
rect 13136 25112 13181 25140
rect 13136 25100 13142 25112
rect 13449 25109 13461 25143
rect 13495 25109 13507 25143
rect 14826 25140 14832 25152
rect 14787 25112 14832 25140
rect 13449 25103 13507 25109
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 18046 25100 18052 25152
rect 18104 25140 18110 25152
rect 19904 25149 19932 25248
rect 20165 25245 20177 25248
rect 20211 25245 20223 25279
rect 20165 25239 20223 25245
rect 20272 25208 20300 25316
rect 21376 25316 21640 25344
rect 21080 25279 21138 25285
rect 21080 25245 21092 25279
rect 21126 25276 21138 25279
rect 21376 25276 21404 25316
rect 21634 25304 21640 25316
rect 21692 25304 21698 25356
rect 21836 25344 21864 25375
rect 21836 25316 22048 25344
rect 21126 25248 21404 25276
rect 21453 25279 21511 25285
rect 21126 25245 21138 25248
rect 21080 25239 21138 25245
rect 21453 25245 21465 25279
rect 21499 25276 21511 25279
rect 21910 25276 21916 25288
rect 21499 25248 21916 25276
rect 21499 25245 21511 25248
rect 21453 25239 21511 25245
rect 21910 25236 21916 25248
rect 21968 25236 21974 25288
rect 22020 25285 22048 25316
rect 22005 25279 22063 25285
rect 22005 25245 22017 25279
rect 22051 25245 22063 25279
rect 22554 25276 22560 25288
rect 22515 25248 22560 25276
rect 22005 25239 22063 25245
rect 22554 25236 22560 25248
rect 22612 25236 22618 25288
rect 22833 25279 22891 25285
rect 22833 25276 22845 25279
rect 22756 25248 22845 25276
rect 21177 25211 21235 25217
rect 21177 25208 21189 25211
rect 20272 25180 21189 25208
rect 21177 25177 21189 25180
rect 21223 25177 21235 25211
rect 21177 25171 21235 25177
rect 21269 25211 21327 25217
rect 21269 25177 21281 25211
rect 21315 25208 21327 25211
rect 21315 25180 22094 25208
rect 21315 25177 21327 25180
rect 21269 25171 21327 25177
rect 22066 25152 22094 25180
rect 18877 25143 18935 25149
rect 18877 25140 18889 25143
rect 18104 25112 18889 25140
rect 18104 25100 18110 25112
rect 18877 25109 18889 25112
rect 18923 25109 18935 25143
rect 18877 25103 18935 25109
rect 19889 25143 19947 25149
rect 19889 25109 19901 25143
rect 19935 25109 19947 25143
rect 22066 25112 22100 25152
rect 19889 25103 19947 25109
rect 22094 25100 22100 25112
rect 22152 25100 22158 25152
rect 22189 25143 22247 25149
rect 22189 25109 22201 25143
rect 22235 25140 22247 25143
rect 22554 25140 22560 25152
rect 22235 25112 22560 25140
rect 22235 25109 22247 25112
rect 22189 25103 22247 25109
rect 22554 25100 22560 25112
rect 22612 25100 22618 25152
rect 22756 25149 22784 25248
rect 22833 25245 22845 25248
rect 22879 25245 22891 25279
rect 24394 25276 24400 25288
rect 24355 25248 24400 25276
rect 22833 25239 22891 25245
rect 24394 25236 24400 25248
rect 24452 25236 24458 25288
rect 22741 25143 22799 25149
rect 22741 25109 22753 25143
rect 22787 25109 22799 25143
rect 22741 25103 22799 25109
rect 1104 25050 29532 25072
rect 1104 24998 10425 25050
rect 10477 24998 10489 25050
rect 10541 24998 10553 25050
rect 10605 24998 10617 25050
rect 10669 24998 10681 25050
rect 10733 24998 19901 25050
rect 19953 24998 19965 25050
rect 20017 24998 20029 25050
rect 20081 24998 20093 25050
rect 20145 24998 20157 25050
rect 20209 24998 29532 25050
rect 1104 24976 29532 24998
rect 9858 24896 9864 24948
rect 9916 24936 9922 24948
rect 10318 24936 10324 24948
rect 9916 24908 10324 24936
rect 9916 24896 9922 24908
rect 10318 24896 10324 24908
rect 10376 24896 10382 24948
rect 12713 24939 12771 24945
rect 12713 24905 12725 24939
rect 12759 24936 12771 24939
rect 13078 24936 13084 24948
rect 12759 24908 13084 24936
rect 12759 24905 12771 24908
rect 12713 24899 12771 24905
rect 13078 24896 13084 24908
rect 13136 24896 13142 24948
rect 16574 24896 16580 24948
rect 16632 24936 16638 24948
rect 16669 24939 16727 24945
rect 16669 24936 16681 24939
rect 16632 24908 16681 24936
rect 16632 24896 16638 24908
rect 16669 24905 16681 24908
rect 16715 24905 16727 24939
rect 16669 24899 16727 24905
rect 19794 24896 19800 24948
rect 19852 24936 19858 24948
rect 22097 24939 22155 24945
rect 22097 24936 22109 24939
rect 19852 24908 22109 24936
rect 19852 24896 19858 24908
rect 22097 24905 22109 24908
rect 22143 24905 22155 24939
rect 22097 24899 22155 24905
rect 2682 24828 2688 24880
rect 2740 24828 2746 24880
rect 4154 24828 4160 24880
rect 4212 24868 4218 24880
rect 4614 24868 4620 24880
rect 4212 24840 4620 24868
rect 4212 24828 4218 24840
rect 4614 24828 4620 24840
rect 4672 24868 4678 24880
rect 4672 24840 5304 24868
rect 4672 24828 4678 24840
rect 3881 24803 3939 24809
rect 3881 24769 3893 24803
rect 3927 24769 3939 24803
rect 3881 24763 3939 24769
rect 4525 24803 4583 24809
rect 4525 24769 4537 24803
rect 4571 24769 4583 24803
rect 5276 24800 5304 24840
rect 8864 24840 9628 24868
rect 5534 24800 5540 24812
rect 5276 24772 5540 24800
rect 4525 24763 4583 24769
rect 1394 24692 1400 24744
rect 1452 24732 1458 24744
rect 1765 24735 1823 24741
rect 1765 24732 1777 24735
rect 1452 24704 1777 24732
rect 1452 24692 1458 24704
rect 1765 24701 1777 24704
rect 1811 24701 1823 24735
rect 1765 24695 1823 24701
rect 2041 24735 2099 24741
rect 2041 24701 2053 24735
rect 2087 24732 2099 24735
rect 3694 24732 3700 24744
rect 2087 24704 3556 24732
rect 3655 24704 3700 24732
rect 2087 24701 2099 24704
rect 2041 24695 2099 24701
rect 3528 24664 3556 24704
rect 3694 24692 3700 24704
rect 3752 24692 3758 24744
rect 3896 24732 3924 24763
rect 3970 24732 3976 24744
rect 3883 24704 3976 24732
rect 3970 24692 3976 24704
rect 4028 24732 4034 24744
rect 4433 24735 4491 24741
rect 4433 24732 4445 24735
rect 4028 24704 4445 24732
rect 4028 24692 4034 24704
rect 4433 24701 4445 24704
rect 4479 24701 4491 24735
rect 4433 24695 4491 24701
rect 4249 24667 4307 24673
rect 4249 24664 4261 24667
rect 3528 24636 4261 24664
rect 4249 24633 4261 24636
rect 4295 24633 4307 24667
rect 4249 24627 4307 24633
rect 3513 24599 3571 24605
rect 3513 24565 3525 24599
rect 3559 24596 3571 24599
rect 3694 24596 3700 24608
rect 3559 24568 3700 24596
rect 3559 24565 3571 24568
rect 3513 24559 3571 24565
rect 3694 24556 3700 24568
rect 3752 24556 3758 24608
rect 4540 24596 4568 24763
rect 5534 24760 5540 24772
rect 5592 24800 5598 24812
rect 6638 24809 6644 24812
rect 6365 24803 6423 24809
rect 6365 24800 6377 24803
rect 5592 24772 6377 24800
rect 5592 24760 5598 24772
rect 6365 24769 6377 24772
rect 6411 24769 6423 24803
rect 6365 24763 6423 24769
rect 6632 24763 6644 24809
rect 6696 24800 6702 24812
rect 6696 24772 6732 24800
rect 6638 24760 6644 24763
rect 6696 24760 6702 24772
rect 6914 24760 6920 24812
rect 6972 24800 6978 24812
rect 8864 24800 8892 24840
rect 6972 24772 8892 24800
rect 8932 24803 8990 24809
rect 6972 24760 6978 24772
rect 8932 24769 8944 24803
rect 8978 24800 8990 24803
rect 9490 24800 9496 24812
rect 8978 24772 9496 24800
rect 8978 24769 8990 24772
rect 8932 24763 8990 24769
rect 9490 24760 9496 24772
rect 9548 24760 9554 24812
rect 9600 24800 9628 24840
rect 12250 24828 12256 24880
rect 12308 24868 12314 24880
rect 12345 24871 12403 24877
rect 12345 24868 12357 24871
rect 12308 24840 12357 24868
rect 12308 24828 12314 24840
rect 12345 24837 12357 24840
rect 12391 24837 12403 24871
rect 12345 24831 12403 24837
rect 13446 24828 13452 24880
rect 13504 24868 13510 24880
rect 14550 24868 14556 24880
rect 13504 24840 14556 24868
rect 13504 24828 13510 24840
rect 14550 24828 14556 24840
rect 14608 24828 14614 24880
rect 14642 24828 14648 24880
rect 14700 24868 14706 24880
rect 14700 24840 14745 24868
rect 14700 24828 14706 24840
rect 14918 24828 14924 24880
rect 14976 24868 14982 24880
rect 14976 24840 15332 24868
rect 14976 24828 14982 24840
rect 10318 24800 10324 24812
rect 9600 24772 9720 24800
rect 10279 24772 10324 24800
rect 8662 24732 8668 24744
rect 8623 24704 8668 24732
rect 8662 24692 8668 24704
rect 8720 24692 8726 24744
rect 9692 24732 9720 24772
rect 10318 24760 10324 24772
rect 10376 24760 10382 24812
rect 14369 24803 14427 24809
rect 10428 24772 12434 24800
rect 10428 24732 10456 24772
rect 9692 24704 10456 24732
rect 11330 24692 11336 24744
rect 11388 24732 11394 24744
rect 12066 24732 12072 24744
rect 11388 24704 12072 24732
rect 11388 24692 11394 24704
rect 12066 24692 12072 24704
rect 12124 24692 12130 24744
rect 12253 24735 12311 24741
rect 12253 24701 12265 24735
rect 12299 24701 12311 24735
rect 12253 24695 12311 24701
rect 7576 24636 8708 24664
rect 7576 24596 7604 24636
rect 7742 24596 7748 24608
rect 4540 24568 7604 24596
rect 7703 24568 7748 24596
rect 7742 24556 7748 24568
rect 7800 24556 7806 24608
rect 8680 24596 8708 24636
rect 9674 24624 9680 24676
rect 9732 24664 9738 24676
rect 10045 24667 10103 24673
rect 10045 24664 10057 24667
rect 9732 24636 10057 24664
rect 9732 24624 9738 24636
rect 10045 24633 10057 24636
rect 10091 24664 10103 24667
rect 10226 24664 10232 24676
rect 10091 24636 10232 24664
rect 10091 24633 10103 24636
rect 10045 24627 10103 24633
rect 10226 24624 10232 24636
rect 10284 24624 10290 24676
rect 10505 24667 10563 24673
rect 10505 24633 10517 24667
rect 10551 24664 10563 24667
rect 10594 24664 10600 24676
rect 10551 24636 10600 24664
rect 10551 24633 10563 24636
rect 10505 24627 10563 24633
rect 10594 24624 10600 24636
rect 10652 24624 10658 24676
rect 11422 24624 11428 24676
rect 11480 24664 11486 24676
rect 12268 24664 12296 24695
rect 11480 24636 12296 24664
rect 12406 24664 12434 24772
rect 14369 24769 14381 24803
rect 14415 24800 14427 24803
rect 14789 24803 14847 24809
rect 14415 24772 14504 24800
rect 14415 24769 14427 24772
rect 14369 24763 14427 24769
rect 14366 24664 14372 24676
rect 12406 24636 14372 24664
rect 11480 24624 11486 24636
rect 14366 24624 14372 24636
rect 14424 24624 14430 24676
rect 8846 24596 8852 24608
rect 8680 24568 8852 24596
rect 8846 24556 8852 24568
rect 8904 24556 8910 24608
rect 14476 24596 14504 24772
rect 14789 24769 14801 24803
rect 14835 24769 14847 24803
rect 14789 24763 14847 24769
rect 14804 24732 14832 24763
rect 15102 24760 15108 24812
rect 15160 24800 15166 24812
rect 15304 24809 15332 24840
rect 15396 24840 15792 24868
rect 15396 24809 15424 24840
rect 15289 24803 15347 24809
rect 15160 24772 15205 24800
rect 15160 24760 15166 24772
rect 15289 24769 15301 24803
rect 15335 24769 15347 24803
rect 15289 24763 15347 24769
rect 15381 24803 15439 24809
rect 15381 24769 15393 24803
rect 15427 24769 15439 24803
rect 15381 24763 15439 24769
rect 15478 24803 15536 24809
rect 15478 24769 15490 24803
rect 15524 24800 15536 24803
rect 15654 24800 15660 24812
rect 15524 24772 15660 24800
rect 15524 24769 15536 24772
rect 15478 24763 15536 24769
rect 15493 24732 15521 24763
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 15764 24800 15792 24840
rect 22554 24828 22560 24880
rect 22612 24868 22618 24880
rect 22612 24840 24440 24868
rect 22612 24828 22618 24840
rect 16206 24800 16212 24812
rect 15764 24772 16212 24800
rect 16206 24760 16212 24772
rect 16264 24760 16270 24812
rect 16666 24760 16672 24812
rect 16724 24800 16730 24812
rect 16853 24803 16911 24809
rect 16853 24800 16865 24803
rect 16724 24772 16865 24800
rect 16724 24760 16730 24772
rect 16853 24769 16865 24772
rect 16899 24769 16911 24803
rect 18046 24800 18052 24812
rect 16853 24763 16911 24769
rect 17788 24772 18052 24800
rect 14804 24704 15521 24732
rect 16224 24732 16252 24760
rect 17788 24732 17816 24772
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 18230 24809 18236 24812
rect 18224 24800 18236 24809
rect 18191 24772 18236 24800
rect 18224 24763 18236 24772
rect 18230 24760 18236 24763
rect 18288 24760 18294 24812
rect 19702 24760 19708 24812
rect 19760 24800 19766 24812
rect 19797 24803 19855 24809
rect 19797 24800 19809 24803
rect 19760 24772 19809 24800
rect 19760 24760 19766 24772
rect 19797 24769 19809 24772
rect 19843 24769 19855 24803
rect 19797 24763 19855 24769
rect 19889 24803 19947 24809
rect 19889 24769 19901 24803
rect 19935 24769 19947 24803
rect 19889 24763 19947 24769
rect 20901 24803 20959 24809
rect 20901 24769 20913 24803
rect 20947 24769 20959 24803
rect 20901 24763 20959 24769
rect 20993 24803 21051 24809
rect 20993 24769 21005 24803
rect 21039 24800 21051 24803
rect 21361 24803 21419 24809
rect 21361 24800 21373 24803
rect 21039 24772 21373 24800
rect 21039 24769 21051 24772
rect 20993 24763 21051 24769
rect 21361 24769 21373 24772
rect 21407 24769 21419 24803
rect 21361 24763 21419 24769
rect 16224 24704 17816 24732
rect 17954 24692 17960 24744
rect 18012 24732 18018 24744
rect 18012 24704 18057 24732
rect 18012 24692 18018 24704
rect 14921 24667 14979 24673
rect 14921 24633 14933 24667
rect 14967 24664 14979 24667
rect 15470 24664 15476 24676
rect 14967 24636 15476 24664
rect 14967 24633 14979 24636
rect 14921 24627 14979 24633
rect 15470 24624 15476 24636
rect 15528 24624 15534 24676
rect 15657 24667 15715 24673
rect 15657 24633 15669 24667
rect 15703 24664 15715 24667
rect 17402 24664 17408 24676
rect 15703 24636 17408 24664
rect 15703 24633 15715 24636
rect 15657 24627 15715 24633
rect 17402 24624 17408 24636
rect 17460 24624 17466 24676
rect 19337 24667 19395 24673
rect 19337 24633 19349 24667
rect 19383 24664 19395 24667
rect 19426 24664 19432 24676
rect 19383 24636 19432 24664
rect 19383 24633 19395 24636
rect 19337 24627 19395 24633
rect 19426 24624 19432 24636
rect 19484 24664 19490 24676
rect 19904 24664 19932 24763
rect 20916 24732 20944 24763
rect 21266 24732 21272 24744
rect 20916 24704 21272 24732
rect 21266 24692 21272 24704
rect 21324 24692 21330 24744
rect 21376 24732 21404 24763
rect 21450 24760 21456 24812
rect 21508 24800 21514 24812
rect 21821 24803 21879 24809
rect 21508 24772 21553 24800
rect 21508 24760 21514 24772
rect 21821 24769 21833 24803
rect 21867 24769 21879 24803
rect 21821 24763 21879 24769
rect 21836 24732 21864 24763
rect 22186 24760 22192 24812
rect 22244 24800 22250 24812
rect 23216 24809 23244 24840
rect 24412 24812 24440 24840
rect 22281 24803 22339 24809
rect 22281 24800 22293 24803
rect 22244 24772 22293 24800
rect 22244 24760 22250 24772
rect 22281 24769 22293 24772
rect 22327 24769 22339 24803
rect 22281 24763 22339 24769
rect 23201 24803 23259 24809
rect 23201 24769 23213 24803
rect 23247 24769 23259 24803
rect 23477 24803 23535 24809
rect 23477 24800 23489 24803
rect 23201 24763 23259 24769
rect 23400 24772 23489 24800
rect 21376 24704 21864 24732
rect 21634 24664 21640 24676
rect 19484 24636 19932 24664
rect 21595 24636 21640 24664
rect 19484 24624 19490 24636
rect 21634 24624 21640 24636
rect 21692 24624 21698 24676
rect 21726 24624 21732 24676
rect 21784 24664 21790 24676
rect 22002 24664 22008 24676
rect 21784 24636 22008 24664
rect 21784 24624 21790 24636
rect 22002 24624 22008 24636
rect 22060 24624 22066 24676
rect 23400 24673 23428 24772
rect 23477 24769 23489 24772
rect 23523 24769 23535 24803
rect 23477 24763 23535 24769
rect 24394 24760 24400 24812
rect 24452 24800 24458 24812
rect 24857 24803 24915 24809
rect 24857 24800 24869 24803
rect 24452 24772 24869 24800
rect 24452 24760 24458 24772
rect 24857 24769 24869 24772
rect 24903 24769 24915 24803
rect 25133 24803 25191 24809
rect 25133 24800 25145 24803
rect 24857 24763 24915 24769
rect 24964 24772 25145 24800
rect 24486 24692 24492 24744
rect 24544 24732 24550 24744
rect 24964 24732 24992 24772
rect 25133 24769 25145 24772
rect 25179 24769 25191 24803
rect 25133 24763 25191 24769
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24769 25743 24803
rect 25685 24763 25743 24769
rect 25700 24732 25728 24763
rect 24544 24704 24992 24732
rect 25056 24704 25728 24732
rect 24544 24692 24550 24704
rect 25056 24673 25084 24704
rect 23385 24667 23443 24673
rect 23385 24633 23397 24667
rect 23431 24633 23443 24667
rect 23385 24627 23443 24633
rect 25041 24667 25099 24673
rect 25041 24633 25053 24667
rect 25087 24633 25099 24667
rect 25041 24627 25099 24633
rect 15010 24596 15016 24608
rect 14476 24568 15016 24596
rect 15010 24556 15016 24568
rect 15068 24556 15074 24608
rect 17678 24556 17684 24608
rect 17736 24596 17742 24608
rect 19242 24596 19248 24608
rect 17736 24568 19248 24596
rect 17736 24556 17742 24568
rect 19242 24556 19248 24568
rect 19300 24596 19306 24608
rect 19613 24599 19671 24605
rect 19613 24596 19625 24599
rect 19300 24568 19625 24596
rect 19300 24556 19306 24568
rect 19613 24565 19625 24568
rect 19659 24565 19671 24599
rect 19613 24559 19671 24565
rect 20073 24599 20131 24605
rect 20073 24565 20085 24599
rect 20119 24596 20131 24599
rect 20254 24596 20260 24608
rect 20119 24568 20260 24596
rect 20119 24565 20131 24568
rect 20073 24559 20131 24565
rect 20254 24556 20260 24568
rect 20312 24556 20318 24608
rect 20898 24556 20904 24608
rect 20956 24596 20962 24608
rect 21177 24599 21235 24605
rect 21177 24596 21189 24599
rect 20956 24568 21189 24596
rect 20956 24556 20962 24568
rect 21177 24565 21189 24568
rect 21223 24565 21235 24599
rect 21177 24559 21235 24565
rect 21910 24556 21916 24608
rect 21968 24596 21974 24608
rect 22373 24599 22431 24605
rect 22373 24596 22385 24599
rect 21968 24568 22385 24596
rect 21968 24556 21974 24568
rect 22373 24565 22385 24568
rect 22419 24565 22431 24599
rect 22373 24559 22431 24565
rect 23661 24599 23719 24605
rect 23661 24565 23673 24599
rect 23707 24596 23719 24599
rect 23750 24596 23756 24608
rect 23707 24568 23756 24596
rect 23707 24565 23719 24568
rect 23661 24559 23719 24565
rect 23750 24556 23756 24568
rect 23808 24556 23814 24608
rect 25314 24596 25320 24608
rect 25275 24568 25320 24596
rect 25314 24556 25320 24568
rect 25372 24556 25378 24608
rect 25866 24596 25872 24608
rect 25827 24568 25872 24596
rect 25866 24556 25872 24568
rect 25924 24556 25930 24608
rect 1104 24506 29532 24528
rect 1104 24454 5688 24506
rect 5740 24454 5752 24506
rect 5804 24454 5816 24506
rect 5868 24454 5880 24506
rect 5932 24454 5944 24506
rect 5996 24454 15163 24506
rect 15215 24454 15227 24506
rect 15279 24454 15291 24506
rect 15343 24454 15355 24506
rect 15407 24454 15419 24506
rect 15471 24454 24639 24506
rect 24691 24454 24703 24506
rect 24755 24454 24767 24506
rect 24819 24454 24831 24506
rect 24883 24454 24895 24506
rect 24947 24454 29532 24506
rect 1104 24432 29532 24454
rect 2682 24392 2688 24404
rect 2643 24364 2688 24392
rect 2682 24352 2688 24364
rect 2740 24352 2746 24404
rect 5813 24395 5871 24401
rect 5813 24361 5825 24395
rect 5859 24392 5871 24395
rect 6086 24392 6092 24404
rect 5859 24364 6092 24392
rect 5859 24361 5871 24364
rect 5813 24355 5871 24361
rect 6086 24352 6092 24364
rect 6144 24352 6150 24404
rect 6362 24392 6368 24404
rect 6323 24364 6368 24392
rect 6362 24352 6368 24364
rect 6420 24352 6426 24404
rect 6549 24395 6607 24401
rect 6549 24361 6561 24395
rect 6595 24392 6607 24395
rect 6638 24392 6644 24404
rect 6595 24364 6644 24392
rect 6595 24361 6607 24364
rect 6549 24355 6607 24361
rect 6638 24352 6644 24364
rect 6696 24352 6702 24404
rect 8294 24352 8300 24404
rect 8352 24392 8358 24404
rect 8665 24395 8723 24401
rect 8665 24392 8677 24395
rect 8352 24364 8677 24392
rect 8352 24352 8358 24364
rect 8665 24361 8677 24364
rect 8711 24392 8723 24395
rect 8757 24395 8815 24401
rect 8757 24392 8769 24395
rect 8711 24364 8769 24392
rect 8711 24361 8723 24364
rect 8665 24355 8723 24361
rect 8757 24361 8769 24364
rect 8803 24361 8815 24395
rect 8757 24355 8815 24361
rect 9490 24352 9496 24404
rect 9548 24392 9554 24404
rect 9585 24395 9643 24401
rect 9585 24392 9597 24395
rect 9548 24364 9597 24392
rect 9548 24352 9554 24364
rect 9585 24361 9597 24364
rect 9631 24361 9643 24395
rect 10042 24392 10048 24404
rect 9955 24364 10048 24392
rect 9585 24355 9643 24361
rect 2409 24327 2467 24333
rect 2409 24293 2421 24327
rect 2455 24293 2467 24327
rect 9766 24324 9772 24336
rect 2409 24287 2467 24293
rect 6196 24296 9772 24324
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2314 24188 2320 24200
rect 2271 24160 2320 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2314 24148 2320 24160
rect 2372 24148 2378 24200
rect 2424 24188 2452 24287
rect 6196 24197 6224 24296
rect 7742 24256 7748 24268
rect 6656 24228 7748 24256
rect 6656 24197 6684 24228
rect 7742 24216 7748 24228
rect 7800 24216 7806 24268
rect 2501 24191 2559 24197
rect 2501 24188 2513 24191
rect 2424 24160 2513 24188
rect 2501 24157 2513 24160
rect 2547 24157 2559 24191
rect 2501 24151 2559 24157
rect 5997 24191 6055 24197
rect 5997 24157 6009 24191
rect 6043 24188 6055 24191
rect 6181 24191 6239 24197
rect 6181 24188 6193 24191
rect 6043 24160 6193 24188
rect 6043 24157 6055 24160
rect 5997 24151 6055 24157
rect 6181 24157 6193 24160
rect 6227 24157 6239 24191
rect 6181 24151 6239 24157
rect 6641 24191 6699 24197
rect 6641 24157 6653 24191
rect 6687 24157 6699 24191
rect 6822 24188 6828 24200
rect 6783 24160 6828 24188
rect 6641 24151 6699 24157
rect 6822 24148 6828 24160
rect 6880 24148 6886 24200
rect 6917 24191 6975 24197
rect 6917 24157 6929 24191
rect 6963 24157 6975 24191
rect 6917 24151 6975 24157
rect 7027 24191 7085 24197
rect 7027 24157 7039 24191
rect 7073 24188 7085 24191
rect 7193 24191 7251 24197
rect 7073 24160 7144 24188
rect 7073 24157 7085 24160
rect 7027 24151 7085 24157
rect 6362 24080 6368 24132
rect 6420 24120 6426 24132
rect 6730 24120 6736 24132
rect 6420 24092 6736 24120
rect 6420 24080 6426 24092
rect 6730 24080 6736 24092
rect 6788 24120 6794 24132
rect 6932 24120 6960 24151
rect 6788 24092 6960 24120
rect 7116 24120 7144 24160
rect 7193 24157 7205 24191
rect 7239 24188 7251 24191
rect 8490 24191 8548 24197
rect 7239 24160 7788 24188
rect 7239 24157 7251 24160
rect 7193 24151 7251 24157
rect 7760 24120 7788 24160
rect 8490 24157 8502 24191
rect 8536 24185 8548 24191
rect 8588 24185 8616 24296
rect 9766 24284 9772 24296
rect 9824 24284 9830 24336
rect 8757 24259 8815 24265
rect 8757 24225 8769 24259
rect 8803 24256 8815 24259
rect 9214 24256 9220 24268
rect 8803 24228 9220 24256
rect 8803 24225 8815 24228
rect 8757 24219 8815 24225
rect 9214 24216 9220 24228
rect 9272 24216 9278 24268
rect 9306 24216 9312 24268
rect 9364 24256 9370 24268
rect 9364 24228 9409 24256
rect 9364 24216 9370 24228
rect 9582 24216 9588 24268
rect 9640 24256 9646 24268
rect 9640 24228 9904 24256
rect 9640 24216 9646 24228
rect 8536 24157 8616 24185
rect 8680 24184 8892 24188
rect 8938 24184 8944 24200
rect 8680 24160 8944 24184
rect 8490 24151 8548 24157
rect 8680 24120 8708 24160
rect 8855 24156 8944 24160
rect 8938 24148 8944 24156
rect 8996 24148 9002 24200
rect 9048 24197 9168 24198
rect 8938 24143 8996 24148
rect 9030 24145 9036 24197
rect 9088 24191 9182 24197
rect 9088 24170 9136 24191
rect 9088 24145 9094 24170
rect 9124 24157 9136 24170
rect 9170 24157 9182 24191
rect 9124 24151 9182 24157
rect 9493 24191 9551 24197
rect 9493 24157 9505 24191
rect 9539 24188 9551 24191
rect 9674 24188 9680 24200
rect 9539 24160 9680 24188
rect 9539 24157 9551 24160
rect 9493 24151 9551 24157
rect 9674 24148 9680 24160
rect 9732 24148 9738 24200
rect 7116 24092 7420 24120
rect 7760 24092 8708 24120
rect 9876 24120 9904 24228
rect 9968 24197 9996 24364
rect 10042 24352 10048 24364
rect 10100 24392 10106 24404
rect 10778 24392 10784 24404
rect 10100 24364 10784 24392
rect 10100 24352 10106 24364
rect 10778 24352 10784 24364
rect 10836 24352 10842 24404
rect 11422 24392 11428 24404
rect 11383 24364 11428 24392
rect 11422 24352 11428 24364
rect 11480 24352 11486 24404
rect 14366 24352 14372 24404
rect 14424 24392 14430 24404
rect 16666 24392 16672 24404
rect 14424 24364 16528 24392
rect 16627 24364 16672 24392
rect 14424 24352 14430 24364
rect 13817 24327 13875 24333
rect 13817 24293 13829 24327
rect 13863 24324 13875 24327
rect 14458 24324 14464 24336
rect 13863 24296 14464 24324
rect 13863 24293 13875 24296
rect 13817 24287 13875 24293
rect 14458 24284 14464 24296
rect 14516 24284 14522 24336
rect 16500 24324 16528 24364
rect 16666 24352 16672 24364
rect 16724 24352 16730 24404
rect 18230 24352 18236 24404
rect 18288 24392 18294 24404
rect 18325 24395 18383 24401
rect 18325 24392 18337 24395
rect 18288 24364 18337 24392
rect 18288 24352 18294 24364
rect 18325 24361 18337 24364
rect 18371 24361 18383 24395
rect 21910 24392 21916 24404
rect 18325 24355 18383 24361
rect 19720 24364 21916 24392
rect 19720 24324 19748 24364
rect 21910 24352 21916 24364
rect 21968 24392 21974 24404
rect 24121 24395 24179 24401
rect 24121 24392 24133 24395
rect 21968 24364 24133 24392
rect 21968 24352 21974 24364
rect 24121 24361 24133 24364
rect 24167 24361 24179 24395
rect 24121 24355 24179 24361
rect 26142 24352 26148 24404
rect 26200 24392 26206 24404
rect 26878 24392 26884 24404
rect 26200 24364 26884 24392
rect 26200 24352 26206 24364
rect 26878 24352 26884 24364
rect 26936 24352 26942 24404
rect 27430 24352 27436 24404
rect 27488 24392 27494 24404
rect 29089 24395 29147 24401
rect 29089 24392 29101 24395
rect 27488 24364 29101 24392
rect 27488 24352 27494 24364
rect 29089 24361 29101 24364
rect 29135 24361 29147 24395
rect 29089 24355 29147 24361
rect 16500 24296 19748 24324
rect 14185 24259 14243 24265
rect 14185 24256 14197 24259
rect 13188 24228 14197 24256
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24157 10011 24191
rect 9953 24151 10011 24157
rect 10045 24191 10103 24197
rect 10045 24157 10057 24191
rect 10091 24188 10103 24191
rect 10594 24188 10600 24200
rect 10091 24160 10600 24188
rect 10091 24157 10103 24160
rect 10045 24151 10103 24157
rect 10060 24120 10088 24151
rect 10594 24148 10600 24160
rect 10652 24188 10658 24200
rect 11609 24191 11667 24197
rect 11609 24188 11621 24191
rect 10652 24160 11621 24188
rect 10652 24148 10658 24160
rect 11609 24157 11621 24160
rect 11655 24157 11667 24191
rect 13188 24188 13216 24228
rect 14185 24225 14197 24228
rect 14231 24225 14243 24259
rect 14918 24256 14924 24268
rect 14185 24219 14243 24225
rect 14384 24228 14924 24256
rect 11609 24151 11667 24157
rect 11716 24160 13216 24188
rect 13265 24191 13323 24197
rect 9876 24092 10088 24120
rect 10312 24123 10370 24129
rect 6788 24080 6794 24092
rect 7392 24064 7420 24092
rect 10312 24089 10324 24123
rect 10358 24120 10370 24123
rect 10778 24120 10784 24132
rect 10358 24092 10784 24120
rect 10358 24089 10370 24092
rect 10312 24083 10370 24089
rect 10778 24080 10784 24092
rect 10836 24080 10842 24132
rect 4062 24012 4068 24064
rect 4120 24052 4126 24064
rect 6914 24052 6920 24064
rect 4120 24024 6920 24052
rect 4120 24012 4126 24024
rect 6914 24012 6920 24024
rect 6972 24012 6978 24064
rect 7374 24052 7380 24064
rect 7335 24024 7380 24052
rect 7374 24012 7380 24024
rect 7432 24012 7438 24064
rect 8389 24055 8447 24061
rect 8389 24021 8401 24055
rect 8435 24052 8447 24055
rect 8478 24052 8484 24064
rect 8435 24024 8484 24052
rect 8435 24021 8447 24024
rect 8389 24015 8447 24021
rect 8478 24012 8484 24024
rect 8536 24012 8542 24064
rect 8846 24012 8852 24064
rect 8904 24052 8910 24064
rect 11716 24052 11744 24160
rect 13265 24157 13277 24191
rect 13311 24157 13323 24191
rect 13446 24188 13452 24200
rect 13407 24160 13452 24188
rect 13265 24151 13323 24157
rect 11876 24123 11934 24129
rect 11876 24089 11888 24123
rect 11922 24120 11934 24123
rect 12158 24120 12164 24132
rect 11922 24092 12164 24120
rect 11922 24089 11934 24092
rect 11876 24083 11934 24089
rect 12158 24080 12164 24092
rect 12216 24080 12222 24132
rect 8904 24024 11744 24052
rect 8904 24012 8910 24024
rect 12250 24012 12256 24064
rect 12308 24052 12314 24064
rect 12989 24055 13047 24061
rect 12989 24052 13001 24055
rect 12308 24024 13001 24052
rect 12308 24012 12314 24024
rect 12989 24021 13001 24024
rect 13035 24021 13047 24055
rect 13280 24052 13308 24151
rect 13446 24148 13452 24160
rect 13504 24148 13510 24200
rect 13685 24191 13743 24197
rect 13685 24157 13697 24191
rect 13731 24188 13743 24191
rect 13906 24188 13912 24200
rect 13731 24160 13912 24188
rect 13731 24157 13743 24160
rect 13685 24151 13743 24157
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 14090 24188 14096 24200
rect 14051 24160 14096 24188
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 14384 24197 14412 24228
rect 14918 24216 14924 24228
rect 14976 24216 14982 24268
rect 18230 24216 18236 24268
rect 18288 24256 18294 24268
rect 18509 24259 18567 24265
rect 18509 24256 18521 24259
rect 18288 24228 18521 24256
rect 18288 24216 18294 24228
rect 18509 24225 18521 24228
rect 18555 24256 18567 24259
rect 19705 24259 19763 24265
rect 19705 24256 19717 24259
rect 18555 24228 19717 24256
rect 18555 24225 18567 24228
rect 18509 24219 18567 24225
rect 19705 24225 19717 24228
rect 19751 24225 19763 24259
rect 19705 24219 19763 24225
rect 14369 24191 14427 24197
rect 14369 24157 14381 24191
rect 14415 24157 14427 24191
rect 14369 24151 14427 24157
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24157 14611 24191
rect 14826 24188 14832 24200
rect 14787 24160 14832 24188
rect 14553 24151 14611 24157
rect 13538 24080 13544 24132
rect 13596 24120 13602 24132
rect 14568 24120 14596 24151
rect 14826 24148 14832 24160
rect 14884 24148 14890 24200
rect 13596 24092 14596 24120
rect 14936 24120 14964 24216
rect 16485 24191 16543 24197
rect 16485 24157 16497 24191
rect 16531 24188 16543 24191
rect 16666 24188 16672 24200
rect 16531 24160 16672 24188
rect 16531 24157 16543 24160
rect 16485 24151 16543 24157
rect 16666 24148 16672 24160
rect 16724 24148 16730 24200
rect 17402 24148 17408 24200
rect 17460 24188 17466 24200
rect 17773 24191 17831 24197
rect 17773 24188 17785 24191
rect 17460 24160 17785 24188
rect 17460 24148 17466 24160
rect 17773 24157 17785 24160
rect 17819 24157 17831 24191
rect 17773 24151 17831 24157
rect 17862 24148 17868 24200
rect 17920 24188 17926 24200
rect 18146 24191 18204 24197
rect 18146 24188 18158 24191
rect 17920 24160 18158 24188
rect 17920 24148 17926 24160
rect 18146 24157 18158 24160
rect 18192 24157 18204 24191
rect 18690 24188 18696 24200
rect 18651 24160 18696 24188
rect 18146 24151 18204 24157
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 19061 24191 19119 24197
rect 19061 24157 19073 24191
rect 19107 24188 19119 24191
rect 19426 24188 19432 24200
rect 19107 24160 19432 24188
rect 19107 24157 19119 24160
rect 19061 24151 19119 24157
rect 19426 24148 19432 24160
rect 19484 24148 19490 24200
rect 21358 24148 21364 24200
rect 21416 24188 21422 24200
rect 21453 24191 21511 24197
rect 21453 24188 21465 24191
rect 21416 24160 21465 24188
rect 21416 24148 21422 24160
rect 21453 24157 21465 24160
rect 21499 24157 21511 24191
rect 21453 24151 21511 24157
rect 21637 24191 21695 24197
rect 21637 24157 21649 24191
rect 21683 24188 21695 24191
rect 21726 24188 21732 24200
rect 21683 24160 21732 24188
rect 21683 24157 21695 24160
rect 21637 24151 21695 24157
rect 21726 24148 21732 24160
rect 21784 24148 21790 24200
rect 17678 24120 17684 24132
rect 14936 24092 17684 24120
rect 13596 24080 13602 24092
rect 17678 24080 17684 24092
rect 17736 24120 17742 24132
rect 17957 24123 18015 24129
rect 17957 24120 17969 24123
rect 17736 24092 17969 24120
rect 17736 24080 17742 24092
rect 17957 24089 17969 24092
rect 18003 24089 18015 24123
rect 17957 24083 18015 24089
rect 18049 24123 18107 24129
rect 18049 24089 18061 24123
rect 18095 24120 18107 24123
rect 18095 24092 18920 24120
rect 18095 24089 18107 24092
rect 18049 24083 18107 24089
rect 14090 24052 14096 24064
rect 13280 24024 14096 24052
rect 12989 24015 13047 24021
rect 14090 24012 14096 24024
rect 14148 24012 14154 24064
rect 14550 24012 14556 24064
rect 14608 24052 14614 24064
rect 18064 24052 18092 24083
rect 18138 24052 18144 24064
rect 14608 24024 18144 24052
rect 14608 24012 14614 24024
rect 18138 24012 18144 24024
rect 18196 24012 18202 24064
rect 18892 24061 18920 24092
rect 19794 24080 19800 24132
rect 19852 24120 19858 24132
rect 19950 24123 20008 24129
rect 19950 24120 19962 24123
rect 19852 24092 19962 24120
rect 19852 24080 19858 24092
rect 19950 24089 19962 24092
rect 19996 24089 20008 24123
rect 21818 24120 21824 24132
rect 21779 24092 21824 24120
rect 19950 24083 20008 24089
rect 21818 24080 21824 24092
rect 21876 24080 21882 24132
rect 21928 24129 21956 24352
rect 22002 24284 22008 24336
rect 22060 24324 22066 24336
rect 22189 24327 22247 24333
rect 22060 24284 22094 24324
rect 22189 24293 22201 24327
rect 22235 24324 22247 24327
rect 26421 24327 26479 24333
rect 26421 24324 26433 24327
rect 22235 24296 22508 24324
rect 22235 24293 22247 24296
rect 22189 24287 22247 24293
rect 22066 24256 22094 24284
rect 22373 24259 22431 24265
rect 22373 24256 22385 24259
rect 22066 24228 22385 24256
rect 22373 24225 22385 24228
rect 22419 24225 22431 24259
rect 22480 24256 22508 24296
rect 26206 24296 26433 24324
rect 22649 24259 22707 24265
rect 22649 24256 22661 24259
rect 22480 24228 22661 24256
rect 22373 24219 22431 24225
rect 22649 24225 22661 24228
rect 22695 24225 22707 24259
rect 22649 24219 22707 24225
rect 23658 24216 23664 24268
rect 23716 24256 23722 24268
rect 24397 24259 24455 24265
rect 24397 24256 24409 24259
rect 23716 24228 24409 24256
rect 23716 24216 23722 24228
rect 24397 24225 24409 24228
rect 24443 24225 24455 24259
rect 24397 24219 24455 24225
rect 25222 24216 25228 24268
rect 25280 24256 25286 24268
rect 26206 24256 26234 24296
rect 26421 24293 26433 24296
rect 26467 24293 26479 24327
rect 26421 24287 26479 24293
rect 25280 24228 26234 24256
rect 25280 24216 25286 24228
rect 22010 24191 22068 24197
rect 22010 24157 22022 24191
rect 22056 24157 22068 24191
rect 22010 24151 22068 24157
rect 21913 24123 21971 24129
rect 21913 24089 21925 24123
rect 21959 24089 21971 24123
rect 21913 24083 21971 24089
rect 18877 24055 18935 24061
rect 18877 24021 18889 24055
rect 18923 24021 18935 24055
rect 19518 24052 19524 24064
rect 19479 24024 19524 24052
rect 18877 24015 18935 24021
rect 19518 24012 19524 24024
rect 19576 24012 19582 24064
rect 19702 24012 19708 24064
rect 19760 24052 19766 24064
rect 20622 24052 20628 24064
rect 19760 24024 20628 24052
rect 19760 24012 19766 24024
rect 20622 24012 20628 24024
rect 20680 24052 20686 24064
rect 21085 24055 21143 24061
rect 21085 24052 21097 24055
rect 20680 24024 21097 24052
rect 20680 24012 20686 24024
rect 21085 24021 21097 24024
rect 21131 24021 21143 24055
rect 21266 24052 21272 24064
rect 21227 24024 21272 24052
rect 21085 24015 21143 24021
rect 21266 24012 21272 24024
rect 21324 24052 21330 24064
rect 21542 24052 21548 24064
rect 21324 24024 21548 24052
rect 21324 24012 21330 24024
rect 21542 24012 21548 24024
rect 21600 24012 21606 24064
rect 21634 24012 21640 24064
rect 21692 24052 21698 24064
rect 22020 24052 22048 24151
rect 23750 24148 23756 24200
rect 23808 24148 23814 24200
rect 26050 24148 26056 24200
rect 26108 24188 26114 24200
rect 26553 24191 26611 24197
rect 26553 24188 26565 24191
rect 26108 24160 26565 24188
rect 26108 24148 26114 24160
rect 26553 24157 26565 24160
rect 26599 24157 26611 24191
rect 26694 24188 26700 24200
rect 26655 24160 26700 24188
rect 26553 24151 26611 24157
rect 26694 24148 26700 24160
rect 26752 24148 26758 24200
rect 26973 24191 27031 24197
rect 26973 24157 26985 24191
rect 27019 24157 27031 24191
rect 27338 24188 27344 24200
rect 27299 24160 27344 24188
rect 26973 24151 27031 24157
rect 24026 24080 24032 24132
rect 24084 24120 24090 24132
rect 24673 24123 24731 24129
rect 24673 24120 24685 24123
rect 24084 24092 24685 24120
rect 24084 24080 24090 24092
rect 24673 24089 24685 24092
rect 24719 24089 24731 24123
rect 24673 24083 24731 24089
rect 25314 24080 25320 24132
rect 25372 24080 25378 24132
rect 26786 24120 26792 24132
rect 25976 24092 26648 24120
rect 26747 24092 26792 24120
rect 21692 24024 22048 24052
rect 21692 24012 21698 24024
rect 25590 24012 25596 24064
rect 25648 24052 25654 24064
rect 25976 24052 26004 24092
rect 26142 24052 26148 24064
rect 25648 24024 26004 24052
rect 26103 24024 26148 24052
rect 25648 24012 25654 24024
rect 26142 24012 26148 24024
rect 26200 24012 26206 24064
rect 26620 24052 26648 24092
rect 26786 24080 26792 24092
rect 26844 24080 26850 24132
rect 26988 24052 27016 24151
rect 27338 24148 27344 24160
rect 27396 24148 27402 24200
rect 27614 24120 27620 24132
rect 27575 24092 27620 24120
rect 27614 24080 27620 24092
rect 27672 24080 27678 24132
rect 28626 24080 28632 24132
rect 28684 24080 28690 24132
rect 26620 24024 27016 24052
rect 27062 24012 27068 24064
rect 27120 24052 27126 24064
rect 27120 24024 27165 24052
rect 27120 24012 27126 24024
rect 1104 23962 29532 23984
rect 1104 23910 10425 23962
rect 10477 23910 10489 23962
rect 10541 23910 10553 23962
rect 10605 23910 10617 23962
rect 10669 23910 10681 23962
rect 10733 23910 19901 23962
rect 19953 23910 19965 23962
rect 20017 23910 20029 23962
rect 20081 23910 20093 23962
rect 20145 23910 20157 23962
rect 20209 23910 29532 23962
rect 1104 23888 29532 23910
rect 1394 23808 1400 23860
rect 1452 23848 1458 23860
rect 4614 23848 4620 23860
rect 1452 23820 4620 23848
rect 1452 23808 1458 23820
rect 4614 23808 4620 23820
rect 4672 23808 4678 23860
rect 5997 23851 6055 23857
rect 5997 23817 6009 23851
rect 6043 23848 6055 23851
rect 6086 23848 6092 23860
rect 6043 23820 6092 23848
rect 6043 23817 6055 23820
rect 5997 23811 6055 23817
rect 6086 23808 6092 23820
rect 6144 23848 6150 23860
rect 7193 23851 7251 23857
rect 7193 23848 7205 23851
rect 6144 23820 7205 23848
rect 6144 23808 6150 23820
rect 7193 23817 7205 23820
rect 7239 23817 7251 23851
rect 7650 23848 7656 23860
rect 7611 23820 7656 23848
rect 7193 23811 7251 23817
rect 7650 23808 7656 23820
rect 7708 23808 7714 23860
rect 8478 23808 8484 23860
rect 8536 23848 8542 23860
rect 9030 23848 9036 23860
rect 8536 23820 9036 23848
rect 8536 23808 8542 23820
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 9214 23808 9220 23860
rect 9272 23848 9278 23860
rect 11790 23848 11796 23860
rect 9272 23820 11796 23848
rect 9272 23808 9278 23820
rect 11790 23808 11796 23820
rect 11848 23808 11854 23860
rect 12158 23848 12164 23860
rect 12119 23820 12164 23848
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 14182 23808 14188 23860
rect 14240 23848 14246 23860
rect 14737 23851 14795 23857
rect 14737 23848 14749 23851
rect 14240 23820 14749 23848
rect 14240 23808 14246 23820
rect 14737 23817 14749 23820
rect 14783 23848 14795 23851
rect 15838 23848 15844 23860
rect 14783 23820 15844 23848
rect 14783 23817 14795 23820
rect 14737 23811 14795 23817
rect 15838 23808 15844 23820
rect 15896 23808 15902 23860
rect 16853 23851 16911 23857
rect 16853 23817 16865 23851
rect 16899 23817 16911 23851
rect 16853 23811 16911 23817
rect 18800 23820 19656 23848
rect 2866 23740 2872 23792
rect 2924 23740 2930 23792
rect 13725 23783 13783 23789
rect 13725 23780 13737 23783
rect 4356 23752 13737 23780
rect 3418 23672 3424 23724
rect 3476 23712 3482 23724
rect 4356 23721 4384 23752
rect 13725 23749 13737 23752
rect 13771 23749 13783 23783
rect 13725 23743 13783 23749
rect 3513 23715 3571 23721
rect 3513 23712 3525 23715
rect 3476 23684 3525 23712
rect 3476 23672 3482 23684
rect 3513 23681 3525 23684
rect 3559 23681 3571 23715
rect 3513 23675 3571 23681
rect 3697 23715 3755 23721
rect 3697 23681 3709 23715
rect 3743 23681 3755 23715
rect 3697 23675 3755 23681
rect 4341 23715 4399 23721
rect 4341 23681 4353 23715
rect 4387 23681 4399 23715
rect 4614 23712 4620 23724
rect 4575 23684 4620 23712
rect 4341 23675 4399 23681
rect 1394 23604 1400 23656
rect 1452 23644 1458 23656
rect 1581 23647 1639 23653
rect 1581 23644 1593 23647
rect 1452 23616 1593 23644
rect 1452 23604 1458 23616
rect 1581 23613 1593 23616
rect 1627 23613 1639 23647
rect 1581 23607 1639 23613
rect 1857 23647 1915 23653
rect 1857 23613 1869 23647
rect 1903 23644 1915 23647
rect 3712 23644 3740 23675
rect 4614 23672 4620 23684
rect 4672 23672 4678 23724
rect 4890 23721 4896 23724
rect 4884 23675 4896 23721
rect 4948 23712 4954 23724
rect 7282 23712 7288 23724
rect 4948 23684 4984 23712
rect 7243 23684 7288 23712
rect 4890 23672 4896 23675
rect 4948 23672 4954 23684
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 9398 23672 9404 23724
rect 9456 23712 9462 23724
rect 9493 23715 9551 23721
rect 9493 23712 9505 23715
rect 9456 23684 9505 23712
rect 9456 23672 9462 23684
rect 9493 23681 9505 23684
rect 9539 23681 9551 23715
rect 9493 23675 9551 23681
rect 9585 23715 9643 23721
rect 9585 23681 9597 23715
rect 9631 23712 9643 23715
rect 9766 23712 9772 23724
rect 9631 23684 9772 23712
rect 9631 23681 9643 23684
rect 9585 23675 9643 23681
rect 9766 23672 9772 23684
rect 9824 23672 9830 23724
rect 10042 23712 10048 23724
rect 10003 23684 10048 23712
rect 10042 23672 10048 23684
rect 10100 23672 10106 23724
rect 10228 23715 10286 23721
rect 10228 23681 10240 23715
rect 10274 23712 10286 23715
rect 10597 23715 10655 23721
rect 10274 23684 10548 23712
rect 10274 23681 10286 23684
rect 10228 23675 10286 23681
rect 3970 23644 3976 23656
rect 1903 23616 3464 23644
rect 3712 23616 3976 23644
rect 1903 23613 1915 23616
rect 1857 23607 1915 23613
rect 3436 23576 3464 23616
rect 3970 23604 3976 23616
rect 4028 23644 4034 23656
rect 4249 23647 4307 23653
rect 4249 23644 4261 23647
rect 4028 23616 4261 23644
rect 4028 23604 4034 23616
rect 4249 23613 4261 23616
rect 4295 23613 4307 23647
rect 4249 23607 4307 23613
rect 7101 23647 7159 23653
rect 7101 23613 7113 23647
rect 7147 23644 7159 23647
rect 7466 23644 7472 23656
rect 7147 23616 7472 23644
rect 7147 23613 7159 23616
rect 7101 23607 7159 23613
rect 7466 23604 7472 23616
rect 7524 23644 7530 23656
rect 9950 23644 9956 23656
rect 7524 23616 9628 23644
rect 7524 23604 7530 23616
rect 9600 23588 9628 23616
rect 9784 23616 9956 23644
rect 9784 23588 9812 23616
rect 9950 23604 9956 23616
rect 10008 23644 10014 23656
rect 10321 23647 10379 23653
rect 10321 23644 10333 23647
rect 10008 23616 10333 23644
rect 10008 23604 10014 23616
rect 10321 23613 10333 23616
rect 10367 23613 10379 23647
rect 10321 23607 10379 23613
rect 10413 23647 10471 23653
rect 10413 23613 10425 23647
rect 10459 23613 10471 23647
rect 10520 23644 10548 23684
rect 10597 23681 10609 23715
rect 10643 23712 10655 23715
rect 11422 23712 11428 23724
rect 10643 23684 11428 23712
rect 10643 23681 10655 23684
rect 10597 23675 10655 23681
rect 11422 23672 11428 23684
rect 11480 23672 11486 23724
rect 11517 23715 11575 23721
rect 11517 23681 11529 23715
rect 11563 23681 11575 23715
rect 11698 23712 11704 23724
rect 11659 23684 11704 23712
rect 11517 23675 11575 23681
rect 10520 23616 11008 23644
rect 10413 23607 10471 23613
rect 4065 23579 4123 23585
rect 4065 23576 4077 23579
rect 3436 23548 4077 23576
rect 4065 23545 4077 23548
rect 4111 23545 4123 23579
rect 4065 23539 4123 23545
rect 9582 23536 9588 23588
rect 9640 23536 9646 23588
rect 9766 23576 9772 23588
rect 9679 23548 9772 23576
rect 9766 23536 9772 23548
rect 9824 23536 9830 23588
rect 9858 23536 9864 23588
rect 9916 23576 9922 23588
rect 10226 23576 10232 23588
rect 9916 23548 10232 23576
rect 9916 23536 9922 23548
rect 10226 23536 10232 23548
rect 10284 23576 10290 23588
rect 10428 23576 10456 23607
rect 10284 23548 10456 23576
rect 10284 23536 10290 23548
rect 10686 23536 10692 23588
rect 10744 23576 10750 23588
rect 10781 23579 10839 23585
rect 10781 23576 10793 23579
rect 10744 23548 10793 23576
rect 10744 23536 10750 23548
rect 10781 23545 10793 23548
rect 10827 23545 10839 23579
rect 10781 23539 10839 23545
rect 10980 23520 11008 23616
rect 11238 23604 11244 23656
rect 11296 23644 11302 23656
rect 11532 23644 11560 23675
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 11882 23712 11888 23724
rect 11843 23684 11888 23712
rect 11882 23672 11888 23684
rect 11940 23672 11946 23724
rect 12069 23715 12127 23721
rect 12069 23681 12081 23715
rect 12115 23712 12127 23715
rect 12250 23712 12256 23724
rect 12115 23684 12256 23712
rect 12115 23681 12127 23684
rect 12069 23675 12127 23681
rect 12250 23672 12256 23684
rect 12308 23672 12314 23724
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23681 13507 23715
rect 13449 23675 13507 23681
rect 13541 23715 13599 23721
rect 13541 23681 13553 23715
rect 13587 23681 13599 23715
rect 13541 23675 13599 23681
rect 11790 23644 11796 23656
rect 11296 23616 11560 23644
rect 11751 23616 11796 23644
rect 11296 23604 11302 23616
rect 11790 23604 11796 23616
rect 11848 23604 11854 23656
rect 3329 23511 3387 23517
rect 3329 23477 3341 23511
rect 3375 23508 3387 23511
rect 3418 23508 3424 23520
rect 3375 23480 3424 23508
rect 3375 23477 3387 23480
rect 3329 23471 3387 23477
rect 3418 23468 3424 23480
rect 3476 23468 3482 23520
rect 8018 23468 8024 23520
rect 8076 23508 8082 23520
rect 9309 23511 9367 23517
rect 9309 23508 9321 23511
rect 8076 23480 9321 23508
rect 8076 23468 8082 23480
rect 9309 23477 9321 23480
rect 9355 23508 9367 23511
rect 10594 23508 10600 23520
rect 9355 23480 10600 23508
rect 9355 23477 9367 23480
rect 9309 23471 9367 23477
rect 10594 23468 10600 23480
rect 10652 23468 10658 23520
rect 10962 23508 10968 23520
rect 10923 23480 10968 23508
rect 10962 23468 10968 23480
rect 11020 23468 11026 23520
rect 11698 23468 11704 23520
rect 11756 23508 11762 23520
rect 12434 23508 12440 23520
rect 11756 23480 12440 23508
rect 11756 23468 11762 23480
rect 12434 23468 12440 23480
rect 12492 23468 12498 23520
rect 13464 23508 13492 23675
rect 13556 23576 13584 23675
rect 13630 23672 13636 23724
rect 13688 23712 13694 23724
rect 13817 23715 13875 23721
rect 13817 23712 13829 23715
rect 13688 23684 13829 23712
rect 13688 23672 13694 23684
rect 13817 23681 13829 23684
rect 13863 23681 13875 23715
rect 13998 23712 14004 23724
rect 13959 23684 14004 23712
rect 13817 23675 13875 23681
rect 13998 23672 14004 23684
rect 14056 23672 14062 23724
rect 14918 23576 14924 23588
rect 13556 23548 14924 23576
rect 14918 23536 14924 23548
rect 14976 23536 14982 23588
rect 14090 23508 14096 23520
rect 13464 23480 14096 23508
rect 14090 23468 14096 23480
rect 14148 23468 14154 23520
rect 15120 23508 15148 23698
rect 16482 23672 16488 23724
rect 16540 23712 16546 23724
rect 16540 23684 16585 23712
rect 16540 23672 16546 23684
rect 16666 23672 16672 23724
rect 16724 23712 16730 23724
rect 16868 23712 16896 23811
rect 18800 23780 18828 23820
rect 17880 23752 18828 23780
rect 17880 23724 17908 23752
rect 19426 23740 19432 23792
rect 19484 23780 19490 23792
rect 19484 23752 19529 23780
rect 19484 23740 19490 23752
rect 17862 23721 17868 23724
rect 17129 23715 17187 23721
rect 17129 23712 17141 23715
rect 16724 23684 16769 23712
rect 16868 23684 17141 23712
rect 16724 23672 16730 23684
rect 17129 23681 17141 23684
rect 17175 23681 17187 23715
rect 17860 23712 17868 23721
rect 17823 23684 17868 23712
rect 17129 23675 17187 23681
rect 17860 23675 17868 23684
rect 17862 23672 17868 23675
rect 17920 23672 17926 23724
rect 17957 23715 18015 23721
rect 17957 23681 17969 23715
rect 18003 23681 18015 23715
rect 17957 23675 18015 23681
rect 18049 23715 18107 23721
rect 18049 23681 18061 23715
rect 18095 23712 18107 23715
rect 18138 23712 18144 23724
rect 18095 23684 18144 23712
rect 18095 23681 18107 23684
rect 18049 23675 18107 23681
rect 16206 23644 16212 23656
rect 16167 23616 16212 23644
rect 16206 23604 16212 23616
rect 16264 23604 16270 23656
rect 17494 23604 17500 23656
rect 17552 23644 17558 23656
rect 17972 23644 18000 23675
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 18230 23672 18236 23724
rect 18288 23712 18294 23724
rect 18506 23712 18512 23724
rect 18288 23684 18333 23712
rect 18467 23684 18512 23712
rect 18288 23672 18294 23684
rect 18506 23672 18512 23684
rect 18564 23672 18570 23724
rect 19334 23721 19340 23724
rect 19291 23715 19340 23721
rect 19291 23681 19303 23715
rect 19337 23681 19340 23715
rect 19291 23675 19340 23681
rect 19334 23672 19340 23675
rect 19392 23672 19398 23724
rect 19628 23721 19656 23820
rect 19794 23808 19800 23860
rect 19852 23857 19858 23860
rect 19852 23848 19863 23857
rect 19852 23820 19897 23848
rect 19852 23811 19863 23820
rect 19852 23808 19858 23811
rect 21082 23808 21088 23860
rect 21140 23848 21146 23860
rect 22002 23848 22008 23860
rect 21140 23820 22008 23848
rect 21140 23808 21146 23820
rect 22002 23808 22008 23820
rect 22060 23848 22066 23860
rect 23109 23851 23167 23857
rect 23109 23848 23121 23851
rect 22060 23820 23121 23848
rect 22060 23808 22066 23820
rect 23109 23817 23121 23820
rect 23155 23848 23167 23851
rect 23658 23848 23664 23860
rect 23155 23820 23664 23848
rect 23155 23817 23167 23820
rect 23109 23811 23167 23817
rect 23658 23808 23664 23820
rect 23716 23808 23722 23860
rect 24486 23808 24492 23860
rect 24544 23848 24550 23860
rect 24673 23851 24731 23857
rect 24673 23848 24685 23851
rect 24544 23820 24685 23848
rect 24544 23808 24550 23820
rect 24673 23817 24685 23820
rect 24719 23817 24731 23851
rect 27338 23848 27344 23860
rect 24673 23811 24731 23817
rect 24964 23820 27344 23848
rect 20254 23740 20260 23792
rect 20312 23780 20318 23792
rect 24854 23780 24860 23792
rect 20312 23752 24860 23780
rect 20312 23740 20318 23752
rect 24854 23740 24860 23752
rect 24912 23740 24918 23792
rect 19521 23715 19579 23721
rect 19521 23681 19533 23715
rect 19567 23681 19579 23715
rect 19521 23675 19579 23681
rect 19618 23715 19676 23721
rect 19618 23681 19630 23715
rect 19664 23681 19676 23715
rect 20162 23712 20168 23724
rect 20123 23684 20168 23712
rect 19618 23675 19676 23681
rect 19536 23644 19564 23675
rect 20162 23672 20168 23684
rect 20220 23712 20226 23724
rect 20533 23715 20591 23721
rect 20533 23712 20545 23715
rect 20220 23684 20545 23712
rect 20220 23672 20226 23684
rect 20533 23681 20545 23684
rect 20579 23681 20591 23715
rect 20533 23675 20591 23681
rect 17552 23616 18000 23644
rect 17552 23604 17558 23616
rect 17972 23576 18000 23616
rect 19352 23616 19564 23644
rect 20548 23644 20576 23675
rect 20622 23672 20628 23724
rect 20680 23712 20686 23724
rect 21085 23715 21143 23721
rect 21085 23712 21097 23715
rect 20680 23684 21097 23712
rect 20680 23672 20686 23684
rect 21085 23681 21097 23684
rect 21131 23681 21143 23715
rect 21085 23675 21143 23681
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23712 22431 23715
rect 22419 23684 22968 23712
rect 22419 23681 22431 23684
rect 22373 23675 22431 23681
rect 22830 23644 22836 23656
rect 20548 23616 22836 23644
rect 18325 23579 18383 23585
rect 18325 23576 18337 23579
rect 17972 23548 18337 23576
rect 18325 23545 18337 23548
rect 18371 23545 18383 23579
rect 18325 23539 18383 23545
rect 16945 23511 17003 23517
rect 16945 23508 16957 23511
rect 15120 23480 16957 23508
rect 16945 23477 16957 23480
rect 16991 23477 17003 23511
rect 17678 23508 17684 23520
rect 17639 23480 17684 23508
rect 16945 23471 17003 23477
rect 17678 23468 17684 23480
rect 17736 23468 17742 23520
rect 19242 23468 19248 23520
rect 19300 23508 19306 23520
rect 19352 23508 19380 23616
rect 22830 23604 22836 23616
rect 22888 23604 22894 23656
rect 22940 23644 22968 23684
rect 23014 23672 23020 23724
rect 23072 23712 23078 23724
rect 23201 23715 23259 23721
rect 23201 23712 23213 23715
rect 23072 23684 23213 23712
rect 23072 23672 23078 23684
rect 23201 23681 23213 23684
rect 23247 23681 23259 23715
rect 23201 23675 23259 23681
rect 24118 23672 24124 23724
rect 24176 23712 24182 23724
rect 24489 23715 24547 23721
rect 24489 23712 24501 23715
rect 24176 23684 24501 23712
rect 24176 23672 24182 23684
rect 24489 23681 24501 23684
rect 24535 23712 24547 23715
rect 24765 23715 24823 23721
rect 24765 23712 24777 23715
rect 24535 23684 24777 23712
rect 24535 23681 24547 23684
rect 24489 23675 24547 23681
rect 24765 23681 24777 23684
rect 24811 23681 24823 23715
rect 24765 23675 24823 23681
rect 23474 23644 23480 23656
rect 22940 23616 23480 23644
rect 23474 23604 23480 23616
rect 23532 23604 23538 23656
rect 23658 23604 23664 23656
rect 23716 23644 23722 23656
rect 24964 23653 24992 23820
rect 27338 23808 27344 23820
rect 27396 23808 27402 23860
rect 27430 23808 27436 23860
rect 27488 23808 27494 23860
rect 28537 23851 28595 23857
rect 28537 23817 28549 23851
rect 28583 23848 28595 23851
rect 28626 23848 28632 23860
rect 28583 23820 28632 23848
rect 28583 23817 28595 23820
rect 28537 23811 28595 23817
rect 28626 23808 28632 23820
rect 28684 23808 28690 23860
rect 25222 23780 25228 23792
rect 25183 23752 25228 23780
rect 25222 23740 25228 23752
rect 25280 23740 25286 23792
rect 25866 23740 25872 23792
rect 25924 23740 25930 23792
rect 26970 23740 26976 23792
rect 27028 23780 27034 23792
rect 27249 23783 27307 23789
rect 27249 23780 27261 23783
rect 27028 23752 27261 23780
rect 27028 23740 27034 23752
rect 27249 23749 27261 23752
rect 27295 23749 27307 23783
rect 27448 23780 27476 23808
rect 27249 23743 27307 23749
rect 27356 23752 27476 23780
rect 26602 23672 26608 23724
rect 26660 23712 26666 23724
rect 27356 23721 27384 23752
rect 27065 23715 27123 23721
rect 27065 23712 27077 23715
rect 26660 23684 27077 23712
rect 26660 23672 26666 23684
rect 27065 23681 27077 23684
rect 27111 23681 27123 23715
rect 27065 23675 27123 23681
rect 27341 23715 27399 23721
rect 27341 23681 27353 23715
rect 27387 23681 27399 23715
rect 27341 23675 27399 23681
rect 27438 23715 27496 23721
rect 27438 23681 27450 23715
rect 27484 23681 27496 23715
rect 27438 23675 27496 23681
rect 28077 23715 28135 23721
rect 28077 23681 28089 23715
rect 28123 23712 28135 23715
rect 28166 23712 28172 23724
rect 28123 23684 28172 23712
rect 28123 23681 28135 23684
rect 28077 23675 28135 23681
rect 24949 23647 25007 23653
rect 24949 23644 24961 23647
rect 23716 23616 24961 23644
rect 23716 23604 23722 23616
rect 24949 23613 24961 23616
rect 24995 23613 25007 23647
rect 26694 23644 26700 23656
rect 24949 23607 25007 23613
rect 25056 23616 26556 23644
rect 26655 23616 26700 23644
rect 19978 23576 19984 23588
rect 19939 23548 19984 23576
rect 19978 23536 19984 23548
rect 20036 23536 20042 23588
rect 21174 23536 21180 23588
rect 21232 23576 21238 23588
rect 21269 23579 21327 23585
rect 21269 23576 21281 23579
rect 21232 23548 21281 23576
rect 21232 23536 21238 23548
rect 21269 23545 21281 23548
rect 21315 23576 21327 23579
rect 22186 23576 22192 23588
rect 21315 23548 22094 23576
rect 22147 23548 22192 23576
rect 21315 23545 21327 23548
rect 21269 23539 21327 23545
rect 19300 23480 19380 23508
rect 19300 23468 19306 23480
rect 19426 23468 19432 23520
rect 19484 23508 19490 23520
rect 20438 23508 20444 23520
rect 19484 23480 20444 23508
rect 19484 23468 19490 23480
rect 20438 23468 20444 23480
rect 20496 23468 20502 23520
rect 22066 23508 22094 23548
rect 22186 23536 22192 23548
rect 22244 23536 22250 23588
rect 24765 23579 24823 23585
rect 24765 23545 24777 23579
rect 24811 23576 24823 23579
rect 25056 23576 25084 23616
rect 24811 23548 25084 23576
rect 26528 23576 26556 23616
rect 26694 23604 26700 23616
rect 26752 23604 26758 23656
rect 27154 23604 27160 23656
rect 27212 23644 27218 23656
rect 27448 23644 27476 23675
rect 28166 23672 28172 23684
rect 28224 23672 28230 23724
rect 28353 23715 28411 23721
rect 28353 23712 28365 23715
rect 28276 23684 28365 23712
rect 27212 23616 27476 23644
rect 27212 23604 27218 23616
rect 27614 23576 27620 23588
rect 26528 23548 27384 23576
rect 27575 23548 27620 23576
rect 24811 23545 24823 23548
rect 24765 23539 24823 23545
rect 26786 23508 26792 23520
rect 22066 23480 26792 23508
rect 26786 23468 26792 23480
rect 26844 23508 26850 23520
rect 27246 23508 27252 23520
rect 26844 23480 27252 23508
rect 26844 23468 26850 23480
rect 27246 23468 27252 23480
rect 27304 23468 27310 23520
rect 27356 23508 27384 23548
rect 27614 23536 27620 23548
rect 27672 23536 27678 23588
rect 28276 23585 28304 23684
rect 28353 23681 28365 23684
rect 28399 23681 28411 23715
rect 28353 23675 28411 23681
rect 28261 23579 28319 23585
rect 28261 23545 28273 23579
rect 28307 23545 28319 23579
rect 28261 23539 28319 23545
rect 28166 23508 28172 23520
rect 27356 23480 28172 23508
rect 28166 23468 28172 23480
rect 28224 23468 28230 23520
rect 1104 23418 29532 23440
rect 1104 23366 5688 23418
rect 5740 23366 5752 23418
rect 5804 23366 5816 23418
rect 5868 23366 5880 23418
rect 5932 23366 5944 23418
rect 5996 23366 15163 23418
rect 15215 23366 15227 23418
rect 15279 23366 15291 23418
rect 15343 23366 15355 23418
rect 15407 23366 15419 23418
rect 15471 23366 24639 23418
rect 24691 23366 24703 23418
rect 24755 23366 24767 23418
rect 24819 23366 24831 23418
rect 24883 23366 24895 23418
rect 24947 23366 29532 23418
rect 1104 23344 29532 23366
rect 2777 23307 2835 23313
rect 2777 23273 2789 23307
rect 2823 23304 2835 23307
rect 2866 23304 2872 23316
rect 2823 23276 2872 23304
rect 2823 23273 2835 23276
rect 2777 23267 2835 23273
rect 2866 23264 2872 23276
rect 2924 23264 2930 23316
rect 3789 23307 3847 23313
rect 3789 23273 3801 23307
rect 3835 23304 3847 23307
rect 3970 23304 3976 23316
rect 3835 23276 3976 23304
rect 3835 23273 3847 23276
rect 3789 23267 3847 23273
rect 3970 23264 3976 23276
rect 4028 23264 4034 23316
rect 4890 23304 4896 23316
rect 4851 23276 4896 23304
rect 4890 23264 4896 23276
rect 4948 23264 4954 23316
rect 6086 23304 6092 23316
rect 5000 23276 6092 23304
rect 2685 23239 2743 23245
rect 2685 23205 2697 23239
rect 2731 23205 2743 23239
rect 2685 23199 2743 23205
rect 2222 23100 2228 23112
rect 2183 23072 2228 23100
rect 2222 23060 2228 23072
rect 2280 23060 2286 23112
rect 2314 23060 2320 23112
rect 2372 23100 2378 23112
rect 2501 23103 2559 23109
rect 2501 23100 2513 23103
rect 2372 23072 2513 23100
rect 2372 23060 2378 23072
rect 2501 23069 2513 23072
rect 2547 23069 2559 23103
rect 2700 23100 2728 23199
rect 2961 23103 3019 23109
rect 2961 23100 2973 23103
rect 2700 23072 2973 23100
rect 2501 23063 2559 23069
rect 2961 23069 2973 23072
rect 3007 23069 3019 23103
rect 2961 23063 3019 23069
rect 3602 23060 3608 23112
rect 3660 23100 3666 23112
rect 5000 23109 5028 23276
rect 6086 23264 6092 23276
rect 6144 23264 6150 23316
rect 9674 23264 9680 23316
rect 9732 23304 9738 23316
rect 10042 23304 10048 23316
rect 9732 23276 10048 23304
rect 9732 23264 9738 23276
rect 10042 23264 10048 23276
rect 10100 23264 10106 23316
rect 10229 23307 10287 23313
rect 10229 23273 10241 23307
rect 10275 23304 10287 23307
rect 12710 23304 12716 23316
rect 10275 23276 12716 23304
rect 10275 23273 10287 23276
rect 10229 23267 10287 23273
rect 12710 23264 12716 23276
rect 12768 23264 12774 23316
rect 15565 23307 15623 23313
rect 15565 23273 15577 23307
rect 15611 23304 15623 23307
rect 16206 23304 16212 23316
rect 15611 23276 16212 23304
rect 15611 23273 15623 23276
rect 15565 23267 15623 23273
rect 16206 23264 16212 23276
rect 16264 23264 16270 23316
rect 17236 23276 18460 23304
rect 5534 23196 5540 23248
rect 5592 23236 5598 23248
rect 5721 23239 5779 23245
rect 5721 23236 5733 23239
rect 5592 23208 5733 23236
rect 5592 23196 5598 23208
rect 5721 23205 5733 23208
rect 5767 23205 5779 23239
rect 5721 23199 5779 23205
rect 5166 23168 5172 23180
rect 5127 23140 5172 23168
rect 5166 23128 5172 23140
rect 5224 23128 5230 23180
rect 5261 23171 5319 23177
rect 5261 23137 5273 23171
rect 5307 23168 5319 23171
rect 5626 23168 5632 23180
rect 5307 23140 5632 23168
rect 5307 23137 5319 23140
rect 5261 23131 5319 23137
rect 5626 23128 5632 23140
rect 5684 23128 5690 23180
rect 5736 23168 5764 23199
rect 9306 23196 9312 23248
rect 9364 23236 9370 23248
rect 9364 23208 10088 23236
rect 9364 23196 9370 23208
rect 6181 23171 6239 23177
rect 6181 23168 6193 23171
rect 5736 23140 6193 23168
rect 6181 23137 6193 23140
rect 6227 23137 6239 23171
rect 6181 23131 6239 23137
rect 8294 23128 8300 23180
rect 8352 23168 8358 23180
rect 9324 23168 9352 23196
rect 8352 23140 8397 23168
rect 8497 23140 9352 23168
rect 8352 23128 8358 23140
rect 3973 23103 4031 23109
rect 3973 23100 3985 23103
rect 3660 23072 3985 23100
rect 3660 23060 3666 23072
rect 3973 23069 3985 23072
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 4985 23103 5043 23109
rect 4985 23069 4997 23103
rect 5031 23069 5043 23103
rect 5350 23100 5356 23112
rect 4985 23063 5043 23069
rect 5092 23072 5356 23100
rect 4709 23035 4767 23041
rect 4709 23001 4721 23035
rect 4755 23032 4767 23035
rect 5092 23032 5120 23072
rect 5350 23060 5356 23072
rect 5408 23060 5414 23112
rect 5537 23103 5595 23109
rect 5537 23069 5549 23103
rect 5583 23100 5595 23103
rect 8018 23100 8024 23112
rect 5583 23072 8024 23100
rect 5583 23069 5595 23072
rect 5537 23063 5595 23069
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 8186 23100 8244 23106
rect 8186 23066 8198 23100
rect 8232 23066 8244 23100
rect 8186 23060 8244 23066
rect 8389 23103 8447 23109
rect 8389 23069 8401 23103
rect 8435 23100 8447 23103
rect 8497 23100 8525 23140
rect 9582 23128 9588 23180
rect 9640 23168 9646 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 9640 23140 9689 23168
rect 9640 23128 9646 23140
rect 9677 23137 9689 23140
rect 9723 23168 9735 23171
rect 9950 23168 9956 23180
rect 9723 23140 9956 23168
rect 9723 23137 9735 23140
rect 9677 23131 9735 23137
rect 9950 23128 9956 23140
rect 10008 23128 10014 23180
rect 10060 23168 10088 23208
rect 10962 23196 10968 23248
rect 11020 23236 11026 23248
rect 17236 23236 17264 23276
rect 11020 23208 17264 23236
rect 18432 23236 18460 23276
rect 18506 23264 18512 23316
rect 18564 23304 18570 23316
rect 18877 23307 18935 23313
rect 18877 23304 18889 23307
rect 18564 23276 18889 23304
rect 18564 23264 18570 23276
rect 18877 23273 18889 23276
rect 18923 23304 18935 23307
rect 19061 23307 19119 23313
rect 19061 23304 19073 23307
rect 18923 23276 19073 23304
rect 18923 23273 18935 23276
rect 18877 23267 18935 23273
rect 19061 23273 19073 23276
rect 19107 23273 19119 23307
rect 19061 23267 19119 23273
rect 19518 23264 19524 23316
rect 19576 23304 19582 23316
rect 19889 23307 19947 23313
rect 19889 23304 19901 23307
rect 19576 23276 19901 23304
rect 19576 23264 19582 23276
rect 19889 23273 19901 23276
rect 19935 23304 19947 23307
rect 20165 23307 20223 23313
rect 20165 23304 20177 23307
rect 19935 23276 20177 23304
rect 19935 23273 19947 23276
rect 19889 23267 19947 23273
rect 20165 23273 20177 23276
rect 20211 23273 20223 23307
rect 27430 23304 27436 23316
rect 20165 23267 20223 23273
rect 20272 23276 27436 23304
rect 20272 23236 20300 23276
rect 27430 23264 27436 23276
rect 27488 23264 27494 23316
rect 29089 23307 29147 23313
rect 29089 23273 29101 23307
rect 29135 23304 29147 23307
rect 29641 23307 29699 23313
rect 29641 23304 29653 23307
rect 29135 23276 29653 23304
rect 29135 23273 29147 23276
rect 29089 23267 29147 23273
rect 29641 23273 29653 23276
rect 29687 23273 29699 23307
rect 29641 23267 29699 23273
rect 18432 23208 20300 23236
rect 11020 23196 11026 23208
rect 22094 23196 22100 23248
rect 22152 23236 22158 23248
rect 22741 23239 22799 23245
rect 22741 23236 22753 23239
rect 22152 23208 22753 23236
rect 22152 23196 22158 23208
rect 22741 23205 22753 23208
rect 22787 23236 22799 23239
rect 24302 23236 24308 23248
rect 22787 23208 24308 23236
rect 22787 23205 22799 23208
rect 22741 23199 22799 23205
rect 24302 23196 24308 23208
rect 24360 23196 24366 23248
rect 25682 23196 25688 23248
rect 25740 23236 25746 23248
rect 26970 23236 26976 23248
rect 25740 23208 26976 23236
rect 25740 23196 25746 23208
rect 26970 23196 26976 23208
rect 27028 23196 27034 23248
rect 27157 23239 27215 23245
rect 27157 23205 27169 23239
rect 27203 23236 27215 23239
rect 27203 23208 27476 23236
rect 27203 23205 27215 23208
rect 27157 23199 27215 23205
rect 11609 23171 11667 23177
rect 11609 23168 11621 23171
rect 10060 23140 11621 23168
rect 11609 23137 11621 23140
rect 11655 23168 11667 23171
rect 11882 23168 11888 23180
rect 11655 23140 11888 23168
rect 11655 23137 11667 23140
rect 11609 23131 11667 23137
rect 11882 23128 11888 23140
rect 11940 23128 11946 23180
rect 12066 23128 12072 23180
rect 12124 23168 12130 23180
rect 14185 23171 14243 23177
rect 14185 23168 14197 23171
rect 12124 23140 14197 23168
rect 12124 23128 12130 23140
rect 14185 23137 14197 23140
rect 14231 23137 14243 23171
rect 17310 23168 17316 23180
rect 14185 23131 14243 23137
rect 14384 23140 17316 23168
rect 8435 23072 8525 23100
rect 8573 23103 8631 23109
rect 8435 23069 8447 23072
rect 8389 23063 8447 23069
rect 8573 23069 8585 23103
rect 8619 23100 8631 23103
rect 9306 23100 9312 23112
rect 8619 23072 9312 23100
rect 8619 23069 8631 23072
rect 8573 23063 8631 23069
rect 9306 23060 9312 23072
rect 9364 23100 9370 23112
rect 9861 23103 9919 23109
rect 9861 23100 9873 23103
rect 9364 23072 9873 23100
rect 9364 23060 9370 23072
rect 9861 23069 9873 23072
rect 9907 23069 9919 23103
rect 9861 23063 9919 23069
rect 10594 23060 10600 23112
rect 10652 23100 10658 23112
rect 11238 23100 11244 23112
rect 10652 23072 11244 23100
rect 10652 23060 10658 23072
rect 11238 23060 11244 23072
rect 11296 23060 11302 23112
rect 11422 23100 11428 23112
rect 11383 23072 11428 23100
rect 11422 23060 11428 23072
rect 11480 23060 11486 23112
rect 11517 23103 11575 23109
rect 11517 23069 11529 23103
rect 11563 23100 11575 23103
rect 11698 23100 11704 23112
rect 11563 23072 11704 23100
rect 11563 23069 11575 23072
rect 11517 23063 11575 23069
rect 11698 23060 11704 23072
rect 11756 23060 11762 23112
rect 11793 23103 11851 23109
rect 11793 23069 11805 23103
rect 11839 23100 11851 23103
rect 12434 23100 12440 23112
rect 11839 23072 12440 23100
rect 11839 23069 11851 23072
rect 11793 23063 11851 23069
rect 12434 23060 12440 23072
rect 12492 23060 12498 23112
rect 14090 23100 14096 23112
rect 14051 23072 14096 23100
rect 14090 23060 14096 23072
rect 14148 23060 14154 23112
rect 14384 23109 14412 23140
rect 17310 23128 17316 23140
rect 17368 23128 17374 23180
rect 19061 23171 19119 23177
rect 19061 23137 19073 23171
rect 19107 23168 19119 23171
rect 19242 23168 19248 23180
rect 19107 23140 19248 23168
rect 19107 23137 19119 23140
rect 19061 23131 19119 23137
rect 19242 23128 19248 23140
rect 19300 23168 19306 23180
rect 19521 23171 19579 23177
rect 19521 23168 19533 23171
rect 19300 23140 19533 23168
rect 19300 23128 19306 23140
rect 19521 23137 19533 23140
rect 19567 23137 19579 23171
rect 19521 23131 19579 23137
rect 14369 23103 14427 23109
rect 14369 23069 14381 23103
rect 14415 23069 14427 23103
rect 14369 23063 14427 23069
rect 14553 23103 14611 23109
rect 14553 23069 14565 23103
rect 14599 23069 14611 23103
rect 14734 23100 14740 23112
rect 14695 23072 14740 23100
rect 14553 23063 14611 23069
rect 4755 23004 5120 23032
rect 4755 23001 4767 23004
rect 4709 22995 4767 23001
rect 5718 22992 5724 23044
rect 5776 23032 5782 23044
rect 6454 23041 6460 23044
rect 5905 23035 5963 23041
rect 5905 23032 5917 23035
rect 5776 23004 5917 23032
rect 5776 22992 5782 23004
rect 5905 23001 5917 23004
rect 5951 23001 5963 23035
rect 5905 22995 5963 23001
rect 6448 22995 6460 23041
rect 6512 23032 6518 23044
rect 8201 23032 8229 23060
rect 6512 23004 6548 23032
rect 7852 23004 8229 23032
rect 9769 23035 9827 23041
rect 6454 22992 6460 22995
rect 6512 22992 6518 23004
rect 7852 22976 7880 23004
rect 9769 23001 9781 23035
rect 9815 23032 9827 23035
rect 10042 23032 10048 23044
rect 9815 23004 10048 23032
rect 9815 23001 9827 23004
rect 9769 22995 9827 23001
rect 10042 22992 10048 23004
rect 10100 22992 10106 23044
rect 11439 23032 11467 23060
rect 12069 23035 12127 23041
rect 12069 23032 12081 23035
rect 11439 23004 12081 23032
rect 12069 23001 12081 23004
rect 12115 23001 12127 23035
rect 12069 22995 12127 23001
rect 13630 22992 13636 23044
rect 13688 23032 13694 23044
rect 14568 23032 14596 23063
rect 14734 23060 14740 23072
rect 14792 23060 14798 23112
rect 15010 23100 15016 23112
rect 14971 23072 15016 23100
rect 15010 23060 15016 23072
rect 15068 23060 15074 23112
rect 15470 23109 15476 23112
rect 15433 23103 15476 23109
rect 15433 23100 15445 23103
rect 15383 23072 15445 23100
rect 15433 23069 15445 23072
rect 15528 23100 15534 23112
rect 15654 23100 15660 23112
rect 15528 23072 15660 23100
rect 15433 23063 15476 23069
rect 15470 23060 15476 23063
rect 15528 23060 15534 23072
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 15838 23060 15844 23112
rect 15896 23060 15902 23112
rect 17497 23103 17555 23109
rect 17497 23069 17509 23103
rect 17543 23100 17555 23103
rect 18138 23100 18144 23112
rect 17543 23072 18144 23100
rect 17543 23069 17555 23072
rect 17497 23063 17555 23069
rect 18138 23060 18144 23072
rect 18196 23060 18202 23112
rect 13688 23004 14596 23032
rect 13688 22992 13694 23004
rect 14918 22992 14924 23044
rect 14976 23032 14982 23044
rect 15197 23035 15255 23041
rect 15197 23032 15209 23035
rect 14976 23004 15209 23032
rect 14976 22992 14982 23004
rect 15197 23001 15209 23004
rect 15243 23001 15255 23035
rect 15197 22995 15255 23001
rect 15289 23035 15347 23041
rect 15289 23001 15301 23035
rect 15335 23032 15347 23035
rect 15856 23032 15884 23060
rect 15335 23004 15884 23032
rect 15335 23001 15347 23004
rect 15289 22995 15347 23001
rect 17678 22992 17684 23044
rect 17736 23041 17742 23044
rect 17736 23035 17800 23041
rect 17736 23001 17754 23035
rect 17788 23001 17800 23035
rect 19536 23032 19564 23131
rect 19702 23128 19708 23180
rect 19760 23168 19766 23180
rect 19889 23171 19947 23177
rect 19889 23168 19901 23171
rect 19760 23140 19901 23168
rect 19760 23128 19766 23140
rect 19889 23137 19901 23140
rect 19935 23168 19947 23171
rect 20257 23171 20315 23177
rect 20257 23168 20269 23171
rect 19935 23140 20269 23168
rect 19935 23137 19947 23140
rect 19889 23131 19947 23137
rect 20257 23137 20269 23140
rect 20303 23137 20315 23171
rect 27338 23168 27344 23180
rect 20257 23131 20315 23137
rect 22204 23140 26234 23168
rect 27299 23140 27344 23168
rect 20162 23060 20168 23112
rect 20220 23100 20226 23112
rect 20717 23103 20775 23109
rect 20717 23100 20729 23103
rect 20220 23072 20265 23100
rect 20364 23072 20729 23100
rect 20220 23060 20226 23072
rect 19536 23004 20116 23032
rect 17736 22995 17800 23001
rect 17736 22992 17742 22995
rect 2406 22964 2412 22976
rect 2367 22936 2412 22964
rect 2406 22924 2412 22936
rect 2464 22924 2470 22976
rect 6638 22924 6644 22976
rect 6696 22964 6702 22976
rect 7282 22964 7288 22976
rect 6696 22936 7288 22964
rect 6696 22924 6702 22936
rect 7282 22924 7288 22936
rect 7340 22964 7346 22976
rect 7561 22967 7619 22973
rect 7561 22964 7573 22967
rect 7340 22936 7573 22964
rect 7340 22924 7346 22936
rect 7561 22933 7573 22936
rect 7607 22933 7619 22967
rect 7834 22964 7840 22976
rect 7795 22936 7840 22964
rect 7561 22927 7619 22933
rect 7834 22924 7840 22936
rect 7892 22924 7898 22976
rect 8202 22924 8208 22976
rect 8260 22964 8266 22976
rect 8665 22967 8723 22973
rect 8665 22964 8677 22967
rect 8260 22936 8677 22964
rect 8260 22924 8266 22936
rect 8665 22933 8677 22936
rect 8711 22933 8723 22967
rect 8665 22927 8723 22933
rect 9401 22967 9459 22973
rect 9401 22933 9413 22967
rect 9447 22964 9459 22967
rect 9582 22964 9588 22976
rect 9447 22936 9588 22964
rect 9447 22933 9459 22936
rect 9401 22927 9459 22933
rect 9582 22924 9588 22936
rect 9640 22924 9646 22976
rect 11882 22964 11888 22976
rect 11843 22936 11888 22964
rect 11882 22924 11888 22936
rect 11940 22924 11946 22976
rect 15838 22964 15844 22976
rect 15751 22936 15844 22964
rect 15838 22924 15844 22936
rect 15896 22964 15902 22976
rect 17218 22964 17224 22976
rect 15896 22936 17224 22964
rect 15896 22924 15902 22936
rect 17218 22924 17224 22936
rect 17276 22924 17282 22976
rect 19334 22924 19340 22976
rect 19392 22964 19398 22976
rect 19705 22967 19763 22973
rect 19705 22964 19717 22967
rect 19392 22936 19717 22964
rect 19392 22924 19398 22936
rect 19705 22933 19717 22936
rect 19751 22933 19763 22967
rect 20088 22964 20116 23004
rect 20364 22964 20392 23072
rect 20717 23069 20729 23072
rect 20763 23069 20775 23103
rect 20717 23063 20775 23069
rect 20993 23103 21051 23109
rect 20993 23069 21005 23103
rect 21039 23100 21051 23103
rect 21082 23100 21088 23112
rect 21039 23072 21088 23100
rect 21039 23069 21051 23072
rect 20993 23063 21051 23069
rect 21082 23060 21088 23072
rect 21140 23060 21146 23112
rect 20806 22992 20812 23044
rect 20864 23032 20870 23044
rect 21238 23035 21296 23041
rect 21238 23032 21250 23035
rect 20864 23004 21250 23032
rect 20864 22992 20870 23004
rect 21238 23001 21250 23004
rect 21284 23001 21296 23035
rect 21238 22995 21296 23001
rect 20088 22936 20392 22964
rect 20533 22967 20591 22973
rect 19705 22927 19763 22933
rect 20533 22933 20545 22967
rect 20579 22964 20591 22967
rect 20622 22964 20628 22976
rect 20579 22936 20628 22964
rect 20579 22933 20591 22936
rect 20533 22927 20591 22933
rect 20622 22924 20628 22936
rect 20680 22924 20686 22976
rect 20901 22967 20959 22973
rect 20901 22933 20913 22967
rect 20947 22964 20959 22967
rect 21634 22964 21640 22976
rect 20947 22936 21640 22964
rect 20947 22933 20959 22936
rect 20901 22927 20959 22933
rect 21634 22924 21640 22936
rect 21692 22964 21698 22976
rect 22204 22964 22232 23140
rect 22557 23103 22615 23109
rect 22557 23100 22569 23103
rect 22388 23072 22569 23100
rect 22388 22976 22416 23072
rect 22557 23069 22569 23072
rect 22603 23069 22615 23103
rect 22557 23063 22615 23069
rect 24486 23060 24492 23112
rect 24544 23100 24550 23112
rect 24581 23103 24639 23109
rect 24581 23100 24593 23103
rect 24544 23072 24593 23100
rect 24544 23060 24550 23072
rect 24581 23069 24593 23072
rect 24627 23069 24639 23103
rect 24581 23063 24639 23069
rect 25038 22992 25044 23044
rect 25096 23032 25102 23044
rect 25317 23035 25375 23041
rect 25317 23032 25329 23035
rect 25096 23004 25329 23032
rect 25096 22992 25102 23004
rect 25317 23001 25329 23004
rect 25363 23032 25375 23035
rect 25682 23032 25688 23044
rect 25363 23004 25688 23032
rect 25363 23001 25375 23004
rect 25317 22995 25375 23001
rect 25682 22992 25688 23004
rect 25740 22992 25746 23044
rect 26206 23032 26234 23140
rect 27338 23128 27344 23140
rect 27396 23128 27402 23180
rect 27448 23168 27476 23208
rect 27617 23171 27675 23177
rect 27617 23168 27629 23171
rect 27448 23140 27629 23168
rect 27617 23137 27629 23140
rect 27663 23137 27675 23171
rect 27617 23131 27675 23137
rect 26602 23100 26608 23112
rect 26563 23072 26608 23100
rect 26602 23060 26608 23072
rect 26660 23060 26666 23112
rect 27025 23103 27083 23109
rect 27025 23069 27037 23103
rect 27071 23100 27083 23103
rect 27154 23100 27160 23112
rect 27071 23072 27160 23100
rect 27071 23069 27083 23072
rect 27025 23063 27083 23069
rect 27154 23060 27160 23072
rect 27212 23060 27218 23112
rect 26786 23032 26792 23044
rect 26206 23004 26792 23032
rect 26786 22992 26792 23004
rect 26844 22992 26850 23044
rect 26881 23035 26939 23041
rect 26881 23001 26893 23035
rect 26927 23001 26939 23035
rect 26881 22995 26939 23001
rect 22370 22964 22376 22976
rect 21692 22936 22232 22964
rect 22331 22936 22376 22964
rect 21692 22924 21698 22936
rect 22370 22924 22376 22936
rect 22428 22924 22434 22976
rect 24670 22924 24676 22976
rect 24728 22964 24734 22976
rect 24765 22967 24823 22973
rect 24765 22964 24777 22967
rect 24728 22936 24777 22964
rect 24728 22924 24734 22936
rect 24765 22933 24777 22936
rect 24811 22933 24823 22967
rect 25498 22964 25504 22976
rect 25459 22936 25504 22964
rect 24765 22927 24823 22933
rect 25498 22924 25504 22936
rect 25556 22924 25562 22976
rect 26896 22964 26924 22995
rect 28626 22992 28632 23044
rect 28684 22992 28690 23044
rect 29104 22964 29132 23267
rect 26896 22936 29132 22964
rect 1104 22874 29532 22896
rect 1104 22822 10425 22874
rect 10477 22822 10489 22874
rect 10541 22822 10553 22874
rect 10605 22822 10617 22874
rect 10669 22822 10681 22874
rect 10733 22822 19901 22874
rect 19953 22822 19965 22874
rect 20017 22822 20029 22874
rect 20081 22822 20093 22874
rect 20145 22822 20157 22874
rect 20209 22822 29532 22874
rect 1104 22800 29532 22822
rect 4893 22763 4951 22769
rect 4893 22729 4905 22763
rect 4939 22729 4951 22763
rect 6454 22760 6460 22772
rect 6415 22732 6460 22760
rect 4893 22723 4951 22729
rect 2406 22652 2412 22704
rect 2464 22652 2470 22704
rect 1394 22624 1400 22636
rect 1355 22596 1400 22624
rect 1394 22584 1400 22596
rect 1452 22584 1458 22636
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22593 4767 22627
rect 4908 22624 4936 22723
rect 6454 22720 6460 22732
rect 6512 22720 6518 22772
rect 6822 22720 6828 22772
rect 6880 22720 6886 22772
rect 9306 22760 9312 22772
rect 9267 22732 9312 22760
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 9490 22720 9496 22772
rect 9548 22760 9554 22772
rect 9548 22732 9674 22760
rect 9548 22720 9554 22732
rect 6840 22692 6868 22720
rect 9646 22692 9674 22732
rect 9950 22720 9956 22772
rect 10008 22760 10014 22772
rect 12158 22760 12164 22772
rect 10008 22732 12164 22760
rect 10008 22720 10014 22732
rect 12158 22720 12164 22732
rect 12216 22720 12222 22772
rect 13630 22720 13636 22772
rect 13688 22760 13694 22772
rect 13725 22763 13783 22769
rect 13725 22760 13737 22763
rect 13688 22732 13737 22760
rect 13688 22720 13694 22732
rect 13725 22729 13737 22732
rect 13771 22729 13783 22763
rect 13725 22723 13783 22729
rect 13817 22763 13875 22769
rect 13817 22729 13829 22763
rect 13863 22760 13875 22763
rect 14090 22760 14096 22772
rect 13863 22732 14096 22760
rect 13863 22729 13875 22732
rect 13817 22723 13875 22729
rect 14090 22720 14096 22732
rect 14148 22720 14154 22772
rect 16853 22763 16911 22769
rect 15212 22732 15976 22760
rect 11784 22695 11842 22701
rect 6473 22664 6868 22692
rect 7944 22664 11560 22692
rect 4985 22627 5043 22633
rect 4985 22624 4997 22627
rect 4908 22596 4997 22624
rect 4709 22587 4767 22593
rect 4985 22593 4997 22596
rect 5031 22593 5043 22627
rect 4985 22587 5043 22593
rect 1670 22556 1676 22568
rect 1631 22528 1676 22556
rect 1670 22516 1676 22528
rect 1728 22516 1734 22568
rect 2314 22516 2320 22568
rect 2372 22556 2378 22568
rect 4724 22556 4752 22587
rect 5074 22556 5080 22568
rect 2372 22528 5080 22556
rect 2372 22516 2378 22528
rect 5074 22516 5080 22528
rect 5132 22516 5138 22568
rect 6473 22556 6501 22664
rect 6549 22627 6607 22633
rect 6549 22593 6561 22627
rect 6595 22624 6607 22627
rect 6638 22624 6644 22636
rect 6595 22596 6644 22624
rect 6595 22593 6607 22596
rect 6549 22587 6607 22593
rect 6638 22584 6644 22596
rect 6696 22584 6702 22636
rect 6822 22624 6828 22636
rect 6783 22596 6828 22624
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 7944 22633 7972 22664
rect 8202 22633 8208 22636
rect 6918 22627 6976 22633
rect 6918 22593 6930 22627
rect 6964 22593 6976 22627
rect 6918 22587 6976 22593
rect 7101 22627 7159 22633
rect 7101 22593 7113 22627
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7929 22627 7987 22633
rect 7929 22593 7941 22627
rect 7975 22593 7987 22627
rect 8196 22624 8208 22633
rect 8163 22596 8208 22624
rect 7929 22587 7987 22593
rect 8196 22587 8208 22596
rect 6733 22559 6791 22565
rect 6733 22556 6745 22559
rect 6473 22528 6745 22556
rect 6733 22525 6745 22528
rect 6779 22525 6791 22559
rect 6733 22519 6791 22525
rect 6181 22491 6239 22497
rect 6181 22457 6193 22491
rect 6227 22488 6239 22491
rect 6270 22488 6276 22500
rect 6227 22460 6276 22488
rect 6227 22457 6239 22460
rect 6181 22451 6239 22457
rect 6270 22448 6276 22460
rect 6328 22488 6334 22500
rect 6932 22488 6960 22587
rect 6328 22460 6960 22488
rect 6328 22448 6334 22460
rect 3050 22380 3056 22432
rect 3108 22420 3114 22432
rect 3145 22423 3203 22429
rect 3145 22420 3157 22423
rect 3108 22392 3157 22420
rect 3108 22380 3114 22392
rect 3145 22389 3157 22392
rect 3191 22389 3203 22423
rect 5166 22420 5172 22432
rect 5127 22392 5172 22420
rect 3145 22383 3203 22389
rect 5166 22380 5172 22392
rect 5224 22380 5230 22432
rect 7116 22420 7144 22587
rect 8202 22584 8208 22587
rect 8260 22584 8266 22636
rect 9493 22627 9551 22633
rect 9493 22593 9505 22627
rect 9539 22593 9551 22627
rect 9493 22587 9551 22593
rect 9508 22556 9536 22587
rect 9582 22584 9588 22636
rect 9640 22624 9646 22636
rect 9676 22627 9734 22633
rect 9676 22624 9688 22627
rect 9640 22596 9688 22624
rect 9640 22584 9646 22596
rect 9676 22593 9688 22596
rect 9722 22593 9734 22627
rect 9676 22587 9734 22593
rect 9766 22584 9772 22636
rect 9824 22624 9830 22636
rect 10042 22624 10048 22636
rect 9824 22596 9869 22624
rect 10003 22596 10048 22624
rect 9824 22584 9830 22596
rect 10042 22584 10048 22596
rect 10100 22584 10106 22636
rect 11532 22633 11560 22664
rect 11784 22661 11796 22695
rect 11830 22692 11842 22695
rect 11882 22692 11888 22704
rect 11830 22664 11888 22692
rect 11830 22661 11842 22664
rect 11784 22655 11842 22661
rect 11882 22652 11888 22664
rect 11940 22652 11946 22704
rect 15212 22701 15240 22732
rect 15197 22695 15255 22701
rect 15197 22661 15209 22695
rect 15243 22661 15255 22695
rect 15197 22655 15255 22661
rect 15289 22695 15347 22701
rect 15289 22661 15301 22695
rect 15335 22692 15347 22695
rect 15838 22692 15844 22704
rect 15335 22664 15844 22692
rect 15335 22661 15347 22664
rect 15289 22655 15347 22661
rect 15838 22652 15844 22664
rect 15896 22652 15902 22704
rect 15948 22701 15976 22732
rect 16853 22729 16865 22763
rect 16899 22729 16911 22763
rect 16853 22723 16911 22729
rect 20165 22763 20223 22769
rect 20165 22729 20177 22763
rect 20211 22760 20223 22763
rect 20254 22760 20260 22772
rect 20211 22732 20260 22760
rect 20211 22729 20223 22732
rect 20165 22723 20223 22729
rect 15933 22695 15991 22701
rect 15933 22661 15945 22695
rect 15979 22661 15991 22695
rect 15933 22655 15991 22661
rect 16025 22695 16083 22701
rect 16025 22661 16037 22695
rect 16071 22692 16083 22695
rect 16482 22692 16488 22704
rect 16071 22664 16488 22692
rect 16071 22661 16083 22664
rect 16025 22655 16083 22661
rect 11517 22627 11575 22633
rect 11517 22593 11529 22627
rect 11563 22593 11575 22627
rect 13538 22624 13544 22636
rect 13499 22596 13544 22624
rect 11517 22587 11575 22593
rect 13538 22584 13544 22596
rect 13596 22584 13602 22636
rect 13998 22624 14004 22636
rect 13959 22596 14004 22624
rect 13998 22584 14004 22596
rect 14056 22584 14062 22636
rect 15010 22624 15016 22636
rect 14971 22596 15016 22624
rect 15010 22584 15016 22596
rect 15068 22584 15074 22636
rect 15470 22633 15476 22636
rect 15433 22627 15476 22633
rect 15433 22593 15445 22627
rect 15433 22587 15476 22593
rect 9861 22559 9919 22565
rect 9508 22528 9720 22556
rect 9692 22500 9720 22528
rect 9861 22525 9873 22559
rect 9907 22556 9919 22559
rect 10226 22556 10232 22568
rect 9907 22528 10232 22556
rect 9907 22525 9919 22528
rect 9861 22519 9919 22525
rect 10226 22516 10232 22528
rect 10284 22516 10290 22568
rect 14826 22516 14832 22568
rect 14884 22556 14890 22568
rect 15448 22556 15476 22587
rect 15528 22584 15534 22636
rect 15654 22584 15660 22636
rect 15712 22624 15718 22636
rect 15749 22627 15807 22633
rect 15749 22624 15761 22627
rect 15712 22596 15761 22624
rect 15712 22584 15718 22596
rect 15749 22593 15761 22596
rect 15795 22593 15807 22627
rect 15749 22587 15807 22593
rect 14884 22528 15476 22556
rect 15948 22556 15976 22655
rect 16482 22652 16488 22664
rect 16540 22652 16546 22704
rect 16114 22584 16120 22636
rect 16172 22633 16178 22636
rect 16172 22624 16180 22633
rect 16666 22624 16672 22636
rect 16172 22596 16217 22624
rect 16627 22596 16672 22624
rect 16172 22587 16180 22596
rect 16172 22584 16178 22587
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 16868 22624 16896 22723
rect 20254 22720 20260 22732
rect 20312 22720 20318 22772
rect 20456 22732 22094 22760
rect 17310 22652 17316 22704
rect 17368 22692 17374 22704
rect 17368 22664 18736 22692
rect 17368 22652 17374 22664
rect 17129 22627 17187 22633
rect 17129 22624 17141 22627
rect 16868 22596 17141 22624
rect 17129 22593 17141 22596
rect 17175 22593 17187 22627
rect 17402 22624 17408 22636
rect 17363 22596 17408 22624
rect 17129 22587 17187 22593
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 17862 22633 17868 22636
rect 17589 22627 17647 22633
rect 17589 22593 17601 22627
rect 17635 22593 17647 22627
rect 17589 22587 17647 22593
rect 17681 22627 17739 22633
rect 17681 22593 17693 22627
rect 17727 22593 17739 22627
rect 17681 22587 17739 22593
rect 17825 22627 17868 22633
rect 17825 22593 17837 22627
rect 17825 22587 17868 22593
rect 17494 22556 17500 22568
rect 15948 22528 17500 22556
rect 14884 22516 14890 22528
rect 17494 22516 17500 22528
rect 17552 22556 17558 22568
rect 17604 22556 17632 22587
rect 17552 22528 17632 22556
rect 17552 22516 17558 22528
rect 9306 22448 9312 22500
rect 9364 22488 9370 22500
rect 9582 22488 9588 22500
rect 9364 22460 9588 22488
rect 9364 22448 9370 22460
rect 9582 22448 9588 22460
rect 9640 22448 9646 22500
rect 9674 22448 9680 22500
rect 9732 22448 9738 22500
rect 14918 22448 14924 22500
rect 14976 22488 14982 22500
rect 17696 22488 17724 22587
rect 17862 22584 17868 22587
rect 17920 22584 17926 22636
rect 18138 22624 18144 22636
rect 18099 22596 18144 22624
rect 18138 22584 18144 22596
rect 18196 22584 18202 22636
rect 18397 22627 18455 22633
rect 18397 22624 18409 22627
rect 18248 22596 18409 22624
rect 18248 22556 18276 22596
rect 18397 22593 18409 22596
rect 18443 22593 18455 22627
rect 18708 22624 18736 22664
rect 19242 22652 19248 22704
rect 19300 22692 19306 22704
rect 19300 22664 20024 22692
rect 19300 22652 19306 22664
rect 19702 22624 19708 22636
rect 18708 22596 19196 22624
rect 19663 22596 19708 22624
rect 18397 22587 18455 22593
rect 17972 22528 18276 22556
rect 19168 22556 19196 22596
rect 19702 22584 19708 22596
rect 19760 22584 19766 22636
rect 19996 22633 20024 22664
rect 19981 22627 20039 22633
rect 19981 22593 19993 22627
rect 20027 22593 20039 22627
rect 19981 22587 20039 22593
rect 19797 22559 19855 22565
rect 19797 22556 19809 22559
rect 19168 22528 19809 22556
rect 17972 22497 18000 22528
rect 19797 22525 19809 22528
rect 19843 22556 19855 22559
rect 20456 22556 20484 22732
rect 22066 22692 22094 22732
rect 22278 22720 22284 22772
rect 22336 22760 22342 22772
rect 22554 22760 22560 22772
rect 22336 22732 22560 22760
rect 22336 22720 22342 22732
rect 22554 22720 22560 22732
rect 22612 22760 22618 22772
rect 22649 22763 22707 22769
rect 22649 22760 22661 22763
rect 22612 22732 22661 22760
rect 22612 22720 22618 22732
rect 22649 22729 22661 22732
rect 22695 22729 22707 22763
rect 26142 22760 26148 22772
rect 22649 22723 22707 22729
rect 23216 22732 26148 22760
rect 22370 22692 22376 22704
rect 22066 22664 22376 22692
rect 20533 22627 20591 22633
rect 20533 22593 20545 22627
rect 20579 22593 20591 22627
rect 22094 22624 22100 22636
rect 22055 22596 22100 22624
rect 20533 22587 20591 22593
rect 19843 22528 20484 22556
rect 19843 22525 19855 22528
rect 19797 22519 19855 22525
rect 14976 22460 17724 22488
rect 14976 22448 14982 22460
rect 9030 22420 9036 22432
rect 7116 22392 9036 22420
rect 9030 22380 9036 22392
rect 9088 22380 9094 22432
rect 10134 22420 10140 22432
rect 10095 22392 10140 22420
rect 10134 22380 10140 22392
rect 10192 22380 10198 22432
rect 12434 22380 12440 22432
rect 12492 22420 12498 22432
rect 12897 22423 12955 22429
rect 12897 22420 12909 22423
rect 12492 22392 12909 22420
rect 12492 22380 12498 22392
rect 12897 22389 12909 22392
rect 12943 22389 12955 22423
rect 12897 22383 12955 22389
rect 15565 22423 15623 22429
rect 15565 22389 15577 22423
rect 15611 22420 15623 22423
rect 16022 22420 16028 22432
rect 15611 22392 16028 22420
rect 15611 22389 15623 22392
rect 15565 22383 15623 22389
rect 16022 22380 16028 22392
rect 16080 22380 16086 22432
rect 16298 22420 16304 22432
rect 16259 22392 16304 22420
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 16945 22423 17003 22429
rect 16945 22389 16957 22423
rect 16991 22420 17003 22423
rect 17034 22420 17040 22432
rect 16991 22392 17040 22420
rect 16991 22389 17003 22392
rect 16945 22383 17003 22389
rect 17034 22380 17040 22392
rect 17092 22380 17098 22432
rect 17696 22420 17724 22460
rect 17957 22491 18015 22497
rect 17957 22457 17969 22491
rect 18003 22457 18015 22491
rect 17957 22451 18015 22457
rect 19076 22460 20116 22488
rect 19076 22420 19104 22460
rect 17696 22392 19104 22420
rect 19521 22423 19579 22429
rect 19521 22389 19533 22423
rect 19567 22420 19579 22423
rect 19978 22420 19984 22432
rect 19567 22392 19984 22420
rect 19567 22389 19579 22392
rect 19521 22383 19579 22389
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 20088 22420 20116 22460
rect 20162 22448 20168 22500
rect 20220 22488 20226 22500
rect 20548 22488 20576 22587
rect 22094 22584 22100 22596
rect 22152 22584 22158 22636
rect 22204 22633 22232 22664
rect 22370 22652 22376 22664
rect 22428 22652 22434 22704
rect 23216 22701 23244 22732
rect 26142 22720 26148 22732
rect 26200 22720 26206 22772
rect 28626 22760 28632 22772
rect 28587 22732 28632 22760
rect 28626 22720 28632 22732
rect 28684 22720 28690 22772
rect 23109 22695 23167 22701
rect 23109 22692 23121 22695
rect 22572 22664 23121 22692
rect 22189 22627 22247 22633
rect 22189 22593 22201 22627
rect 22235 22593 22247 22627
rect 22189 22587 22247 22593
rect 22465 22627 22523 22633
rect 22465 22593 22477 22627
rect 22511 22593 22523 22627
rect 22465 22587 22523 22593
rect 22112 22556 22140 22584
rect 22480 22556 22508 22587
rect 22112 22528 22508 22556
rect 22572 22488 22600 22664
rect 23109 22661 23121 22664
rect 23155 22661 23167 22695
rect 23109 22655 23167 22661
rect 23201 22695 23259 22701
rect 23201 22661 23213 22695
rect 23247 22661 23259 22695
rect 23201 22655 23259 22661
rect 24670 22652 24676 22704
rect 24728 22652 24734 22704
rect 25498 22652 25504 22704
rect 25556 22692 25562 22704
rect 25869 22695 25927 22701
rect 25869 22692 25881 22695
rect 25556 22664 25881 22692
rect 25556 22652 25562 22664
rect 25869 22661 25881 22664
rect 25915 22661 25927 22695
rect 25869 22655 25927 22661
rect 22925 22627 22983 22633
rect 22925 22593 22937 22627
rect 22971 22593 22983 22627
rect 22925 22587 22983 22593
rect 22940 22556 22968 22587
rect 23290 22584 23296 22636
rect 23348 22633 23354 22636
rect 23348 22624 23356 22633
rect 23658 22624 23664 22636
rect 23348 22596 23393 22624
rect 23619 22596 23664 22624
rect 23348 22587 23356 22596
rect 23348 22584 23354 22587
rect 23658 22584 23664 22596
rect 23716 22584 23722 22636
rect 25590 22624 25596 22636
rect 25551 22596 25596 22624
rect 25590 22584 25596 22596
rect 25648 22584 25654 22636
rect 25682 22584 25688 22636
rect 25740 22624 25746 22636
rect 26050 22633 26056 22636
rect 25777 22627 25835 22633
rect 25777 22624 25789 22627
rect 25740 22596 25789 22624
rect 25740 22584 25746 22596
rect 25777 22593 25789 22596
rect 25823 22593 25835 22627
rect 25777 22587 25835 22593
rect 26013 22627 26056 22633
rect 26013 22593 26025 22627
rect 26013 22587 26056 22593
rect 26050 22584 26056 22587
rect 26108 22584 26114 22636
rect 26510 22624 26516 22636
rect 26471 22596 26516 22624
rect 26510 22584 26516 22596
rect 26568 22584 26574 22636
rect 28077 22627 28135 22633
rect 28077 22593 28089 22627
rect 28123 22624 28135 22627
rect 28166 22624 28172 22636
rect 28123 22596 28172 22624
rect 28123 22593 28135 22596
rect 28077 22587 28135 22593
rect 28166 22584 28172 22596
rect 28224 22584 28230 22636
rect 28445 22627 28503 22633
rect 28445 22624 28457 22627
rect 28276 22596 28457 22624
rect 23198 22556 23204 22568
rect 22940 22528 23204 22556
rect 23198 22516 23204 22528
rect 23256 22516 23262 22568
rect 23934 22556 23940 22568
rect 23895 22528 23940 22556
rect 23934 22516 23940 22528
rect 23992 22516 23998 22568
rect 25406 22556 25412 22568
rect 25367 22528 25412 22556
rect 25406 22516 25412 22528
rect 25464 22516 25470 22568
rect 28276 22497 28304 22596
rect 28445 22593 28457 22596
rect 28491 22593 28503 22627
rect 28445 22587 28503 22593
rect 20220 22460 20576 22488
rect 20640 22460 22094 22488
rect 20220 22448 20226 22460
rect 20346 22420 20352 22432
rect 20088 22392 20352 22420
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 20530 22380 20536 22432
rect 20588 22420 20594 22432
rect 20640 22420 20668 22460
rect 20588 22392 20668 22420
rect 20588 22380 20594 22392
rect 20714 22380 20720 22432
rect 20772 22420 20778 22432
rect 21910 22420 21916 22432
rect 20772 22392 21916 22420
rect 20772 22380 20778 22392
rect 21910 22380 21916 22392
rect 21968 22380 21974 22432
rect 22066 22420 22094 22460
rect 22388 22460 22600 22488
rect 28261 22491 28319 22497
rect 22388 22429 22416 22460
rect 28261 22457 28273 22491
rect 28307 22457 28319 22491
rect 28261 22451 28319 22457
rect 22373 22423 22431 22429
rect 22373 22420 22385 22423
rect 22066 22392 22385 22420
rect 22373 22389 22385 22392
rect 22419 22389 22431 22423
rect 22373 22383 22431 22389
rect 23477 22423 23535 22429
rect 23477 22389 23489 22423
rect 23523 22420 23535 22423
rect 24026 22420 24032 22432
rect 23523 22392 24032 22420
rect 23523 22389 23535 22392
rect 23477 22383 23535 22389
rect 24026 22380 24032 22392
rect 24084 22380 24090 22432
rect 26142 22420 26148 22432
rect 26103 22392 26148 22420
rect 26142 22380 26148 22392
rect 26200 22380 26206 22432
rect 26326 22420 26332 22432
rect 26287 22392 26332 22420
rect 26326 22380 26332 22392
rect 26384 22380 26390 22432
rect 1104 22330 29532 22352
rect 1104 22278 5688 22330
rect 5740 22278 5752 22330
rect 5804 22278 5816 22330
rect 5868 22278 5880 22330
rect 5932 22278 5944 22330
rect 5996 22278 15163 22330
rect 15215 22278 15227 22330
rect 15279 22278 15291 22330
rect 15343 22278 15355 22330
rect 15407 22278 15419 22330
rect 15471 22278 24639 22330
rect 24691 22278 24703 22330
rect 24755 22278 24767 22330
rect 24819 22278 24831 22330
rect 24883 22278 24895 22330
rect 24947 22278 29532 22330
rect 1104 22256 29532 22278
rect 1670 22176 1676 22228
rect 1728 22216 1734 22228
rect 1857 22219 1915 22225
rect 1857 22216 1869 22219
rect 1728 22188 1869 22216
rect 1728 22176 1734 22188
rect 1857 22185 1869 22188
rect 1903 22185 1915 22219
rect 1857 22179 1915 22185
rect 2133 22219 2191 22225
rect 2133 22185 2145 22219
rect 2179 22216 2191 22219
rect 2222 22216 2228 22228
rect 2179 22188 2228 22216
rect 2179 22185 2191 22188
rect 2133 22179 2191 22185
rect 2222 22176 2228 22188
rect 2280 22176 2286 22228
rect 3970 22176 3976 22228
rect 4028 22216 4034 22228
rect 4028 22188 17816 22216
rect 4028 22176 4034 22188
rect 6365 22151 6423 22157
rect 6365 22117 6377 22151
rect 6411 22117 6423 22151
rect 6365 22111 6423 22117
rect 7101 22151 7159 22157
rect 7101 22117 7113 22151
rect 7147 22148 7159 22151
rect 8202 22148 8208 22160
rect 7147 22120 8208 22148
rect 7147 22117 7159 22120
rect 7101 22111 7159 22117
rect 1394 22040 1400 22092
rect 1452 22080 1458 22092
rect 3804 22089 3924 22094
rect 3804 22083 3939 22089
rect 3804 22080 3893 22083
rect 1452 22066 3893 22080
rect 1452 22052 3832 22066
rect 1452 22040 1458 22052
rect 3881 22049 3893 22066
rect 3927 22049 3939 22083
rect 3881 22043 3939 22049
rect 5460 22052 6316 22080
rect 2041 22015 2099 22021
rect 2041 21981 2053 22015
rect 2087 21981 2099 22015
rect 2314 22012 2320 22024
rect 2275 21984 2320 22012
rect 2041 21975 2099 21981
rect 2056 21944 2084 21975
rect 2314 21972 2320 21984
rect 2372 21972 2378 22024
rect 3237 22015 3295 22021
rect 3237 21981 3249 22015
rect 3283 22012 3295 22015
rect 3283 21984 3832 22012
rect 3283 21981 3295 21984
rect 3237 21975 3295 21981
rect 2943 21947 3001 21953
rect 2943 21944 2955 21947
rect 2056 21916 2955 21944
rect 2943 21913 2955 21916
rect 2989 21913 3001 21947
rect 2943 21907 3001 21913
rect 3513 21947 3571 21953
rect 3513 21913 3525 21947
rect 3559 21944 3571 21947
rect 3602 21944 3608 21956
rect 3559 21916 3608 21944
rect 3559 21913 3571 21916
rect 3513 21907 3571 21913
rect 3602 21904 3608 21916
rect 3660 21904 3666 21956
rect 3050 21836 3056 21888
rect 3108 21876 3114 21888
rect 3421 21879 3479 21885
rect 3421 21876 3433 21879
rect 3108 21848 3433 21876
rect 3108 21836 3114 21848
rect 3421 21845 3433 21848
rect 3467 21845 3479 21879
rect 3804 21876 3832 21984
rect 4154 21944 4160 21956
rect 4115 21916 4160 21944
rect 4154 21904 4160 21916
rect 4212 21904 4218 21956
rect 5166 21904 5172 21956
rect 5224 21904 5230 21956
rect 5460 21876 5488 22052
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 21981 6239 22015
rect 6181 21975 6239 21981
rect 6196 21888 6224 21975
rect 6288 21944 6316 22052
rect 6380 22012 6408 22111
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 12158 22108 12164 22160
rect 12216 22148 12222 22160
rect 12216 22120 12664 22148
rect 12216 22108 12222 22120
rect 6546 22080 6552 22092
rect 6507 22052 6552 22080
rect 6546 22040 6552 22052
rect 6604 22040 6610 22092
rect 12636 22089 12664 22120
rect 14826 22108 14832 22160
rect 14884 22148 14890 22160
rect 15105 22151 15163 22157
rect 15105 22148 15117 22151
rect 14884 22120 15117 22148
rect 14884 22108 14890 22120
rect 15105 22117 15117 22120
rect 15151 22117 15163 22151
rect 17218 22148 17224 22160
rect 17131 22120 17224 22148
rect 15105 22111 15163 22117
rect 17218 22108 17224 22120
rect 17276 22148 17282 22160
rect 17678 22148 17684 22160
rect 17276 22120 17684 22148
rect 17276 22108 17282 22120
rect 17678 22108 17684 22120
rect 17736 22108 17742 22160
rect 17788 22148 17816 22188
rect 20070 22176 20076 22228
rect 20128 22216 20134 22228
rect 20530 22216 20536 22228
rect 20128 22188 20536 22216
rect 20128 22176 20134 22188
rect 20530 22176 20536 22188
rect 20588 22176 20594 22228
rect 20717 22219 20775 22225
rect 20717 22185 20729 22219
rect 20763 22216 20775 22219
rect 20806 22216 20812 22228
rect 20763 22188 20812 22216
rect 20763 22185 20775 22188
rect 20717 22179 20775 22185
rect 20806 22176 20812 22188
rect 20864 22176 20870 22228
rect 22094 22176 22100 22228
rect 22152 22216 22158 22228
rect 22557 22219 22615 22225
rect 22557 22216 22569 22219
rect 22152 22188 22569 22216
rect 22152 22176 22158 22188
rect 22557 22185 22569 22188
rect 22603 22185 22615 22219
rect 23934 22216 23940 22228
rect 23895 22188 23940 22216
rect 22557 22179 22615 22185
rect 23934 22176 23940 22188
rect 23992 22176 23998 22228
rect 24486 22176 24492 22228
rect 24544 22216 24550 22228
rect 24581 22219 24639 22225
rect 24581 22216 24593 22219
rect 24544 22188 24593 22216
rect 24544 22176 24550 22188
rect 24581 22185 24593 22188
rect 24627 22185 24639 22219
rect 24581 22179 24639 22185
rect 26142 22176 26148 22228
rect 26200 22216 26206 22228
rect 26893 22219 26951 22225
rect 26893 22216 26905 22219
rect 26200 22188 26905 22216
rect 26200 22176 26206 22188
rect 26893 22185 26905 22188
rect 26939 22185 26951 22219
rect 26893 22179 26951 22185
rect 25409 22151 25467 22157
rect 25409 22148 25421 22151
rect 17788 22120 21036 22148
rect 7193 22083 7251 22089
rect 7193 22049 7205 22083
rect 7239 22049 7251 22083
rect 7193 22043 7251 22049
rect 12621 22083 12679 22089
rect 12621 22049 12633 22083
rect 12667 22049 12679 22083
rect 13173 22083 13231 22089
rect 13173 22080 13185 22083
rect 12621 22043 12679 22049
rect 12912 22052 13185 22080
rect 6638 22012 6644 22024
rect 6380 21984 6644 22012
rect 6638 21972 6644 21984
rect 6696 22012 6702 22024
rect 7208 22012 7236 22043
rect 6696 21984 7236 22012
rect 7285 22015 7343 22021
rect 6696 21972 6702 21984
rect 7285 21981 7297 22015
rect 7331 22012 7343 22015
rect 7331 21984 9536 22012
rect 7331 21981 7343 21984
rect 7285 21975 7343 21981
rect 9214 21944 9220 21956
rect 6288 21916 9220 21944
rect 9214 21904 9220 21916
rect 9272 21904 9278 21956
rect 9508 21944 9536 21984
rect 9582 21972 9588 22024
rect 9640 22012 9646 22024
rect 10413 22015 10471 22021
rect 10413 22012 10425 22015
rect 9640 21984 10425 22012
rect 9640 21972 9646 21984
rect 10413 21981 10425 21984
rect 10459 22012 10471 22015
rect 10505 22015 10563 22021
rect 10505 22012 10517 22015
rect 10459 21984 10517 22012
rect 10459 21981 10471 21984
rect 10413 21975 10471 21981
rect 10505 21981 10517 21984
rect 10551 21981 10563 22015
rect 12912 22012 12940 22052
rect 13173 22049 13185 22052
rect 13219 22049 13231 22083
rect 13998 22080 14004 22092
rect 13173 22043 13231 22049
rect 13280 22052 14004 22080
rect 10505 21975 10563 21981
rect 10612 21984 12940 22012
rect 13081 22015 13139 22021
rect 10134 21944 10140 21956
rect 10192 21953 10198 21956
rect 9508 21916 9996 21944
rect 10104 21916 10140 21944
rect 5626 21876 5632 21888
rect 3804 21848 5488 21876
rect 5587 21848 5632 21876
rect 3421 21839 3479 21845
rect 5626 21836 5632 21848
rect 5684 21836 5690 21888
rect 6178 21876 6184 21888
rect 6091 21848 6184 21876
rect 6178 21836 6184 21848
rect 6236 21876 6242 21888
rect 8662 21876 8668 21888
rect 6236 21848 8668 21876
rect 6236 21836 6242 21848
rect 8662 21836 8668 21848
rect 8720 21836 8726 21888
rect 9033 21879 9091 21885
rect 9033 21845 9045 21879
rect 9079 21876 9091 21879
rect 9766 21876 9772 21888
rect 9079 21848 9772 21876
rect 9079 21845 9091 21848
rect 9033 21839 9091 21845
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 9968 21876 9996 21916
rect 10134 21904 10140 21916
rect 10192 21907 10204 21953
rect 10192 21904 10198 21907
rect 10612 21876 10640 21984
rect 13081 21981 13093 22015
rect 13127 22012 13139 22015
rect 13280 22012 13308 22052
rect 13998 22040 14004 22052
rect 14056 22040 14062 22092
rect 14734 22080 14740 22092
rect 14695 22052 14740 22080
rect 14734 22040 14740 22052
rect 14792 22040 14798 22092
rect 15396 22052 17356 22080
rect 13127 21984 13308 22012
rect 13357 22015 13415 22021
rect 13127 21981 13139 21984
rect 13081 21975 13139 21981
rect 13357 21981 13369 22015
rect 13403 21981 13415 22015
rect 13538 22012 13544 22024
rect 13499 21984 13544 22012
rect 13357 21975 13415 21981
rect 10778 21953 10784 21956
rect 10772 21907 10784 21953
rect 10836 21944 10842 21956
rect 12529 21947 12587 21953
rect 12529 21944 12541 21947
rect 10836 21916 10872 21944
rect 11900 21916 12541 21944
rect 10778 21904 10784 21907
rect 10836 21904 10842 21916
rect 11900 21888 11928 21916
rect 12529 21913 12541 21916
rect 12575 21913 12587 21947
rect 13372 21944 13400 21975
rect 13538 21972 13544 21984
rect 13596 21972 13602 22024
rect 13814 22012 13820 22024
rect 13775 21984 13820 22012
rect 13814 21972 13820 21984
rect 13872 21972 13878 22024
rect 14458 22012 14464 22024
rect 14419 21984 14464 22012
rect 14458 21972 14464 21984
rect 14516 21972 14522 22024
rect 15286 22012 15292 22024
rect 15247 21984 15292 22012
rect 15286 21972 15292 21984
rect 15344 21972 15350 22024
rect 15396 21944 15424 22052
rect 15473 22015 15531 22021
rect 15473 21981 15485 22015
rect 15519 21981 15531 22015
rect 17328 22012 17356 22052
rect 17402 22040 17408 22092
rect 17460 22080 17466 22092
rect 18230 22080 18236 22092
rect 17460 22052 18236 22080
rect 17460 22040 17466 22052
rect 18230 22040 18236 22052
rect 18288 22080 18294 22092
rect 18874 22080 18880 22092
rect 18288 22052 18880 22080
rect 18288 22040 18294 22052
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 19794 22040 19800 22092
rect 19852 22080 19858 22092
rect 20070 22080 20076 22092
rect 19852 22052 20076 22080
rect 19852 22040 19858 22052
rect 20070 22040 20076 22052
rect 20128 22080 20134 22092
rect 20128 22052 20484 22080
rect 20128 22040 20134 22052
rect 19702 22012 19708 22024
rect 17328 21984 19708 22012
rect 15473 21975 15531 21981
rect 13372 21916 15424 21944
rect 12529 21907 12587 21913
rect 11882 21876 11888 21888
rect 9968 21848 10640 21876
rect 11843 21848 11888 21876
rect 11882 21836 11888 21848
rect 11940 21836 11946 21888
rect 12069 21879 12127 21885
rect 12069 21845 12081 21879
rect 12115 21876 12127 21879
rect 12342 21876 12348 21888
rect 12115 21848 12348 21876
rect 12115 21845 12127 21848
rect 12069 21839 12127 21845
rect 12342 21836 12348 21848
rect 12400 21836 12406 21888
rect 12434 21836 12440 21888
rect 12492 21876 12498 21888
rect 12492 21848 12537 21876
rect 12492 21836 12498 21848
rect 13998 21836 14004 21888
rect 14056 21876 14062 21888
rect 14093 21879 14151 21885
rect 14093 21876 14105 21879
rect 14056 21848 14105 21876
rect 14056 21836 14062 21848
rect 14093 21845 14105 21848
rect 14139 21845 14151 21879
rect 14093 21839 14151 21845
rect 14553 21879 14611 21885
rect 14553 21845 14565 21879
rect 14599 21876 14611 21879
rect 14642 21876 14648 21888
rect 14599 21848 14648 21876
rect 14599 21845 14611 21848
rect 14553 21839 14611 21845
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 15488 21876 15516 21975
rect 19702 21972 19708 21984
rect 19760 21972 19766 22024
rect 19886 22012 19892 22024
rect 19847 21984 19892 22012
rect 19886 21972 19892 21984
rect 19944 21972 19950 22024
rect 20165 22015 20223 22021
rect 20165 21981 20177 22015
rect 20211 21981 20223 22015
rect 20346 22012 20352 22024
rect 20307 21984 20352 22012
rect 20165 21975 20223 21981
rect 15749 21947 15807 21953
rect 15749 21913 15761 21947
rect 15795 21944 15807 21947
rect 16022 21944 16028 21956
rect 15795 21916 16028 21944
rect 15795 21913 15807 21916
rect 15749 21907 15807 21913
rect 16022 21904 16028 21916
rect 16080 21904 16086 21956
rect 17034 21944 17040 21956
rect 16974 21916 17040 21944
rect 17034 21904 17040 21916
rect 17092 21904 17098 21956
rect 20180 21944 20208 21975
rect 20346 21972 20352 21984
rect 20404 21972 20410 22024
rect 20456 22021 20484 22052
rect 20441 22015 20499 22021
rect 20441 21981 20453 22015
rect 20487 21981 20499 22015
rect 20441 21975 20499 21981
rect 20530 21972 20536 22024
rect 20588 22021 20594 22024
rect 20588 22012 20596 22021
rect 21008 22012 21036 22120
rect 22204 22120 25421 22148
rect 21082 22040 21088 22092
rect 21140 22080 21146 22092
rect 21177 22083 21235 22089
rect 21177 22080 21189 22083
rect 21140 22052 21189 22080
rect 21140 22040 21146 22052
rect 21177 22049 21189 22052
rect 21223 22049 21235 22083
rect 21177 22043 21235 22049
rect 22204 22012 22232 22120
rect 25409 22117 25421 22120
rect 25455 22148 25467 22151
rect 25498 22148 25504 22160
rect 25455 22120 25504 22148
rect 25455 22117 25467 22120
rect 25409 22111 25467 22117
rect 25498 22108 25504 22120
rect 25556 22108 25562 22160
rect 23290 22040 23296 22092
rect 23348 22080 23354 22092
rect 23348 22052 23704 22080
rect 23348 22040 23354 22052
rect 22830 22012 22836 22024
rect 20588 21984 20633 22012
rect 21008 21984 22232 22012
rect 22791 21984 22836 22012
rect 20588 21975 20596 21984
rect 20588 21972 20594 21975
rect 22830 21972 22836 21984
rect 22888 22012 22894 22024
rect 23109 22015 23167 22021
rect 23109 22012 23121 22015
rect 22888 21984 23121 22012
rect 22888 21972 22894 21984
rect 23109 21981 23121 21984
rect 23155 21981 23167 22015
rect 23109 21975 23167 21981
rect 23198 21972 23204 22024
rect 23256 22012 23262 22024
rect 23385 22015 23443 22021
rect 23385 22012 23397 22015
rect 23256 21984 23397 22012
rect 23256 21972 23262 21984
rect 23385 21981 23397 21984
rect 23431 21981 23443 22015
rect 23676 22012 23704 22052
rect 23758 22015 23816 22021
rect 23758 22012 23770 22015
rect 23676 21984 23770 22012
rect 23385 21975 23443 21981
rect 23758 21981 23770 21984
rect 23804 21981 23816 22015
rect 23758 21975 23816 21981
rect 24397 22015 24455 22021
rect 24397 21981 24409 22015
rect 24443 22012 24455 22015
rect 24486 22012 24492 22024
rect 24443 21984 24492 22012
rect 24443 21981 24455 21984
rect 24397 21975 24455 21981
rect 24486 21972 24492 21984
rect 24544 21972 24550 22024
rect 27154 21972 27160 22024
rect 27212 22012 27218 22024
rect 27212 21984 27257 22012
rect 27212 21972 27218 21984
rect 20254 21944 20260 21956
rect 20180 21916 20260 21944
rect 20254 21904 20260 21916
rect 20312 21904 20318 21956
rect 20990 21904 20996 21956
rect 21048 21944 21054 21956
rect 21422 21947 21480 21953
rect 21422 21944 21434 21947
rect 21048 21916 21434 21944
rect 21048 21904 21054 21916
rect 21422 21913 21434 21916
rect 21468 21913 21480 21947
rect 21422 21907 21480 21913
rect 21910 21904 21916 21956
rect 21968 21944 21974 21956
rect 23014 21944 23020 21956
rect 21968 21916 22876 21944
rect 22975 21916 23020 21944
rect 21968 21904 21974 21916
rect 15838 21876 15844 21888
rect 15488 21848 15844 21876
rect 15838 21836 15844 21848
rect 15896 21876 15902 21888
rect 17954 21876 17960 21888
rect 15896 21848 17960 21876
rect 15896 21836 15902 21848
rect 17954 21836 17960 21848
rect 18012 21836 18018 21888
rect 19610 21836 19616 21888
rect 19668 21876 19674 21888
rect 20073 21879 20131 21885
rect 20073 21876 20085 21879
rect 19668 21848 20085 21876
rect 19668 21836 19674 21848
rect 20073 21845 20085 21848
rect 20119 21876 20131 21879
rect 22646 21876 22652 21888
rect 20119 21848 22652 21876
rect 20119 21845 20131 21848
rect 20073 21839 20131 21845
rect 22646 21836 22652 21848
rect 22704 21836 22710 21888
rect 22848 21876 22876 21916
rect 23014 21904 23020 21916
rect 23072 21904 23078 21956
rect 23569 21947 23627 21953
rect 23569 21913 23581 21947
rect 23615 21913 23627 21947
rect 23569 21907 23627 21913
rect 23661 21947 23719 21953
rect 23661 21913 23673 21947
rect 23707 21944 23719 21947
rect 25406 21944 25412 21956
rect 23707 21916 25412 21944
rect 23707 21913 23719 21916
rect 23661 21907 23719 21913
rect 23584 21876 23612 21907
rect 25406 21904 25412 21916
rect 25464 21904 25470 21956
rect 26326 21904 26332 21956
rect 26384 21904 26390 21956
rect 22848 21848 23612 21876
rect 24026 21836 24032 21888
rect 24084 21876 24090 21888
rect 24302 21876 24308 21888
rect 24084 21848 24308 21876
rect 24084 21836 24090 21848
rect 24302 21836 24308 21848
rect 24360 21836 24366 21888
rect 25958 21836 25964 21888
rect 26016 21876 26022 21888
rect 26510 21876 26516 21888
rect 26016 21848 26516 21876
rect 26016 21836 26022 21848
rect 26510 21836 26516 21848
rect 26568 21836 26574 21888
rect 1104 21786 29532 21808
rect 1104 21734 10425 21786
rect 10477 21734 10489 21786
rect 10541 21734 10553 21786
rect 10605 21734 10617 21786
rect 10669 21734 10681 21786
rect 10733 21734 19901 21786
rect 19953 21734 19965 21786
rect 20017 21734 20029 21786
rect 20081 21734 20093 21786
rect 20145 21734 20157 21786
rect 20209 21734 29532 21786
rect 1104 21712 29532 21734
rect 3418 21672 3424 21684
rect 3379 21644 3424 21672
rect 3418 21632 3424 21644
rect 3476 21632 3482 21684
rect 4154 21632 4160 21684
rect 4212 21672 4218 21684
rect 4433 21675 4491 21681
rect 4433 21672 4445 21675
rect 4212 21644 4445 21672
rect 4212 21632 4218 21644
rect 4433 21641 4445 21644
rect 4479 21641 4491 21675
rect 4433 21635 4491 21641
rect 5074 21632 5080 21684
rect 5132 21672 5138 21684
rect 5721 21675 5779 21681
rect 5721 21672 5733 21675
rect 5132 21644 5733 21672
rect 5132 21632 5138 21644
rect 5721 21641 5733 21644
rect 5767 21641 5779 21675
rect 10505 21675 10563 21681
rect 5721 21635 5779 21641
rect 5828 21644 10456 21672
rect 4522 21564 4528 21616
rect 4580 21604 4586 21616
rect 5445 21607 5503 21613
rect 5445 21604 5457 21607
rect 4580 21576 5457 21604
rect 4580 21564 4586 21576
rect 5445 21573 5457 21576
rect 5491 21604 5503 21607
rect 5626 21604 5632 21616
rect 5491 21576 5632 21604
rect 5491 21573 5503 21576
rect 5445 21567 5503 21573
rect 5626 21564 5632 21576
rect 5684 21564 5690 21616
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21536 4675 21539
rect 4967 21539 5025 21545
rect 4967 21536 4979 21539
rect 4663 21508 4979 21536
rect 4663 21505 4675 21508
rect 4617 21499 4675 21505
rect 4967 21505 4979 21508
rect 5013 21505 5025 21539
rect 4967 21499 5025 21505
rect 5261 21539 5319 21545
rect 5261 21505 5273 21539
rect 5307 21536 5319 21539
rect 5828 21536 5856 21644
rect 7558 21564 7564 21616
rect 7616 21564 7622 21616
rect 8386 21564 8392 21616
rect 8444 21604 8450 21616
rect 9585 21607 9643 21613
rect 8444 21576 8892 21604
rect 8444 21564 8450 21576
rect 5307 21508 5856 21536
rect 5905 21539 5963 21545
rect 5307 21505 5319 21508
rect 5261 21499 5319 21505
rect 5905 21505 5917 21539
rect 5951 21536 5963 21539
rect 6089 21539 6147 21545
rect 6089 21536 6101 21539
rect 5951 21508 6101 21536
rect 5951 21505 5963 21508
rect 5905 21499 5963 21505
rect 6089 21505 6101 21508
rect 6135 21536 6147 21539
rect 7006 21536 7012 21548
rect 6135 21508 7012 21536
rect 6135 21505 6147 21508
rect 6089 21499 6147 21505
rect 7006 21496 7012 21508
rect 7064 21496 7070 21548
rect 8864 21545 8892 21576
rect 9585 21573 9597 21607
rect 9631 21604 9643 21607
rect 10318 21604 10324 21616
rect 9631 21576 10324 21604
rect 9631 21573 9643 21576
rect 9585 21567 9643 21573
rect 10318 21564 10324 21576
rect 10376 21564 10382 21616
rect 10428 21604 10456 21644
rect 10505 21641 10517 21675
rect 10551 21672 10563 21675
rect 10778 21672 10784 21684
rect 10551 21644 10784 21672
rect 10551 21641 10563 21644
rect 10505 21635 10563 21641
rect 10778 21632 10784 21644
rect 10836 21632 10842 21684
rect 15286 21632 15292 21684
rect 15344 21672 15350 21684
rect 16206 21672 16212 21684
rect 15344 21644 16212 21672
rect 15344 21632 15350 21644
rect 16206 21632 16212 21644
rect 16264 21632 16270 21684
rect 16666 21632 16672 21684
rect 16724 21672 16730 21684
rect 17773 21675 17831 21681
rect 17773 21672 17785 21675
rect 16724 21644 17785 21672
rect 16724 21632 16730 21644
rect 17773 21641 17785 21644
rect 17819 21641 17831 21675
rect 17773 21635 17831 21641
rect 13998 21604 14004 21616
rect 10428 21576 14004 21604
rect 13998 21564 14004 21576
rect 14056 21564 14062 21616
rect 15378 21604 15384 21616
rect 15339 21576 15384 21604
rect 15378 21564 15384 21576
rect 15436 21564 15442 21616
rect 15473 21607 15531 21613
rect 15473 21573 15485 21607
rect 15519 21604 15531 21607
rect 17788 21604 17816 21635
rect 17862 21632 17868 21684
rect 17920 21672 17926 21684
rect 19429 21675 19487 21681
rect 19429 21672 19441 21675
rect 17920 21644 19441 21672
rect 17920 21632 17926 21644
rect 19429 21641 19441 21644
rect 19475 21641 19487 21675
rect 19429 21635 19487 21641
rect 19702 21632 19708 21684
rect 19760 21672 19766 21684
rect 22094 21672 22100 21684
rect 19760 21644 22100 21672
rect 19760 21632 19766 21644
rect 22094 21632 22100 21644
rect 22152 21632 22158 21684
rect 22646 21632 22652 21684
rect 22704 21672 22710 21684
rect 27338 21672 27344 21684
rect 22704 21644 27344 21672
rect 22704 21632 22710 21644
rect 15519 21576 15608 21604
rect 17788 21576 18092 21604
rect 15519 21573 15531 21576
rect 15473 21567 15531 21573
rect 8849 21539 8907 21545
rect 8849 21505 8861 21539
rect 8895 21505 8907 21539
rect 8849 21499 8907 21505
rect 9122 21496 9128 21548
rect 9180 21536 9186 21548
rect 9217 21539 9275 21545
rect 9217 21536 9229 21539
rect 9180 21508 9229 21536
rect 9180 21496 9186 21508
rect 9217 21505 9229 21508
rect 9263 21505 9275 21539
rect 9398 21536 9404 21548
rect 9359 21508 9404 21536
rect 9217 21499 9275 21505
rect 9398 21496 9404 21508
rect 9456 21496 9462 21548
rect 9858 21536 9864 21548
rect 9819 21508 9864 21536
rect 9858 21496 9864 21508
rect 9916 21496 9922 21548
rect 10026 21539 10084 21545
rect 10026 21536 10038 21539
rect 9968 21508 10038 21536
rect 3142 21468 3148 21480
rect 3103 21440 3148 21468
rect 3142 21428 3148 21440
rect 3200 21428 3206 21480
rect 3234 21428 3240 21480
rect 3292 21468 3298 21480
rect 3329 21471 3387 21477
rect 3329 21468 3341 21471
rect 3292 21440 3341 21468
rect 3292 21428 3298 21440
rect 3329 21437 3341 21440
rect 3375 21437 3387 21471
rect 3329 21431 3387 21437
rect 3602 21428 3608 21480
rect 3660 21468 3666 21480
rect 5537 21471 5595 21477
rect 5537 21468 5549 21471
rect 3660 21440 5549 21468
rect 3660 21428 3666 21440
rect 5537 21437 5549 21440
rect 5583 21468 5595 21471
rect 6178 21468 6184 21480
rect 5583 21440 6184 21468
rect 5583 21437 5595 21440
rect 5537 21431 5595 21437
rect 6178 21428 6184 21440
rect 6236 21428 6242 21480
rect 8294 21468 8300 21480
rect 8255 21440 8300 21468
rect 8294 21428 8300 21440
rect 8352 21428 8358 21480
rect 8570 21468 8576 21480
rect 8531 21440 8576 21468
rect 8570 21428 8576 21440
rect 8628 21428 8634 21480
rect 8938 21428 8944 21480
rect 8996 21468 9002 21480
rect 9677 21471 9735 21477
rect 9677 21468 9689 21471
rect 8996 21440 9689 21468
rect 8996 21428 9002 21440
rect 9677 21437 9689 21440
rect 9723 21468 9735 21471
rect 9968 21468 9996 21508
rect 10026 21505 10038 21508
rect 10072 21505 10084 21539
rect 10226 21536 10232 21548
rect 10187 21508 10232 21536
rect 10026 21499 10084 21505
rect 10226 21496 10232 21508
rect 10284 21496 10290 21548
rect 10413 21539 10471 21545
rect 10413 21505 10425 21539
rect 10459 21536 10471 21539
rect 11882 21536 11888 21548
rect 10459 21508 11888 21536
rect 10459 21505 10471 21508
rect 10413 21499 10471 21505
rect 11882 21496 11888 21508
rect 11940 21496 11946 21548
rect 12437 21539 12495 21545
rect 12437 21505 12449 21539
rect 12483 21536 12495 21539
rect 12526 21536 12532 21548
rect 12483 21508 12532 21536
rect 12483 21505 12495 21508
rect 12437 21499 12495 21505
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 12618 21496 12624 21548
rect 12676 21536 12682 21548
rect 12713 21539 12771 21545
rect 12713 21536 12725 21539
rect 12676 21508 12725 21536
rect 12676 21496 12682 21508
rect 12713 21505 12725 21508
rect 12759 21505 12771 21539
rect 12713 21499 12771 21505
rect 13078 21496 13084 21548
rect 13136 21536 13142 21548
rect 13265 21539 13323 21545
rect 13265 21536 13277 21539
rect 13136 21508 13277 21536
rect 13136 21496 13142 21508
rect 13265 21505 13277 21508
rect 13311 21536 13323 21539
rect 13538 21536 13544 21548
rect 13311 21508 13544 21536
rect 13311 21505 13323 21508
rect 13265 21499 13323 21505
rect 13538 21496 13544 21508
rect 13596 21496 13602 21548
rect 14090 21536 14096 21548
rect 14003 21508 14096 21536
rect 14090 21496 14096 21508
rect 14148 21536 14154 21548
rect 14458 21536 14464 21548
rect 14148 21508 14464 21536
rect 14148 21496 14154 21508
rect 14458 21496 14464 21508
rect 14516 21496 14522 21548
rect 14734 21496 14740 21548
rect 14792 21536 14798 21548
rect 15580 21536 15608 21576
rect 15930 21536 15936 21548
rect 14792 21508 15516 21536
rect 15580 21508 15936 21536
rect 14792 21496 14798 21508
rect 10134 21468 10140 21480
rect 9723 21440 9996 21468
rect 10095 21440 10140 21468
rect 9723 21437 9735 21440
rect 9677 21431 9735 21437
rect 10134 21428 10140 21440
rect 10192 21428 10198 21480
rect 10502 21428 10508 21480
rect 10560 21468 10566 21480
rect 15488 21468 15516 21508
rect 15930 21496 15936 21508
rect 15988 21496 15994 21548
rect 17126 21536 17132 21548
rect 17087 21508 17132 21536
rect 17126 21496 17132 21508
rect 17184 21496 17190 21548
rect 18064 21545 18092 21576
rect 18138 21564 18144 21616
rect 18196 21604 18202 21616
rect 19794 21604 19800 21616
rect 18196 21576 19800 21604
rect 18196 21564 18202 21576
rect 19794 21564 19800 21576
rect 19852 21604 19858 21616
rect 20625 21607 20683 21613
rect 20625 21604 20637 21607
rect 19852 21576 20637 21604
rect 19852 21564 19858 21576
rect 20625 21573 20637 21576
rect 20671 21573 20683 21607
rect 20625 21567 20683 21573
rect 23014 21564 23020 21616
rect 23072 21604 23078 21616
rect 24029 21607 24087 21613
rect 24029 21604 24041 21607
rect 23072 21576 24041 21604
rect 23072 21564 23078 21576
rect 24029 21573 24041 21576
rect 24075 21573 24087 21607
rect 24029 21567 24087 21573
rect 25590 21564 25596 21616
rect 25648 21604 25654 21616
rect 25648 21576 26188 21604
rect 25648 21564 25654 21576
rect 17957 21539 18015 21545
rect 17957 21505 17969 21539
rect 18003 21505 18015 21539
rect 17957 21499 18015 21505
rect 18049 21539 18107 21545
rect 18049 21505 18061 21539
rect 18095 21505 18107 21539
rect 18049 21499 18107 21505
rect 19613 21539 19671 21545
rect 19613 21505 19625 21539
rect 19659 21536 19671 21539
rect 19659 21508 20208 21536
rect 19659 21505 19671 21508
rect 19613 21499 19671 21505
rect 15657 21471 15715 21477
rect 15657 21468 15669 21471
rect 10560 21440 15148 21468
rect 15488 21440 15669 21468
rect 10560 21428 10566 21440
rect 1486 21360 1492 21412
rect 1544 21400 1550 21412
rect 12342 21400 12348 21412
rect 1544 21372 7328 21400
rect 1544 21360 1550 21372
rect 3510 21292 3516 21344
rect 3568 21332 3574 21344
rect 3789 21335 3847 21341
rect 3789 21332 3801 21335
rect 3568 21304 3801 21332
rect 3568 21292 3574 21304
rect 3789 21301 3801 21304
rect 3835 21301 3847 21335
rect 3789 21295 3847 21301
rect 6730 21292 6736 21344
rect 6788 21332 6794 21344
rect 6825 21335 6883 21341
rect 6825 21332 6837 21335
rect 6788 21304 6837 21332
rect 6788 21292 6794 21304
rect 6825 21301 6837 21304
rect 6871 21301 6883 21335
rect 7300 21332 7328 21372
rect 8496 21372 12348 21400
rect 8496 21332 8524 21372
rect 12342 21360 12348 21372
rect 12400 21360 12406 21412
rect 12618 21400 12624 21412
rect 12579 21372 12624 21400
rect 12618 21360 12624 21372
rect 12676 21360 12682 21412
rect 15013 21403 15071 21409
rect 15013 21400 15025 21403
rect 12728 21372 15025 21400
rect 8662 21332 8668 21344
rect 7300 21304 8524 21332
rect 8623 21304 8668 21332
rect 6825 21295 6883 21301
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 9030 21332 9036 21344
rect 8991 21304 9036 21332
rect 9030 21292 9036 21304
rect 9088 21292 9094 21344
rect 9214 21292 9220 21344
rect 9272 21332 9278 21344
rect 12728 21332 12756 21372
rect 15013 21369 15025 21372
rect 15059 21369 15071 21403
rect 15120 21400 15148 21440
rect 15657 21437 15669 21440
rect 15703 21468 15715 21471
rect 16114 21468 16120 21480
rect 15703 21440 16120 21468
rect 15703 21437 15715 21440
rect 15657 21431 15715 21437
rect 16114 21428 16120 21440
rect 16172 21428 16178 21480
rect 17972 21468 18000 21499
rect 18138 21468 18144 21480
rect 17972 21440 18144 21468
rect 18138 21428 18144 21440
rect 18196 21428 18202 21480
rect 19794 21400 19800 21412
rect 15120 21372 19800 21400
rect 15013 21363 15071 21369
rect 19794 21360 19800 21372
rect 19852 21360 19858 21412
rect 12894 21332 12900 21344
rect 9272 21304 12756 21332
rect 12855 21304 12900 21332
rect 9272 21292 9278 21304
rect 12894 21292 12900 21304
rect 12952 21292 12958 21344
rect 13262 21292 13268 21344
rect 13320 21332 13326 21344
rect 13449 21335 13507 21341
rect 13449 21332 13461 21335
rect 13320 21304 13461 21332
rect 13320 21292 13326 21304
rect 13449 21301 13461 21304
rect 13495 21301 13507 21335
rect 13449 21295 13507 21301
rect 14277 21335 14335 21341
rect 14277 21301 14289 21335
rect 14323 21332 14335 21335
rect 14918 21332 14924 21344
rect 14323 21304 14924 21332
rect 14323 21301 14335 21304
rect 14277 21295 14335 21301
rect 14918 21292 14924 21304
rect 14976 21332 14982 21344
rect 15654 21332 15660 21344
rect 14976 21304 15660 21332
rect 14976 21292 14982 21304
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 16850 21292 16856 21344
rect 16908 21332 16914 21344
rect 16945 21335 17003 21341
rect 16945 21332 16957 21335
rect 16908 21304 16957 21332
rect 16908 21292 16914 21304
rect 16945 21301 16957 21304
rect 16991 21301 17003 21335
rect 16945 21295 17003 21301
rect 18233 21335 18291 21341
rect 18233 21301 18245 21335
rect 18279 21332 18291 21335
rect 18966 21332 18972 21344
rect 18279 21304 18972 21332
rect 18279 21301 18291 21304
rect 18233 21295 18291 21301
rect 18966 21292 18972 21304
rect 19024 21292 19030 21344
rect 20180 21332 20208 21508
rect 20254 21496 20260 21548
rect 20312 21536 20318 21548
rect 20441 21539 20499 21545
rect 20441 21536 20453 21539
rect 20312 21508 20453 21536
rect 20312 21496 20318 21508
rect 20441 21505 20453 21508
rect 20487 21505 20499 21539
rect 20441 21499 20499 21505
rect 20714 21496 20720 21548
rect 20772 21536 20778 21548
rect 20861 21539 20919 21545
rect 20772 21508 20817 21536
rect 20772 21496 20778 21508
rect 20861 21505 20873 21539
rect 20907 21536 20919 21539
rect 22830 21536 22836 21548
rect 20907 21505 20944 21536
rect 22791 21508 22836 21536
rect 20861 21499 20944 21505
rect 20346 21428 20352 21480
rect 20404 21468 20410 21480
rect 20530 21468 20536 21480
rect 20404 21440 20536 21468
rect 20404 21428 20410 21440
rect 20530 21428 20536 21440
rect 20588 21468 20594 21480
rect 20916 21468 20944 21499
rect 22830 21496 22836 21508
rect 22888 21496 22894 21548
rect 24210 21496 24216 21548
rect 24268 21536 24274 21548
rect 24305 21539 24363 21545
rect 24305 21536 24317 21539
rect 24268 21508 24317 21536
rect 24268 21496 24274 21508
rect 24305 21505 24317 21508
rect 24351 21505 24363 21539
rect 24305 21499 24363 21505
rect 24486 21496 24492 21548
rect 24544 21536 24550 21548
rect 26160 21545 26188 21576
rect 26234 21564 26240 21616
rect 26292 21564 26298 21616
rect 26344 21613 26372 21644
rect 27338 21632 27344 21644
rect 27396 21632 27402 21684
rect 28810 21672 28816 21684
rect 27724 21644 28816 21672
rect 26329 21607 26387 21613
rect 26329 21573 26341 21607
rect 26375 21573 26387 21607
rect 26329 21567 26387 21573
rect 26421 21607 26479 21613
rect 26421 21573 26433 21607
rect 26467 21604 26479 21607
rect 27724 21604 27752 21644
rect 28810 21632 28816 21644
rect 28868 21632 28874 21684
rect 26467 21576 27752 21604
rect 26467 21573 26479 21576
rect 26421 21567 26479 21573
rect 27982 21564 27988 21616
rect 28040 21564 28046 21616
rect 24581 21539 24639 21545
rect 24581 21536 24593 21539
rect 24544 21508 24593 21536
rect 24544 21496 24550 21508
rect 24581 21505 24593 21508
rect 24627 21505 24639 21539
rect 24581 21499 24639 21505
rect 25869 21539 25927 21545
rect 25869 21505 25881 21539
rect 25915 21505 25927 21539
rect 25869 21499 25927 21505
rect 26145 21539 26203 21545
rect 26145 21505 26157 21539
rect 26191 21505 26203 21539
rect 26252 21536 26280 21564
rect 26518 21539 26576 21545
rect 26518 21536 26530 21539
rect 26252 21508 26530 21536
rect 26145 21499 26203 21505
rect 26518 21505 26530 21508
rect 26564 21505 26576 21539
rect 26518 21499 26576 21505
rect 20588 21440 20944 21468
rect 20588 21428 20594 21440
rect 20990 21400 20996 21412
rect 20951 21372 20996 21400
rect 20990 21360 20996 21372
rect 21048 21360 21054 21412
rect 24213 21403 24271 21409
rect 24213 21369 24225 21403
rect 24259 21400 24271 21403
rect 24302 21400 24308 21412
rect 24259 21372 24308 21400
rect 24259 21369 24271 21372
rect 24213 21363 24271 21369
rect 24302 21360 24308 21372
rect 24360 21360 24366 21412
rect 21082 21332 21088 21344
rect 20180 21304 21088 21332
rect 21082 21292 21088 21304
rect 21140 21292 21146 21344
rect 22646 21332 22652 21344
rect 22607 21304 22652 21332
rect 22646 21292 22652 21304
rect 22704 21292 22710 21344
rect 24486 21332 24492 21344
rect 24447 21304 24492 21332
rect 24486 21292 24492 21304
rect 24544 21292 24550 21344
rect 24765 21335 24823 21341
rect 24765 21301 24777 21335
rect 24811 21332 24823 21335
rect 25038 21332 25044 21344
rect 24811 21304 25044 21332
rect 24811 21301 24823 21304
rect 24765 21295 24823 21301
rect 25038 21292 25044 21304
rect 25096 21292 25102 21344
rect 25884 21332 25912 21499
rect 25958 21428 25964 21480
rect 26016 21468 26022 21480
rect 26016 21440 26096 21468
rect 26016 21428 26022 21440
rect 26068 21409 26096 21440
rect 26234 21428 26240 21480
rect 26292 21468 26298 21480
rect 27062 21468 27068 21480
rect 26292 21440 27068 21468
rect 26292 21428 26298 21440
rect 27062 21428 27068 21440
rect 27120 21428 27126 21480
rect 27341 21471 27399 21477
rect 27341 21468 27353 21471
rect 27172 21440 27353 21468
rect 26053 21403 26111 21409
rect 26053 21369 26065 21403
rect 26099 21369 26111 21403
rect 26053 21363 26111 21369
rect 26697 21403 26755 21409
rect 26697 21369 26709 21403
rect 26743 21400 26755 21403
rect 27172 21400 27200 21440
rect 27341 21437 27353 21440
rect 27387 21437 27399 21471
rect 27341 21431 27399 21437
rect 26743 21372 27200 21400
rect 26743 21369 26755 21372
rect 26697 21363 26755 21369
rect 26326 21332 26332 21344
rect 25884 21304 26332 21332
rect 26326 21292 26332 21304
rect 26384 21292 26390 21344
rect 1104 21242 29532 21264
rect 1104 21190 5688 21242
rect 5740 21190 5752 21242
rect 5804 21190 5816 21242
rect 5868 21190 5880 21242
rect 5932 21190 5944 21242
rect 5996 21190 15163 21242
rect 15215 21190 15227 21242
rect 15279 21190 15291 21242
rect 15343 21190 15355 21242
rect 15407 21190 15419 21242
rect 15471 21190 24639 21242
rect 24691 21190 24703 21242
rect 24755 21190 24767 21242
rect 24819 21190 24831 21242
rect 24883 21190 24895 21242
rect 24947 21190 29532 21242
rect 1104 21168 29532 21190
rect 4062 21088 4068 21140
rect 4120 21128 4126 21140
rect 4120 21100 8524 21128
rect 4120 21088 4126 21100
rect 2777 21063 2835 21069
rect 2777 21029 2789 21063
rect 2823 21060 2835 21063
rect 3234 21060 3240 21072
rect 2823 21032 3240 21060
rect 2823 21029 2835 21032
rect 2777 21023 2835 21029
rect 3234 21020 3240 21032
rect 3292 21020 3298 21072
rect 7193 21063 7251 21069
rect 7193 21029 7205 21063
rect 7239 21060 7251 21063
rect 8294 21060 8300 21072
rect 7239 21032 8300 21060
rect 7239 21029 7251 21032
rect 7193 21023 7251 21029
rect 8294 21020 8300 21032
rect 8352 21020 8358 21072
rect 8496 21060 8524 21100
rect 8570 21088 8576 21140
rect 8628 21128 8634 21140
rect 9582 21128 9588 21140
rect 8628 21100 9588 21128
rect 8628 21088 8634 21100
rect 9582 21088 9588 21100
rect 9640 21128 9646 21140
rect 10321 21131 10379 21137
rect 10321 21128 10333 21131
rect 9640 21100 10333 21128
rect 9640 21088 9646 21100
rect 10321 21097 10333 21100
rect 10367 21097 10379 21131
rect 10321 21091 10379 21097
rect 11149 21131 11207 21137
rect 11149 21097 11161 21131
rect 11195 21128 11207 21131
rect 12434 21128 12440 21140
rect 11195 21100 12440 21128
rect 11195 21097 11207 21100
rect 11149 21091 11207 21097
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 16482 21128 16488 21140
rect 15396 21100 16488 21128
rect 8938 21060 8944 21072
rect 8496 21032 8944 21060
rect 8938 21020 8944 21032
rect 8996 21020 9002 21072
rect 9122 21060 9128 21072
rect 9083 21032 9128 21060
rect 9122 21020 9128 21032
rect 9180 21060 9186 21072
rect 9309 21063 9367 21069
rect 9309 21060 9321 21063
rect 9180 21032 9321 21060
rect 9180 21020 9186 21032
rect 9309 21029 9321 21032
rect 9355 21029 9367 21063
rect 9309 21023 9367 21029
rect 10778 21020 10784 21072
rect 10836 21060 10842 21072
rect 11241 21063 11299 21069
rect 11241 21060 11253 21063
rect 10836 21032 11253 21060
rect 10836 21020 10842 21032
rect 11241 21029 11253 21032
rect 11287 21029 11299 21063
rect 11241 21023 11299 21029
rect 3418 20952 3424 21004
rect 3476 20992 3482 21004
rect 3513 20995 3571 21001
rect 3513 20992 3525 20995
rect 3476 20964 3525 20992
rect 3476 20952 3482 20964
rect 3513 20961 3525 20964
rect 3559 20961 3571 20995
rect 5997 20995 6055 21001
rect 5997 20992 6009 20995
rect 3513 20955 3571 20961
rect 5000 20964 6009 20992
rect 1394 20924 1400 20936
rect 1355 20896 1400 20924
rect 1394 20884 1400 20896
rect 1452 20884 1458 20936
rect 3234 20924 3240 20936
rect 3195 20896 3240 20924
rect 3234 20884 3240 20896
rect 3292 20884 3298 20936
rect 3326 20884 3332 20936
rect 3384 20924 3390 20936
rect 3602 20924 3608 20936
rect 3384 20896 3429 20924
rect 3563 20896 3608 20924
rect 3384 20884 3390 20896
rect 3602 20884 3608 20896
rect 3660 20884 3666 20936
rect 3789 20927 3847 20933
rect 3789 20893 3801 20927
rect 3835 20924 3847 20927
rect 4614 20924 4620 20936
rect 3835 20896 4620 20924
rect 3835 20893 3847 20896
rect 3789 20887 3847 20893
rect 4614 20884 4620 20896
rect 4672 20884 4678 20936
rect 4062 20865 4068 20868
rect 1664 20859 1722 20865
rect 1664 20825 1676 20859
rect 1710 20856 1722 20859
rect 3053 20859 3111 20865
rect 3053 20856 3065 20859
rect 1710 20828 3065 20856
rect 1710 20825 1722 20828
rect 1664 20819 1722 20825
rect 3053 20825 3065 20828
rect 3099 20825 3111 20859
rect 4056 20856 4068 20865
rect 4023 20828 4068 20856
rect 3053 20819 3111 20825
rect 4056 20819 4068 20828
rect 4062 20816 4068 20819
rect 4120 20816 4126 20868
rect 3878 20748 3884 20800
rect 3936 20788 3942 20800
rect 5000 20788 5028 20964
rect 5997 20961 6009 20964
rect 6043 20961 6055 20995
rect 6730 20992 6736 21004
rect 5997 20955 6055 20961
rect 6380 20964 6736 20992
rect 5813 20927 5871 20933
rect 5813 20893 5825 20927
rect 5859 20924 5871 20927
rect 6380 20924 6408 20964
rect 6730 20952 6736 20964
rect 6788 20952 6794 21004
rect 7377 20995 7435 21001
rect 7377 20992 7389 20995
rect 6932 20964 7389 20992
rect 6638 20924 6644 20936
rect 5859 20896 6408 20924
rect 6551 20896 6644 20924
rect 5859 20893 5871 20896
rect 5813 20887 5871 20893
rect 6638 20884 6644 20896
rect 6696 20924 6702 20936
rect 6932 20924 6960 20964
rect 7377 20961 7389 20964
rect 7423 20961 7435 20995
rect 7377 20955 7435 20961
rect 8864 20964 10640 20992
rect 6696 20896 6960 20924
rect 7285 20927 7343 20933
rect 6696 20884 6702 20896
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 8864 20924 8892 20964
rect 7331 20896 8892 20924
rect 8941 20927 8999 20933
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 8941 20893 8953 20927
rect 8987 20924 8999 20927
rect 9122 20924 9128 20936
rect 8987 20896 9128 20924
rect 8987 20893 8999 20896
rect 8941 20887 8999 20893
rect 9122 20884 9128 20896
rect 9180 20884 9186 20936
rect 9766 20924 9772 20936
rect 9679 20896 9772 20924
rect 9766 20884 9772 20896
rect 9824 20924 9830 20936
rect 10229 20927 10287 20933
rect 9824 20896 10189 20924
rect 9824 20884 9830 20896
rect 5905 20859 5963 20865
rect 5905 20856 5917 20859
rect 5184 20828 5917 20856
rect 5184 20800 5212 20828
rect 5905 20825 5917 20828
rect 5951 20825 5963 20859
rect 5905 20819 5963 20825
rect 9398 20816 9404 20868
rect 9456 20856 9462 20868
rect 10161 20856 10189 20896
rect 10229 20893 10241 20927
rect 10275 20924 10287 20927
rect 10318 20924 10324 20936
rect 10275 20896 10324 20924
rect 10275 20893 10287 20896
rect 10229 20887 10287 20893
rect 10318 20884 10324 20896
rect 10376 20884 10382 20936
rect 10502 20884 10508 20936
rect 10560 20884 10566 20936
rect 10520 20856 10548 20884
rect 9456 20828 9904 20856
rect 10161 20828 10548 20856
rect 10612 20856 10640 20964
rect 11330 20952 11336 21004
rect 11388 20992 11394 21004
rect 12069 20995 12127 21001
rect 12069 20992 12081 20995
rect 11388 20964 12081 20992
rect 11388 20952 11394 20964
rect 12069 20961 12081 20964
rect 12115 20961 12127 20995
rect 12069 20955 12127 20961
rect 13262 20952 13268 21004
rect 13320 20992 13326 21004
rect 14826 20992 14832 21004
rect 13320 20964 14832 20992
rect 13320 20952 13326 20964
rect 14826 20952 14832 20964
rect 14884 20992 14890 21004
rect 15396 20992 15424 21100
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 19794 21088 19800 21140
rect 19852 21128 19858 21140
rect 22186 21128 22192 21140
rect 19852 21100 22192 21128
rect 19852 21088 19858 21100
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 23290 21088 23296 21140
rect 23348 21128 23354 21140
rect 23845 21131 23903 21137
rect 23845 21128 23857 21131
rect 23348 21100 23857 21128
rect 23348 21088 23354 21100
rect 23845 21097 23857 21100
rect 23891 21097 23903 21131
rect 24118 21128 24124 21140
rect 24079 21100 24124 21128
rect 23845 21091 23903 21097
rect 24118 21088 24124 21100
rect 24176 21088 24182 21140
rect 24394 21088 24400 21140
rect 24452 21128 24458 21140
rect 24452 21100 26372 21128
rect 24452 21088 24458 21100
rect 15654 21060 15660 21072
rect 15615 21032 15660 21060
rect 15654 21020 15660 21032
rect 15712 21020 15718 21072
rect 17954 21020 17960 21072
rect 18012 21060 18018 21072
rect 18322 21060 18328 21072
rect 18012 21032 18328 21060
rect 18012 21020 18018 21032
rect 18322 21020 18328 21032
rect 18380 21060 18386 21072
rect 18417 21063 18475 21069
rect 18417 21060 18429 21063
rect 18380 21032 18429 21060
rect 18380 21020 18386 21032
rect 18417 21029 18429 21032
rect 18463 21060 18475 21063
rect 19242 21060 19248 21072
rect 18463 21032 19248 21060
rect 18463 21029 18475 21032
rect 18417 21023 18475 21029
rect 19242 21020 19248 21032
rect 19300 21020 19306 21072
rect 20530 21060 20536 21072
rect 20180 21032 20392 21060
rect 20491 21032 20536 21060
rect 15838 20992 15844 21004
rect 14884 20964 15424 20992
rect 15799 20964 15844 20992
rect 14884 20952 14890 20964
rect 10689 20927 10747 20933
rect 10689 20893 10701 20927
rect 10735 20924 10747 20927
rect 10962 20924 10968 20936
rect 10735 20896 10968 20924
rect 10735 20893 10747 20896
rect 10689 20887 10747 20893
rect 10962 20884 10968 20896
rect 11020 20884 11026 20936
rect 11054 20884 11060 20936
rect 11112 20924 11118 20936
rect 11425 20927 11483 20933
rect 11425 20924 11437 20927
rect 11112 20896 11437 20924
rect 11112 20884 11118 20896
rect 11425 20893 11437 20896
rect 11471 20893 11483 20927
rect 11425 20887 11483 20893
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 12492 20896 12537 20924
rect 12492 20884 12498 20896
rect 14918 20884 14924 20936
rect 14976 20924 14982 20936
rect 15102 20924 15108 20936
rect 14976 20896 15108 20924
rect 14976 20884 14982 20896
rect 15102 20884 15108 20896
rect 15160 20884 15166 20936
rect 15396 20933 15424 20964
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 16117 20995 16175 21001
rect 16117 20961 16129 20995
rect 16163 20992 16175 20995
rect 16482 20992 16488 21004
rect 16163 20964 16488 20992
rect 16163 20961 16175 20964
rect 16117 20955 16175 20961
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 17310 20952 17316 21004
rect 17368 20992 17374 21004
rect 17678 20992 17684 21004
rect 17368 20964 17684 20992
rect 17368 20952 17374 20964
rect 17678 20952 17684 20964
rect 17736 20952 17742 21004
rect 20180 20992 20208 21032
rect 18156 20964 20208 20992
rect 20364 20992 20392 21032
rect 20530 21020 20536 21032
rect 20588 21020 20594 21072
rect 24210 21060 24216 21072
rect 23501 21032 24216 21060
rect 22002 20992 22008 21004
rect 20364 20964 22008 20992
rect 18156 20936 18184 20964
rect 22002 20952 22008 20964
rect 22060 20992 22066 21004
rect 23501 20992 23529 21032
rect 24210 21020 24216 21032
rect 24268 21020 24274 21072
rect 22060 20964 23529 20992
rect 23569 20995 23627 21001
rect 22060 20952 22066 20964
rect 23569 20961 23581 20995
rect 23615 20992 23627 20995
rect 24302 20992 24308 21004
rect 23615 20964 24308 20992
rect 23615 20961 23627 20964
rect 23569 20955 23627 20961
rect 24302 20952 24308 20964
rect 24360 20992 24366 21004
rect 26234 20992 26240 21004
rect 24360 20964 26240 20992
rect 24360 20952 24366 20964
rect 26234 20952 26240 20964
rect 26292 20952 26298 21004
rect 15381 20927 15439 20933
rect 15381 20893 15393 20927
rect 15427 20893 15439 20927
rect 15381 20887 15439 20893
rect 15525 20927 15583 20933
rect 15525 20893 15537 20927
rect 15571 20924 15583 20927
rect 15746 20924 15752 20936
rect 15571 20896 15752 20924
rect 15571 20893 15583 20896
rect 15525 20887 15583 20893
rect 15746 20884 15752 20896
rect 15804 20884 15810 20936
rect 18049 20927 18107 20933
rect 18049 20893 18061 20927
rect 18095 20924 18107 20927
rect 18138 20924 18144 20936
rect 18095 20896 18144 20924
rect 18095 20893 18107 20896
rect 18049 20887 18107 20893
rect 18138 20884 18144 20896
rect 18196 20884 18202 20936
rect 18601 20927 18659 20933
rect 18601 20893 18613 20927
rect 18647 20924 18659 20927
rect 18690 20924 18696 20936
rect 18647 20896 18696 20924
rect 18647 20893 18659 20896
rect 18601 20887 18659 20893
rect 18690 20884 18696 20896
rect 18748 20884 18754 20936
rect 18966 20924 18972 20936
rect 18927 20896 18972 20924
rect 18966 20884 18972 20896
rect 19024 20884 19030 20936
rect 19426 20924 19432 20936
rect 19387 20896 19432 20924
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 19794 20924 19800 20936
rect 19755 20896 19800 20924
rect 19794 20884 19800 20896
rect 19852 20884 19858 20936
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20924 20039 20927
rect 20070 20924 20076 20936
rect 20027 20896 20076 20924
rect 20027 20893 20039 20896
rect 19981 20887 20039 20893
rect 20070 20884 20076 20896
rect 20128 20884 20134 20936
rect 20162 20884 20168 20936
rect 20220 20924 20226 20936
rect 20220 20896 20265 20924
rect 20220 20884 20226 20896
rect 20346 20884 20352 20936
rect 20404 20933 20410 20936
rect 20404 20924 20412 20933
rect 20901 20927 20959 20933
rect 20404 20896 20449 20924
rect 20404 20887 20412 20896
rect 20901 20893 20913 20927
rect 20947 20924 20959 20927
rect 21082 20924 21088 20936
rect 20947 20896 21088 20924
rect 20947 20893 20959 20896
rect 20901 20887 20959 20893
rect 20404 20884 20410 20887
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 23658 20924 23664 20936
rect 23619 20896 23664 20924
rect 23658 20884 23664 20896
rect 23716 20884 23722 20936
rect 23937 20927 23995 20933
rect 23937 20893 23949 20927
rect 23983 20924 23995 20927
rect 24213 20927 24271 20933
rect 24213 20924 24225 20927
rect 23983 20896 24225 20924
rect 23983 20893 23995 20896
rect 23937 20887 23995 20893
rect 24213 20893 24225 20896
rect 24259 20893 24271 20927
rect 26344 20924 26372 21100
rect 26602 21088 26608 21140
rect 26660 21128 26666 21140
rect 26789 21131 26847 21137
rect 26789 21128 26801 21131
rect 26660 21100 26801 21128
rect 26660 21088 26666 21100
rect 26789 21097 26801 21100
rect 26835 21097 26847 21131
rect 27982 21128 27988 21140
rect 27943 21100 27988 21128
rect 26789 21091 26847 21097
rect 27982 21088 27988 21100
rect 28040 21088 28046 21140
rect 27525 21063 27583 21069
rect 27525 21029 27537 21063
rect 27571 21029 27583 21063
rect 27525 21023 27583 21029
rect 26418 20952 26424 21004
rect 26476 20992 26482 21004
rect 26476 20964 27384 20992
rect 26476 20952 26482 20964
rect 26510 20924 26516 20936
rect 26344 20896 26516 20924
rect 24213 20887 24271 20893
rect 26510 20884 26516 20896
rect 26568 20884 26574 20936
rect 27356 20933 27384 20964
rect 26605 20927 26663 20933
rect 26605 20893 26617 20927
rect 26651 20893 26663 20927
rect 26605 20887 26663 20893
rect 27341 20927 27399 20933
rect 27341 20893 27353 20927
rect 27387 20893 27399 20927
rect 27540 20924 27568 21023
rect 27801 20927 27859 20933
rect 27801 20924 27813 20927
rect 27540 20896 27813 20924
rect 27341 20887 27399 20893
rect 27801 20893 27813 20896
rect 27847 20893 27859 20927
rect 27801 20887 27859 20893
rect 12066 20856 12072 20868
rect 10612 20828 12072 20856
rect 9456 20816 9462 20828
rect 9876 20800 9904 20828
rect 12066 20816 12072 20828
rect 12124 20816 12130 20868
rect 12894 20816 12900 20868
rect 12952 20816 12958 20868
rect 13814 20816 13820 20868
rect 13872 20856 13878 20868
rect 13909 20859 13967 20865
rect 13909 20856 13921 20859
rect 13872 20828 13921 20856
rect 13872 20816 13878 20828
rect 13909 20825 13921 20828
rect 13955 20856 13967 20859
rect 14366 20856 14372 20868
rect 13955 20828 14372 20856
rect 13955 20825 13967 20828
rect 13909 20819 13967 20825
rect 14366 20816 14372 20828
rect 14424 20816 14430 20868
rect 15289 20859 15347 20865
rect 15289 20825 15301 20859
rect 15335 20856 15347 20859
rect 15838 20856 15844 20868
rect 15335 20828 15844 20856
rect 15335 20825 15347 20828
rect 15289 20819 15347 20825
rect 15838 20816 15844 20828
rect 15896 20856 15902 20868
rect 15896 20828 15976 20856
rect 15896 20816 15902 20828
rect 5166 20788 5172 20800
rect 3936 20760 5028 20788
rect 5127 20760 5172 20788
rect 3936 20748 3942 20760
rect 5166 20748 5172 20760
rect 5224 20748 5230 20800
rect 5445 20791 5503 20797
rect 5445 20757 5457 20791
rect 5491 20788 5503 20791
rect 5626 20788 5632 20800
rect 5491 20760 5632 20788
rect 5491 20757 5503 20760
rect 5445 20751 5503 20757
rect 5626 20748 5632 20760
rect 5684 20748 5690 20800
rect 9490 20748 9496 20800
rect 9548 20788 9554 20800
rect 9585 20791 9643 20797
rect 9585 20788 9597 20791
rect 9548 20760 9597 20788
rect 9548 20748 9554 20760
rect 9585 20757 9597 20760
rect 9631 20757 9643 20791
rect 9858 20788 9864 20800
rect 9819 20760 9864 20788
rect 9585 20751 9643 20757
rect 9858 20748 9864 20760
rect 9916 20748 9922 20800
rect 10226 20748 10232 20800
rect 10284 20788 10290 20800
rect 10505 20791 10563 20797
rect 10505 20788 10517 20791
rect 10284 20760 10517 20788
rect 10284 20748 10290 20760
rect 10505 20757 10517 20760
rect 10551 20757 10563 20791
rect 10505 20751 10563 20757
rect 12342 20748 12348 20800
rect 12400 20788 12406 20800
rect 15746 20788 15752 20800
rect 12400 20760 15752 20788
rect 12400 20748 12406 20760
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 15948 20788 15976 20828
rect 16850 20816 16856 20868
rect 16908 20816 16914 20868
rect 20257 20859 20315 20865
rect 17420 20828 20116 20856
rect 17420 20788 17448 20828
rect 15948 20760 17448 20788
rect 17494 20748 17500 20800
rect 17552 20788 17558 20800
rect 17589 20791 17647 20797
rect 17589 20788 17601 20791
rect 17552 20760 17601 20788
rect 17552 20748 17558 20760
rect 17589 20757 17601 20760
rect 17635 20757 17647 20791
rect 17862 20788 17868 20800
rect 17823 20760 17868 20788
rect 17589 20751 17647 20757
rect 17862 20748 17868 20760
rect 17920 20748 17926 20800
rect 18690 20748 18696 20800
rect 18748 20788 18754 20800
rect 18785 20791 18843 20797
rect 18785 20788 18797 20791
rect 18748 20760 18797 20788
rect 18748 20748 18754 20760
rect 18785 20757 18797 20760
rect 18831 20757 18843 20791
rect 18785 20751 18843 20757
rect 18874 20748 18880 20800
rect 18932 20788 18938 20800
rect 19245 20791 19303 20797
rect 19245 20788 19257 20791
rect 18932 20760 19257 20788
rect 18932 20748 18938 20760
rect 19245 20757 19257 20760
rect 19291 20757 19303 20791
rect 19245 20751 19303 20757
rect 19518 20748 19524 20800
rect 19576 20788 19582 20800
rect 19613 20791 19671 20797
rect 19613 20788 19625 20791
rect 19576 20760 19625 20788
rect 19576 20748 19582 20760
rect 19613 20757 19625 20760
rect 19659 20757 19671 20791
rect 20088 20788 20116 20828
rect 20257 20825 20269 20859
rect 20303 20856 20315 20859
rect 21174 20856 21180 20868
rect 20303 20828 21180 20856
rect 20303 20825 20315 20828
rect 20257 20819 20315 20825
rect 20272 20788 20300 20819
rect 21174 20816 21180 20828
rect 21232 20816 21238 20868
rect 22646 20816 22652 20868
rect 22704 20816 22710 20868
rect 23293 20859 23351 20865
rect 23293 20825 23305 20859
rect 23339 20856 23351 20859
rect 23382 20856 23388 20868
rect 23339 20828 23388 20856
rect 23339 20825 23351 20828
rect 23293 20819 23351 20825
rect 23382 20816 23388 20828
rect 23440 20816 23446 20868
rect 23676 20856 23704 20884
rect 24394 20856 24400 20868
rect 23676 20828 24400 20856
rect 24394 20816 24400 20828
rect 24452 20816 24458 20868
rect 24946 20816 24952 20868
rect 25004 20816 25010 20868
rect 25961 20859 26019 20865
rect 25961 20825 25973 20859
rect 26007 20825 26019 20859
rect 26620 20856 26648 20887
rect 25961 20819 26019 20825
rect 26436 20828 26648 20856
rect 20088 20760 20300 20788
rect 19613 20751 19671 20757
rect 20346 20748 20352 20800
rect 20404 20788 20410 20800
rect 20717 20791 20775 20797
rect 20717 20788 20729 20791
rect 20404 20760 20729 20788
rect 20404 20748 20410 20760
rect 20717 20757 20729 20760
rect 20763 20757 20775 20791
rect 20717 20751 20775 20757
rect 21821 20791 21879 20797
rect 21821 20757 21833 20791
rect 21867 20788 21879 20791
rect 22370 20788 22376 20800
rect 21867 20760 22376 20788
rect 21867 20757 21879 20760
rect 21821 20751 21879 20757
rect 22370 20748 22376 20760
rect 22428 20748 22434 20800
rect 23842 20748 23848 20800
rect 23900 20788 23906 20800
rect 24489 20791 24547 20797
rect 24489 20788 24501 20791
rect 23900 20760 24501 20788
rect 23900 20748 23906 20760
rect 24489 20757 24501 20760
rect 24535 20757 24547 20791
rect 24489 20751 24547 20757
rect 24578 20748 24584 20800
rect 24636 20788 24642 20800
rect 25976 20788 26004 20819
rect 26436 20800 26464 20828
rect 26418 20788 26424 20800
rect 24636 20760 26004 20788
rect 26379 20760 26424 20788
rect 24636 20748 24642 20760
rect 26418 20748 26424 20760
rect 26476 20748 26482 20800
rect 1104 20698 29532 20720
rect 1104 20646 10425 20698
rect 10477 20646 10489 20698
rect 10541 20646 10553 20698
rect 10605 20646 10617 20698
rect 10669 20646 10681 20698
rect 10733 20646 19901 20698
rect 19953 20646 19965 20698
rect 20017 20646 20029 20698
rect 20081 20646 20093 20698
rect 20145 20646 20157 20698
rect 20209 20646 29532 20698
rect 1104 20624 29532 20646
rect 3050 20584 3056 20596
rect 3011 20556 3056 20584
rect 3050 20544 3056 20556
rect 3108 20544 3114 20596
rect 3421 20587 3479 20593
rect 3421 20553 3433 20587
rect 3467 20584 3479 20587
rect 3602 20584 3608 20596
rect 3467 20556 3608 20584
rect 3467 20553 3479 20556
rect 3421 20547 3479 20553
rect 3602 20544 3608 20556
rect 3660 20544 3666 20596
rect 4062 20584 4068 20596
rect 4023 20556 4068 20584
rect 4062 20544 4068 20556
rect 4120 20544 4126 20596
rect 7009 20587 7067 20593
rect 7009 20553 7021 20587
rect 7055 20584 7067 20587
rect 9398 20584 9404 20596
rect 7055 20556 9404 20584
rect 7055 20553 7067 20556
rect 7009 20547 7067 20553
rect 3326 20476 3332 20528
rect 3384 20516 3390 20528
rect 5258 20516 5264 20528
rect 3384 20488 5264 20516
rect 3384 20476 3390 20488
rect 3510 20448 3516 20460
rect 3471 20420 3516 20448
rect 3510 20408 3516 20420
rect 3568 20408 3574 20460
rect 3804 20457 3832 20488
rect 5258 20476 5264 20488
rect 5316 20476 5322 20528
rect 5353 20519 5411 20525
rect 5353 20485 5365 20519
rect 5399 20516 5411 20519
rect 5534 20516 5540 20528
rect 5399 20488 5540 20516
rect 5399 20485 5411 20488
rect 5353 20479 5411 20485
rect 5534 20476 5540 20488
rect 5592 20516 5598 20528
rect 6549 20519 6607 20525
rect 6549 20516 6561 20519
rect 5592 20488 6561 20516
rect 5592 20476 5598 20488
rect 6549 20485 6561 20488
rect 6595 20485 6607 20519
rect 6549 20479 6607 20485
rect 6733 20519 6791 20525
rect 6733 20485 6745 20519
rect 6779 20516 6791 20519
rect 7024 20516 7052 20547
rect 9398 20544 9404 20556
rect 9456 20544 9462 20596
rect 10134 20544 10140 20596
rect 10192 20584 10198 20596
rect 11054 20584 11060 20596
rect 10192 20556 11060 20584
rect 10192 20544 10198 20556
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 12434 20544 12440 20596
rect 12492 20584 12498 20596
rect 12805 20587 12863 20593
rect 12805 20584 12817 20587
rect 12492 20556 12817 20584
rect 12492 20544 12498 20556
rect 12805 20553 12817 20556
rect 12851 20553 12863 20587
rect 12805 20547 12863 20553
rect 15010 20544 15016 20596
rect 15068 20584 15074 20596
rect 15105 20587 15163 20593
rect 15105 20584 15117 20587
rect 15068 20556 15117 20584
rect 15068 20544 15074 20556
rect 15105 20553 15117 20556
rect 15151 20553 15163 20587
rect 15105 20547 15163 20553
rect 17037 20587 17095 20593
rect 17037 20553 17049 20587
rect 17083 20584 17095 20587
rect 17126 20584 17132 20596
rect 17083 20556 17132 20584
rect 17083 20553 17095 20556
rect 17037 20547 17095 20553
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 17770 20544 17776 20596
rect 17828 20584 17834 20596
rect 19794 20584 19800 20596
rect 17828 20556 19661 20584
rect 19707 20556 19800 20584
rect 17828 20544 17834 20556
rect 10778 20516 10784 20528
rect 6779 20488 7052 20516
rect 10626 20488 10784 20516
rect 6779 20485 6791 20488
rect 6733 20479 6791 20485
rect 10778 20476 10784 20488
rect 10836 20476 10842 20528
rect 13538 20476 13544 20528
rect 13596 20516 13602 20528
rect 14829 20519 14887 20525
rect 14829 20516 14841 20519
rect 13596 20488 14841 20516
rect 13596 20476 13602 20488
rect 14829 20485 14841 20488
rect 14875 20485 14887 20519
rect 15933 20519 15991 20525
rect 15933 20516 15945 20519
rect 14829 20479 14887 20485
rect 15764 20488 15945 20516
rect 15764 20460 15792 20488
rect 15933 20485 15945 20488
rect 15979 20516 15991 20519
rect 16393 20519 16451 20525
rect 16393 20516 16405 20519
rect 15979 20488 16405 20516
rect 15979 20485 15991 20488
rect 15933 20479 15991 20485
rect 16393 20485 16405 20488
rect 16439 20516 16451 20519
rect 17494 20516 17500 20528
rect 16439 20488 17500 20516
rect 16439 20485 16451 20488
rect 16393 20479 16451 20485
rect 17494 20476 17500 20488
rect 17552 20476 17558 20528
rect 18690 20476 18696 20528
rect 18748 20476 18754 20528
rect 19242 20476 19248 20528
rect 19300 20516 19306 20528
rect 19633 20516 19661 20556
rect 19794 20544 19800 20556
rect 19852 20584 19858 20596
rect 20254 20584 20260 20596
rect 19852 20556 20260 20584
rect 19852 20544 19858 20556
rect 20254 20544 20260 20556
rect 20312 20544 20318 20596
rect 22002 20584 22008 20596
rect 21963 20556 22008 20584
rect 22002 20544 22008 20556
rect 22060 20544 22066 20596
rect 22649 20587 22707 20593
rect 22649 20553 22661 20587
rect 22695 20584 22707 20587
rect 22830 20584 22836 20596
rect 22695 20556 22836 20584
rect 22695 20553 22707 20556
rect 22649 20547 22707 20553
rect 22830 20544 22836 20556
rect 22888 20544 22894 20596
rect 23474 20584 23480 20596
rect 23032 20556 23480 20584
rect 20432 20519 20490 20525
rect 19300 20488 19472 20516
rect 19633 20488 19748 20516
rect 19300 20476 19306 20488
rect 3789 20451 3847 20457
rect 3789 20417 3801 20451
rect 3835 20417 3847 20451
rect 3789 20411 3847 20417
rect 3881 20451 3939 20457
rect 3881 20417 3893 20451
rect 3927 20448 3939 20451
rect 5166 20448 5172 20460
rect 3927 20420 5172 20448
rect 3927 20417 3939 20420
rect 3881 20411 3939 20417
rect 5166 20408 5172 20420
rect 5224 20408 5230 20460
rect 7282 20448 7288 20460
rect 7243 20420 7288 20448
rect 7282 20408 7288 20420
rect 7340 20408 7346 20460
rect 7742 20448 7748 20460
rect 7703 20420 7748 20448
rect 7742 20408 7748 20420
rect 7800 20408 7806 20460
rect 8941 20451 8999 20457
rect 8941 20417 8953 20451
rect 8987 20448 8999 20451
rect 9122 20448 9128 20460
rect 8987 20420 9128 20448
rect 8987 20417 8999 20420
rect 8941 20411 8999 20417
rect 9122 20408 9128 20420
rect 9180 20448 9186 20460
rect 9217 20451 9275 20457
rect 9217 20448 9229 20451
rect 9180 20420 9229 20448
rect 9180 20408 9186 20420
rect 9217 20417 9229 20420
rect 9263 20417 9275 20451
rect 9217 20411 9275 20417
rect 11885 20451 11943 20457
rect 11885 20417 11897 20451
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 2777 20383 2835 20389
rect 2777 20349 2789 20383
rect 2823 20349 2835 20383
rect 2958 20380 2964 20392
rect 2919 20352 2964 20380
rect 2777 20343 2835 20349
rect 2792 20312 2820 20343
rect 2958 20340 2964 20352
rect 3016 20340 3022 20392
rect 9766 20380 9772 20392
rect 9646 20352 9772 20380
rect 3142 20312 3148 20324
rect 2792 20284 3148 20312
rect 3142 20272 3148 20284
rect 3200 20312 3206 20324
rect 3878 20312 3884 20324
rect 3200 20284 3884 20312
rect 3200 20272 3206 20284
rect 3878 20272 3884 20284
rect 3936 20272 3942 20324
rect 4614 20272 4620 20324
rect 4672 20312 4678 20324
rect 5169 20315 5227 20321
rect 5169 20312 5181 20315
rect 4672 20284 5181 20312
rect 4672 20272 4678 20284
rect 5169 20281 5181 20284
rect 5215 20281 5227 20315
rect 5169 20275 5227 20281
rect 7469 20315 7527 20321
rect 7469 20281 7481 20315
rect 7515 20312 7527 20315
rect 8754 20312 8760 20324
rect 7515 20284 8760 20312
rect 7515 20281 7527 20284
rect 7469 20275 7527 20281
rect 8754 20272 8760 20284
rect 8812 20272 8818 20324
rect 9125 20315 9183 20321
rect 9125 20281 9137 20315
rect 9171 20312 9183 20315
rect 9646 20312 9674 20352
rect 9766 20340 9772 20352
rect 9824 20340 9830 20392
rect 11054 20380 11060 20392
rect 11015 20352 11060 20380
rect 11054 20340 11060 20352
rect 11112 20340 11118 20392
rect 11330 20380 11336 20392
rect 11291 20352 11336 20380
rect 11330 20340 11336 20352
rect 11388 20340 11394 20392
rect 9171 20284 9674 20312
rect 9171 20281 9183 20284
rect 9125 20275 9183 20281
rect 3510 20204 3516 20256
rect 3568 20244 3574 20256
rect 3605 20247 3663 20253
rect 3605 20244 3617 20247
rect 3568 20216 3617 20244
rect 3568 20204 3574 20216
rect 3605 20213 3617 20216
rect 3651 20213 3663 20247
rect 7558 20244 7564 20256
rect 7519 20216 7564 20244
rect 3605 20207 3663 20213
rect 7558 20204 7564 20216
rect 7616 20204 7622 20256
rect 9401 20247 9459 20253
rect 9401 20213 9413 20247
rect 9447 20244 9459 20247
rect 9490 20244 9496 20256
rect 9447 20216 9496 20244
rect 9447 20213 9459 20216
rect 9401 20207 9459 20213
rect 9490 20204 9496 20216
rect 9548 20204 9554 20256
rect 9585 20247 9643 20253
rect 9585 20213 9597 20247
rect 9631 20244 9643 20247
rect 11900 20244 11928 20411
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 12492 20420 12537 20448
rect 12492 20408 12498 20420
rect 12894 20408 12900 20460
rect 12952 20448 12958 20460
rect 12989 20451 13047 20457
rect 12989 20448 13001 20451
rect 12952 20420 13001 20448
rect 12952 20408 12958 20420
rect 12989 20417 13001 20420
rect 13035 20417 13047 20451
rect 14093 20451 14151 20457
rect 14093 20448 14105 20451
rect 12989 20411 13047 20417
rect 13648 20420 14105 20448
rect 12250 20380 12256 20392
rect 12211 20352 12256 20380
rect 12250 20340 12256 20352
rect 12308 20340 12314 20392
rect 12452 20380 12480 20408
rect 13648 20380 13676 20420
rect 14093 20417 14105 20420
rect 14139 20448 14151 20451
rect 14645 20451 14703 20457
rect 14645 20448 14657 20451
rect 14139 20420 14657 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 14645 20417 14657 20420
rect 14691 20448 14703 20451
rect 14734 20448 14740 20460
rect 14691 20420 14740 20448
rect 14691 20417 14703 20420
rect 14645 20411 14703 20417
rect 14734 20408 14740 20420
rect 14792 20408 14798 20460
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 15289 20451 15347 20457
rect 15289 20448 15301 20451
rect 14976 20420 15301 20448
rect 14976 20408 14982 20420
rect 15289 20417 15301 20420
rect 15335 20417 15347 20451
rect 15289 20411 15347 20417
rect 15657 20451 15715 20457
rect 15657 20417 15669 20451
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 12452 20352 13676 20380
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 14185 20383 14243 20389
rect 14185 20380 14197 20383
rect 13872 20352 14197 20380
rect 13872 20340 13878 20352
rect 14185 20349 14197 20352
rect 14231 20349 14243 20383
rect 15010 20380 15016 20392
rect 14971 20352 15016 20380
rect 14185 20343 14243 20349
rect 15010 20340 15016 20352
rect 15068 20340 15074 20392
rect 15672 20380 15700 20411
rect 15746 20408 15752 20460
rect 15804 20408 15810 20460
rect 15841 20451 15899 20457
rect 15841 20444 15853 20451
rect 15887 20444 15899 20451
rect 16022 20448 16028 20460
rect 16080 20457 16086 20460
rect 15838 20392 15844 20444
rect 15896 20392 15902 20444
rect 15988 20420 16028 20448
rect 16022 20408 16028 20420
rect 16080 20411 16088 20457
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20448 17279 20451
rect 17402 20448 17408 20460
rect 17267 20420 17408 20448
rect 17267 20417 17279 20420
rect 17221 20411 17279 20417
rect 16080 20408 16086 20411
rect 17402 20408 17408 20420
rect 17460 20448 17466 20460
rect 17862 20448 17868 20460
rect 17460 20420 17868 20448
rect 17460 20408 17466 20420
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 19444 20457 19472 20488
rect 19429 20451 19487 20457
rect 19429 20417 19441 20451
rect 19475 20417 19487 20451
rect 19429 20411 19487 20417
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20448 19579 20451
rect 19613 20451 19671 20457
rect 19613 20448 19625 20451
rect 19567 20420 19625 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 19613 20417 19625 20420
rect 19659 20417 19671 20451
rect 19720 20448 19748 20488
rect 20432 20485 20444 20519
rect 20478 20516 20490 20519
rect 20530 20516 20536 20528
rect 20478 20488 20536 20516
rect 20478 20485 20490 20488
rect 20432 20479 20490 20485
rect 20530 20476 20536 20488
rect 20588 20476 20594 20528
rect 23032 20516 23060 20556
rect 23474 20544 23480 20556
rect 23532 20584 23538 20596
rect 24486 20584 24492 20596
rect 23532 20556 24492 20584
rect 23532 20544 23538 20556
rect 24486 20544 24492 20556
rect 24544 20544 24550 20596
rect 24946 20544 24952 20596
rect 25004 20584 25010 20596
rect 25041 20587 25099 20593
rect 25041 20584 25053 20587
rect 25004 20556 25053 20584
rect 25004 20544 25010 20556
rect 25041 20553 25053 20556
rect 25087 20553 25099 20587
rect 25041 20547 25099 20553
rect 26697 20587 26755 20593
rect 26697 20553 26709 20587
rect 26743 20584 26755 20587
rect 27246 20584 27252 20596
rect 26743 20556 27252 20584
rect 26743 20553 26755 20556
rect 26697 20547 26755 20553
rect 27246 20544 27252 20556
rect 27304 20544 27310 20596
rect 22480 20488 23060 20516
rect 22186 20448 22192 20460
rect 19720 20420 21220 20448
rect 22147 20420 22192 20448
rect 19613 20411 19671 20417
rect 19150 20380 19156 20392
rect 15672 20352 15792 20380
rect 19111 20352 19156 20380
rect 15764 20324 15792 20352
rect 19150 20340 19156 20352
rect 19208 20340 19214 20392
rect 19444 20380 19472 20411
rect 20165 20383 20223 20389
rect 20165 20380 20177 20383
rect 19444 20352 20177 20380
rect 20165 20349 20177 20352
rect 20211 20349 20223 20383
rect 21192 20380 21220 20420
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 22480 20457 22508 20488
rect 23106 20476 23112 20528
rect 23164 20516 23170 20528
rect 23164 20488 23209 20516
rect 23308 20488 24072 20516
rect 23164 20476 23170 20488
rect 23308 20460 23336 20488
rect 22465 20451 22523 20457
rect 22465 20417 22477 20451
rect 22511 20417 22523 20451
rect 22465 20411 22523 20417
rect 22833 20451 22891 20457
rect 22833 20417 22845 20451
rect 22879 20417 22891 20451
rect 22833 20411 22891 20417
rect 22554 20380 22560 20392
rect 21192 20352 22560 20380
rect 20165 20343 20223 20349
rect 22554 20340 22560 20352
rect 22612 20340 22618 20392
rect 11977 20315 12035 20321
rect 11977 20281 11989 20315
rect 12023 20312 12035 20315
rect 12342 20312 12348 20324
rect 12023 20284 12348 20312
rect 12023 20281 12035 20284
rect 11977 20275 12035 20281
rect 12342 20272 12348 20284
rect 12400 20312 12406 20324
rect 12400 20284 14136 20312
rect 12400 20272 12406 20284
rect 12526 20244 12532 20256
rect 9631 20216 12532 20244
rect 9631 20213 9643 20216
rect 9585 20207 9643 20213
rect 12526 20204 12532 20216
rect 12584 20204 12590 20256
rect 12621 20247 12679 20253
rect 12621 20213 12633 20247
rect 12667 20244 12679 20247
rect 12710 20244 12716 20256
rect 12667 20216 12716 20244
rect 12667 20213 12679 20216
rect 12621 20207 12679 20213
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 14108 20253 14136 20284
rect 15746 20272 15752 20324
rect 15804 20272 15810 20324
rect 16209 20315 16267 20321
rect 16209 20281 16221 20315
rect 16255 20312 16267 20315
rect 16482 20312 16488 20324
rect 16255 20284 16488 20312
rect 16255 20281 16267 20284
rect 16209 20275 16267 20281
rect 16482 20272 16488 20284
rect 16540 20272 16546 20324
rect 17604 20284 18000 20312
rect 14093 20247 14151 20253
rect 14093 20213 14105 20247
rect 14139 20213 14151 20247
rect 14093 20207 14151 20213
rect 14461 20247 14519 20253
rect 14461 20213 14473 20247
rect 14507 20244 14519 20247
rect 17604 20244 17632 20284
rect 14507 20216 17632 20244
rect 14507 20213 14519 20216
rect 14461 20207 14519 20213
rect 17678 20204 17684 20256
rect 17736 20244 17742 20256
rect 17972 20244 18000 20284
rect 19426 20272 19432 20324
rect 19484 20312 19490 20324
rect 19521 20315 19579 20321
rect 19521 20312 19533 20315
rect 19484 20284 19533 20312
rect 19484 20272 19490 20284
rect 19521 20281 19533 20284
rect 19567 20281 19579 20315
rect 22848 20312 22876 20411
rect 23014 20408 23020 20460
rect 23072 20448 23078 20460
rect 23290 20457 23296 20460
rect 23253 20451 23296 20457
rect 23072 20420 23117 20448
rect 23072 20408 23078 20420
rect 23253 20417 23265 20451
rect 23253 20411 23296 20417
rect 23290 20408 23296 20411
rect 23348 20408 23354 20460
rect 23569 20451 23627 20457
rect 23569 20417 23581 20451
rect 23615 20417 23627 20451
rect 23750 20448 23756 20460
rect 23711 20420 23756 20448
rect 23569 20411 23627 20417
rect 23584 20380 23612 20411
rect 23750 20408 23756 20420
rect 23808 20408 23814 20460
rect 23842 20408 23848 20460
rect 23900 20448 23906 20460
rect 24044 20457 24072 20488
rect 26786 20476 26792 20528
rect 26844 20516 26850 20528
rect 27157 20519 27215 20525
rect 27157 20516 27169 20519
rect 26844 20488 27169 20516
rect 26844 20476 26850 20488
rect 27157 20485 27169 20488
rect 27203 20485 27215 20519
rect 27709 20519 27767 20525
rect 27709 20516 27721 20519
rect 27157 20479 27215 20485
rect 27264 20488 27721 20516
rect 23989 20451 24072 20457
rect 23900 20420 23945 20448
rect 23900 20408 23906 20420
rect 23989 20417 24001 20451
rect 24035 20420 24072 20451
rect 24857 20451 24915 20457
rect 24035 20417 24047 20420
rect 23989 20411 24047 20417
rect 24857 20417 24869 20451
rect 24903 20448 24915 20451
rect 25038 20448 25044 20460
rect 24903 20420 25044 20448
rect 24903 20417 24915 20420
rect 24857 20411 24915 20417
rect 25038 20408 25044 20420
rect 25096 20408 25102 20460
rect 25590 20408 25596 20460
rect 25648 20408 25654 20460
rect 25961 20451 26019 20457
rect 25961 20417 25973 20451
rect 26007 20448 26019 20451
rect 26418 20448 26424 20460
rect 26007 20420 26424 20448
rect 26007 20417 26019 20420
rect 25961 20411 26019 20417
rect 26418 20408 26424 20420
rect 26476 20408 26482 20460
rect 26510 20408 26516 20460
rect 26568 20448 26574 20460
rect 26973 20451 27031 20457
rect 26568 20420 26613 20448
rect 26568 20408 26574 20420
rect 26973 20417 26985 20451
rect 27019 20417 27031 20451
rect 26973 20411 27031 20417
rect 22986 20352 24716 20380
rect 22986 20312 23014 20352
rect 23216 20324 23244 20352
rect 22848 20284 23014 20312
rect 19521 20275 19579 20281
rect 23198 20272 23204 20324
rect 23256 20272 23262 20324
rect 23382 20312 23388 20324
rect 23343 20284 23388 20312
rect 23382 20272 23388 20284
rect 23440 20272 23446 20324
rect 24121 20315 24179 20321
rect 24121 20281 24133 20315
rect 24167 20312 24179 20315
rect 24578 20312 24584 20324
rect 24167 20284 24584 20312
rect 24167 20281 24179 20284
rect 24121 20275 24179 20281
rect 24578 20272 24584 20284
rect 24636 20272 24642 20324
rect 21358 20244 21364 20256
rect 17736 20216 17781 20244
rect 17972 20216 21364 20244
rect 17736 20204 17742 20216
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 21450 20204 21456 20256
rect 21508 20244 21514 20256
rect 21545 20247 21603 20253
rect 21545 20244 21557 20247
rect 21508 20216 21557 20244
rect 21508 20204 21514 20216
rect 21545 20213 21557 20216
rect 21591 20213 21603 20247
rect 22370 20244 22376 20256
rect 22283 20216 22376 20244
rect 21545 20207 21603 20213
rect 22370 20204 22376 20216
rect 22428 20244 22434 20256
rect 23106 20244 23112 20256
rect 22428 20216 23112 20244
rect 22428 20204 22434 20216
rect 23106 20204 23112 20216
rect 23164 20204 23170 20256
rect 23842 20204 23848 20256
rect 23900 20244 23906 20256
rect 24305 20247 24363 20253
rect 24305 20244 24317 20247
rect 23900 20216 24317 20244
rect 23900 20204 23906 20216
rect 24305 20213 24317 20216
rect 24351 20213 24363 20247
rect 24688 20244 24716 20352
rect 25314 20340 25320 20392
rect 25372 20380 25378 20392
rect 25608 20380 25636 20408
rect 26988 20380 27016 20411
rect 27062 20408 27068 20460
rect 27120 20448 27126 20460
rect 27264 20457 27292 20488
rect 27709 20485 27721 20488
rect 27755 20485 27767 20519
rect 27709 20479 27767 20485
rect 27249 20451 27307 20457
rect 27249 20448 27261 20451
rect 27120 20420 27261 20448
rect 27120 20408 27126 20420
rect 27249 20417 27261 20420
rect 27295 20417 27307 20451
rect 27249 20411 27307 20417
rect 27346 20451 27404 20457
rect 27346 20417 27358 20451
rect 27392 20417 27404 20451
rect 27346 20411 27404 20417
rect 25372 20352 27016 20380
rect 25372 20340 25378 20352
rect 25590 20272 25596 20324
rect 25648 20312 25654 20324
rect 26050 20312 26056 20324
rect 25648 20284 26056 20312
rect 25648 20272 25654 20284
rect 26050 20272 26056 20284
rect 26108 20312 26114 20324
rect 27356 20312 27384 20411
rect 26108 20284 27384 20312
rect 26108 20272 26114 20284
rect 25777 20247 25835 20253
rect 25777 20244 25789 20247
rect 24688 20216 25789 20244
rect 24305 20207 24363 20213
rect 25777 20213 25789 20216
rect 25823 20213 25835 20247
rect 25777 20207 25835 20213
rect 26878 20204 26884 20256
rect 26936 20244 26942 20256
rect 27525 20247 27583 20253
rect 27525 20244 27537 20247
rect 26936 20216 27537 20244
rect 26936 20204 26942 20216
rect 27525 20213 27537 20216
rect 27571 20213 27583 20247
rect 27525 20207 27583 20213
rect 1104 20154 29532 20176
rect 1104 20102 5688 20154
rect 5740 20102 5752 20154
rect 5804 20102 5816 20154
rect 5868 20102 5880 20154
rect 5932 20102 5944 20154
rect 5996 20102 15163 20154
rect 15215 20102 15227 20154
rect 15279 20102 15291 20154
rect 15343 20102 15355 20154
rect 15407 20102 15419 20154
rect 15471 20102 24639 20154
rect 24691 20102 24703 20154
rect 24755 20102 24767 20154
rect 24819 20102 24831 20154
rect 24883 20102 24895 20154
rect 24947 20102 29532 20154
rect 1104 20080 29532 20102
rect 6546 20000 6552 20052
rect 6604 20040 6610 20052
rect 6733 20043 6791 20049
rect 6733 20040 6745 20043
rect 6604 20012 6745 20040
rect 6604 20000 6610 20012
rect 6733 20009 6745 20012
rect 6779 20009 6791 20043
rect 6733 20003 6791 20009
rect 9766 20000 9772 20052
rect 9824 20040 9830 20052
rect 10962 20040 10968 20052
rect 9824 20012 10968 20040
rect 9824 20000 9830 20012
rect 10962 20000 10968 20012
rect 11020 20000 11026 20052
rect 13722 20040 13728 20052
rect 13683 20012 13728 20040
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 16022 20000 16028 20052
rect 16080 20040 16086 20052
rect 16117 20043 16175 20049
rect 16117 20040 16129 20043
rect 16080 20012 16129 20040
rect 16080 20000 16086 20012
rect 16117 20009 16129 20012
rect 16163 20009 16175 20043
rect 17678 20040 17684 20052
rect 17639 20012 17684 20040
rect 16117 20003 16175 20009
rect 17678 20000 17684 20012
rect 17736 20000 17742 20052
rect 18325 20043 18383 20049
rect 18325 20009 18337 20043
rect 18371 20040 18383 20043
rect 19150 20040 19156 20052
rect 18371 20012 19156 20040
rect 18371 20009 18383 20012
rect 18325 20003 18383 20009
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 19242 20000 19248 20052
rect 19300 20040 19306 20052
rect 19300 20012 20852 20040
rect 19300 20000 19306 20012
rect 11054 19932 11060 19984
rect 11112 19972 11118 19984
rect 15105 19975 15163 19981
rect 11112 19944 12664 19972
rect 11112 19932 11118 19944
rect 8202 19904 8208 19916
rect 8163 19876 8208 19904
rect 8202 19864 8208 19876
rect 8260 19864 8266 19916
rect 8481 19907 8539 19913
rect 8481 19873 8493 19907
rect 8527 19904 8539 19907
rect 8570 19904 8576 19916
rect 8527 19876 8576 19904
rect 8527 19873 8539 19876
rect 8481 19867 8539 19873
rect 8570 19864 8576 19876
rect 8628 19904 8634 19916
rect 8938 19904 8944 19916
rect 8628 19876 8944 19904
rect 8628 19864 8634 19876
rect 8938 19864 8944 19876
rect 8996 19904 9002 19916
rect 10781 19907 10839 19913
rect 10781 19904 10793 19907
rect 8996 19876 10793 19904
rect 8996 19864 9002 19876
rect 10781 19873 10793 19876
rect 10827 19904 10839 19907
rect 11330 19904 11336 19916
rect 10827 19876 11336 19904
rect 10827 19873 10839 19876
rect 10781 19867 10839 19873
rect 11330 19864 11336 19876
rect 11388 19864 11394 19916
rect 12636 19913 12664 19944
rect 15105 19941 15117 19975
rect 15151 19941 15163 19975
rect 15105 19935 15163 19941
rect 12621 19907 12679 19913
rect 12621 19873 12633 19907
rect 12667 19873 12679 19907
rect 13538 19904 13544 19916
rect 12621 19867 12679 19873
rect 13004 19876 13544 19904
rect 13004 19848 13032 19876
rect 13538 19864 13544 19876
rect 13596 19904 13602 19916
rect 14185 19907 14243 19913
rect 14185 19904 14197 19907
rect 13596 19876 14197 19904
rect 13596 19864 13602 19876
rect 14185 19873 14197 19876
rect 14231 19873 14243 19907
rect 15120 19904 15148 19935
rect 15746 19904 15752 19916
rect 15120 19876 15752 19904
rect 14185 19867 14243 19873
rect 15746 19864 15752 19876
rect 15804 19904 15810 19916
rect 17696 19904 17724 20000
rect 20254 19932 20260 19984
rect 20312 19972 20318 19984
rect 20441 19975 20499 19981
rect 20441 19972 20453 19975
rect 20312 19944 20453 19972
rect 20312 19932 20318 19944
rect 20441 19941 20453 19944
rect 20487 19941 20499 19975
rect 20441 19935 20499 19941
rect 17862 19904 17868 19916
rect 15804 19876 16712 19904
rect 17696 19876 17868 19904
rect 15804 19864 15810 19876
rect 16684 19848 16712 19876
rect 17862 19864 17868 19876
rect 17920 19904 17926 19916
rect 20714 19904 20720 19916
rect 17920 19876 18092 19904
rect 17920 19864 17926 19876
rect 4614 19836 4620 19848
rect 4575 19808 4620 19836
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 8754 19836 8760 19848
rect 8715 19808 8760 19836
rect 8754 19796 8760 19808
rect 8812 19796 8818 19848
rect 12342 19836 12348 19848
rect 12303 19808 12348 19836
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19805 12587 19839
rect 12529 19799 12587 19805
rect 4884 19771 4942 19777
rect 4884 19737 4896 19771
rect 4930 19768 4942 19771
rect 4982 19768 4988 19780
rect 4930 19740 4988 19768
rect 4930 19737 4942 19740
rect 4884 19731 4942 19737
rect 4982 19728 4988 19740
rect 5040 19728 5046 19780
rect 5994 19700 6000 19712
rect 5955 19672 6000 19700
rect 5994 19660 6000 19672
rect 6052 19660 6058 19712
rect 7760 19700 7788 19754
rect 10042 19728 10048 19780
rect 10100 19728 10106 19780
rect 10505 19771 10563 19777
rect 10505 19737 10517 19771
rect 10551 19768 10563 19771
rect 11698 19768 11704 19780
rect 10551 19740 11704 19768
rect 10551 19737 10563 19740
rect 10505 19731 10563 19737
rect 11698 19728 11704 19740
rect 11756 19728 11762 19780
rect 12544 19768 12572 19799
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 12805 19839 12863 19845
rect 12805 19836 12817 19839
rect 12768 19808 12817 19836
rect 12768 19796 12774 19808
rect 12805 19805 12817 19808
rect 12851 19805 12863 19839
rect 12986 19836 12992 19848
rect 12947 19808 12992 19836
rect 12805 19799 12863 19805
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 14093 19839 14151 19845
rect 14093 19836 14105 19839
rect 13832 19808 14105 19836
rect 13832 19780 13860 19808
rect 14093 19805 14105 19808
rect 14139 19805 14151 19839
rect 14918 19836 14924 19848
rect 14879 19808 14924 19836
rect 14093 19799 14151 19805
rect 14918 19796 14924 19808
rect 14976 19796 14982 19848
rect 15010 19796 15016 19848
rect 15068 19836 15074 19848
rect 15197 19839 15255 19845
rect 15197 19836 15209 19839
rect 15068 19808 15209 19836
rect 15068 19796 15074 19808
rect 15197 19805 15209 19808
rect 15243 19805 15255 19839
rect 15470 19836 15476 19848
rect 15431 19808 15476 19836
rect 15197 19799 15255 19805
rect 12406 19740 12572 19768
rect 8573 19703 8631 19709
rect 8573 19700 8585 19703
rect 7760 19672 8585 19700
rect 8573 19669 8585 19672
rect 8619 19669 8631 19703
rect 8573 19663 8631 19669
rect 9033 19703 9091 19709
rect 9033 19669 9045 19703
rect 9079 19700 9091 19703
rect 10778 19700 10784 19712
rect 9079 19672 10784 19700
rect 9079 19669 9091 19672
rect 9033 19663 9091 19669
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 11054 19660 11060 19712
rect 11112 19700 11118 19712
rect 11882 19700 11888 19712
rect 11112 19672 11888 19700
rect 11112 19660 11118 19672
rect 11882 19660 11888 19672
rect 11940 19700 11946 19712
rect 12406 19700 12434 19740
rect 12618 19728 12624 19780
rect 12676 19768 12682 19780
rect 13449 19771 13507 19777
rect 13449 19768 13461 19771
rect 12676 19740 13461 19768
rect 12676 19728 12682 19740
rect 13449 19737 13461 19740
rect 13495 19737 13507 19771
rect 13449 19731 13507 19737
rect 13633 19771 13691 19777
rect 13633 19737 13645 19771
rect 13679 19768 13691 19771
rect 13814 19768 13820 19780
rect 13679 19740 13820 19768
rect 13679 19737 13691 19740
rect 13633 19731 13691 19737
rect 13814 19728 13820 19740
rect 13872 19728 13878 19780
rect 11940 19672 12434 19700
rect 15212 19700 15240 19799
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 15562 19796 15568 19848
rect 15620 19845 15626 19848
rect 15620 19836 15628 19845
rect 15620 19808 15665 19836
rect 15620 19799 15628 19808
rect 15620 19796 15626 19799
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 15896 19808 15945 19836
rect 15896 19796 15902 19808
rect 15933 19805 15945 19808
rect 15979 19836 15991 19839
rect 16206 19836 16212 19848
rect 15979 19808 16212 19836
rect 15979 19805 15991 19808
rect 15933 19799 15991 19805
rect 16206 19796 16212 19808
rect 16264 19796 16270 19848
rect 16666 19796 16672 19848
rect 16724 19836 16730 19848
rect 18064 19845 18092 19876
rect 20088 19876 20720 19904
rect 17773 19839 17831 19845
rect 17773 19836 17785 19839
rect 16724 19808 17785 19836
rect 16724 19796 16730 19808
rect 17773 19805 17785 19808
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 18050 19839 18108 19845
rect 18050 19805 18062 19839
rect 18096 19805 18108 19839
rect 18050 19799 18108 19805
rect 15381 19771 15439 19777
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 16850 19768 16856 19780
rect 15427 19740 16856 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 16850 19728 16856 19740
rect 16908 19728 16914 19780
rect 15562 19700 15568 19712
rect 15212 19672 15568 19700
rect 11940 19660 11946 19672
rect 15562 19660 15568 19672
rect 15620 19660 15626 19712
rect 15746 19700 15752 19712
rect 15804 19709 15810 19712
rect 15715 19672 15752 19700
rect 15746 19660 15752 19672
rect 15804 19663 15815 19709
rect 16577 19703 16635 19709
rect 16577 19669 16589 19703
rect 16623 19700 16635 19703
rect 17126 19700 17132 19712
rect 16623 19672 17132 19700
rect 16623 19669 16635 19672
rect 16577 19663 16635 19669
rect 15804 19660 15810 19663
rect 17126 19660 17132 19672
rect 17184 19660 17190 19712
rect 17788 19700 17816 19799
rect 18138 19796 18144 19848
rect 18196 19845 18202 19848
rect 18196 19836 18204 19845
rect 18782 19836 18788 19848
rect 18196 19808 18241 19836
rect 18524 19808 18788 19836
rect 18196 19799 18204 19808
rect 18196 19796 18202 19799
rect 17954 19728 17960 19780
rect 18012 19768 18018 19780
rect 18012 19740 18057 19768
rect 18012 19728 18018 19740
rect 18524 19700 18552 19808
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 19794 19796 19800 19848
rect 19852 19836 19858 19848
rect 19889 19839 19947 19845
rect 19889 19836 19901 19839
rect 19852 19808 19901 19836
rect 19852 19796 19858 19808
rect 19889 19805 19901 19808
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 18598 19728 18604 19780
rect 18656 19768 18662 19780
rect 20088 19777 20116 19876
rect 20714 19864 20720 19876
rect 20772 19864 20778 19916
rect 20824 19904 20852 20012
rect 21174 20000 21180 20052
rect 21232 20040 21238 20052
rect 21269 20043 21327 20049
rect 21269 20040 21281 20043
rect 21232 20012 21281 20040
rect 21232 20000 21238 20012
rect 21269 20009 21281 20012
rect 21315 20040 21327 20043
rect 23014 20040 23020 20052
rect 21315 20012 23020 20040
rect 21315 20009 21327 20012
rect 21269 20003 21327 20009
rect 23014 20000 23020 20012
rect 23072 20000 23078 20052
rect 25314 20040 25320 20052
rect 25275 20012 25320 20040
rect 25314 20000 25320 20012
rect 25372 20000 25378 20052
rect 25590 20040 25596 20052
rect 25551 20012 25596 20040
rect 25590 20000 25596 20012
rect 25648 20000 25654 20052
rect 26326 20040 26332 20052
rect 26287 20012 26332 20040
rect 26326 20000 26332 20012
rect 26384 20000 26390 20052
rect 22741 19975 22799 19981
rect 22741 19941 22753 19975
rect 22787 19972 22799 19975
rect 23382 19972 23388 19984
rect 22787 19944 23388 19972
rect 22787 19941 22799 19944
rect 22741 19935 22799 19941
rect 23382 19932 23388 19944
rect 23440 19972 23446 19984
rect 23440 19944 25544 19972
rect 23440 19932 23446 19944
rect 23290 19904 23296 19916
rect 20824 19876 23296 19904
rect 23290 19864 23296 19876
rect 23348 19864 23354 19916
rect 25056 19876 25452 19904
rect 25056 19848 25084 19876
rect 20346 19845 20352 19848
rect 20309 19839 20352 19845
rect 20309 19805 20321 19839
rect 20309 19799 20352 19805
rect 20346 19796 20352 19799
rect 20404 19796 20410 19848
rect 21450 19836 21456 19848
rect 21411 19808 21456 19836
rect 21450 19796 21456 19808
rect 21508 19796 21514 19848
rect 22186 19796 22192 19848
rect 22244 19836 22250 19848
rect 22557 19839 22615 19845
rect 22557 19836 22569 19839
rect 22244 19808 22569 19836
rect 22244 19796 22250 19808
rect 22557 19805 22569 19808
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 22738 19796 22744 19848
rect 22796 19796 22802 19848
rect 25038 19836 25044 19848
rect 24999 19808 25044 19836
rect 25038 19796 25044 19808
rect 25096 19796 25102 19848
rect 25424 19845 25452 19876
rect 25133 19839 25191 19845
rect 25133 19805 25145 19839
rect 25179 19805 25191 19839
rect 25133 19799 25191 19805
rect 25409 19839 25467 19845
rect 25409 19805 25421 19839
rect 25455 19805 25467 19839
rect 25516 19836 25544 19944
rect 26234 19864 26240 19916
rect 26292 19904 26298 19916
rect 26605 19907 26663 19913
rect 26605 19904 26617 19907
rect 26292 19876 26617 19904
rect 26292 19864 26298 19876
rect 26605 19873 26617 19876
rect 26651 19873 26663 19907
rect 26878 19904 26884 19916
rect 26839 19876 26884 19904
rect 26605 19867 26663 19873
rect 26878 19864 26884 19876
rect 26936 19864 26942 19916
rect 26145 19839 26203 19845
rect 26145 19836 26157 19839
rect 25516 19808 26157 19836
rect 25409 19799 25467 19805
rect 26145 19805 26157 19808
rect 26191 19805 26203 19839
rect 26145 19799 26203 19805
rect 20073 19771 20131 19777
rect 20073 19768 20085 19771
rect 18656 19740 20085 19768
rect 18656 19728 18662 19740
rect 20073 19737 20085 19740
rect 20119 19737 20131 19771
rect 20073 19731 20131 19737
rect 20165 19771 20223 19777
rect 20165 19737 20177 19771
rect 20211 19768 20223 19771
rect 20714 19768 20720 19780
rect 20211 19740 20720 19768
rect 20211 19737 20223 19740
rect 20165 19731 20223 19737
rect 20714 19728 20720 19740
rect 20772 19728 20778 19780
rect 22094 19728 22100 19780
rect 22152 19768 22158 19780
rect 22462 19768 22468 19780
rect 22152 19740 22468 19768
rect 22152 19728 22158 19740
rect 22462 19728 22468 19740
rect 22520 19768 22526 19780
rect 22756 19768 22784 19796
rect 22520 19740 22784 19768
rect 22520 19728 22526 19740
rect 25148 19712 25176 19799
rect 28166 19796 28172 19848
rect 28224 19836 28230 19848
rect 28721 19839 28779 19845
rect 28721 19836 28733 19839
rect 28224 19808 28733 19836
rect 28224 19796 28230 19808
rect 28721 19805 28733 19808
rect 28767 19805 28779 19839
rect 28721 19799 28779 19805
rect 27614 19728 27620 19780
rect 27672 19728 27678 19780
rect 17788 19672 18552 19700
rect 18690 19660 18696 19712
rect 18748 19700 18754 19712
rect 21542 19700 21548 19712
rect 18748 19672 21548 19700
rect 18748 19660 18754 19672
rect 21542 19660 21548 19672
rect 21600 19660 21606 19712
rect 21818 19660 21824 19712
rect 21876 19700 21882 19712
rect 22002 19700 22008 19712
rect 21876 19672 22008 19700
rect 21876 19660 21882 19672
rect 22002 19660 22008 19672
rect 22060 19700 22066 19712
rect 22278 19700 22284 19712
rect 22060 19672 22284 19700
rect 22060 19660 22066 19672
rect 22278 19660 22284 19672
rect 22336 19660 22342 19712
rect 24949 19703 25007 19709
rect 24949 19669 24961 19703
rect 24995 19700 25007 19703
rect 25130 19700 25136 19712
rect 24995 19672 25136 19700
rect 24995 19669 25007 19672
rect 24949 19663 25007 19669
rect 25130 19660 25136 19672
rect 25188 19660 25194 19712
rect 26970 19660 26976 19712
rect 27028 19700 27034 19712
rect 28353 19703 28411 19709
rect 28353 19700 28365 19703
rect 27028 19672 28365 19700
rect 27028 19660 27034 19672
rect 28353 19669 28365 19672
rect 28399 19669 28411 19703
rect 28534 19700 28540 19712
rect 28495 19672 28540 19700
rect 28353 19663 28411 19669
rect 28534 19660 28540 19672
rect 28592 19660 28598 19712
rect 1104 19610 29532 19632
rect 1104 19558 10425 19610
rect 10477 19558 10489 19610
rect 10541 19558 10553 19610
rect 10605 19558 10617 19610
rect 10669 19558 10681 19610
rect 10733 19558 19901 19610
rect 19953 19558 19965 19610
rect 20017 19558 20029 19610
rect 20081 19558 20093 19610
rect 20145 19558 20157 19610
rect 20209 19558 29532 19610
rect 1104 19536 29532 19558
rect 2777 19499 2835 19505
rect 2777 19465 2789 19499
rect 2823 19496 2835 19499
rect 2958 19496 2964 19508
rect 2823 19468 2964 19496
rect 2823 19465 2835 19468
rect 2777 19459 2835 19465
rect 2958 19456 2964 19468
rect 3016 19456 3022 19508
rect 4065 19499 4123 19505
rect 4065 19465 4077 19499
rect 4111 19496 4123 19499
rect 4522 19496 4528 19508
rect 4111 19468 4528 19496
rect 4111 19465 4123 19468
rect 4065 19459 4123 19465
rect 4522 19456 4528 19468
rect 4580 19456 4586 19508
rect 4982 19496 4988 19508
rect 4943 19468 4988 19496
rect 4982 19456 4988 19468
rect 5040 19456 5046 19508
rect 5994 19456 6000 19508
rect 6052 19496 6058 19508
rect 6825 19499 6883 19505
rect 6825 19496 6837 19499
rect 6052 19468 6837 19496
rect 6052 19456 6058 19468
rect 6825 19465 6837 19468
rect 6871 19465 6883 19499
rect 6825 19459 6883 19465
rect 7282 19456 7288 19508
rect 7340 19496 7346 19508
rect 7469 19499 7527 19505
rect 7469 19496 7481 19499
rect 7340 19468 7481 19496
rect 7340 19456 7346 19468
rect 7469 19465 7481 19468
rect 7515 19465 7527 19499
rect 7742 19496 7748 19508
rect 7703 19468 7748 19496
rect 7469 19459 7527 19465
rect 2976 19428 3004 19456
rect 6012 19428 6040 19456
rect 2976 19400 3280 19428
rect 3252 19369 3280 19400
rect 5184 19400 6040 19428
rect 1664 19363 1722 19369
rect 1664 19329 1676 19363
rect 1710 19360 1722 19363
rect 3053 19363 3111 19369
rect 3053 19360 3065 19363
rect 1710 19332 3065 19360
rect 1710 19329 1722 19332
rect 1664 19323 1722 19329
rect 3053 19329 3065 19332
rect 3099 19329 3111 19363
rect 3053 19323 3111 19329
rect 3237 19363 3295 19369
rect 3237 19329 3249 19363
rect 3283 19329 3295 19363
rect 3237 19323 3295 19329
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 4062 19360 4068 19372
rect 3375 19332 4068 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 5184 19369 5212 19400
rect 6546 19388 6552 19440
rect 6604 19428 6610 19440
rect 6733 19431 6791 19437
rect 6733 19428 6745 19431
rect 6604 19400 6745 19428
rect 6604 19388 6610 19400
rect 6733 19397 6745 19400
rect 6779 19397 6791 19431
rect 6733 19391 6791 19397
rect 5169 19363 5227 19369
rect 5169 19329 5181 19363
rect 5215 19329 5227 19363
rect 5169 19323 5227 19329
rect 5258 19320 5264 19372
rect 5316 19360 5322 19372
rect 5316 19332 5361 19360
rect 5316 19320 5322 19332
rect 7006 19320 7012 19372
rect 7064 19360 7070 19372
rect 7285 19363 7343 19369
rect 7285 19360 7297 19363
rect 7064 19332 7297 19360
rect 7064 19320 7070 19332
rect 7285 19329 7297 19332
rect 7331 19329 7343 19363
rect 7484 19360 7512 19459
rect 7742 19456 7748 19468
rect 7800 19456 7806 19508
rect 9493 19499 9551 19505
rect 9493 19465 9505 19499
rect 9539 19465 9551 19499
rect 9493 19459 9551 19465
rect 7926 19428 7932 19440
rect 7887 19400 7932 19428
rect 7926 19388 7932 19400
rect 7984 19388 7990 19440
rect 9508 19428 9536 19459
rect 9582 19456 9588 19508
rect 9640 19496 9646 19508
rect 9769 19499 9827 19505
rect 9769 19496 9781 19499
rect 9640 19468 9781 19496
rect 9640 19456 9646 19468
rect 9769 19465 9781 19468
rect 9815 19465 9827 19499
rect 9769 19459 9827 19465
rect 10042 19456 10048 19508
rect 10100 19496 10106 19508
rect 10137 19499 10195 19505
rect 10137 19496 10149 19499
rect 10100 19468 10149 19496
rect 10100 19456 10106 19468
rect 10137 19465 10149 19468
rect 10183 19465 10195 19499
rect 12894 19496 12900 19508
rect 12855 19468 12900 19496
rect 10137 19459 10195 19465
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 13449 19499 13507 19505
rect 13449 19496 13461 19499
rect 13320 19468 13461 19496
rect 13320 19456 13326 19468
rect 13449 19465 13461 19468
rect 13495 19496 13507 19499
rect 14918 19496 14924 19508
rect 13495 19468 14924 19496
rect 13495 19465 13507 19468
rect 13449 19459 13507 19465
rect 14918 19456 14924 19468
rect 14976 19456 14982 19508
rect 16022 19456 16028 19508
rect 16080 19496 16086 19508
rect 18138 19496 18144 19508
rect 16080 19468 18144 19496
rect 16080 19456 16086 19468
rect 9508 19400 10364 19428
rect 7558 19360 7564 19372
rect 7471 19332 7564 19360
rect 7285 19323 7343 19329
rect 1394 19292 1400 19304
rect 1355 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19252 1458 19304
rect 3605 19295 3663 19301
rect 3605 19261 3617 19295
rect 3651 19261 3663 19295
rect 4154 19292 4160 19304
rect 4115 19264 4160 19292
rect 3605 19255 3663 19261
rect 3620 19224 3648 19255
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 4249 19295 4307 19301
rect 4249 19261 4261 19295
rect 4295 19261 4307 19295
rect 5534 19292 5540 19304
rect 5495 19264 5540 19292
rect 4249 19255 4307 19261
rect 3697 19227 3755 19233
rect 3697 19224 3709 19227
rect 3620 19196 3709 19224
rect 3697 19193 3709 19196
rect 3743 19193 3755 19227
rect 3697 19187 3755 19193
rect 3878 19184 3884 19236
rect 3936 19224 3942 19236
rect 4264 19224 4292 19255
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 6917 19295 6975 19301
rect 6917 19261 6929 19295
rect 6963 19261 6975 19295
rect 7300 19292 7328 19323
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 7944 19292 7972 19388
rect 9309 19363 9367 19369
rect 9309 19329 9321 19363
rect 9355 19360 9367 19363
rect 9490 19360 9496 19372
rect 9355 19332 9496 19360
rect 9355 19329 9367 19332
rect 9309 19323 9367 19329
rect 9490 19320 9496 19332
rect 9548 19320 9554 19372
rect 9585 19363 9643 19369
rect 9585 19329 9597 19363
rect 9631 19329 9643 19363
rect 9585 19323 9643 19329
rect 7300 19264 7972 19292
rect 9600 19292 9628 19323
rect 9674 19320 9680 19372
rect 9732 19360 9738 19372
rect 9861 19363 9919 19369
rect 9861 19360 9873 19363
rect 9732 19332 9873 19360
rect 9732 19320 9738 19332
rect 9861 19329 9873 19332
rect 9907 19329 9919 19363
rect 9861 19323 9919 19329
rect 9950 19320 9956 19372
rect 10008 19320 10014 19372
rect 10134 19360 10140 19372
rect 10060 19332 10140 19360
rect 9766 19292 9772 19304
rect 9600 19264 9772 19292
rect 6917 19255 6975 19261
rect 6546 19224 6552 19236
rect 3936 19196 6552 19224
rect 3936 19184 3942 19196
rect 6546 19184 6552 19196
rect 6604 19224 6610 19236
rect 6932 19224 6960 19255
rect 9766 19252 9772 19264
rect 9824 19292 9830 19304
rect 9968 19292 9996 19320
rect 9824 19264 9996 19292
rect 9824 19252 9830 19264
rect 10060 19233 10088 19332
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 10336 19369 10364 19400
rect 10778 19388 10784 19440
rect 10836 19428 10842 19440
rect 11974 19428 11980 19440
rect 10836 19400 11980 19428
rect 10836 19388 10842 19400
rect 11164 19369 11192 19400
rect 11974 19388 11980 19400
rect 12032 19428 12038 19440
rect 12158 19428 12164 19440
rect 12032 19400 12164 19428
rect 12032 19388 12038 19400
rect 12158 19388 12164 19400
rect 12216 19388 12222 19440
rect 16850 19428 16856 19440
rect 16811 19400 16856 19428
rect 16850 19388 16856 19400
rect 16908 19388 16914 19440
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19329 10379 19363
rect 10321 19323 10379 19329
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19329 11207 19363
rect 11149 19323 11207 19329
rect 11609 19363 11667 19369
rect 11609 19329 11621 19363
rect 11655 19329 11667 19363
rect 11609 19323 11667 19329
rect 6604 19196 6960 19224
rect 10045 19227 10103 19233
rect 6604 19184 6610 19196
rect 10045 19193 10057 19227
rect 10091 19193 10103 19227
rect 10045 19187 10103 19193
rect 11241 19227 11299 19233
rect 11241 19193 11253 19227
rect 11287 19224 11299 19227
rect 11514 19224 11520 19236
rect 11287 19196 11520 19224
rect 11287 19193 11299 19196
rect 11241 19187 11299 19193
rect 11514 19184 11520 19196
rect 11572 19224 11578 19236
rect 11624 19224 11652 19323
rect 11698 19320 11704 19372
rect 11756 19320 11762 19372
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19360 11851 19363
rect 11882 19360 11888 19372
rect 11839 19332 11888 19360
rect 11839 19329 11851 19332
rect 11793 19323 11851 19329
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 12066 19360 12072 19372
rect 12027 19332 12072 19360
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 12253 19363 12311 19369
rect 12253 19329 12265 19363
rect 12299 19360 12311 19363
rect 12342 19360 12348 19372
rect 12299 19332 12348 19360
rect 12299 19329 12311 19332
rect 12253 19323 12311 19329
rect 12342 19320 12348 19332
rect 12400 19320 12406 19372
rect 12618 19320 12624 19372
rect 12676 19360 12682 19372
rect 13265 19363 13323 19369
rect 13265 19360 13277 19363
rect 12676 19332 13277 19360
rect 12676 19320 12682 19332
rect 13265 19329 13277 19332
rect 13311 19329 13323 19363
rect 13265 19323 13323 19329
rect 13354 19320 13360 19372
rect 13412 19360 13418 19372
rect 14185 19363 14243 19369
rect 13412 19332 13457 19360
rect 13412 19320 13418 19332
rect 14185 19329 14197 19363
rect 14231 19360 14243 19363
rect 14366 19360 14372 19372
rect 14231 19332 14372 19360
rect 14231 19329 14243 19332
rect 14185 19323 14243 19329
rect 14366 19320 14372 19332
rect 14424 19360 14430 19372
rect 14921 19363 14979 19369
rect 14921 19360 14933 19363
rect 14424 19332 14933 19360
rect 14424 19320 14430 19332
rect 14921 19329 14933 19332
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 15930 19320 15936 19372
rect 15988 19360 15994 19372
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 15988 19332 16129 19360
rect 15988 19320 15994 19332
rect 16117 19329 16129 19332
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 16393 19363 16451 19369
rect 16393 19329 16405 19363
rect 16439 19360 16451 19363
rect 16666 19360 16672 19372
rect 16439 19332 16528 19360
rect 16627 19332 16672 19360
rect 16439 19329 16451 19332
rect 16393 19323 16451 19329
rect 11716 19292 11744 19320
rect 11977 19295 12035 19301
rect 11977 19292 11989 19295
rect 11716 19264 11989 19292
rect 11977 19261 11989 19264
rect 12023 19261 12035 19295
rect 11977 19255 12035 19261
rect 13173 19295 13231 19301
rect 13173 19261 13185 19295
rect 13219 19292 13231 19295
rect 13446 19292 13452 19304
rect 13219 19264 13452 19292
rect 13219 19261 13231 19264
rect 13173 19255 13231 19261
rect 13446 19252 13452 19264
rect 13504 19252 13510 19304
rect 14274 19292 14280 19304
rect 14235 19264 14280 19292
rect 14274 19252 14280 19264
rect 14332 19252 14338 19304
rect 16022 19292 16028 19304
rect 15983 19264 16028 19292
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 16500 19292 16528 19332
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 17052 19369 17080 19468
rect 18138 19456 18144 19468
rect 18196 19496 18202 19508
rect 18196 19468 18267 19496
rect 18196 19456 18202 19468
rect 17238 19431 17296 19437
rect 17238 19397 17250 19431
rect 17284 19428 17296 19431
rect 18046 19428 18052 19440
rect 17284 19400 18052 19428
rect 17284 19397 17296 19400
rect 17238 19391 17296 19397
rect 18046 19388 18052 19400
rect 18104 19388 18110 19440
rect 18239 19428 18267 19468
rect 18506 19456 18512 19508
rect 18564 19496 18570 19508
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 18564 19468 20453 19496
rect 18564 19456 18570 19468
rect 20441 19465 20453 19468
rect 20487 19465 20499 19499
rect 20441 19459 20499 19465
rect 20714 19456 20720 19508
rect 20772 19496 20778 19508
rect 21177 19499 21235 19505
rect 21177 19496 21189 19499
rect 20772 19468 21189 19496
rect 20772 19456 20778 19468
rect 21177 19465 21189 19468
rect 21223 19465 21235 19499
rect 21177 19459 21235 19465
rect 21637 19499 21695 19505
rect 21637 19465 21649 19499
rect 21683 19496 21695 19499
rect 22094 19496 22100 19508
rect 21683 19468 22100 19496
rect 21683 19465 21695 19468
rect 21637 19459 21695 19465
rect 18598 19428 18604 19440
rect 18239 19400 18368 19428
rect 18559 19400 18604 19428
rect 16945 19363 17003 19369
rect 16945 19329 16957 19363
rect 16991 19329 17003 19363
rect 16945 19323 17003 19329
rect 17042 19363 17100 19369
rect 17042 19329 17054 19363
rect 17088 19329 17100 19363
rect 17678 19360 17684 19372
rect 17639 19332 17684 19360
rect 17042 19323 17100 19329
rect 16960 19292 16988 19323
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 18340 19369 18368 19400
rect 18598 19388 18604 19400
rect 18656 19388 18662 19440
rect 21192 19428 21220 19459
rect 22094 19456 22100 19468
rect 22152 19456 22158 19508
rect 23474 19496 23480 19508
rect 22204 19468 23480 19496
rect 21726 19428 21732 19440
rect 21192 19400 21732 19428
rect 21726 19388 21732 19400
rect 21784 19428 21790 19440
rect 21784 19400 21864 19428
rect 21784 19388 21790 19400
rect 18340 19363 18423 19369
rect 18340 19332 18377 19363
rect 18365 19329 18377 19332
rect 18411 19329 18423 19363
rect 18365 19323 18423 19329
rect 18509 19363 18567 19369
rect 18509 19329 18521 19363
rect 18555 19329 18567 19363
rect 18782 19360 18788 19372
rect 18743 19332 18788 19360
rect 18509 19323 18567 19329
rect 17126 19292 17132 19304
rect 16500 19264 16620 19292
rect 16960 19264 17132 19292
rect 14292 19224 14320 19252
rect 14550 19224 14556 19236
rect 11572 19196 14320 19224
rect 14511 19196 14556 19224
rect 11572 19184 11578 19196
rect 14550 19184 14556 19196
rect 14608 19184 14614 19236
rect 14734 19224 14740 19236
rect 14695 19196 14740 19224
rect 14734 19184 14740 19196
rect 14792 19184 14798 19236
rect 16592 19224 16620 19264
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 18524 19292 18552 19323
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19360 20315 19363
rect 20714 19360 20720 19372
rect 20303 19332 20720 19360
rect 20303 19329 20315 19332
rect 20257 19323 20315 19329
rect 20714 19320 20720 19332
rect 20772 19320 20778 19372
rect 21358 19360 21364 19372
rect 21319 19332 21364 19360
rect 21358 19320 21364 19332
rect 21416 19320 21422 19372
rect 21450 19320 21456 19372
rect 21508 19360 21514 19372
rect 21836 19369 21864 19400
rect 21821 19363 21879 19369
rect 21508 19332 21553 19360
rect 21508 19320 21514 19332
rect 21821 19329 21833 19363
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 22002 19320 22008 19372
rect 22060 19360 22066 19372
rect 22094 19360 22100 19372
rect 22060 19332 22100 19360
rect 22060 19320 22066 19332
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 22204 19360 22232 19468
rect 23474 19456 23480 19468
rect 23532 19456 23538 19508
rect 26053 19499 26111 19505
rect 26053 19496 26065 19499
rect 23860 19468 26065 19496
rect 22278 19388 22284 19440
rect 22336 19428 22342 19440
rect 23860 19437 23888 19468
rect 26053 19465 26065 19468
rect 26099 19496 26111 19499
rect 26418 19496 26424 19508
rect 26099 19468 26424 19496
rect 26099 19465 26111 19468
rect 26053 19459 26111 19465
rect 26418 19456 26424 19468
rect 26476 19456 26482 19508
rect 27341 19499 27399 19505
rect 27341 19465 27353 19499
rect 27387 19465 27399 19499
rect 27614 19496 27620 19508
rect 27575 19468 27620 19496
rect 27341 19459 27399 19465
rect 23753 19431 23811 19437
rect 23753 19428 23765 19431
rect 22336 19400 23765 19428
rect 22336 19388 22342 19400
rect 23753 19397 23765 19400
rect 23799 19397 23811 19431
rect 23753 19391 23811 19397
rect 23845 19431 23903 19437
rect 23845 19397 23857 19431
rect 23891 19397 23903 19431
rect 23845 19391 23903 19397
rect 25222 19388 25228 19440
rect 25280 19388 25286 19440
rect 22413 19363 22471 19369
rect 22413 19360 22425 19363
rect 22204 19332 22425 19360
rect 22413 19329 22425 19332
rect 22459 19329 22471 19363
rect 22556 19363 22614 19369
rect 22556 19360 22568 19363
rect 22535 19332 22568 19360
rect 22413 19323 22471 19329
rect 22556 19329 22568 19332
rect 22602 19329 22614 19363
rect 22556 19323 22614 19329
rect 22649 19363 22707 19369
rect 22649 19329 22661 19363
rect 22695 19360 22707 19363
rect 22738 19360 22744 19372
rect 22695 19332 22744 19360
rect 22695 19329 22707 19332
rect 22649 19323 22707 19329
rect 20622 19292 20628 19304
rect 18524 19264 19012 19292
rect 20583 19264 20628 19292
rect 17770 19224 17776 19236
rect 16592 19196 17776 19224
rect 17770 19184 17776 19196
rect 17828 19184 17834 19236
rect 3510 19156 3516 19168
rect 3471 19128 3516 19156
rect 3510 19116 3516 19128
rect 3568 19116 3574 19168
rect 5445 19159 5503 19165
rect 5445 19125 5457 19159
rect 5491 19156 5503 19159
rect 5534 19156 5540 19168
rect 5491 19128 5540 19156
rect 5491 19125 5503 19128
rect 5445 19119 5503 19125
rect 5534 19116 5540 19128
rect 5592 19116 5598 19168
rect 6362 19156 6368 19168
rect 6323 19128 6368 19156
rect 6362 19116 6368 19128
rect 6420 19116 6426 19168
rect 13262 19156 13268 19168
rect 13223 19128 13268 19156
rect 13262 19116 13268 19128
rect 13320 19116 13326 19168
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 14185 19159 14243 19165
rect 14185 19156 14197 19159
rect 13780 19128 14197 19156
rect 13780 19116 13786 19128
rect 14185 19125 14197 19128
rect 14231 19125 14243 19159
rect 17494 19156 17500 19168
rect 17455 19128 17500 19156
rect 14185 19119 14243 19125
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18414 19156 18420 19168
rect 18279 19128 18420 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18414 19116 18420 19128
rect 18472 19116 18478 19168
rect 18984 19165 19012 19264
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 22020 19233 22048 19320
rect 22571 19306 22600 19323
rect 22738 19320 22744 19332
rect 22796 19320 22802 19372
rect 22833 19363 22891 19369
rect 22833 19329 22845 19363
rect 22879 19360 22891 19363
rect 22922 19360 22928 19372
rect 22879 19332 22928 19360
rect 22879 19329 22891 19332
rect 22833 19323 22891 19329
rect 22922 19320 22928 19332
rect 22980 19360 22986 19372
rect 23290 19360 23296 19372
rect 22980 19332 23152 19360
rect 23251 19332 23296 19360
rect 22980 19320 22986 19332
rect 22571 19236 22599 19306
rect 23124 19292 23152 19332
rect 23290 19320 23296 19332
rect 23348 19320 23354 19372
rect 23569 19363 23627 19369
rect 23569 19360 23581 19363
rect 23400 19332 23581 19360
rect 23400 19292 23428 19332
rect 23569 19329 23581 19332
rect 23615 19360 23627 19363
rect 23658 19360 23664 19372
rect 23615 19332 23664 19360
rect 23615 19329 23627 19332
rect 23569 19323 23627 19329
rect 23658 19320 23664 19332
rect 23716 19320 23722 19372
rect 23942 19363 24000 19369
rect 23942 19360 23954 19363
rect 23768 19332 23954 19360
rect 23768 19292 23796 19332
rect 23942 19329 23954 19332
rect 23988 19329 24000 19363
rect 24302 19360 24308 19372
rect 24263 19332 24308 19360
rect 23942 19323 24000 19329
rect 24302 19320 24308 19332
rect 24360 19320 24366 19372
rect 26326 19320 26332 19372
rect 26384 19360 26390 19372
rect 26513 19363 26571 19369
rect 26513 19360 26525 19363
rect 26384 19332 26525 19360
rect 26384 19320 26390 19332
rect 26513 19329 26525 19332
rect 26559 19360 26571 19363
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 26559 19332 27169 19360
rect 26559 19329 26571 19332
rect 26513 19323 26571 19329
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27356 19360 27384 19459
rect 27614 19456 27620 19468
rect 27672 19456 27678 19508
rect 27433 19363 27491 19369
rect 27433 19360 27445 19363
rect 27356 19332 27445 19360
rect 27157 19323 27215 19329
rect 27433 19329 27445 19332
rect 27479 19329 27491 19363
rect 27433 19323 27491 19329
rect 28261 19363 28319 19369
rect 28261 19329 28273 19363
rect 28307 19360 28319 19363
rect 28534 19360 28540 19372
rect 28307 19332 28540 19360
rect 28307 19329 28319 19332
rect 28261 19323 28319 19329
rect 28534 19320 28540 19332
rect 28592 19320 28598 19372
rect 24581 19295 24639 19301
rect 24581 19292 24593 19295
rect 23124 19264 23428 19292
rect 23676 19264 23796 19292
rect 24136 19264 24593 19292
rect 22005 19227 22063 19233
rect 22005 19193 22017 19227
rect 22051 19193 22063 19227
rect 22554 19224 22560 19236
rect 22467 19196 22560 19224
rect 22005 19187 22063 19193
rect 22554 19184 22560 19196
rect 22612 19224 22618 19236
rect 22612 19196 23060 19224
rect 22612 19184 22618 19196
rect 18969 19159 19027 19165
rect 18969 19125 18981 19159
rect 19015 19156 19027 19159
rect 19058 19156 19064 19168
rect 19015 19128 19064 19156
rect 19015 19125 19027 19128
rect 18969 19119 19027 19125
rect 19058 19116 19064 19128
rect 19116 19116 19122 19168
rect 20809 19159 20867 19165
rect 20809 19125 20821 19159
rect 20855 19156 20867 19159
rect 21082 19156 21088 19168
rect 20855 19128 21088 19156
rect 20855 19125 20867 19128
rect 20809 19119 20867 19125
rect 21082 19116 21088 19128
rect 21140 19156 21146 19168
rect 21450 19156 21456 19168
rect 21140 19128 21456 19156
rect 21140 19116 21146 19128
rect 21450 19116 21456 19128
rect 21508 19116 21514 19168
rect 22281 19159 22339 19165
rect 22281 19125 22293 19159
rect 22327 19156 22339 19159
rect 22370 19156 22376 19168
rect 22327 19128 22376 19156
rect 22327 19125 22339 19128
rect 22281 19119 22339 19125
rect 22370 19116 22376 19128
rect 22428 19116 22434 19168
rect 23032 19165 23060 19196
rect 23676 19168 23704 19264
rect 24136 19233 24164 19264
rect 24581 19261 24593 19264
rect 24627 19261 24639 19295
rect 24581 19255 24639 19261
rect 24121 19227 24179 19233
rect 24121 19193 24133 19227
rect 24167 19193 24179 19227
rect 24121 19187 24179 19193
rect 23017 19159 23075 19165
rect 23017 19125 23029 19159
rect 23063 19156 23075 19159
rect 23382 19156 23388 19168
rect 23063 19128 23388 19156
rect 23063 19125 23075 19128
rect 23017 19119 23075 19125
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 23474 19116 23480 19168
rect 23532 19156 23538 19168
rect 23658 19156 23664 19168
rect 23532 19128 23664 19156
rect 23532 19116 23538 19128
rect 23658 19116 23664 19128
rect 23716 19116 23722 19168
rect 24026 19116 24032 19168
rect 24084 19156 24090 19168
rect 25774 19156 25780 19168
rect 24084 19128 25780 19156
rect 24084 19116 24090 19128
rect 25774 19116 25780 19128
rect 25832 19116 25838 19168
rect 26329 19159 26387 19165
rect 26329 19125 26341 19159
rect 26375 19156 26387 19159
rect 26418 19156 26424 19168
rect 26375 19128 26424 19156
rect 26375 19125 26387 19128
rect 26329 19119 26387 19125
rect 26418 19116 26424 19128
rect 26476 19116 26482 19168
rect 28350 19116 28356 19168
rect 28408 19156 28414 19168
rect 28445 19159 28503 19165
rect 28445 19156 28457 19159
rect 28408 19128 28457 19156
rect 28408 19116 28414 19128
rect 28445 19125 28457 19128
rect 28491 19125 28503 19159
rect 28445 19119 28503 19125
rect 1104 19066 29532 19088
rect 1104 19014 5688 19066
rect 5740 19014 5752 19066
rect 5804 19014 5816 19066
rect 5868 19014 5880 19066
rect 5932 19014 5944 19066
rect 5996 19014 15163 19066
rect 15215 19014 15227 19066
rect 15279 19014 15291 19066
rect 15343 19014 15355 19066
rect 15407 19014 15419 19066
rect 15471 19014 24639 19066
rect 24691 19014 24703 19066
rect 24755 19014 24767 19066
rect 24819 19014 24831 19066
rect 24883 19014 24895 19066
rect 24947 19014 29532 19066
rect 1104 18992 29532 19014
rect 3510 18912 3516 18964
rect 3568 18952 3574 18964
rect 3881 18955 3939 18961
rect 3881 18952 3893 18955
rect 3568 18924 3893 18952
rect 3568 18912 3574 18924
rect 3881 18921 3893 18924
rect 3927 18921 3939 18955
rect 3881 18915 3939 18921
rect 6454 18912 6460 18964
rect 6512 18952 6518 18964
rect 25222 18952 25228 18964
rect 6512 18924 25084 18952
rect 25183 18924 25228 18952
rect 6512 18912 6518 18924
rect 12986 18884 12992 18896
rect 12452 18856 12992 18884
rect 3237 18819 3295 18825
rect 3237 18785 3249 18819
rect 3283 18816 3295 18819
rect 3789 18819 3847 18825
rect 3789 18816 3801 18819
rect 3283 18788 3801 18816
rect 3283 18785 3295 18788
rect 3237 18779 3295 18785
rect 3789 18785 3801 18788
rect 3835 18785 3847 18819
rect 3789 18779 3847 18785
rect 9214 18776 9220 18828
rect 9272 18816 9278 18828
rect 11149 18819 11207 18825
rect 11149 18816 11161 18819
rect 9272 18788 11161 18816
rect 9272 18776 9278 18788
rect 11149 18785 11161 18788
rect 11195 18785 11207 18819
rect 11149 18779 11207 18785
rect 11977 18819 12035 18825
rect 11977 18785 11989 18819
rect 12023 18816 12035 18819
rect 12342 18816 12348 18828
rect 12023 18788 12348 18816
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 12342 18776 12348 18788
rect 12400 18776 12406 18828
rect 12452 18825 12480 18856
rect 12986 18844 12992 18856
rect 13044 18844 13050 18896
rect 13262 18884 13268 18896
rect 13175 18856 13268 18884
rect 13262 18844 13268 18856
rect 13320 18884 13326 18896
rect 15838 18884 15844 18896
rect 13320 18856 15844 18884
rect 13320 18844 13326 18856
rect 15838 18844 15844 18856
rect 15896 18844 15902 18896
rect 21542 18884 21548 18896
rect 21503 18856 21548 18884
rect 21542 18844 21548 18856
rect 21600 18844 21606 18896
rect 23382 18844 23388 18896
rect 23440 18884 23446 18896
rect 23845 18887 23903 18893
rect 23845 18884 23857 18887
rect 23440 18856 23857 18884
rect 23440 18844 23446 18856
rect 23845 18853 23857 18856
rect 23891 18853 23903 18887
rect 25056 18884 25084 18924
rect 25222 18912 25228 18924
rect 25280 18912 25286 18964
rect 26326 18884 26332 18896
rect 25056 18856 26332 18884
rect 23845 18847 23903 18853
rect 26326 18844 26332 18856
rect 26384 18844 26390 18896
rect 12437 18819 12495 18825
rect 12437 18785 12449 18819
rect 12483 18785 12495 18819
rect 12437 18779 12495 18785
rect 12529 18819 12587 18825
rect 12529 18785 12541 18819
rect 12575 18816 12587 18819
rect 12618 18816 12624 18828
rect 12575 18788 12624 18816
rect 12575 18785 12587 18788
rect 12529 18779 12587 18785
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 13722 18816 13728 18828
rect 12768 18788 13728 18816
rect 12768 18776 12774 18788
rect 13722 18776 13728 18788
rect 13780 18816 13786 18828
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 13780 18788 14105 18816
rect 13780 18776 13786 18788
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 14274 18776 14280 18828
rect 14332 18816 14338 18828
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 14332 18788 14381 18816
rect 14332 18776 14338 18788
rect 14369 18785 14381 18788
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 14553 18819 14611 18825
rect 14553 18785 14565 18819
rect 14599 18816 14611 18819
rect 14826 18816 14832 18828
rect 14599 18788 14832 18816
rect 14599 18785 14611 18788
rect 14553 18779 14611 18785
rect 14826 18776 14832 18788
rect 14884 18776 14890 18828
rect 15933 18819 15991 18825
rect 15933 18785 15945 18819
rect 15979 18816 15991 18819
rect 16114 18816 16120 18828
rect 15979 18788 16120 18816
rect 15979 18785 15991 18788
rect 15933 18779 15991 18785
rect 16114 18776 16120 18788
rect 16172 18776 16178 18828
rect 18046 18816 18052 18828
rect 18007 18788 18052 18816
rect 18046 18776 18052 18788
rect 18104 18776 18110 18828
rect 18322 18816 18328 18828
rect 18283 18788 18328 18816
rect 18322 18776 18328 18788
rect 18380 18816 18386 18828
rect 19981 18819 20039 18825
rect 19981 18816 19993 18819
rect 18380 18788 19993 18816
rect 18380 18776 18386 18788
rect 19981 18785 19993 18788
rect 20027 18785 20039 18819
rect 19981 18779 20039 18785
rect 22097 18819 22155 18825
rect 22097 18785 22109 18819
rect 22143 18816 22155 18819
rect 24302 18816 24308 18828
rect 22143 18788 24308 18816
rect 22143 18785 22155 18788
rect 22097 18779 22155 18785
rect 24302 18776 24308 18788
rect 24360 18776 24366 18828
rect 25130 18816 25136 18828
rect 24688 18788 25136 18816
rect 3421 18751 3479 18757
rect 3421 18717 3433 18751
rect 3467 18717 3479 18751
rect 3421 18711 3479 18717
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18748 3663 18751
rect 3694 18748 3700 18760
rect 3651 18720 3700 18748
rect 3651 18717 3663 18720
rect 3605 18711 3663 18717
rect 3436 18680 3464 18711
rect 3694 18708 3700 18720
rect 3752 18708 3758 18760
rect 4062 18748 4068 18760
rect 4023 18720 4068 18748
rect 4062 18708 4068 18720
rect 4120 18708 4126 18760
rect 4154 18708 4160 18760
rect 4212 18748 4218 18760
rect 4212 18720 4257 18748
rect 4212 18708 4218 18720
rect 4614 18708 4620 18760
rect 4672 18748 4678 18760
rect 4890 18748 4896 18760
rect 4672 18720 4896 18748
rect 4672 18708 4678 18720
rect 4890 18708 4896 18720
rect 4948 18708 4954 18760
rect 7466 18748 7472 18760
rect 7427 18720 7472 18748
rect 7466 18708 7472 18720
rect 7524 18708 7530 18760
rect 9674 18748 9680 18760
rect 9635 18720 9680 18748
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 10778 18748 10784 18760
rect 10739 18720 10784 18748
rect 10778 18708 10784 18720
rect 10836 18708 10842 18760
rect 11054 18748 11060 18760
rect 11015 18720 11060 18748
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 11238 18708 11244 18760
rect 11296 18748 11302 18760
rect 11333 18751 11391 18757
rect 11333 18748 11345 18751
rect 11296 18720 11345 18748
rect 11296 18708 11302 18720
rect 11333 18717 11345 18720
rect 11379 18717 11391 18751
rect 11514 18748 11520 18760
rect 11475 18720 11520 18748
rect 11333 18711 11391 18717
rect 3970 18680 3976 18692
rect 3436 18652 3976 18680
rect 3970 18640 3976 18652
rect 4028 18640 4034 18692
rect 5160 18683 5218 18689
rect 5160 18649 5172 18683
rect 5206 18680 5218 18683
rect 5258 18680 5264 18692
rect 5206 18652 5264 18680
rect 5206 18649 5218 18652
rect 5160 18643 5218 18649
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 11348 18680 11376 18711
rect 11514 18708 11520 18720
rect 11572 18708 11578 18760
rect 11882 18708 11888 18760
rect 11940 18748 11946 18760
rect 12161 18751 12219 18757
rect 12161 18748 12173 18751
rect 11940 18720 12173 18748
rect 11940 18708 11946 18720
rect 12161 18717 12173 18720
rect 12207 18717 12219 18751
rect 12161 18711 12219 18717
rect 12250 18708 12256 18760
rect 12308 18748 12314 18760
rect 12802 18748 12808 18760
rect 12308 18720 12353 18748
rect 12763 18720 12808 18748
rect 12308 18708 12314 18720
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 12986 18748 12992 18760
rect 12947 18720 12992 18748
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18748 13139 18751
rect 13354 18748 13360 18760
rect 13127 18720 13360 18748
rect 13127 18717 13139 18720
rect 13081 18711 13139 18717
rect 11793 18683 11851 18689
rect 11793 18680 11805 18683
rect 11348 18652 11805 18680
rect 11793 18649 11805 18652
rect 11839 18680 11851 18683
rect 12066 18680 12072 18692
rect 11839 18652 12072 18680
rect 11839 18649 11851 18652
rect 11793 18643 11851 18649
rect 12066 18640 12072 18652
rect 12124 18640 12130 18692
rect 12894 18640 12900 18692
rect 12952 18680 12958 18692
rect 13096 18680 13124 18711
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 15654 18748 15660 18760
rect 15615 18720 15660 18748
rect 15654 18708 15660 18720
rect 15712 18708 15718 18760
rect 15749 18751 15807 18757
rect 15749 18717 15761 18751
rect 15795 18748 15807 18751
rect 16022 18748 16028 18760
rect 15795 18720 16028 18748
rect 15795 18717 15807 18720
rect 15749 18711 15807 18717
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 20254 18757 20260 18760
rect 18417 18751 18475 18757
rect 18417 18748 18429 18751
rect 18340 18720 18429 18748
rect 12952 18652 13124 18680
rect 14829 18683 14887 18689
rect 12952 18640 12958 18652
rect 14829 18649 14841 18683
rect 14875 18680 14887 18683
rect 15010 18680 15016 18692
rect 14875 18652 15016 18680
rect 14875 18649 14887 18652
rect 14829 18643 14887 18649
rect 15010 18640 15016 18652
rect 15068 18640 15074 18692
rect 17494 18640 17500 18692
rect 17552 18640 17558 18692
rect 4338 18612 4344 18624
rect 4299 18584 4344 18612
rect 4338 18572 4344 18584
rect 4396 18572 4402 18624
rect 6273 18615 6331 18621
rect 6273 18581 6285 18615
rect 6319 18612 6331 18615
rect 6454 18612 6460 18624
rect 6319 18584 6460 18612
rect 6319 18581 6331 18584
rect 6273 18575 6331 18581
rect 6454 18572 6460 18584
rect 6512 18572 6518 18624
rect 7650 18612 7656 18624
rect 7611 18584 7656 18612
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 9861 18615 9919 18621
rect 9861 18581 9873 18615
rect 9907 18612 9919 18615
rect 9950 18612 9956 18624
rect 9907 18584 9956 18612
rect 9907 18581 9919 18584
rect 9861 18575 9919 18581
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 12342 18572 12348 18624
rect 12400 18612 12406 18624
rect 13262 18612 13268 18624
rect 12400 18584 13268 18612
rect 12400 18572 12406 18584
rect 13262 18572 13268 18584
rect 13320 18572 13326 18624
rect 13538 18572 13544 18624
rect 13596 18612 13602 18624
rect 14461 18615 14519 18621
rect 14461 18612 14473 18615
rect 13596 18584 14473 18612
rect 13596 18572 13602 18584
rect 14461 18581 14473 18584
rect 14507 18581 14519 18615
rect 14461 18575 14519 18581
rect 15289 18615 15347 18621
rect 15289 18581 15301 18615
rect 15335 18612 15347 18615
rect 16298 18612 16304 18624
rect 15335 18584 16304 18612
rect 15335 18581 15347 18584
rect 15289 18575 15347 18581
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 16577 18615 16635 18621
rect 16577 18581 16589 18615
rect 16623 18612 16635 18615
rect 17126 18612 17132 18624
rect 16623 18584 17132 18612
rect 16623 18581 16635 18584
rect 16577 18575 16635 18581
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 17402 18572 17408 18624
rect 17460 18612 17466 18624
rect 18340 18612 18368 18720
rect 18417 18717 18429 18720
rect 18463 18717 18475 18751
rect 18785 18751 18843 18757
rect 18785 18748 18797 18751
rect 18417 18711 18475 18717
rect 18616 18720 18797 18748
rect 18616 18621 18644 18720
rect 18785 18717 18797 18720
rect 18831 18717 18843 18751
rect 20248 18748 20260 18757
rect 20215 18720 20260 18748
rect 18785 18711 18843 18717
rect 20248 18711 20260 18720
rect 20254 18708 20260 18711
rect 20312 18708 20318 18760
rect 21726 18748 21732 18760
rect 21687 18720 21732 18748
rect 21726 18708 21732 18720
rect 21784 18708 21790 18760
rect 23658 18708 23664 18760
rect 23716 18748 23722 18760
rect 24486 18748 24492 18760
rect 23716 18720 24492 18748
rect 23716 18708 23722 18720
rect 24486 18708 24492 18720
rect 24544 18708 24550 18760
rect 24688 18757 24716 18788
rect 25130 18776 25136 18788
rect 25188 18776 25194 18828
rect 26234 18776 26240 18828
rect 26292 18816 26298 18828
rect 27341 18819 27399 18825
rect 27341 18816 27353 18819
rect 26292 18788 27353 18816
rect 26292 18776 26298 18788
rect 27341 18785 27353 18788
rect 27387 18785 27399 18819
rect 27341 18779 27399 18785
rect 24673 18751 24731 18757
rect 24673 18717 24685 18751
rect 24719 18717 24731 18751
rect 24673 18711 24731 18717
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18717 24823 18751
rect 25041 18751 25099 18757
rect 25041 18748 25053 18751
rect 24765 18711 24823 18717
rect 24964 18720 25053 18748
rect 22370 18680 22376 18692
rect 22331 18652 22376 18680
rect 22370 18640 22376 18652
rect 22428 18640 22434 18692
rect 23382 18640 23388 18692
rect 23440 18640 23446 18692
rect 24394 18640 24400 18692
rect 24452 18680 24458 18692
rect 24780 18680 24808 18711
rect 24452 18652 24808 18680
rect 24452 18640 24458 18652
rect 17460 18584 18368 18612
rect 18601 18615 18659 18621
rect 17460 18572 17466 18584
rect 18601 18581 18613 18615
rect 18647 18581 18659 18615
rect 18966 18612 18972 18624
rect 18927 18584 18972 18612
rect 18601 18575 18659 18581
rect 18966 18572 18972 18584
rect 19024 18572 19030 18624
rect 20714 18572 20720 18624
rect 20772 18612 20778 18624
rect 21358 18612 21364 18624
rect 20772 18584 21364 18612
rect 20772 18572 20778 18584
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 23750 18572 23756 18624
rect 23808 18612 23814 18624
rect 24964 18621 24992 18720
rect 25041 18717 25053 18720
rect 25087 18717 25099 18751
rect 26418 18748 26424 18760
rect 26379 18720 26424 18748
rect 25041 18711 25099 18717
rect 26418 18708 26424 18720
rect 26476 18708 26482 18760
rect 27617 18683 27675 18689
rect 27617 18649 27629 18683
rect 27663 18680 27675 18683
rect 27706 18680 27712 18692
rect 27663 18652 27712 18680
rect 27663 18649 27675 18652
rect 27617 18643 27675 18649
rect 27706 18640 27712 18652
rect 27764 18640 27770 18692
rect 28350 18640 28356 18692
rect 28408 18640 28414 18692
rect 24489 18615 24547 18621
rect 24489 18612 24501 18615
rect 23808 18584 24501 18612
rect 23808 18572 23814 18584
rect 24489 18581 24501 18584
rect 24535 18581 24547 18615
rect 24489 18575 24547 18581
rect 24949 18615 25007 18621
rect 24949 18581 24961 18615
rect 24995 18581 25007 18615
rect 26234 18612 26240 18624
rect 26195 18584 26240 18612
rect 24949 18575 25007 18581
rect 26234 18572 26240 18584
rect 26292 18572 26298 18624
rect 27798 18572 27804 18624
rect 27856 18612 27862 18624
rect 29089 18615 29147 18621
rect 29089 18612 29101 18615
rect 27856 18584 29101 18612
rect 27856 18572 27862 18584
rect 29089 18581 29101 18584
rect 29135 18581 29147 18615
rect 29089 18575 29147 18581
rect 1104 18522 29532 18544
rect 1104 18470 10425 18522
rect 10477 18470 10489 18522
rect 10541 18470 10553 18522
rect 10605 18470 10617 18522
rect 10669 18470 10681 18522
rect 10733 18470 19901 18522
rect 19953 18470 19965 18522
rect 20017 18470 20029 18522
rect 20081 18470 20093 18522
rect 20145 18470 20157 18522
rect 20209 18470 29532 18522
rect 1104 18448 29532 18470
rect 2593 18411 2651 18417
rect 2593 18377 2605 18411
rect 2639 18408 2651 18411
rect 3510 18408 3516 18420
rect 2639 18380 3516 18408
rect 2639 18377 2651 18380
rect 2593 18371 2651 18377
rect 3510 18368 3516 18380
rect 3568 18368 3574 18420
rect 4065 18411 4123 18417
rect 4065 18377 4077 18411
rect 4111 18408 4123 18411
rect 4154 18408 4160 18420
rect 4111 18380 4160 18408
rect 4111 18377 4123 18380
rect 4065 18371 4123 18377
rect 4154 18368 4160 18380
rect 4212 18368 4218 18420
rect 4525 18411 4583 18417
rect 4525 18377 4537 18411
rect 4571 18408 4583 18411
rect 5074 18408 5080 18420
rect 4571 18380 5080 18408
rect 4571 18377 4583 18380
rect 4525 18371 4583 18377
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 5258 18408 5264 18420
rect 5219 18380 5264 18408
rect 5258 18368 5264 18380
rect 5316 18368 5322 18420
rect 11146 18368 11152 18420
rect 11204 18408 11210 18420
rect 12434 18408 12440 18420
rect 11204 18380 12440 18408
rect 11204 18368 11210 18380
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 12526 18368 12532 18420
rect 12584 18408 12590 18420
rect 15381 18411 15439 18417
rect 15381 18408 15393 18411
rect 12584 18380 15393 18408
rect 12584 18368 12590 18380
rect 15381 18377 15393 18380
rect 15427 18377 15439 18411
rect 15746 18408 15752 18420
rect 15707 18380 15752 18408
rect 15381 18371 15439 18377
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 17589 18411 17647 18417
rect 17589 18377 17601 18411
rect 17635 18408 17647 18411
rect 17678 18408 17684 18420
rect 17635 18380 17684 18408
rect 17635 18377 17647 18380
rect 17589 18371 17647 18377
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 17770 18368 17776 18420
rect 17828 18408 17834 18420
rect 20901 18411 20959 18417
rect 20901 18408 20913 18411
rect 17828 18380 20913 18408
rect 17828 18368 17834 18380
rect 20901 18377 20913 18380
rect 20947 18377 20959 18411
rect 20901 18371 20959 18377
rect 23293 18411 23351 18417
rect 23293 18377 23305 18411
rect 23339 18377 23351 18411
rect 23293 18371 23351 18377
rect 1394 18300 1400 18352
rect 1452 18340 1458 18352
rect 4890 18340 4896 18352
rect 1452 18312 4896 18340
rect 1452 18300 1458 18312
rect 2700 18281 2728 18312
rect 4890 18300 4896 18312
rect 4948 18300 4954 18352
rect 6454 18340 6460 18352
rect 5460 18312 6460 18340
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18272 2467 18275
rect 2685 18275 2743 18281
rect 2455 18244 2645 18272
rect 2455 18241 2467 18244
rect 2409 18235 2467 18241
rect 2617 18068 2645 18244
rect 2685 18241 2697 18275
rect 2731 18241 2743 18275
rect 2685 18235 2743 18241
rect 2952 18275 3010 18281
rect 2952 18241 2964 18275
rect 2998 18272 3010 18275
rect 4338 18272 4344 18284
rect 2998 18244 4344 18272
rect 2998 18241 3010 18244
rect 2952 18235 3010 18241
rect 4338 18232 4344 18244
rect 4396 18232 4402 18284
rect 4706 18272 4712 18284
rect 4667 18244 4712 18272
rect 4706 18232 4712 18244
rect 4764 18232 4770 18284
rect 5460 18281 5488 18312
rect 6454 18300 6460 18312
rect 6512 18300 6518 18352
rect 7650 18300 7656 18352
rect 7708 18300 7714 18352
rect 9214 18340 9220 18352
rect 9175 18312 9220 18340
rect 9214 18300 9220 18312
rect 9272 18300 9278 18352
rect 9950 18300 9956 18352
rect 10008 18300 10014 18352
rect 12802 18300 12808 18352
rect 12860 18340 12866 18352
rect 13081 18343 13139 18349
rect 13081 18340 13093 18343
rect 12860 18312 13093 18340
rect 12860 18300 12866 18312
rect 13081 18309 13093 18312
rect 13127 18340 13139 18343
rect 13170 18340 13176 18352
rect 13127 18312 13176 18340
rect 13127 18309 13139 18312
rect 13081 18303 13139 18309
rect 13170 18300 13176 18312
rect 13228 18300 13234 18352
rect 14366 18340 14372 18352
rect 14327 18312 14372 18340
rect 14366 18300 14372 18312
rect 14424 18300 14430 18352
rect 18322 18340 18328 18352
rect 18156 18312 18328 18340
rect 18156 18284 18184 18312
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 18414 18300 18420 18352
rect 18472 18340 18478 18352
rect 18472 18312 18517 18340
rect 18472 18300 18478 18312
rect 18966 18300 18972 18352
rect 19024 18300 19030 18352
rect 5445 18275 5503 18281
rect 5445 18241 5457 18275
rect 5491 18241 5503 18275
rect 5445 18235 5503 18241
rect 5537 18275 5595 18281
rect 5537 18241 5549 18275
rect 5583 18241 5595 18275
rect 5537 18235 5595 18241
rect 5813 18275 5871 18281
rect 5813 18241 5825 18275
rect 5859 18272 5871 18275
rect 6362 18272 6368 18284
rect 5859 18244 6368 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 5074 18164 5080 18216
rect 5132 18204 5138 18216
rect 5552 18204 5580 18235
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 10965 18275 11023 18281
rect 10965 18241 10977 18275
rect 11011 18241 11023 18275
rect 10965 18235 11023 18241
rect 6638 18204 6644 18216
rect 5132 18176 5580 18204
rect 6599 18176 6644 18204
rect 5132 18164 5138 18176
rect 6638 18164 6644 18176
rect 6696 18164 6702 18216
rect 6914 18204 6920 18216
rect 6875 18176 6920 18204
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 8938 18204 8944 18216
rect 8899 18176 8944 18204
rect 8938 18164 8944 18176
rect 8996 18164 9002 18216
rect 10689 18207 10747 18213
rect 10689 18173 10701 18207
rect 10735 18204 10747 18207
rect 10980 18204 11008 18235
rect 11974 18232 11980 18284
rect 12032 18272 12038 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 12032 18244 12173 18272
rect 12032 18232 12038 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18272 12403 18275
rect 12710 18272 12716 18284
rect 12391 18244 12716 18272
rect 12391 18241 12403 18244
rect 12345 18235 12403 18241
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 13265 18275 13323 18281
rect 13265 18241 13277 18275
rect 13311 18272 13323 18275
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13311 18244 14013 18272
rect 13311 18241 13323 18244
rect 13265 18235 13323 18241
rect 14001 18241 14013 18244
rect 14047 18241 14059 18275
rect 14001 18235 14059 18241
rect 14185 18275 14243 18281
rect 14185 18241 14197 18275
rect 14231 18272 14243 18275
rect 14274 18272 14280 18284
rect 14231 18244 14280 18272
rect 14231 18241 14243 18244
rect 14185 18235 14243 18241
rect 14016 18204 14044 18235
rect 14274 18232 14280 18244
rect 14332 18232 14338 18284
rect 14734 18272 14740 18284
rect 14695 18244 14740 18272
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 17402 18272 17408 18284
rect 17363 18244 17408 18272
rect 17402 18232 17408 18244
rect 17460 18272 17466 18284
rect 17681 18275 17739 18281
rect 17681 18272 17693 18275
rect 17460 18244 17693 18272
rect 17460 18232 17466 18244
rect 17681 18241 17693 18244
rect 17727 18241 17739 18275
rect 18138 18272 18144 18284
rect 18051 18244 18144 18272
rect 17681 18235 17739 18241
rect 18138 18232 18144 18244
rect 18196 18232 18202 18284
rect 20714 18272 20720 18284
rect 20675 18244 20720 18272
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 21082 18272 21088 18284
rect 21043 18244 21088 18272
rect 21082 18232 21088 18244
rect 21140 18232 21146 18284
rect 23109 18275 23167 18281
rect 23109 18241 23121 18275
rect 23155 18241 23167 18275
rect 23308 18272 23336 18371
rect 23382 18368 23388 18420
rect 23440 18408 23446 18420
rect 23440 18380 23485 18408
rect 23440 18368 23446 18380
rect 24302 18368 24308 18420
rect 24360 18368 24366 18420
rect 24026 18300 24032 18352
rect 24084 18340 24090 18352
rect 24320 18340 24348 18368
rect 24084 18312 24256 18340
rect 24320 18312 24992 18340
rect 24084 18300 24090 18312
rect 23569 18275 23627 18281
rect 23569 18272 23581 18275
rect 23308 18244 23581 18272
rect 23109 18235 23167 18241
rect 23569 18241 23581 18244
rect 23615 18241 23627 18275
rect 23569 18235 23627 18241
rect 14752 18204 14780 18232
rect 15838 18204 15844 18216
rect 10735 18176 12388 18204
rect 14016 18176 14780 18204
rect 15799 18176 15844 18204
rect 10735 18173 10747 18176
rect 10689 18167 10747 18173
rect 5534 18096 5540 18148
rect 5592 18136 5598 18148
rect 5721 18139 5779 18145
rect 5721 18136 5733 18139
rect 5592 18108 5733 18136
rect 5592 18096 5598 18108
rect 5721 18105 5733 18108
rect 5767 18105 5779 18139
rect 5721 18099 5779 18105
rect 12360 18136 12388 18176
rect 15838 18164 15844 18176
rect 15896 18164 15902 18216
rect 16025 18207 16083 18213
rect 16025 18173 16037 18207
rect 16071 18204 16083 18207
rect 16114 18204 16120 18216
rect 16071 18176 16120 18204
rect 16071 18173 16083 18176
rect 16025 18167 16083 18173
rect 16114 18164 16120 18176
rect 16172 18164 16178 18216
rect 23124 18204 23152 18235
rect 23750 18232 23756 18284
rect 23808 18272 23814 18284
rect 24121 18275 24179 18281
rect 24121 18272 24133 18275
rect 23808 18244 24133 18272
rect 23808 18232 23814 18244
rect 24121 18241 24133 18244
rect 24167 18241 24179 18275
rect 24228 18272 24256 18312
rect 24305 18275 24363 18281
rect 24305 18272 24317 18275
rect 24228 18244 24317 18272
rect 24121 18235 24179 18241
rect 24305 18241 24317 18244
rect 24351 18241 24363 18275
rect 24305 18235 24363 18241
rect 24397 18275 24455 18281
rect 24397 18241 24409 18275
rect 24443 18241 24455 18275
rect 24397 18235 24455 18241
rect 23474 18204 23480 18216
rect 23124 18176 23480 18204
rect 23474 18164 23480 18176
rect 23532 18164 23538 18216
rect 24412 18204 24440 18235
rect 24486 18232 24492 18284
rect 24544 18281 24550 18284
rect 24964 18281 24992 18312
rect 26234 18300 26240 18352
rect 26292 18300 26298 18352
rect 27246 18300 27252 18352
rect 27304 18340 27310 18352
rect 27304 18312 27568 18340
rect 27304 18300 27310 18312
rect 24544 18272 24552 18281
rect 24949 18275 25007 18281
rect 24544 18244 24589 18272
rect 24544 18235 24552 18244
rect 24949 18241 24961 18275
rect 24995 18241 25007 18275
rect 24949 18235 25007 18241
rect 24544 18232 24550 18235
rect 26602 18232 26608 18284
rect 26660 18272 26666 18284
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 26660 18244 27169 18272
rect 26660 18232 26666 18244
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27338 18272 27344 18284
rect 27299 18244 27344 18272
rect 27157 18235 27215 18241
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 27540 18281 27568 18312
rect 27433 18275 27491 18281
rect 27433 18241 27445 18275
rect 27479 18241 27491 18275
rect 27433 18235 27491 18241
rect 27530 18275 27588 18281
rect 27530 18241 27542 18275
rect 27576 18241 27588 18275
rect 27530 18235 27588 18241
rect 25225 18207 25283 18213
rect 25225 18204 25237 18207
rect 24412 18176 24532 18204
rect 13538 18136 13544 18148
rect 12360 18108 13544 18136
rect 3602 18068 3608 18080
rect 2617 18040 3608 18068
rect 3602 18028 3608 18040
rect 3660 18028 3666 18080
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 8389 18071 8447 18077
rect 8389 18068 8401 18071
rect 8352 18040 8401 18068
rect 8352 18028 8358 18040
rect 8389 18037 8401 18040
rect 8435 18037 8447 18071
rect 8389 18031 8447 18037
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 11057 18071 11115 18077
rect 11057 18068 11069 18071
rect 10836 18040 11069 18068
rect 10836 18028 10842 18040
rect 11057 18037 11069 18040
rect 11103 18037 11115 18071
rect 11974 18068 11980 18080
rect 11935 18040 11980 18068
rect 11057 18031 11115 18037
rect 11974 18028 11980 18040
rect 12032 18028 12038 18080
rect 12360 18077 12388 18108
rect 13538 18096 13544 18108
rect 13596 18096 13602 18148
rect 12345 18071 12403 18077
rect 12345 18037 12357 18071
rect 12391 18037 12403 18071
rect 12345 18031 12403 18037
rect 12894 18028 12900 18080
rect 12952 18068 12958 18080
rect 12989 18071 13047 18077
rect 12989 18068 13001 18071
rect 12952 18040 13001 18068
rect 12952 18028 12958 18040
rect 12989 18037 13001 18040
rect 13035 18037 13047 18071
rect 14826 18068 14832 18080
rect 14787 18040 14832 18068
rect 12989 18031 13047 18037
rect 14826 18028 14832 18040
rect 14884 18028 14890 18080
rect 17865 18071 17923 18077
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 18230 18068 18236 18080
rect 17911 18040 18236 18068
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 19058 18028 19064 18080
rect 19116 18068 19122 18080
rect 19889 18071 19947 18077
rect 19889 18068 19901 18071
rect 19116 18040 19901 18068
rect 19116 18028 19122 18040
rect 19889 18037 19901 18040
rect 19935 18068 19947 18071
rect 20346 18068 20352 18080
rect 19935 18040 20352 18068
rect 19935 18037 19947 18040
rect 19889 18031 19947 18037
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 20622 18068 20628 18080
rect 20583 18040 20628 18068
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 24504 18068 24532 18176
rect 24688 18176 25237 18204
rect 24688 18145 24716 18176
rect 25225 18173 25237 18176
rect 25271 18173 25283 18207
rect 25225 18167 25283 18173
rect 27062 18164 27068 18216
rect 27120 18204 27126 18216
rect 27356 18204 27384 18232
rect 27120 18176 27384 18204
rect 27448 18204 27476 18235
rect 27448 18176 27844 18204
rect 27120 18164 27126 18176
rect 24673 18139 24731 18145
rect 24673 18105 24685 18139
rect 24719 18105 24731 18139
rect 27706 18136 27712 18148
rect 27667 18108 27712 18136
rect 24673 18099 24731 18105
rect 27706 18096 27712 18108
rect 27764 18096 27770 18148
rect 27816 18080 27844 18176
rect 25038 18068 25044 18080
rect 24504 18040 25044 18068
rect 25038 18028 25044 18040
rect 25096 18068 25102 18080
rect 26697 18071 26755 18077
rect 26697 18068 26709 18071
rect 25096 18040 26709 18068
rect 25096 18028 25102 18040
rect 26697 18037 26709 18040
rect 26743 18037 26755 18071
rect 26697 18031 26755 18037
rect 27798 18028 27804 18080
rect 27856 18068 27862 18080
rect 27893 18071 27951 18077
rect 27893 18068 27905 18071
rect 27856 18040 27905 18068
rect 27856 18028 27862 18040
rect 27893 18037 27905 18040
rect 27939 18037 27951 18071
rect 27893 18031 27951 18037
rect 1104 17978 29532 18000
rect 1104 17926 5688 17978
rect 5740 17926 5752 17978
rect 5804 17926 5816 17978
rect 5868 17926 5880 17978
rect 5932 17926 5944 17978
rect 5996 17926 15163 17978
rect 15215 17926 15227 17978
rect 15279 17926 15291 17978
rect 15343 17926 15355 17978
rect 15407 17926 15419 17978
rect 15471 17926 24639 17978
rect 24691 17926 24703 17978
rect 24755 17926 24767 17978
rect 24819 17926 24831 17978
rect 24883 17926 24895 17978
rect 24947 17926 29532 17978
rect 1104 17904 29532 17926
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 3878 17864 3884 17876
rect 3476 17836 3884 17864
rect 3476 17824 3482 17836
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4246 17864 4252 17876
rect 4120 17836 4252 17864
rect 4120 17824 4126 17836
rect 4246 17824 4252 17836
rect 4304 17824 4310 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7193 17867 7251 17873
rect 7193 17864 7205 17867
rect 6972 17836 7205 17864
rect 6972 17824 6978 17836
rect 7193 17833 7205 17836
rect 7239 17833 7251 17867
rect 7466 17864 7472 17876
rect 7427 17836 7472 17864
rect 7193 17827 7251 17833
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 12345 17867 12403 17873
rect 12345 17864 12357 17867
rect 11112 17836 12357 17864
rect 11112 17824 11118 17836
rect 12345 17833 12357 17836
rect 12391 17833 12403 17867
rect 12345 17827 12403 17833
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 24486 17864 24492 17876
rect 12492 17836 24492 17864
rect 12492 17824 12498 17836
rect 24486 17824 24492 17836
rect 24544 17824 24550 17876
rect 4080 17796 4108 17824
rect 3436 17768 4108 17796
rect 7837 17799 7895 17805
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 3234 17660 3240 17672
rect 3195 17632 3240 17660
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 3329 17663 3387 17669
rect 3329 17629 3341 17663
rect 3375 17660 3387 17663
rect 3436 17660 3464 17768
rect 7837 17765 7849 17799
rect 7883 17765 7895 17799
rect 12526 17796 12532 17808
rect 7837 17759 7895 17765
rect 8220 17768 12532 17796
rect 3513 17731 3571 17737
rect 3513 17697 3525 17731
rect 3559 17728 3571 17731
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 3559 17700 4077 17728
rect 3559 17697 3571 17700
rect 3513 17691 3571 17697
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 6454 17728 6460 17740
rect 6415 17700 6460 17728
rect 4065 17691 4123 17697
rect 6454 17688 6460 17700
rect 6512 17688 6518 17740
rect 6546 17688 6552 17740
rect 6604 17728 6610 17740
rect 7852 17728 7880 17759
rect 8220 17737 8248 17768
rect 12526 17756 12532 17768
rect 12584 17756 12590 17808
rect 19702 17756 19708 17808
rect 19760 17796 19766 17808
rect 20073 17799 20131 17805
rect 20073 17796 20085 17799
rect 19760 17768 20085 17796
rect 19760 17756 19766 17768
rect 20073 17765 20085 17768
rect 20119 17765 20131 17799
rect 21266 17796 21272 17808
rect 20073 17759 20131 17765
rect 20364 17768 21272 17796
rect 6604 17700 6649 17728
rect 7392 17700 7880 17728
rect 8205 17731 8263 17737
rect 6604 17688 6610 17700
rect 3602 17660 3608 17672
rect 3375 17632 3464 17660
rect 3563 17632 3608 17660
rect 3375 17629 3387 17632
rect 3329 17623 3387 17629
rect 3602 17620 3608 17632
rect 3660 17620 3666 17672
rect 3789 17663 3847 17669
rect 3789 17629 3801 17663
rect 3835 17629 3847 17663
rect 3970 17660 3976 17672
rect 3931 17632 3976 17660
rect 3789 17623 3847 17629
rect 1664 17595 1722 17601
rect 1664 17561 1676 17595
rect 1710 17592 1722 17595
rect 3053 17595 3111 17601
rect 3053 17592 3065 17595
rect 1710 17564 3065 17592
rect 1710 17561 1722 17564
rect 1664 17555 1722 17561
rect 3053 17561 3065 17564
rect 3099 17561 3111 17595
rect 3053 17555 3111 17561
rect 3252 17592 3280 17620
rect 3804 17592 3832 17623
rect 3970 17620 3976 17632
rect 4028 17620 4034 17672
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 4706 17660 4712 17672
rect 4479 17632 4712 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 7392 17669 7420 17700
rect 8205 17697 8217 17731
rect 8251 17697 8263 17731
rect 8205 17691 8263 17697
rect 11790 17688 11796 17740
rect 11848 17728 11854 17740
rect 12713 17731 12771 17737
rect 12713 17728 12725 17731
rect 11848 17700 12725 17728
rect 11848 17688 11854 17700
rect 12713 17697 12725 17700
rect 12759 17728 12771 17731
rect 14550 17728 14556 17740
rect 12759 17700 14556 17728
rect 12759 17697 12771 17700
rect 12713 17691 12771 17697
rect 14550 17688 14556 17700
rect 14608 17688 14614 17740
rect 14737 17731 14795 17737
rect 14737 17697 14749 17731
rect 14783 17728 14795 17731
rect 15654 17728 15660 17740
rect 14783 17700 15660 17728
rect 14783 17697 14795 17700
rect 14737 17691 14795 17697
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 16209 17731 16267 17737
rect 16209 17697 16221 17731
rect 16255 17728 16267 17731
rect 18138 17728 18144 17740
rect 16255 17700 18144 17728
rect 16255 17697 16267 17700
rect 16209 17691 16267 17697
rect 18138 17688 18144 17700
rect 18196 17688 18202 17740
rect 19610 17688 19616 17740
rect 19668 17728 19674 17740
rect 20162 17728 20168 17740
rect 19668 17700 20168 17728
rect 19668 17688 19674 17700
rect 20162 17688 20168 17700
rect 20220 17688 20226 17740
rect 7377 17663 7435 17669
rect 7377 17629 7389 17663
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 7558 17620 7564 17672
rect 7616 17660 7622 17672
rect 7653 17663 7711 17669
rect 7653 17660 7665 17663
rect 7616 17632 7665 17660
rect 7616 17620 7622 17632
rect 7653 17629 7665 17632
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17660 9551 17663
rect 9582 17660 9588 17672
rect 9539 17632 9588 17660
rect 9539 17629 9551 17632
rect 9493 17623 9551 17629
rect 9582 17620 9588 17632
rect 9640 17660 9646 17672
rect 9953 17663 10011 17669
rect 9953 17660 9965 17663
rect 9640 17632 9965 17660
rect 9640 17620 9646 17632
rect 9953 17629 9965 17632
rect 9999 17629 10011 17663
rect 12437 17663 12495 17669
rect 12437 17650 12449 17663
rect 12483 17650 12495 17663
rect 9953 17623 10011 17629
rect 3252 17564 3832 17592
rect 6365 17595 6423 17601
rect 2777 17527 2835 17533
rect 2777 17493 2789 17527
rect 2823 17524 2835 17527
rect 3252 17524 3280 17564
rect 6365 17561 6377 17595
rect 6411 17592 6423 17595
rect 8294 17592 8300 17604
rect 6411 17564 8300 17592
rect 6411 17561 6423 17564
rect 6365 17555 6423 17561
rect 8294 17552 8300 17564
rect 8352 17552 8358 17604
rect 8386 17552 8392 17604
rect 8444 17592 8450 17604
rect 12434 17598 12440 17650
rect 12492 17598 12498 17650
rect 12526 17619 12532 17671
rect 12584 17669 12590 17671
rect 12584 17663 12633 17669
rect 12584 17629 12587 17663
rect 12621 17660 12633 17663
rect 12806 17663 12864 17669
rect 12806 17660 12818 17663
rect 12621 17631 12664 17660
rect 12728 17632 12818 17660
rect 12621 17629 12633 17631
rect 12584 17623 12633 17629
rect 12584 17619 12590 17623
rect 12728 17604 12756 17632
rect 12806 17629 12818 17632
rect 12852 17629 12864 17663
rect 12986 17660 12992 17672
rect 12947 17632 12992 17660
rect 12806 17623 12864 17629
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13170 17660 13176 17672
rect 13127 17632 13176 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 13170 17620 13176 17632
rect 13228 17620 13234 17672
rect 13538 17620 13544 17672
rect 13596 17669 13602 17672
rect 13596 17663 13645 17669
rect 13596 17629 13599 17663
rect 13633 17629 13645 17663
rect 13817 17663 13875 17669
rect 13817 17660 13829 17663
rect 13596 17623 13645 17629
rect 13740 17632 13829 17660
rect 13596 17620 13602 17623
rect 13740 17604 13768 17632
rect 13817 17629 13829 17632
rect 13863 17629 13875 17663
rect 13817 17623 13875 17629
rect 13998 17620 14004 17672
rect 14056 17660 14062 17672
rect 14323 17663 14381 17669
rect 14323 17660 14335 17663
rect 14056 17632 14335 17660
rect 14056 17620 14062 17632
rect 14323 17629 14335 17632
rect 14369 17629 14381 17663
rect 14323 17623 14381 17629
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17660 14519 17663
rect 14918 17660 14924 17672
rect 14507 17632 14924 17660
rect 14507 17629 14519 17632
rect 14461 17623 14519 17629
rect 8444 17564 8489 17592
rect 8444 17552 8450 17564
rect 12710 17552 12716 17604
rect 12768 17552 12774 17604
rect 13722 17552 13728 17604
rect 13780 17552 13786 17604
rect 13909 17595 13967 17601
rect 13909 17561 13921 17595
rect 13955 17592 13967 17595
rect 14476 17592 14504 17623
rect 14918 17620 14924 17632
rect 14976 17620 14982 17672
rect 18230 17620 18236 17672
rect 18288 17660 18294 17672
rect 18325 17663 18383 17669
rect 18325 17660 18337 17663
rect 18288 17632 18337 17660
rect 18288 17620 18294 17632
rect 18325 17629 18337 17632
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 20252 17663 20310 17669
rect 20252 17629 20264 17663
rect 20298 17660 20310 17663
rect 20364 17660 20392 17768
rect 21266 17756 21272 17768
rect 21324 17756 21330 17808
rect 22741 17799 22799 17805
rect 22741 17765 22753 17799
rect 22787 17796 22799 17799
rect 23566 17796 23572 17808
rect 22787 17768 23572 17796
rect 22787 17765 22799 17768
rect 22741 17759 22799 17765
rect 23566 17756 23572 17768
rect 23624 17756 23630 17808
rect 27338 17796 27344 17808
rect 27299 17768 27344 17796
rect 27338 17756 27344 17768
rect 27396 17756 27402 17808
rect 22830 17728 22836 17740
rect 22204 17700 22836 17728
rect 20298 17632 20392 17660
rect 20625 17663 20683 17669
rect 20298 17629 20310 17632
rect 20252 17623 20310 17629
rect 20625 17629 20637 17663
rect 20671 17660 20683 17663
rect 20714 17660 20720 17672
rect 20671 17632 20720 17660
rect 20671 17629 20683 17632
rect 20625 17623 20683 17629
rect 20714 17620 20720 17632
rect 20772 17660 20778 17672
rect 20898 17660 20904 17672
rect 20772 17632 20904 17660
rect 20772 17620 20778 17632
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 22204 17669 22232 17700
rect 22830 17688 22836 17700
rect 22888 17688 22894 17740
rect 23658 17728 23664 17740
rect 23032 17700 23664 17728
rect 22189 17663 22247 17669
rect 22189 17629 22201 17663
rect 22235 17629 22247 17663
rect 22189 17623 22247 17629
rect 22609 17663 22667 17669
rect 22609 17629 22621 17663
rect 22655 17660 22667 17663
rect 23032 17660 23060 17700
rect 23658 17688 23664 17700
rect 23716 17688 23722 17740
rect 26418 17688 26424 17740
rect 26476 17728 26482 17740
rect 27430 17728 27436 17740
rect 26476 17700 27436 17728
rect 26476 17688 26482 17700
rect 22655 17632 23060 17660
rect 23109 17663 23167 17669
rect 22655 17629 22667 17632
rect 22609 17623 22667 17629
rect 23109 17629 23121 17663
rect 23155 17629 23167 17663
rect 23382 17660 23388 17672
rect 23343 17632 23388 17660
rect 23109 17623 23167 17629
rect 13955 17564 14504 17592
rect 13955 17561 13967 17564
rect 13909 17555 13967 17561
rect 14550 17552 14556 17604
rect 14608 17592 14614 17604
rect 14829 17595 14887 17601
rect 14829 17592 14841 17595
rect 14608 17564 14841 17592
rect 14608 17552 14614 17564
rect 14829 17561 14841 17564
rect 14875 17561 14887 17595
rect 14829 17555 14887 17561
rect 15286 17552 15292 17604
rect 15344 17592 15350 17604
rect 16485 17595 16543 17601
rect 16485 17592 16497 17595
rect 15344 17564 16497 17592
rect 15344 17552 15350 17564
rect 16485 17561 16497 17564
rect 16531 17561 16543 17595
rect 20349 17595 20407 17601
rect 20349 17592 20361 17595
rect 17710 17564 18184 17592
rect 16485 17555 16543 17561
rect 2823 17496 3280 17524
rect 5997 17527 6055 17533
rect 2823 17493 2835 17496
rect 2777 17487 2835 17493
rect 5997 17493 6009 17527
rect 6043 17524 6055 17527
rect 6086 17524 6092 17536
rect 6043 17496 6092 17524
rect 6043 17493 6055 17496
rect 5997 17487 6055 17493
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 9766 17524 9772 17536
rect 9727 17496 9772 17524
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 12158 17484 12164 17536
rect 12216 17524 12222 17536
rect 13265 17527 13323 17533
rect 13265 17524 13277 17527
rect 12216 17496 13277 17524
rect 12216 17484 12222 17496
rect 13265 17493 13277 17496
rect 13311 17524 13323 17527
rect 13998 17524 14004 17536
rect 13311 17496 14004 17524
rect 13311 17493 13323 17496
rect 13265 17487 13323 17493
rect 13998 17484 14004 17496
rect 14056 17484 14062 17536
rect 14182 17524 14188 17536
rect 14143 17496 14188 17524
rect 14182 17484 14188 17496
rect 14240 17484 14246 17536
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 16666 17524 16672 17536
rect 14700 17496 16672 17524
rect 14700 17484 14706 17496
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 17954 17524 17960 17536
rect 17915 17496 17960 17524
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 18156 17533 18184 17564
rect 19812 17564 20361 17592
rect 18141 17527 18199 17533
rect 18141 17493 18153 17527
rect 18187 17493 18199 17527
rect 18141 17487 18199 17493
rect 18230 17484 18236 17536
rect 18288 17524 18294 17536
rect 19812 17533 19840 17564
rect 20349 17561 20361 17564
rect 20395 17561 20407 17595
rect 20349 17555 20407 17561
rect 20441 17595 20499 17601
rect 20441 17561 20453 17595
rect 20487 17561 20499 17595
rect 22370 17592 22376 17604
rect 22331 17564 22376 17592
rect 20441 17555 20499 17561
rect 19797 17527 19855 17533
rect 19797 17524 19809 17527
rect 18288 17496 19809 17524
rect 18288 17484 18294 17496
rect 19797 17493 19809 17496
rect 19843 17493 19855 17527
rect 19797 17487 19855 17493
rect 20254 17484 20260 17536
rect 20312 17524 20318 17536
rect 20456 17524 20484 17555
rect 22370 17552 22376 17564
rect 22428 17552 22434 17604
rect 22465 17595 22523 17601
rect 22465 17561 22477 17595
rect 22511 17561 22523 17595
rect 23124 17592 23152 17623
rect 23382 17620 23388 17632
rect 23440 17620 23446 17672
rect 24394 17620 24400 17672
rect 24452 17660 24458 17672
rect 24673 17663 24731 17669
rect 24673 17660 24685 17663
rect 24452 17632 24685 17660
rect 24452 17620 24458 17632
rect 24673 17629 24685 17632
rect 24719 17629 24731 17663
rect 25317 17663 25375 17669
rect 25317 17660 25329 17663
rect 24673 17623 24731 17629
rect 24872 17632 25329 17660
rect 23474 17592 23480 17604
rect 23124 17564 23480 17592
rect 22465 17555 22523 17561
rect 20312 17496 20484 17524
rect 20312 17484 20318 17496
rect 20622 17484 20628 17536
rect 20680 17524 20686 17536
rect 20717 17527 20775 17533
rect 20717 17524 20729 17527
rect 20680 17496 20729 17524
rect 20680 17484 20686 17496
rect 20717 17493 20729 17496
rect 20763 17493 20775 17527
rect 20898 17524 20904 17536
rect 20859 17496 20904 17524
rect 20717 17487 20775 17493
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 22094 17484 22100 17536
rect 22152 17524 22158 17536
rect 22480 17524 22508 17555
rect 23474 17552 23480 17564
rect 23532 17592 23538 17604
rect 23532 17564 23612 17592
rect 23532 17552 23538 17564
rect 23290 17524 23296 17536
rect 22152 17496 22508 17524
rect 23251 17496 23296 17524
rect 22152 17484 22158 17496
rect 23290 17484 23296 17496
rect 23348 17484 23354 17536
rect 23584 17533 23612 17564
rect 23569 17527 23627 17533
rect 23569 17493 23581 17527
rect 23615 17524 23627 17527
rect 24412 17524 24440 17620
rect 24872 17533 24900 17632
rect 25317 17629 25329 17632
rect 25363 17629 25375 17663
rect 25317 17623 25375 17629
rect 26602 17620 26608 17672
rect 26660 17660 26666 17672
rect 26988 17669 27016 17700
rect 27430 17688 27436 17700
rect 27488 17688 27494 17740
rect 27246 17669 27252 17672
rect 26789 17663 26847 17669
rect 26789 17660 26801 17663
rect 26660 17632 26801 17660
rect 26660 17620 26666 17632
rect 26789 17629 26801 17632
rect 26835 17629 26847 17663
rect 26789 17623 26847 17629
rect 26973 17663 27031 17669
rect 26973 17629 26985 17663
rect 27019 17629 27031 17663
rect 26973 17623 27031 17629
rect 27209 17663 27252 17669
rect 27209 17629 27221 17663
rect 27209 17623 27252 17629
rect 27246 17620 27252 17623
rect 27304 17620 27310 17672
rect 27065 17595 27123 17601
rect 27065 17561 27077 17595
rect 27111 17561 27123 17595
rect 27065 17555 27123 17561
rect 23615 17496 24440 17524
rect 24857 17527 24915 17533
rect 23615 17493 23627 17496
rect 23569 17487 23627 17493
rect 24857 17493 24869 17527
rect 24903 17493 24915 17527
rect 25038 17524 25044 17536
rect 24999 17496 25044 17524
rect 24857 17487 24915 17493
rect 25038 17484 25044 17496
rect 25096 17484 25102 17536
rect 25133 17527 25191 17533
rect 25133 17493 25145 17527
rect 25179 17524 25191 17527
rect 25222 17524 25228 17536
rect 25179 17496 25228 17524
rect 25179 17493 25191 17496
rect 25133 17487 25191 17493
rect 25222 17484 25228 17496
rect 25280 17484 25286 17536
rect 27080 17524 27108 17555
rect 27617 17527 27675 17533
rect 27617 17524 27629 17527
rect 27080 17496 27629 17524
rect 27617 17493 27629 17496
rect 27663 17524 27675 17527
rect 29641 17527 29699 17533
rect 29641 17524 29653 17527
rect 27663 17496 29653 17524
rect 27663 17493 27675 17496
rect 27617 17487 27675 17493
rect 29641 17493 29653 17496
rect 29687 17493 29699 17527
rect 29641 17487 29699 17493
rect 1104 17434 29532 17456
rect 1104 17382 10425 17434
rect 10477 17382 10489 17434
rect 10541 17382 10553 17434
rect 10605 17382 10617 17434
rect 10669 17382 10681 17434
rect 10733 17382 19901 17434
rect 19953 17382 19965 17434
rect 20017 17382 20029 17434
rect 20081 17382 20093 17434
rect 20145 17382 20157 17434
rect 20209 17382 29532 17434
rect 1104 17360 29532 17382
rect 7653 17323 7711 17329
rect 7653 17289 7665 17323
rect 7699 17289 7711 17323
rect 7653 17283 7711 17289
rect 12897 17323 12955 17329
rect 12897 17289 12909 17323
rect 12943 17320 12955 17323
rect 12986 17320 12992 17332
rect 12943 17292 12992 17320
rect 12943 17289 12955 17292
rect 12897 17283 12955 17289
rect 4890 17252 4896 17264
rect 4724 17224 4896 17252
rect 4361 17187 4419 17193
rect 4361 17153 4373 17187
rect 4407 17184 4419 17187
rect 4522 17184 4528 17196
rect 4407 17156 4528 17184
rect 4407 17153 4419 17156
rect 4361 17147 4419 17153
rect 4522 17144 4528 17156
rect 4580 17144 4586 17196
rect 4724 17193 4752 17224
rect 4890 17212 4896 17224
rect 4948 17252 4954 17264
rect 6638 17252 6644 17264
rect 4948 17224 6644 17252
rect 4948 17212 4954 17224
rect 6638 17212 6644 17224
rect 6696 17212 6702 17264
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17184 4675 17187
rect 4709 17187 4767 17193
rect 4709 17184 4721 17187
rect 4663 17156 4721 17184
rect 4663 17153 4675 17156
rect 4617 17147 4675 17153
rect 4709 17153 4721 17156
rect 4755 17153 4767 17187
rect 4709 17147 4767 17153
rect 4976 17187 5034 17193
rect 4976 17153 4988 17187
rect 5022 17184 5034 17187
rect 5350 17184 5356 17196
rect 5022 17156 5356 17184
rect 5022 17153 5034 17156
rect 4976 17147 5034 17153
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17184 7527 17187
rect 7558 17184 7564 17196
rect 7515 17156 7564 17184
rect 7515 17153 7527 17156
rect 7469 17147 7527 17153
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 7668 17184 7696 17283
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 13078 17280 13084 17332
rect 13136 17320 13142 17332
rect 13633 17323 13691 17329
rect 13633 17320 13645 17323
rect 13136 17292 13645 17320
rect 13136 17280 13142 17292
rect 13633 17289 13645 17292
rect 13679 17289 13691 17323
rect 13633 17283 13691 17289
rect 14936 17292 15884 17320
rect 9950 17212 9956 17264
rect 10008 17212 10014 17264
rect 11977 17255 12035 17261
rect 11977 17221 11989 17255
rect 12023 17252 12035 17255
rect 14274 17252 14280 17264
rect 12023 17224 14280 17252
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 7837 17187 7895 17193
rect 7837 17184 7849 17187
rect 7668 17156 7849 17184
rect 7837 17153 7849 17156
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9033 17187 9091 17193
rect 9033 17184 9045 17187
rect 8996 17156 9045 17184
rect 8996 17144 9002 17156
rect 9033 17153 9045 17156
rect 9079 17153 9091 17187
rect 9033 17147 9091 17153
rect 12066 17144 12072 17196
rect 12124 17184 12130 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12124 17156 12449 17184
rect 12124 17144 12130 17156
rect 12437 17153 12449 17156
rect 12483 17184 12495 17187
rect 12710 17184 12716 17196
rect 12483 17156 12716 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 12986 17184 12992 17196
rect 12820 17156 12992 17184
rect 9309 17119 9367 17125
rect 9309 17085 9321 17119
rect 9355 17116 9367 17119
rect 10962 17116 10968 17128
rect 9355 17088 10968 17116
rect 9355 17085 9367 17088
rect 9309 17079 9367 17085
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 11885 17119 11943 17125
rect 11885 17085 11897 17119
rect 11931 17085 11943 17119
rect 12158 17116 12164 17128
rect 12119 17088 12164 17116
rect 11885 17079 11943 17085
rect 11900 17048 11928 17079
rect 12158 17076 12164 17088
rect 12216 17076 12222 17128
rect 12820 17048 12848 17156
rect 12986 17144 12992 17156
rect 13044 17184 13050 17196
rect 13556 17193 13584 17224
rect 14274 17212 14280 17224
rect 14332 17252 14338 17264
rect 14645 17255 14703 17261
rect 14645 17252 14657 17255
rect 14332 17224 14657 17252
rect 14332 17212 14338 17224
rect 14645 17221 14657 17224
rect 14691 17252 14703 17255
rect 14691 17224 14872 17252
rect 14691 17221 14703 17224
rect 14645 17215 14703 17221
rect 13265 17187 13323 17193
rect 13265 17184 13277 17187
rect 13044 17156 13277 17184
rect 13044 17144 13050 17156
rect 13265 17153 13277 17156
rect 13311 17153 13323 17187
rect 13265 17147 13323 17153
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17153 13599 17187
rect 13814 17184 13820 17196
rect 13775 17156 13820 17184
rect 13541 17147 13599 17153
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 14844 17193 14872 17224
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17184 14519 17187
rect 14737 17187 14795 17193
rect 14507 17156 14596 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 13078 17116 13084 17128
rect 13039 17088 13084 17116
rect 13078 17076 13084 17088
rect 13136 17076 13142 17128
rect 13173 17119 13231 17125
rect 13173 17085 13185 17119
rect 13219 17085 13231 17119
rect 13173 17079 13231 17085
rect 13357 17119 13415 17125
rect 13357 17085 13369 17119
rect 13403 17085 13415 17119
rect 13357 17079 13415 17085
rect 11900 17020 12848 17048
rect 3237 16983 3295 16989
rect 3237 16949 3249 16983
rect 3283 16980 3295 16983
rect 4338 16980 4344 16992
rect 3283 16952 4344 16980
rect 3283 16949 3295 16952
rect 3237 16943 3295 16949
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 6089 16983 6147 16989
rect 6089 16949 6101 16983
rect 6135 16980 6147 16983
rect 6454 16980 6460 16992
rect 6135 16952 6460 16980
rect 6135 16949 6147 16952
rect 6089 16943 6147 16949
rect 6454 16940 6460 16952
rect 6512 16940 6518 16992
rect 8021 16983 8079 16989
rect 8021 16949 8033 16983
rect 8067 16980 8079 16983
rect 8294 16980 8300 16992
rect 8067 16952 8300 16980
rect 8067 16949 8079 16952
rect 8021 16943 8079 16949
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 10318 16940 10324 16992
rect 10376 16980 10382 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 10376 16952 10793 16980
rect 10376 16940 10382 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 10781 16943 10839 16949
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 11204 16952 11713 16980
rect 11204 16940 11210 16952
rect 11701 16949 11713 16952
rect 11747 16949 11759 16983
rect 11701 16943 11759 16949
rect 11790 16940 11796 16992
rect 11848 16980 11854 16992
rect 12253 16983 12311 16989
rect 12253 16980 12265 16983
rect 11848 16952 12265 16980
rect 11848 16940 11854 16952
rect 12253 16949 12265 16952
rect 12299 16949 12311 16983
rect 13188 16980 13216 17079
rect 13372 17048 13400 17079
rect 13630 17048 13636 17060
rect 13372 17020 13636 17048
rect 13630 17008 13636 17020
rect 13688 17048 13694 17060
rect 14277 17051 14335 17057
rect 14277 17048 14289 17051
rect 13688 17020 14289 17048
rect 13688 17008 13694 17020
rect 14277 17017 14289 17020
rect 14323 17017 14335 17051
rect 14568 17048 14596 17156
rect 14737 17153 14749 17187
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 14829 17187 14887 17193
rect 14829 17153 14841 17187
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 14642 17076 14648 17128
rect 14700 17116 14706 17128
rect 14752 17116 14780 17147
rect 14936 17116 14964 17292
rect 15856 17252 15884 17292
rect 15930 17280 15936 17332
rect 15988 17320 15994 17332
rect 16301 17323 16359 17329
rect 16301 17320 16313 17323
rect 15988 17292 16313 17320
rect 15988 17280 15994 17292
rect 16301 17289 16313 17292
rect 16347 17289 16359 17323
rect 16666 17320 16672 17332
rect 16627 17292 16672 17320
rect 16301 17283 16359 17289
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 18322 17280 18328 17332
rect 18380 17320 18386 17332
rect 20622 17320 20628 17332
rect 18380 17292 20628 17320
rect 18380 17280 18386 17292
rect 17954 17252 17960 17264
rect 15120 17224 15792 17252
rect 15856 17224 17960 17252
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 15120 17193 15148 17224
rect 15105 17187 15163 17193
rect 15105 17184 15117 17187
rect 15068 17156 15117 17184
rect 15068 17144 15074 17156
rect 15105 17153 15117 17156
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17184 15439 17187
rect 15470 17184 15476 17196
rect 15427 17156 15476 17184
rect 15427 17153 15439 17156
rect 15381 17147 15439 17153
rect 15470 17144 15476 17156
rect 15528 17144 15534 17196
rect 15565 17187 15623 17193
rect 15565 17153 15577 17187
rect 15611 17184 15623 17187
rect 15654 17184 15660 17196
rect 15611 17156 15660 17184
rect 15611 17153 15623 17156
rect 15565 17147 15623 17153
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 15764 17193 15792 17224
rect 16040 17193 16068 17224
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 19242 17212 19248 17264
rect 19300 17212 19306 17264
rect 19702 17252 19708 17264
rect 19663 17224 19708 17252
rect 19702 17212 19708 17224
rect 19760 17212 19766 17264
rect 19794 17212 19800 17264
rect 19852 17252 19858 17264
rect 19852 17224 20024 17252
rect 19852 17212 19858 17224
rect 15749 17187 15807 17193
rect 15749 17153 15761 17187
rect 15795 17153 15807 17187
rect 15749 17147 15807 17153
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17153 16083 17187
rect 16206 17184 16212 17196
rect 16167 17156 16212 17184
rect 16025 17147 16083 17153
rect 16206 17144 16212 17156
rect 16264 17184 16270 17196
rect 19996 17193 20024 17224
rect 20088 17193 20116 17292
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 21910 17280 21916 17332
rect 21968 17320 21974 17332
rect 22646 17320 22652 17332
rect 21968 17292 22652 17320
rect 21968 17280 21974 17292
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 23937 17323 23995 17329
rect 23937 17320 23949 17323
rect 23124 17292 23949 17320
rect 20901 17255 20959 17261
rect 20901 17221 20913 17255
rect 20947 17252 20959 17255
rect 21634 17252 21640 17264
rect 20947 17224 21640 17252
rect 20947 17221 20959 17224
rect 20901 17215 20959 17221
rect 21634 17212 21640 17224
rect 21692 17212 21698 17264
rect 23124 17238 23152 17292
rect 23937 17289 23949 17292
rect 23983 17289 23995 17323
rect 24486 17320 24492 17332
rect 24447 17292 24492 17320
rect 23937 17283 23995 17289
rect 24486 17280 24492 17292
rect 24544 17280 24550 17332
rect 23290 17212 23296 17264
rect 23348 17252 23354 17264
rect 23348 17224 24164 17252
rect 23348 17212 23354 17224
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16264 17156 16865 17184
rect 16264 17144 16270 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17153 20131 17187
rect 20441 17187 20499 17193
rect 20441 17184 20453 17187
rect 20073 17147 20131 17153
rect 20272 17156 20453 17184
rect 15286 17116 15292 17128
rect 14700 17088 14964 17116
rect 15247 17088 15292 17116
rect 14700 17076 14706 17088
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 16114 17116 16120 17128
rect 16075 17088 16120 17116
rect 16114 17076 16120 17088
rect 16172 17076 16178 17128
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19610 17116 19616 17128
rect 19392 17088 19616 17116
rect 19392 17076 19398 17088
rect 19610 17076 19616 17088
rect 19668 17076 19674 17128
rect 14826 17048 14832 17060
rect 14568 17020 14832 17048
rect 14277 17011 14335 17017
rect 14826 17008 14832 17020
rect 14884 17048 14890 17060
rect 15562 17048 15568 17060
rect 14884 17020 15568 17048
rect 14884 17008 14890 17020
rect 15562 17008 15568 17020
rect 15620 17008 15626 17060
rect 20272 17057 20300 17156
rect 20441 17153 20453 17156
rect 20487 17153 20499 17187
rect 20714 17184 20720 17196
rect 20675 17156 20720 17184
rect 20441 17147 20499 17153
rect 20714 17144 20720 17156
rect 20772 17144 20778 17196
rect 20990 17144 20996 17196
rect 21048 17184 21054 17196
rect 21137 17187 21195 17193
rect 21048 17156 21093 17184
rect 21048 17144 21054 17156
rect 21137 17153 21149 17187
rect 21183 17184 21195 17187
rect 21266 17184 21272 17196
rect 21183 17156 21272 17184
rect 21183 17153 21195 17156
rect 21137 17147 21195 17153
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 24136 17193 24164 17224
rect 25222 17212 25228 17264
rect 25280 17212 25286 17264
rect 27249 17255 27307 17261
rect 27249 17221 27261 17255
rect 27295 17252 27307 17255
rect 27338 17252 27344 17264
rect 27295 17224 27344 17252
rect 27295 17221 27307 17224
rect 27249 17215 27307 17221
rect 27338 17212 27344 17224
rect 27396 17212 27402 17264
rect 27982 17212 27988 17264
rect 28040 17212 28046 17264
rect 24121 17187 24179 17193
rect 24121 17153 24133 17187
rect 24167 17153 24179 17187
rect 24121 17147 24179 17153
rect 23566 17116 23572 17128
rect 23527 17088 23572 17116
rect 23566 17076 23572 17088
rect 23624 17076 23630 17128
rect 23845 17119 23903 17125
rect 23845 17085 23857 17119
rect 23891 17085 23903 17119
rect 25958 17116 25964 17128
rect 25919 17088 25964 17116
rect 23845 17079 23903 17085
rect 20257 17051 20315 17057
rect 20257 17017 20269 17051
rect 20303 17017 20315 17051
rect 20257 17011 20315 17017
rect 14642 16980 14648 16992
rect 13188 16952 14648 16980
rect 12253 16943 12311 16949
rect 14642 16940 14648 16952
rect 14700 16940 14706 16992
rect 18138 16940 18144 16992
rect 18196 16980 18202 16992
rect 18233 16983 18291 16989
rect 18233 16980 18245 16983
rect 18196 16952 18245 16980
rect 18196 16940 18202 16952
rect 18233 16949 18245 16952
rect 18279 16949 18291 16983
rect 18233 16943 18291 16949
rect 20530 16940 20536 16992
rect 20588 16980 20594 16992
rect 20625 16983 20683 16989
rect 20625 16980 20637 16983
rect 20588 16952 20637 16980
rect 20588 16940 20594 16952
rect 20625 16949 20637 16952
rect 20671 16949 20683 16983
rect 20625 16943 20683 16949
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 21542 16980 21548 16992
rect 21315 16952 21548 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21542 16940 21548 16952
rect 21600 16940 21606 16992
rect 22094 16940 22100 16992
rect 22152 16980 22158 16992
rect 22152 16952 22197 16980
rect 22152 16940 22158 16952
rect 22554 16940 22560 16992
rect 22612 16980 22618 16992
rect 23860 16980 23888 17079
rect 25958 17076 25964 17088
rect 26016 17076 26022 17128
rect 26234 17116 26240 17128
rect 26195 17088 26240 17116
rect 26234 17076 26240 17088
rect 26292 17116 26298 17128
rect 26973 17119 27031 17125
rect 26973 17116 26985 17119
rect 26292 17088 26985 17116
rect 26292 17076 26298 17088
rect 26973 17085 26985 17088
rect 27019 17085 27031 17119
rect 26973 17079 27031 17085
rect 22612 16952 23888 16980
rect 22612 16940 22618 16952
rect 24394 16940 24400 16992
rect 24452 16980 24458 16992
rect 26326 16980 26332 16992
rect 24452 16952 26332 16980
rect 24452 16940 24458 16952
rect 26326 16940 26332 16952
rect 26384 16940 26390 16992
rect 28721 16983 28779 16989
rect 28721 16949 28733 16983
rect 28767 16980 28779 16983
rect 29641 16983 29699 16989
rect 29641 16980 29653 16983
rect 28767 16952 29653 16980
rect 28767 16949 28779 16952
rect 28721 16943 28779 16949
rect 29641 16949 29653 16952
rect 29687 16949 29699 16983
rect 29641 16943 29699 16949
rect 1104 16890 29532 16912
rect 1104 16838 5688 16890
rect 5740 16838 5752 16890
rect 5804 16838 5816 16890
rect 5868 16838 5880 16890
rect 5932 16838 5944 16890
rect 5996 16838 15163 16890
rect 15215 16838 15227 16890
rect 15279 16838 15291 16890
rect 15343 16838 15355 16890
rect 15407 16838 15419 16890
rect 15471 16838 24639 16890
rect 24691 16838 24703 16890
rect 24755 16838 24767 16890
rect 24819 16838 24831 16890
rect 24883 16838 24895 16890
rect 24947 16838 29532 16890
rect 1104 16816 29532 16838
rect 4522 16736 4528 16788
rect 4580 16776 4586 16788
rect 4617 16779 4675 16785
rect 4617 16776 4629 16779
rect 4580 16748 4629 16776
rect 4580 16736 4586 16748
rect 4617 16745 4629 16748
rect 4663 16745 4675 16779
rect 5350 16776 5356 16788
rect 5311 16748 5356 16776
rect 4617 16739 4675 16745
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 5813 16779 5871 16785
rect 5813 16776 5825 16779
rect 5592 16748 5825 16776
rect 5592 16736 5598 16748
rect 5813 16745 5825 16748
rect 5859 16745 5871 16779
rect 5813 16739 5871 16745
rect 6638 16736 6644 16788
rect 6696 16776 6702 16788
rect 9950 16776 9956 16788
rect 6696 16748 6960 16776
rect 9911 16748 9956 16776
rect 6696 16736 6702 16748
rect 4985 16711 5043 16717
rect 4985 16677 4997 16711
rect 5031 16708 5043 16711
rect 5552 16708 5580 16736
rect 5031 16680 5580 16708
rect 5644 16680 6500 16708
rect 5031 16677 5043 16680
rect 4985 16671 5043 16677
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 5000 16640 5028 16671
rect 5644 16640 5672 16680
rect 6472 16652 6500 16680
rect 4724 16612 5028 16640
rect 5552 16612 5672 16640
rect 5905 16643 5963 16649
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 3234 16572 3240 16584
rect 3007 16544 3240 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 3234 16532 3240 16544
rect 3292 16572 3298 16584
rect 3694 16572 3700 16584
rect 3292 16544 3700 16572
rect 3292 16532 3298 16544
rect 3694 16532 3700 16544
rect 3752 16532 3758 16584
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16572 4123 16575
rect 4154 16572 4160 16584
rect 4111 16544 4160 16572
rect 4111 16541 4123 16544
rect 4065 16535 4123 16541
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 4338 16572 4344 16584
rect 4299 16544 4344 16572
rect 4338 16532 4344 16544
rect 4396 16532 4402 16584
rect 4485 16575 4543 16581
rect 4485 16541 4497 16575
rect 4531 16572 4543 16575
rect 4724 16572 4752 16612
rect 5552 16581 5580 16612
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 6086 16640 6092 16652
rect 5951 16612 6092 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 6454 16640 6460 16652
rect 6415 16612 6460 16640
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 6932 16649 6960 16748
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 11701 16779 11759 16785
rect 11701 16745 11713 16779
rect 11747 16776 11759 16779
rect 11974 16776 11980 16788
rect 11747 16748 11980 16776
rect 11747 16745 11759 16748
rect 11701 16739 11759 16745
rect 11974 16736 11980 16748
rect 12032 16736 12038 16788
rect 12066 16736 12072 16788
rect 12124 16776 12130 16788
rect 15473 16779 15531 16785
rect 15473 16776 15485 16779
rect 12124 16748 12169 16776
rect 12406 16748 15485 16776
rect 12124 16736 12130 16748
rect 9858 16668 9864 16720
rect 9916 16708 9922 16720
rect 12406 16708 12434 16748
rect 15473 16745 15485 16748
rect 15519 16776 15531 16779
rect 19334 16776 19340 16788
rect 15519 16748 19340 16776
rect 15519 16745 15531 16748
rect 15473 16739 15531 16745
rect 19334 16736 19340 16748
rect 19392 16736 19398 16788
rect 21726 16736 21732 16788
rect 21784 16776 21790 16788
rect 25041 16779 25099 16785
rect 21784 16748 24992 16776
rect 21784 16736 21790 16748
rect 9916 16680 12434 16708
rect 9916 16668 9922 16680
rect 12526 16668 12532 16720
rect 12584 16708 12590 16720
rect 13354 16708 13360 16720
rect 12584 16680 13360 16708
rect 12584 16668 12590 16680
rect 13354 16668 13360 16680
rect 13412 16668 13418 16720
rect 18322 16668 18328 16720
rect 18380 16708 18386 16720
rect 18601 16711 18659 16717
rect 18601 16708 18613 16711
rect 18380 16680 18613 16708
rect 18380 16668 18386 16680
rect 18601 16677 18613 16680
rect 18647 16677 18659 16711
rect 19242 16708 19248 16720
rect 19203 16680 19248 16708
rect 18601 16671 18659 16677
rect 6917 16643 6975 16649
rect 6604 16612 6649 16640
rect 6604 16600 6610 16612
rect 6917 16609 6929 16643
rect 6963 16609 6975 16643
rect 10962 16640 10968 16652
rect 10923 16612 10968 16640
rect 6917 16603 6975 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 11609 16643 11667 16649
rect 11609 16640 11621 16643
rect 11348 16612 11621 16640
rect 11348 16584 11376 16612
rect 11609 16609 11621 16612
rect 11655 16609 11667 16643
rect 11609 16603 11667 16609
rect 12161 16643 12219 16649
rect 12161 16609 12173 16643
rect 12207 16640 12219 16643
rect 12434 16640 12440 16652
rect 12207 16612 12440 16640
rect 12207 16609 12219 16612
rect 12161 16603 12219 16609
rect 12434 16600 12440 16612
rect 12492 16640 12498 16652
rect 12710 16640 12716 16652
rect 12492 16612 12716 16640
rect 12492 16600 12498 16612
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 16816 16612 17264 16640
rect 16816 16600 16822 16612
rect 4531 16544 4752 16572
rect 4801 16575 4859 16581
rect 4531 16541 4543 16544
rect 4485 16535 4543 16541
rect 4801 16541 4813 16575
rect 4847 16541 4859 16575
rect 4801 16535 4859 16541
rect 5537 16575 5595 16581
rect 5537 16541 5549 16575
rect 5583 16541 5595 16575
rect 5537 16535 5595 16541
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16541 5687 16575
rect 5629 16535 5687 16541
rect 1664 16507 1722 16513
rect 1664 16473 1676 16507
rect 1710 16504 1722 16507
rect 2314 16504 2320 16516
rect 1710 16476 2320 16504
rect 1710 16473 1722 16476
rect 1664 16467 1722 16473
rect 2314 16464 2320 16476
rect 2372 16464 2378 16516
rect 3145 16507 3203 16513
rect 3145 16473 3157 16507
rect 3191 16473 3203 16507
rect 3145 16467 3203 16473
rect 3329 16507 3387 16513
rect 3329 16473 3341 16507
rect 3375 16504 3387 16507
rect 3970 16504 3976 16516
rect 3375 16476 3976 16504
rect 3375 16473 3387 16476
rect 3329 16467 3387 16473
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 3160 16436 3188 16467
rect 3970 16464 3976 16476
rect 4028 16464 4034 16516
rect 4246 16504 4252 16516
rect 4207 16476 4252 16504
rect 4246 16464 4252 16476
rect 4304 16464 4310 16516
rect 4614 16464 4620 16516
rect 4672 16504 4678 16516
rect 4816 16504 4844 16535
rect 4672 16476 4844 16504
rect 4672 16464 4678 16476
rect 5074 16464 5080 16516
rect 5132 16504 5138 16516
rect 5644 16504 5672 16535
rect 8294 16532 8300 16584
rect 8352 16532 8358 16584
rect 9766 16572 9772 16584
rect 9727 16544 9772 16572
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 10689 16575 10747 16581
rect 10689 16541 10701 16575
rect 10735 16572 10747 16575
rect 10778 16572 10784 16584
rect 10735 16544 10784 16572
rect 10735 16541 10747 16544
rect 10689 16535 10747 16541
rect 10778 16532 10784 16544
rect 10836 16532 10842 16584
rect 10873 16575 10931 16581
rect 10873 16541 10885 16575
rect 10919 16541 10931 16575
rect 11146 16572 11152 16584
rect 11107 16544 11152 16572
rect 10873 16535 10931 16541
rect 5132 16476 5672 16504
rect 6365 16507 6423 16513
rect 5132 16464 5138 16476
rect 6365 16473 6377 16507
rect 6411 16504 6423 16507
rect 7190 16504 7196 16516
rect 6411 16476 7052 16504
rect 7151 16476 7196 16504
rect 6411 16473 6423 16476
rect 6365 16467 6423 16473
rect 2832 16408 3188 16436
rect 2832 16396 2838 16408
rect 5350 16396 5356 16448
rect 5408 16436 5414 16448
rect 5997 16439 6055 16445
rect 5997 16436 6009 16439
rect 5408 16408 6009 16436
rect 5408 16396 5414 16408
rect 5997 16405 6009 16408
rect 6043 16405 6055 16439
rect 7024 16436 7052 16476
rect 7190 16464 7196 16476
rect 7248 16464 7254 16516
rect 10888 16504 10916 16535
rect 11146 16532 11152 16544
rect 11204 16532 11210 16584
rect 11330 16572 11336 16584
rect 11291 16544 11336 16572
rect 11330 16532 11336 16544
rect 11388 16532 11394 16584
rect 11514 16572 11520 16584
rect 11475 16544 11520 16572
rect 11514 16532 11520 16544
rect 11572 16572 11578 16584
rect 11882 16572 11888 16584
rect 11572 16544 11888 16572
rect 11572 16532 11578 16544
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 11974 16532 11980 16584
rect 12032 16572 12038 16584
rect 12069 16575 12127 16581
rect 12069 16572 12081 16575
rect 12032 16544 12081 16572
rect 12032 16532 12038 16544
rect 12069 16541 12081 16544
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16572 12679 16575
rect 13814 16572 13820 16584
rect 12667 16544 13820 16572
rect 12667 16541 12679 16544
rect 12621 16535 12679 16541
rect 13814 16532 13820 16544
rect 13872 16532 13878 16584
rect 16574 16532 16580 16584
rect 16632 16572 16638 16584
rect 17236 16581 17264 16612
rect 17129 16575 17187 16581
rect 17129 16572 17141 16575
rect 16632 16544 17141 16572
rect 16632 16532 16638 16544
rect 17129 16541 17141 16544
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16572 17279 16575
rect 17770 16572 17776 16584
rect 17267 16544 17776 16572
rect 17267 16541 17279 16544
rect 17221 16535 17279 16541
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 18616 16572 18644 16671
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 24486 16668 24492 16720
rect 24544 16668 24550 16720
rect 24964 16708 24992 16748
rect 25041 16745 25053 16779
rect 25087 16776 25099 16779
rect 25958 16776 25964 16788
rect 25087 16748 25964 16776
rect 25087 16745 25099 16748
rect 25041 16739 25099 16745
rect 25958 16736 25964 16748
rect 26016 16736 26022 16788
rect 27982 16736 27988 16788
rect 28040 16776 28046 16788
rect 28077 16779 28135 16785
rect 28077 16776 28089 16779
rect 28040 16748 28089 16776
rect 28040 16736 28046 16748
rect 28077 16745 28089 16748
rect 28123 16745 28135 16779
rect 28077 16739 28135 16745
rect 25498 16708 25504 16720
rect 24964 16680 25504 16708
rect 25498 16668 25504 16680
rect 25556 16668 25562 16720
rect 21542 16640 21548 16652
rect 21503 16612 21548 16640
rect 21542 16600 21548 16612
rect 21600 16600 21606 16652
rect 21821 16643 21879 16649
rect 21821 16609 21833 16643
rect 21867 16640 21879 16643
rect 22646 16640 22652 16652
rect 21867 16612 22652 16640
rect 21867 16609 21879 16612
rect 21821 16603 21879 16609
rect 22646 16600 22652 16612
rect 22704 16600 22710 16652
rect 24504 16640 24532 16668
rect 25225 16643 25283 16649
rect 25225 16640 25237 16643
rect 24504 16612 25237 16640
rect 18785 16575 18843 16581
rect 18785 16572 18797 16575
rect 18616 16544 18797 16572
rect 18785 16541 18797 16544
rect 18831 16541 18843 16575
rect 19429 16575 19487 16581
rect 19429 16572 19441 16575
rect 18785 16535 18843 16541
rect 18984 16544 19441 16572
rect 11238 16504 11244 16516
rect 10888 16476 11244 16504
rect 11238 16464 11244 16476
rect 11296 16464 11302 16516
rect 12342 16504 12348 16516
rect 11900 16476 12348 16504
rect 8478 16436 8484 16448
rect 7024 16408 8484 16436
rect 5997 16399 6055 16405
rect 8478 16396 8484 16408
rect 8536 16436 8542 16448
rect 11900 16445 11928 16476
rect 12342 16464 12348 16476
rect 12400 16504 12406 16516
rect 15286 16504 15292 16516
rect 12400 16476 15292 16504
rect 12400 16464 12406 16476
rect 15286 16464 15292 16476
rect 15344 16464 15350 16516
rect 16761 16507 16819 16513
rect 16761 16473 16773 16507
rect 16807 16473 16819 16507
rect 16761 16467 16819 16473
rect 8665 16439 8723 16445
rect 8665 16436 8677 16439
rect 8536 16408 8677 16436
rect 8536 16396 8542 16408
rect 8665 16405 8677 16408
rect 8711 16405 8723 16439
rect 8665 16399 8723 16405
rect 11885 16439 11943 16445
rect 11885 16405 11897 16439
rect 11931 16405 11943 16439
rect 11885 16399 11943 16405
rect 12437 16439 12495 16445
rect 12437 16405 12449 16439
rect 12483 16436 12495 16439
rect 12618 16436 12624 16448
rect 12483 16408 12624 16436
rect 12483 16405 12495 16408
rect 12437 16399 12495 16405
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 12710 16396 12716 16448
rect 12768 16436 12774 16448
rect 13170 16436 13176 16448
rect 12768 16408 13176 16436
rect 12768 16396 12774 16408
rect 13170 16396 13176 16408
rect 13228 16436 13234 16448
rect 15194 16436 15200 16448
rect 13228 16408 15200 16436
rect 13228 16396 13234 16408
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 16776 16436 16804 16467
rect 16850 16436 16856 16448
rect 16776 16408 16856 16436
rect 16850 16396 16856 16408
rect 16908 16396 16914 16448
rect 17034 16396 17040 16448
rect 17092 16436 17098 16448
rect 18506 16436 18512 16448
rect 17092 16408 18512 16436
rect 17092 16396 17098 16408
rect 18506 16396 18512 16408
rect 18564 16396 18570 16448
rect 18984 16445 19012 16544
rect 19429 16541 19441 16544
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16572 23719 16575
rect 23750 16572 23756 16584
rect 23707 16544 23756 16572
rect 23707 16541 23719 16544
rect 23661 16535 23719 16541
rect 23750 16532 23756 16544
rect 23808 16532 23814 16584
rect 24486 16572 24492 16584
rect 24447 16544 24492 16572
rect 24486 16532 24492 16544
rect 24544 16532 24550 16584
rect 24780 16581 24808 16612
rect 25225 16609 25237 16612
rect 25271 16609 25283 16643
rect 25225 16603 25283 16609
rect 24765 16575 24823 16581
rect 24765 16541 24777 16575
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 24909 16575 24967 16581
rect 24909 16541 24921 16575
rect 24955 16572 24967 16575
rect 25314 16572 25320 16584
rect 24955 16544 25320 16572
rect 24955 16541 24967 16544
rect 24909 16535 24967 16541
rect 25314 16532 25320 16544
rect 25372 16532 25378 16584
rect 26697 16575 26755 16581
rect 26697 16541 26709 16575
rect 26743 16541 26755 16575
rect 27154 16572 27160 16584
rect 27115 16544 27160 16572
rect 26697 16535 26755 16541
rect 20530 16464 20536 16516
rect 20588 16464 20594 16516
rect 24673 16507 24731 16513
rect 24673 16473 24685 16507
rect 24719 16504 24731 16507
rect 26418 16504 26424 16516
rect 24719 16476 26424 16504
rect 24719 16473 24731 16476
rect 24673 16467 24731 16473
rect 26418 16464 26424 16476
rect 26476 16464 26482 16516
rect 18969 16439 19027 16445
rect 18969 16405 18981 16439
rect 19015 16405 19027 16439
rect 18969 16399 19027 16405
rect 20073 16439 20131 16445
rect 20073 16405 20085 16439
rect 20119 16436 20131 16439
rect 20898 16436 20904 16448
rect 20119 16408 20904 16436
rect 20119 16405 20131 16408
rect 20073 16399 20131 16405
rect 20898 16396 20904 16408
rect 20956 16396 20962 16448
rect 23845 16439 23903 16445
rect 23845 16405 23857 16439
rect 23891 16436 23903 16439
rect 23934 16436 23940 16448
rect 23891 16408 23940 16436
rect 23891 16405 23903 16408
rect 23845 16399 23903 16405
rect 23934 16396 23940 16408
rect 23992 16396 23998 16448
rect 24026 16396 24032 16448
rect 24084 16436 24090 16448
rect 26712 16436 26740 16535
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 27522 16572 27528 16584
rect 27580 16581 27586 16584
rect 27488 16544 27528 16572
rect 27522 16532 27528 16544
rect 27580 16535 27588 16581
rect 27893 16575 27951 16581
rect 27893 16572 27905 16575
rect 27632 16544 27905 16572
rect 27580 16532 27586 16535
rect 27062 16464 27068 16516
rect 27120 16504 27126 16516
rect 27341 16507 27399 16513
rect 27341 16504 27353 16507
rect 27120 16476 27353 16504
rect 27120 16464 27126 16476
rect 27341 16473 27353 16476
rect 27387 16473 27399 16507
rect 27341 16467 27399 16473
rect 27430 16464 27436 16516
rect 27488 16504 27494 16516
rect 27488 16476 27533 16504
rect 27488 16464 27494 16476
rect 24084 16408 26740 16436
rect 26881 16439 26939 16445
rect 24084 16396 24090 16408
rect 26881 16405 26893 16439
rect 26927 16436 26939 16439
rect 27632 16436 27660 16544
rect 27893 16541 27905 16544
rect 27939 16541 27951 16575
rect 27893 16535 27951 16541
rect 26927 16408 27660 16436
rect 26927 16405 26939 16408
rect 26881 16399 26939 16405
rect 27706 16396 27712 16448
rect 27764 16445 27770 16448
rect 27764 16436 27775 16445
rect 27764 16408 27809 16436
rect 27764 16399 27775 16408
rect 27764 16396 27770 16399
rect 1104 16346 29532 16368
rect 1104 16294 10425 16346
rect 10477 16294 10489 16346
rect 10541 16294 10553 16346
rect 10605 16294 10617 16346
rect 10669 16294 10681 16346
rect 10733 16294 19901 16346
rect 19953 16294 19965 16346
rect 20017 16294 20029 16346
rect 20081 16294 20093 16346
rect 20145 16294 20157 16346
rect 20209 16294 29532 16346
rect 1104 16272 29532 16294
rect 2866 16232 2872 16244
rect 2827 16204 2872 16232
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 4062 16192 4068 16244
rect 4120 16232 4126 16244
rect 5074 16232 5080 16244
rect 4120 16204 4844 16232
rect 5035 16204 5080 16232
rect 4120 16192 4126 16204
rect 2314 16164 2320 16176
rect 2275 16136 2320 16164
rect 2314 16124 2320 16136
rect 2372 16124 2378 16176
rect 3605 16167 3663 16173
rect 3605 16164 3617 16167
rect 2792 16136 3617 16164
rect 2792 16108 2820 16136
rect 3605 16133 3617 16136
rect 3651 16133 3663 16167
rect 3605 16127 3663 16133
rect 3694 16124 3700 16176
rect 3752 16164 3758 16176
rect 4706 16164 4712 16176
rect 3752 16136 3797 16164
rect 4356 16136 4712 16164
rect 3752 16124 3758 16136
rect 2774 16105 2780 16108
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16065 2559 16099
rect 2501 16059 2559 16065
rect 2757 16099 2780 16105
rect 2757 16065 2769 16099
rect 2757 16059 2780 16065
rect 2516 15960 2544 16059
rect 2774 16056 2780 16059
rect 2832 16056 2838 16108
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16096 3019 16099
rect 3237 16099 3295 16105
rect 3237 16096 3249 16099
rect 3007 16068 3249 16096
rect 3007 16065 3019 16068
rect 2961 16059 3019 16065
rect 3237 16065 3249 16068
rect 3283 16065 3295 16099
rect 3237 16059 3295 16065
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16065 3479 16099
rect 3970 16096 3976 16108
rect 3931 16068 3976 16096
rect 3421 16059 3479 16065
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 16028 3111 16031
rect 3142 16028 3148 16040
rect 3099 16000 3148 16028
rect 3099 15997 3111 16000
rect 3053 15991 3111 15997
rect 3142 15988 3148 16000
rect 3200 15988 3206 16040
rect 3326 15988 3332 16040
rect 3384 16028 3390 16040
rect 3436 16028 3464 16059
rect 3970 16056 3976 16068
rect 4028 16056 4034 16108
rect 4356 16105 4384 16136
rect 4706 16124 4712 16136
rect 4764 16124 4770 16176
rect 4816 16164 4844 16204
rect 5074 16192 5080 16204
rect 5132 16192 5138 16244
rect 7190 16192 7196 16244
rect 7248 16232 7254 16244
rect 7469 16235 7527 16241
rect 7469 16232 7481 16235
rect 7248 16204 7481 16232
rect 7248 16192 7254 16204
rect 7469 16201 7481 16204
rect 7515 16201 7527 16235
rect 8478 16232 8484 16244
rect 8439 16204 8484 16232
rect 7469 16195 7527 16201
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 10962 16232 10968 16244
rect 8588 16204 10968 16232
rect 8588 16164 8616 16204
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 11057 16235 11115 16241
rect 11057 16201 11069 16235
rect 11103 16232 11115 16235
rect 11330 16232 11336 16244
rect 11103 16204 11336 16232
rect 11103 16201 11115 16204
rect 11057 16195 11115 16201
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 12894 16192 12900 16244
rect 12952 16192 12958 16244
rect 14001 16235 14059 16241
rect 14001 16201 14013 16235
rect 14047 16232 14059 16235
rect 14182 16232 14188 16244
rect 14047 16204 14188 16232
rect 14047 16201 14059 16204
rect 14001 16195 14059 16201
rect 14182 16192 14188 16204
rect 14240 16192 14246 16244
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 16022 16232 16028 16244
rect 14599 16204 16028 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 4816 16136 8616 16164
rect 9309 16167 9367 16173
rect 9309 16133 9321 16167
rect 9355 16133 9367 16167
rect 9309 16127 9367 16133
rect 9401 16167 9459 16173
rect 9401 16133 9413 16167
rect 9447 16164 9459 16167
rect 11882 16164 11888 16176
rect 9447 16136 11888 16164
rect 9447 16133 9459 16136
rect 9401 16127 9459 16133
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16065 4399 16099
rect 4614 16096 4620 16108
rect 4575 16068 4620 16096
rect 4341 16059 4399 16065
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 4890 16056 4896 16108
rect 4948 16096 4954 16108
rect 7653 16099 7711 16105
rect 4948 16068 4993 16096
rect 4948 16056 4954 16068
rect 7653 16065 7665 16099
rect 7699 16096 7711 16099
rect 7699 16068 8064 16096
rect 7699 16065 7711 16068
rect 7653 16059 7711 16065
rect 3881 16031 3939 16037
rect 3881 16028 3893 16031
rect 3384 16000 3893 16028
rect 3384 15988 3390 16000
rect 3881 15997 3893 16000
rect 3927 15997 3939 16031
rect 3881 15991 3939 15997
rect 3602 15960 3608 15972
rect 2516 15932 3608 15960
rect 3602 15920 3608 15932
rect 3660 15960 3666 15972
rect 8036 15969 8064 16068
rect 8386 16056 8392 16108
rect 8444 16096 8450 16108
rect 8573 16099 8631 16105
rect 8573 16096 8585 16099
rect 8444 16068 8585 16096
rect 8444 16056 8450 16068
rect 8573 16065 8585 16068
rect 8619 16096 8631 16099
rect 9122 16096 9128 16108
rect 8619 16068 9128 16096
rect 8619 16065 8631 16068
rect 8573 16059 8631 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 8478 16028 8484 16040
rect 8439 16000 8484 16028
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 9214 16028 9220 16040
rect 9175 16000 9220 16028
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 8021 15963 8079 15969
rect 3660 15932 4844 15960
rect 3660 15920 3666 15932
rect 3050 15852 3056 15904
rect 3108 15892 3114 15904
rect 4433 15895 4491 15901
rect 4433 15892 4445 15895
rect 3108 15864 4445 15892
rect 3108 15852 3114 15864
rect 4433 15861 4445 15864
rect 4479 15892 4491 15895
rect 4614 15892 4620 15904
rect 4479 15864 4620 15892
rect 4479 15861 4491 15864
rect 4433 15855 4491 15861
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 4816 15901 4844 15932
rect 8021 15929 8033 15963
rect 8067 15929 8079 15963
rect 9324 15960 9352 16127
rect 11882 16124 11888 16136
rect 11940 16124 11946 16176
rect 12710 16164 12716 16176
rect 11992 16136 12716 16164
rect 10226 16056 10232 16108
rect 10284 16096 10290 16108
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 10284 16068 10517 16096
rect 10284 16056 10290 16068
rect 10505 16065 10517 16068
rect 10551 16065 10563 16099
rect 10965 16099 11023 16105
rect 10965 16096 10977 16099
rect 10505 16059 10563 16065
rect 10888 16068 10977 16096
rect 10318 15988 10324 16040
rect 10376 16028 10382 16040
rect 10888 16028 10916 16068
rect 10965 16065 10977 16068
rect 11011 16065 11023 16099
rect 10965 16059 11023 16065
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11992 16096 12020 16136
rect 12710 16124 12716 16136
rect 12768 16124 12774 16176
rect 12066 16105 12072 16108
rect 11112 16068 12020 16096
rect 12049 16099 12072 16105
rect 11112 16056 11118 16068
rect 12049 16065 12061 16099
rect 12049 16059 12072 16065
rect 12066 16056 12072 16059
rect 12124 16056 12130 16108
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16065 12219 16099
rect 12161 16059 12219 16065
rect 10376 16000 10916 16028
rect 10376 15988 10382 16000
rect 12176 15960 12204 16059
rect 12342 16056 12348 16108
rect 12400 16096 12406 16108
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 12400 16068 12449 16096
rect 12400 16056 12406 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12618 16096 12624 16108
rect 12579 16068 12624 16096
rect 12437 16059 12495 16065
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 12912 16105 12940 16192
rect 13004 16136 14504 16164
rect 13004 16105 13032 16136
rect 12804 16099 12862 16105
rect 12804 16065 12816 16099
rect 12850 16065 12862 16099
rect 12804 16059 12862 16065
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16065 12955 16099
rect 12897 16059 12955 16065
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13173 16099 13231 16105
rect 13173 16065 13185 16099
rect 13219 16096 13231 16099
rect 13446 16096 13452 16108
rect 13219 16068 13452 16096
rect 13219 16065 13231 16068
rect 13173 16059 13231 16065
rect 12526 16028 12532 16040
rect 12487 16000 12532 16028
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 12434 15960 12440 15972
rect 9324 15932 12020 15960
rect 12176 15932 12440 15960
rect 8021 15923 8079 15929
rect 4801 15895 4859 15901
rect 4801 15861 4813 15895
rect 4847 15892 4859 15895
rect 5534 15892 5540 15904
rect 4847 15864 5540 15892
rect 4847 15861 4859 15864
rect 4801 15855 4859 15861
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 8110 15852 8116 15904
rect 8168 15892 8174 15904
rect 8849 15895 8907 15901
rect 8849 15892 8861 15895
rect 8168 15864 8861 15892
rect 8168 15852 8174 15864
rect 8849 15861 8861 15864
rect 8895 15861 8907 15895
rect 8849 15855 8907 15861
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 10778 15892 10784 15904
rect 10735 15864 10784 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 10962 15852 10968 15904
rect 11020 15892 11026 15904
rect 11885 15895 11943 15901
rect 11885 15892 11897 15895
rect 11020 15864 11897 15892
rect 11020 15852 11026 15864
rect 11885 15861 11897 15864
rect 11931 15861 11943 15895
rect 11992 15892 12020 15932
rect 12434 15920 12440 15932
rect 12492 15920 12498 15972
rect 12819 15960 12847 16059
rect 13446 16056 13452 16068
rect 13504 16056 13510 16108
rect 14093 16099 14151 16105
rect 14093 16065 14105 16099
rect 14139 16096 14151 16099
rect 14274 16096 14280 16108
rect 14139 16068 14280 16096
rect 14139 16065 14151 16068
rect 14093 16059 14151 16065
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 14366 16056 14372 16108
rect 14424 16096 14430 16108
rect 14476 16105 14504 16136
rect 14461 16099 14519 16105
rect 14461 16096 14473 16099
rect 14424 16068 14473 16096
rect 14424 16056 14430 16068
rect 14461 16065 14473 16068
rect 14507 16065 14519 16099
rect 14461 16059 14519 16065
rect 14185 16031 14243 16037
rect 14185 15997 14197 16031
rect 14231 16028 14243 16031
rect 14568 16028 14596 16195
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 16758 16192 16764 16244
rect 16816 16232 16822 16244
rect 16853 16235 16911 16241
rect 16853 16232 16865 16235
rect 16816 16204 16865 16232
rect 16816 16192 16822 16204
rect 16853 16201 16865 16204
rect 16899 16201 16911 16235
rect 16853 16195 16911 16201
rect 16942 16192 16948 16244
rect 17000 16232 17006 16244
rect 19242 16232 19248 16244
rect 17000 16204 17045 16232
rect 17144 16204 19248 16232
rect 17000 16192 17006 16204
rect 16114 16164 16120 16176
rect 15764 16136 16120 16164
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14231 16000 14596 16028
rect 14844 16068 14933 16096
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 14844 15972 14872 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 15286 16096 15292 16108
rect 15247 16068 15292 16096
rect 14921 16059 14979 16065
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15764 16105 15792 16136
rect 16114 16124 16120 16136
rect 16172 16164 16178 16176
rect 17144 16164 17172 16204
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 19518 16192 19524 16244
rect 19576 16232 19582 16244
rect 20257 16235 20315 16241
rect 20257 16232 20269 16235
rect 19576 16204 20269 16232
rect 19576 16192 19582 16204
rect 20257 16201 20269 16204
rect 20303 16201 20315 16235
rect 22186 16232 22192 16244
rect 20257 16195 20315 16201
rect 22112 16204 22192 16232
rect 16172 16136 17172 16164
rect 17221 16167 17279 16173
rect 16172 16124 16178 16136
rect 17221 16133 17233 16167
rect 17267 16164 17279 16167
rect 17678 16164 17684 16176
rect 17267 16136 17684 16164
rect 17267 16133 17279 16136
rect 17221 16127 17279 16133
rect 17678 16124 17684 16136
rect 17736 16124 17742 16176
rect 18322 16124 18328 16176
rect 18380 16124 18386 16176
rect 18874 16124 18880 16176
rect 18932 16164 18938 16176
rect 19536 16164 19564 16192
rect 18932 16136 19564 16164
rect 18932 16124 18938 16136
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 15930 16056 15936 16108
rect 15988 16096 15994 16108
rect 16025 16099 16083 16105
rect 16025 16096 16037 16099
rect 15988 16068 16037 16096
rect 15988 16056 15994 16068
rect 16025 16065 16037 16068
rect 16071 16096 16083 16099
rect 16390 16096 16396 16108
rect 16071 16068 16396 16096
rect 16071 16065 16083 16068
rect 16025 16059 16083 16065
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 16666 16096 16672 16108
rect 16627 16068 16672 16096
rect 16666 16056 16672 16068
rect 16724 16056 16730 16108
rect 16758 16056 16764 16108
rect 16816 16096 16822 16108
rect 17034 16096 17040 16108
rect 16816 16068 17040 16096
rect 16816 16056 16822 16068
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 20272 16096 20300 16195
rect 22112 16173 22140 16204
rect 22186 16192 22192 16204
rect 22244 16192 22250 16244
rect 22646 16192 22652 16244
rect 22704 16232 22710 16244
rect 26234 16232 26240 16244
rect 22704 16204 26240 16232
rect 22704 16192 22710 16204
rect 22097 16167 22155 16173
rect 22097 16133 22109 16167
rect 22143 16133 22155 16167
rect 22097 16127 22155 16133
rect 23934 16124 23940 16176
rect 23992 16124 23998 16176
rect 20441 16099 20499 16105
rect 20441 16096 20453 16099
rect 20272 16068 20453 16096
rect 20441 16065 20453 16068
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 21174 16056 21180 16108
rect 21232 16096 21238 16108
rect 21913 16099 21971 16105
rect 21913 16096 21925 16099
rect 21232 16068 21925 16096
rect 21232 16056 21238 16068
rect 21913 16065 21925 16068
rect 21959 16065 21971 16099
rect 21913 16059 21971 16065
rect 22189 16099 22247 16105
rect 22189 16065 22201 16099
rect 22235 16065 22247 16099
rect 22189 16059 22247 16065
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 15997 15071 16031
rect 15194 16028 15200 16040
rect 15155 16000 15200 16028
rect 15013 15991 15071 15997
rect 12894 15960 12900 15972
rect 12819 15932 12900 15960
rect 12894 15920 12900 15932
rect 12952 15920 12958 15972
rect 13633 15963 13691 15969
rect 13633 15960 13645 15963
rect 13004 15932 13645 15960
rect 13004 15892 13032 15932
rect 13633 15929 13645 15932
rect 13679 15929 13691 15963
rect 13633 15923 13691 15929
rect 14550 15920 14556 15972
rect 14608 15960 14614 15972
rect 14826 15960 14832 15972
rect 14608 15932 14832 15960
rect 14608 15920 14614 15932
rect 14826 15920 14832 15932
rect 14884 15920 14890 15972
rect 15028 15960 15056 15991
rect 15194 15988 15200 16000
rect 15252 15988 15258 16040
rect 16114 16028 16120 16040
rect 15764 16000 16120 16028
rect 15764 15960 15792 16000
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 17313 16031 17371 16037
rect 17313 15997 17325 16031
rect 17359 15997 17371 16031
rect 17586 16028 17592 16040
rect 17547 16000 17592 16028
rect 17313 15991 17371 15997
rect 15930 15960 15936 15972
rect 15028 15932 15792 15960
rect 15891 15932 15936 15960
rect 15930 15920 15936 15932
rect 15988 15960 15994 15972
rect 15988 15932 16068 15960
rect 15988 15920 15994 15932
rect 11992 15864 13032 15892
rect 13265 15895 13323 15901
rect 11885 15855 11943 15861
rect 13265 15861 13277 15895
rect 13311 15892 13323 15895
rect 13538 15892 13544 15904
rect 13311 15864 13544 15892
rect 13311 15861 13323 15864
rect 13265 15855 13323 15861
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 15654 15892 15660 15904
rect 15615 15864 15660 15892
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 16040 15901 16068 15932
rect 16025 15895 16083 15901
rect 16025 15861 16037 15895
rect 16071 15861 16083 15895
rect 16025 15855 16083 15861
rect 16393 15895 16451 15901
rect 16393 15861 16405 15895
rect 16439 15892 16451 15895
rect 16666 15892 16672 15904
rect 16439 15864 16672 15892
rect 16439 15861 16451 15864
rect 16393 15855 16451 15861
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 17328 15892 17356 15991
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 17770 15892 17776 15904
rect 17328 15864 17776 15892
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 19058 15892 19064 15904
rect 19019 15864 19064 15892
rect 19058 15852 19064 15864
rect 19116 15852 19122 15904
rect 20625 15895 20683 15901
rect 20625 15861 20637 15895
rect 20671 15892 20683 15895
rect 21082 15892 21088 15904
rect 20671 15864 21088 15892
rect 20671 15861 20683 15864
rect 20625 15855 20683 15861
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 22204 15892 22232 16059
rect 22278 16056 22284 16108
rect 22336 16105 22342 16108
rect 22336 16096 22344 16105
rect 22646 16096 22652 16108
rect 22336 16068 22381 16096
rect 22607 16068 22652 16096
rect 22336 16059 22344 16068
rect 22336 16056 22342 16059
rect 22646 16056 22652 16068
rect 22704 16056 22710 16108
rect 24302 16056 24308 16108
rect 24360 16096 24366 16108
rect 24581 16099 24639 16105
rect 24581 16096 24593 16099
rect 24360 16068 24593 16096
rect 24360 16056 24366 16068
rect 24581 16065 24593 16068
rect 24627 16065 24639 16099
rect 24872 16096 24900 16204
rect 26234 16192 26240 16204
rect 26292 16232 26298 16244
rect 26292 16204 27384 16232
rect 26292 16192 26298 16204
rect 26602 16164 26608 16176
rect 26450 16136 26608 16164
rect 26602 16124 26608 16136
rect 26660 16124 26666 16176
rect 24946 16096 24952 16108
rect 24859 16068 24952 16096
rect 24581 16059 24639 16065
rect 24946 16056 24952 16068
rect 25004 16056 25010 16108
rect 27356 16105 27384 16204
rect 27617 16167 27675 16173
rect 27617 16133 27629 16167
rect 27663 16164 27675 16167
rect 27706 16164 27712 16176
rect 27663 16136 27712 16164
rect 27663 16133 27675 16136
rect 27617 16127 27675 16133
rect 27706 16124 27712 16136
rect 27764 16124 27770 16176
rect 28626 16124 28632 16176
rect 28684 16124 28690 16176
rect 27341 16099 27399 16105
rect 27341 16065 27353 16099
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 22925 16031 22983 16037
rect 22925 16028 22937 16031
rect 22480 16000 22937 16028
rect 22480 15969 22508 16000
rect 22925 15997 22937 16000
rect 22971 15997 22983 16031
rect 24394 16028 24400 16040
rect 24355 16000 24400 16028
rect 22925 15991 22983 15997
rect 24394 15988 24400 16000
rect 24452 15988 24458 16040
rect 25222 16028 25228 16040
rect 25183 16000 25228 16028
rect 25222 15988 25228 16000
rect 25280 15988 25286 16040
rect 22465 15963 22523 15969
rect 22465 15929 22477 15963
rect 22511 15929 22523 15963
rect 22465 15923 22523 15929
rect 24412 15892 24440 15988
rect 22204 15864 24440 15892
rect 24765 15895 24823 15901
rect 24765 15861 24777 15895
rect 24811 15892 24823 15895
rect 25314 15892 25320 15904
rect 24811 15864 25320 15892
rect 24811 15861 24823 15864
rect 24765 15855 24823 15861
rect 25314 15852 25320 15864
rect 25372 15852 25378 15904
rect 25406 15852 25412 15904
rect 25464 15892 25470 15904
rect 26697 15895 26755 15901
rect 26697 15892 26709 15895
rect 25464 15864 26709 15892
rect 25464 15852 25470 15864
rect 26697 15861 26709 15864
rect 26743 15861 26755 15895
rect 26697 15855 26755 15861
rect 27338 15852 27344 15904
rect 27396 15892 27402 15904
rect 29089 15895 29147 15901
rect 29089 15892 29101 15895
rect 27396 15864 29101 15892
rect 27396 15852 27402 15864
rect 29089 15861 29101 15864
rect 29135 15861 29147 15895
rect 29089 15855 29147 15861
rect 1104 15802 29532 15824
rect 1104 15750 5688 15802
rect 5740 15750 5752 15802
rect 5804 15750 5816 15802
rect 5868 15750 5880 15802
rect 5932 15750 5944 15802
rect 5996 15750 15163 15802
rect 15215 15750 15227 15802
rect 15279 15750 15291 15802
rect 15343 15750 15355 15802
rect 15407 15750 15419 15802
rect 15471 15750 24639 15802
rect 24691 15750 24703 15802
rect 24755 15750 24767 15802
rect 24819 15750 24831 15802
rect 24883 15750 24895 15802
rect 24947 15750 29532 15802
rect 1104 15728 29532 15750
rect 3970 15648 3976 15700
rect 4028 15688 4034 15700
rect 4525 15691 4583 15697
rect 4525 15688 4537 15691
rect 4028 15660 4537 15688
rect 4028 15648 4034 15660
rect 3878 15620 3884 15632
rect 2884 15592 3884 15620
rect 2884 15561 2912 15592
rect 3878 15580 3884 15592
rect 3936 15580 3942 15632
rect 2869 15555 2927 15561
rect 2869 15521 2881 15555
rect 2915 15521 2927 15555
rect 3050 15552 3056 15564
rect 3011 15524 3056 15552
rect 2869 15515 2927 15521
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 3234 15512 3240 15564
rect 3292 15552 3298 15564
rect 4157 15555 4215 15561
rect 3292 15524 3372 15552
rect 3292 15512 3298 15524
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 3016 15456 3061 15484
rect 3016 15444 3022 15456
rect 3142 15444 3148 15496
rect 3200 15484 3206 15496
rect 3344 15493 3372 15524
rect 4157 15521 4169 15555
rect 4203 15552 4215 15555
rect 4246 15552 4252 15564
rect 4203 15524 4252 15552
rect 4203 15521 4215 15524
rect 4157 15515 4215 15521
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 4376 15561 4404 15660
rect 4525 15657 4537 15660
rect 4571 15657 4583 15691
rect 4525 15651 4583 15657
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 14366 15688 14372 15700
rect 8536 15660 12434 15688
rect 14327 15660 14372 15688
rect 8536 15648 8542 15660
rect 5721 15623 5779 15629
rect 5721 15589 5733 15623
rect 5767 15589 5779 15623
rect 5721 15583 5779 15589
rect 9217 15623 9275 15629
rect 9217 15589 9229 15623
rect 9263 15589 9275 15623
rect 12406 15620 12434 15660
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 16298 15688 16304 15700
rect 14476 15660 16304 15688
rect 14476 15620 14504 15660
rect 16298 15648 16304 15660
rect 16356 15648 16362 15700
rect 17221 15691 17279 15697
rect 17221 15657 17233 15691
rect 17267 15688 17279 15691
rect 17586 15688 17592 15700
rect 17267 15660 17592 15688
rect 17267 15657 17279 15660
rect 17221 15651 17279 15657
rect 17586 15648 17592 15660
rect 17644 15648 17650 15700
rect 18322 15648 18328 15700
rect 18380 15688 18386 15700
rect 18417 15691 18475 15697
rect 18417 15688 18429 15691
rect 18380 15660 18429 15688
rect 18380 15648 18386 15660
rect 18417 15657 18429 15660
rect 18463 15657 18475 15691
rect 18417 15651 18475 15657
rect 19337 15691 19395 15697
rect 19337 15657 19349 15691
rect 19383 15688 19395 15691
rect 19518 15688 19524 15700
rect 19383 15660 19524 15688
rect 19383 15657 19395 15660
rect 19337 15651 19395 15657
rect 19518 15648 19524 15660
rect 19576 15648 19582 15700
rect 21361 15691 21419 15697
rect 21361 15688 21373 15691
rect 19812 15660 21373 15688
rect 12406 15592 14504 15620
rect 16025 15623 16083 15629
rect 9217 15583 9275 15589
rect 16025 15589 16037 15623
rect 16071 15620 16083 15623
rect 16206 15620 16212 15632
rect 16071 15592 16212 15620
rect 16071 15589 16083 15592
rect 16025 15583 16083 15589
rect 4341 15555 4404 15561
rect 4341 15521 4353 15555
rect 4387 15524 4404 15555
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 3329 15487 3387 15493
rect 3200 15456 3293 15484
rect 3200 15444 3206 15456
rect 3329 15453 3341 15487
rect 3375 15453 3387 15487
rect 4433 15487 4491 15493
rect 4433 15484 4445 15487
rect 3329 15447 3387 15453
rect 4376 15456 4445 15484
rect 3160 15416 3188 15444
rect 4376 15416 4404 15456
rect 4433 15453 4445 15456
rect 4479 15453 4491 15487
rect 4522 15478 4528 15530
rect 4580 15478 4586 15530
rect 4433 15447 4491 15453
rect 4525 15453 4537 15478
rect 4571 15453 4583 15478
rect 4525 15447 4583 15453
rect 4614 15444 4620 15496
rect 4672 15484 4678 15496
rect 4672 15456 4717 15484
rect 4672 15444 4678 15456
rect 5074 15444 5080 15496
rect 5132 15484 5138 15496
rect 5169 15487 5227 15493
rect 5169 15484 5181 15487
rect 5132 15456 5181 15484
rect 5132 15444 5138 15456
rect 5169 15453 5181 15456
rect 5215 15453 5227 15487
rect 5350 15484 5356 15496
rect 5311 15456 5356 15484
rect 5169 15447 5227 15453
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 5534 15484 5540 15496
rect 5592 15493 5598 15496
rect 5500 15456 5540 15484
rect 5534 15444 5540 15456
rect 5592 15447 5600 15493
rect 5736 15484 5764 15583
rect 7110 15487 7168 15493
rect 7110 15484 7122 15487
rect 5736 15456 7122 15484
rect 7110 15453 7122 15456
rect 7156 15453 7168 15487
rect 7374 15484 7380 15496
rect 7335 15456 7380 15484
rect 7110 15447 7168 15453
rect 5592 15444 5598 15447
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 8110 15484 8116 15496
rect 8071 15456 8116 15484
rect 8110 15444 8116 15456
rect 8168 15444 8174 15496
rect 9033 15487 9091 15493
rect 9033 15453 9045 15487
rect 9079 15453 9091 15487
rect 9232 15484 9260 15583
rect 16206 15580 16212 15592
rect 16264 15580 16270 15632
rect 19812 15620 19840 15660
rect 21361 15657 21373 15660
rect 21407 15688 21419 15691
rect 21542 15688 21548 15700
rect 21407 15660 21548 15688
rect 21407 15657 21419 15660
rect 21361 15651 21419 15657
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 22646 15648 22652 15700
rect 22704 15688 22710 15700
rect 23750 15688 23756 15700
rect 22704 15660 23244 15688
rect 23711 15660 23756 15688
rect 22704 15648 22710 15660
rect 16592 15592 19840 15620
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15552 10011 15555
rect 10962 15552 10968 15564
rect 9999 15524 10968 15552
rect 9999 15521 10011 15524
rect 9953 15515 10011 15521
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 11425 15555 11483 15561
rect 11425 15521 11437 15555
rect 11471 15552 11483 15555
rect 11471 15524 12434 15552
rect 11471 15521 11483 15524
rect 11425 15515 11483 15521
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 9232 15456 9505 15484
rect 9033 15447 9091 15453
rect 9493 15453 9505 15456
rect 9539 15453 9551 15487
rect 9674 15484 9680 15496
rect 9635 15456 9680 15484
rect 9493 15447 9551 15453
rect 4632 15416 4660 15444
rect 5092 15416 5120 15444
rect 3160 15388 4108 15416
rect 4376 15388 4660 15416
rect 4724 15388 5120 15416
rect 2038 15308 2044 15360
rect 2096 15348 2102 15360
rect 2685 15351 2743 15357
rect 2685 15348 2697 15351
rect 2096 15320 2697 15348
rect 2096 15308 2102 15320
rect 2685 15317 2697 15320
rect 2731 15317 2743 15351
rect 2685 15311 2743 15317
rect 3878 15308 3884 15360
rect 3936 15348 3942 15360
rect 3973 15351 4031 15357
rect 3973 15348 3985 15351
rect 3936 15320 3985 15348
rect 3936 15308 3942 15320
rect 3973 15317 3985 15320
rect 4019 15317 4031 15351
rect 4080 15348 4108 15388
rect 4724 15348 4752 15388
rect 5442 15376 5448 15428
rect 5500 15425 5506 15428
rect 5500 15416 5508 15425
rect 9048 15416 9076 15447
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 11054 15444 11060 15496
rect 11112 15444 11118 15496
rect 12406 15484 12434 15524
rect 12710 15512 12716 15564
rect 12768 15552 12774 15564
rect 12768 15524 15792 15552
rect 12768 15512 12774 15524
rect 13814 15484 13820 15496
rect 12406 15456 13820 15484
rect 13814 15444 13820 15456
rect 13872 15484 13878 15496
rect 15764 15484 15792 15524
rect 15838 15512 15844 15564
rect 15896 15552 15902 15564
rect 16117 15555 16175 15561
rect 16117 15552 16129 15555
rect 15896 15524 16129 15552
rect 15896 15512 15902 15524
rect 16117 15521 16129 15524
rect 16163 15521 16175 15555
rect 16592 15552 16620 15592
rect 16117 15515 16175 15521
rect 16224 15524 16620 15552
rect 16224 15484 16252 15524
rect 16666 15512 16672 15564
rect 16724 15552 16730 15564
rect 16724 15524 17540 15552
rect 16724 15512 16730 15524
rect 13872 15456 14320 15484
rect 15764 15456 16252 15484
rect 16301 15487 16359 15493
rect 13872 15444 13878 15456
rect 5500 15388 6040 15416
rect 9048 15388 9812 15416
rect 5500 15379 5508 15388
rect 5500 15376 5506 15379
rect 4890 15348 4896 15360
rect 4080 15320 4752 15348
rect 4851 15320 4896 15348
rect 3973 15311 4031 15317
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 6012 15357 6040 15388
rect 9784 15360 9812 15388
rect 12342 15376 12348 15428
rect 12400 15416 12406 15428
rect 13630 15416 13636 15428
rect 12400 15388 13636 15416
rect 12400 15376 12406 15388
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 14090 15416 14096 15428
rect 14051 15388 14096 15416
rect 14090 15376 14096 15388
rect 14148 15376 14154 15428
rect 14292 15425 14320 15456
rect 16301 15453 16313 15487
rect 16347 15484 16359 15487
rect 16390 15484 16396 15496
rect 16347 15456 16396 15484
rect 16347 15453 16359 15456
rect 16301 15447 16359 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 16485 15487 16543 15493
rect 16485 15453 16497 15487
rect 16531 15484 16543 15487
rect 16574 15484 16580 15496
rect 16531 15456 16580 15484
rect 16531 15453 16543 15456
rect 16485 15447 16543 15453
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 16942 15444 16948 15496
rect 17000 15484 17006 15496
rect 17512 15493 17540 15524
rect 17678 15512 17684 15564
rect 17736 15552 17742 15564
rect 17773 15555 17831 15561
rect 17773 15552 17785 15555
rect 17736 15524 17785 15552
rect 17736 15512 17742 15524
rect 17773 15521 17785 15524
rect 17819 15521 17831 15555
rect 17773 15515 17831 15521
rect 17865 15555 17923 15561
rect 17865 15521 17877 15555
rect 17911 15552 17923 15555
rect 19058 15552 19064 15564
rect 17911 15524 19064 15552
rect 17911 15521 17923 15524
rect 17865 15515 17923 15521
rect 17359 15487 17417 15493
rect 17359 15484 17371 15487
rect 17000 15456 17371 15484
rect 17000 15444 17006 15456
rect 17359 15453 17371 15456
rect 17405 15453 17417 15487
rect 17359 15447 17417 15453
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15453 17555 15487
rect 17880 15484 17908 15515
rect 19058 15512 19064 15524
rect 19116 15512 19122 15564
rect 19242 15512 19248 15564
rect 19300 15552 19306 15564
rect 22830 15552 22836 15564
rect 19300 15524 22836 15552
rect 19300 15512 19306 15524
rect 22830 15512 22836 15524
rect 22888 15512 22894 15564
rect 23109 15555 23167 15561
rect 23109 15521 23121 15555
rect 23155 15552 23167 15555
rect 23216 15552 23244 15660
rect 23750 15648 23756 15660
rect 23808 15648 23814 15700
rect 25133 15691 25191 15697
rect 25133 15657 25145 15691
rect 25179 15688 25191 15691
rect 25222 15688 25228 15700
rect 25179 15660 25228 15688
rect 25179 15657 25191 15660
rect 25133 15651 25191 15657
rect 25222 15648 25228 15660
rect 25280 15648 25286 15700
rect 25682 15648 25688 15700
rect 25740 15688 25746 15700
rect 26602 15688 26608 15700
rect 25740 15660 26464 15688
rect 26563 15660 26608 15688
rect 25740 15648 25746 15660
rect 25406 15580 25412 15632
rect 25464 15620 25470 15632
rect 25777 15623 25835 15629
rect 25777 15620 25789 15623
rect 25464 15592 25789 15620
rect 25464 15580 25470 15592
rect 25777 15589 25789 15592
rect 25823 15589 25835 15623
rect 26436 15620 26464 15660
rect 26602 15648 26608 15660
rect 26660 15648 26666 15700
rect 28626 15688 28632 15700
rect 28587 15660 28632 15688
rect 28626 15648 28632 15660
rect 28684 15648 28690 15700
rect 26881 15623 26939 15629
rect 26881 15620 26893 15623
rect 26436 15592 26893 15620
rect 25777 15583 25835 15589
rect 26881 15589 26893 15592
rect 26927 15620 26939 15623
rect 26973 15623 27031 15629
rect 26973 15620 26985 15623
rect 26927 15592 26985 15620
rect 26927 15589 26939 15592
rect 26881 15583 26939 15589
rect 26973 15589 26985 15592
rect 27019 15589 27031 15623
rect 26973 15583 27031 15589
rect 27614 15580 27620 15632
rect 27672 15620 27678 15632
rect 27709 15623 27767 15629
rect 27709 15620 27721 15623
rect 27672 15592 27721 15620
rect 27672 15580 27678 15592
rect 27709 15589 27721 15592
rect 27755 15589 27767 15623
rect 27709 15583 27767 15589
rect 28261 15623 28319 15629
rect 28261 15589 28273 15623
rect 28307 15589 28319 15623
rect 28261 15583 28319 15589
rect 23155 15524 23244 15552
rect 25608 15524 27568 15552
rect 23155 15521 23167 15524
rect 23109 15515 23167 15521
rect 17497 15447 17555 15453
rect 17604 15456 17908 15484
rect 18233 15487 18291 15493
rect 14277 15419 14335 15425
rect 14277 15385 14289 15419
rect 14323 15416 14335 15419
rect 15010 15416 15016 15428
rect 14323 15388 15016 15416
rect 14323 15385 14335 15388
rect 14277 15379 14335 15385
rect 15010 15376 15016 15388
rect 15068 15376 15074 15428
rect 15562 15376 15568 15428
rect 15620 15416 15626 15428
rect 15657 15419 15715 15425
rect 15657 15416 15669 15419
rect 15620 15388 15669 15416
rect 15620 15376 15626 15388
rect 15657 15385 15669 15388
rect 15703 15385 15715 15419
rect 15657 15379 15715 15385
rect 15841 15419 15899 15425
rect 15841 15385 15853 15419
rect 15887 15416 15899 15419
rect 17604 15416 17632 15456
rect 18233 15453 18245 15487
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 18693 15487 18751 15493
rect 18693 15453 18705 15487
rect 18739 15484 18751 15487
rect 18782 15484 18788 15496
rect 18739 15456 18788 15484
rect 18739 15453 18751 15456
rect 18693 15447 18751 15453
rect 15887 15388 17632 15416
rect 18248 15416 18276 15447
rect 18782 15444 18788 15456
rect 18840 15444 18846 15496
rect 18966 15484 18972 15496
rect 18927 15456 18972 15484
rect 18966 15444 18972 15456
rect 19024 15444 19030 15496
rect 19702 15444 19708 15496
rect 19760 15444 19766 15496
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15453 21143 15487
rect 23382 15484 23388 15496
rect 23343 15456 23388 15484
rect 21085 15447 21143 15453
rect 20806 15416 20812 15428
rect 18248 15388 18828 15416
rect 20767 15388 20812 15416
rect 15887 15385 15899 15388
rect 15841 15379 15899 15385
rect 5997 15351 6055 15357
rect 5997 15317 6009 15351
rect 6043 15317 6055 15351
rect 5997 15311 6055 15317
rect 7742 15308 7748 15360
rect 7800 15348 7806 15360
rect 7929 15351 7987 15357
rect 7929 15348 7941 15351
rect 7800 15320 7941 15348
rect 7800 15308 7806 15320
rect 7929 15317 7941 15320
rect 7975 15317 7987 15351
rect 9306 15348 9312 15360
rect 9267 15320 9312 15348
rect 7929 15311 7987 15317
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 9766 15308 9772 15360
rect 9824 15308 9830 15360
rect 10318 15308 10324 15360
rect 10376 15348 10382 15360
rect 10962 15348 10968 15360
rect 10376 15320 10968 15348
rect 10376 15308 10382 15320
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 13538 15348 13544 15360
rect 12768 15320 13544 15348
rect 12768 15308 12774 15320
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 15672 15348 15700 15379
rect 16022 15348 16028 15360
rect 15672 15320 16028 15348
rect 16022 15308 16028 15320
rect 16080 15308 16086 15360
rect 18506 15348 18512 15360
rect 18467 15320 18512 15348
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 18800 15357 18828 15388
rect 20806 15376 20812 15388
rect 20864 15376 20870 15428
rect 18785 15351 18843 15357
rect 18785 15317 18797 15351
rect 18831 15317 18843 15351
rect 18785 15311 18843 15317
rect 20530 15308 20536 15360
rect 20588 15348 20594 15360
rect 21100 15348 21128 15447
rect 23382 15444 23388 15456
rect 23440 15444 23446 15496
rect 23566 15444 23572 15496
rect 23624 15484 23630 15496
rect 24026 15484 24032 15496
rect 23624 15456 24032 15484
rect 23624 15444 23630 15456
rect 24026 15444 24032 15456
rect 24084 15444 24090 15496
rect 24394 15444 24400 15496
rect 24452 15484 24458 15496
rect 25314 15493 25320 15496
rect 24489 15487 24547 15493
rect 24489 15484 24501 15487
rect 24452 15456 24501 15484
rect 24452 15444 24458 15456
rect 24489 15453 24501 15456
rect 24535 15453 24547 15487
rect 25312 15484 25320 15493
rect 25227 15456 25320 15484
rect 24489 15447 24547 15453
rect 25312 15447 25320 15456
rect 25372 15484 25378 15496
rect 25608 15484 25636 15524
rect 27540 15496 27568 15524
rect 25372 15456 25636 15484
rect 25685 15487 25743 15493
rect 25314 15444 25320 15447
rect 25372 15444 25378 15456
rect 25685 15453 25697 15487
rect 25731 15453 25743 15487
rect 26326 15484 26332 15496
rect 26287 15456 26332 15484
rect 25685 15447 25743 15453
rect 22830 15416 22836 15428
rect 20588 15320 21128 15348
rect 22388 15348 22416 15402
rect 22791 15388 22836 15416
rect 22830 15376 22836 15388
rect 22888 15376 22894 15428
rect 22922 15376 22928 15428
rect 22980 15416 22986 15428
rect 24302 15416 24308 15428
rect 22980 15388 24308 15416
rect 22980 15376 22986 15388
rect 24302 15376 24308 15388
rect 24360 15376 24366 15428
rect 25406 15416 25412 15428
rect 25367 15388 25412 15416
rect 25406 15376 25412 15388
rect 25464 15376 25470 15428
rect 25498 15376 25504 15428
rect 25556 15416 25562 15428
rect 25700 15416 25728 15447
rect 26326 15444 26332 15456
rect 26384 15444 26390 15496
rect 26789 15463 26847 15469
rect 26789 15429 26801 15463
rect 26835 15429 26847 15463
rect 26878 15444 26884 15496
rect 26936 15484 26942 15496
rect 27154 15484 27160 15496
rect 26936 15456 27160 15484
rect 26936 15444 26942 15456
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 27522 15444 27528 15496
rect 27580 15493 27586 15496
rect 27580 15484 27588 15493
rect 28077 15487 28135 15493
rect 27580 15456 27625 15484
rect 27580 15447 27588 15456
rect 28077 15453 28089 15487
rect 28123 15453 28135 15487
rect 28276 15484 28304 15583
rect 28445 15487 28503 15493
rect 28445 15484 28457 15487
rect 28276 15456 28457 15484
rect 28077 15447 28135 15453
rect 28445 15453 28457 15456
rect 28491 15453 28503 15487
rect 28445 15447 28503 15453
rect 27580 15444 27586 15447
rect 26694 15416 26700 15428
rect 25556 15388 25601 15416
rect 25700 15388 26700 15416
rect 25556 15376 25562 15388
rect 23201 15351 23259 15357
rect 23201 15348 23213 15351
rect 22388 15320 23213 15348
rect 20588 15308 20594 15320
rect 23201 15317 23213 15320
rect 23247 15317 23259 15351
rect 23201 15311 23259 15317
rect 24486 15308 24492 15360
rect 24544 15348 24550 15360
rect 24673 15351 24731 15357
rect 24673 15348 24685 15351
rect 24544 15320 24685 15348
rect 24544 15308 24550 15320
rect 24673 15317 24685 15320
rect 24719 15348 24731 15351
rect 25700 15348 25728 15388
rect 26694 15376 26700 15388
rect 26752 15376 26758 15428
rect 26789 15423 26847 15429
rect 24719 15320 25728 15348
rect 26513 15351 26571 15357
rect 24719 15317 24731 15320
rect 24673 15311 24731 15317
rect 26513 15317 26525 15351
rect 26559 15348 26571 15351
rect 26804 15348 26832 15423
rect 27341 15419 27399 15425
rect 27341 15385 27353 15419
rect 27387 15385 27399 15419
rect 27341 15379 27399 15385
rect 26559 15320 26832 15348
rect 26881 15351 26939 15357
rect 26559 15317 26571 15320
rect 26513 15311 26571 15317
rect 26881 15317 26893 15351
rect 26927 15348 26939 15351
rect 27356 15348 27384 15379
rect 27430 15376 27436 15428
rect 27488 15416 27494 15428
rect 27488 15388 27533 15416
rect 27488 15376 27494 15388
rect 26927 15320 27384 15348
rect 26927 15317 26939 15320
rect 26881 15311 26939 15317
rect 27522 15308 27528 15360
rect 27580 15348 27586 15360
rect 28092 15348 28120 15447
rect 27580 15320 28120 15348
rect 27580 15308 27586 15320
rect 1104 15258 29532 15280
rect 1104 15206 10425 15258
rect 10477 15206 10489 15258
rect 10541 15206 10553 15258
rect 10605 15206 10617 15258
rect 10669 15206 10681 15258
rect 10733 15206 19901 15258
rect 19953 15206 19965 15258
rect 20017 15206 20029 15258
rect 20081 15206 20093 15258
rect 20145 15206 20157 15258
rect 20209 15206 29532 15258
rect 1104 15184 29532 15206
rect 2958 15104 2964 15156
rect 3016 15144 3022 15156
rect 3053 15147 3111 15153
rect 3053 15144 3065 15147
rect 3016 15116 3065 15144
rect 3016 15104 3022 15116
rect 3053 15113 3065 15116
rect 3099 15113 3111 15147
rect 3053 15107 3111 15113
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 4249 15147 4307 15153
rect 4249 15144 4261 15147
rect 4212 15116 4261 15144
rect 4212 15104 4218 15116
rect 4249 15113 4261 15116
rect 4295 15113 4307 15147
rect 4249 15107 4307 15113
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 4755 15116 5764 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 2774 15076 2780 15088
rect 1412 15048 2780 15076
rect 1412 15017 1440 15048
rect 2774 15036 2780 15048
rect 2832 15036 2838 15088
rect 4614 15076 4620 15088
rect 3620 15048 4620 15076
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 1664 15011 1722 15017
rect 1664 14977 1676 15011
rect 1710 15008 1722 15011
rect 1946 15008 1952 15020
rect 1710 14980 1952 15008
rect 1710 14977 1722 14980
rect 1664 14971 1722 14977
rect 1946 14968 1952 14980
rect 2004 14968 2010 15020
rect 3234 15008 3240 15020
rect 3195 14980 3240 15008
rect 3234 14968 3240 14980
rect 3292 14968 3298 15020
rect 3326 14968 3332 15020
rect 3384 15008 3390 15020
rect 3620 15017 3648 15048
rect 4614 15036 4620 15048
rect 4672 15036 4678 15088
rect 3605 15011 3663 15017
rect 3384 14980 3429 15008
rect 3384 14968 3390 14980
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3878 15008 3884 15020
rect 3839 14980 3884 15008
rect 3605 14971 3663 14977
rect 2777 14875 2835 14881
rect 2777 14841 2789 14875
rect 2823 14872 2835 14875
rect 3142 14872 3148 14884
rect 2823 14844 3148 14872
rect 2823 14841 2835 14844
rect 2777 14835 2835 14841
rect 3142 14832 3148 14844
rect 3200 14872 3206 14884
rect 3620 14872 3648 14971
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 3786 14900 3792 14952
rect 3844 14940 3850 14952
rect 3973 14943 4031 14949
rect 3973 14940 3985 14943
rect 3844 14912 3985 14940
rect 3844 14900 3850 14912
rect 3973 14909 3985 14912
rect 4019 14909 4031 14943
rect 3973 14903 4031 14909
rect 4430 14900 4436 14952
rect 4488 14940 4494 14952
rect 4724 14940 4752 15107
rect 5442 15076 5448 15088
rect 5403 15048 5448 15076
rect 5442 15036 5448 15048
rect 5500 15036 5506 15088
rect 4890 15008 4896 15020
rect 4851 14980 4896 15008
rect 4890 14968 4896 14980
rect 4948 14968 4954 15020
rect 5736 15017 5764 15116
rect 10226 15104 10232 15156
rect 10284 15144 10290 15156
rect 10689 15147 10747 15153
rect 10689 15144 10701 15147
rect 10284 15116 10701 15144
rect 10284 15104 10290 15116
rect 10689 15113 10701 15116
rect 10735 15113 10747 15147
rect 10689 15107 10747 15113
rect 10965 15147 11023 15153
rect 10965 15113 10977 15147
rect 11011 15144 11023 15147
rect 11054 15144 11060 15156
rect 11011 15116 11060 15144
rect 11011 15113 11023 15116
rect 10965 15107 11023 15113
rect 7742 15076 7748 15088
rect 7703 15048 7748 15076
rect 7742 15036 7748 15048
rect 7800 15036 7806 15088
rect 9306 15076 9312 15088
rect 8970 15048 9312 15076
rect 9306 15036 9312 15048
rect 9364 15036 9370 15088
rect 10704 15076 10732 15107
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 11940 15116 12173 15144
rect 11940 15104 11946 15116
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 15473 15147 15531 15153
rect 15473 15144 15485 15147
rect 12161 15107 12219 15113
rect 13464 15116 15485 15144
rect 12526 15076 12532 15088
rect 10704 15048 12532 15076
rect 12526 15036 12532 15048
rect 12584 15036 12590 15088
rect 13464 15076 13492 15116
rect 15473 15113 15485 15116
rect 15519 15113 15531 15147
rect 15473 15107 15531 15113
rect 16114 15104 16120 15156
rect 16172 15144 16178 15156
rect 16761 15147 16819 15153
rect 16761 15144 16773 15147
rect 16172 15116 16773 15144
rect 16172 15104 16178 15116
rect 16761 15113 16773 15116
rect 16807 15113 16819 15147
rect 16761 15107 16819 15113
rect 17770 15104 17776 15156
rect 17828 15144 17834 15156
rect 19794 15144 19800 15156
rect 17828 15116 19800 15144
rect 17828 15104 17834 15116
rect 19794 15104 19800 15116
rect 19852 15144 19858 15156
rect 19981 15147 20039 15153
rect 19981 15144 19993 15147
rect 19852 15116 19993 15144
rect 19852 15104 19858 15116
rect 19981 15113 19993 15116
rect 20027 15144 20039 15147
rect 20530 15144 20536 15156
rect 20027 15116 20536 15144
rect 20027 15113 20039 15116
rect 19981 15107 20039 15113
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 21174 15104 21180 15156
rect 21232 15144 21238 15156
rect 21453 15147 21511 15153
rect 21453 15144 21465 15147
rect 21232 15116 21465 15144
rect 21232 15104 21238 15116
rect 21453 15113 21465 15116
rect 21499 15113 21511 15147
rect 21453 15107 21511 15113
rect 21542 15104 21548 15156
rect 21600 15144 21606 15156
rect 22741 15147 22799 15153
rect 21600 15116 22094 15144
rect 21600 15104 21606 15116
rect 12820 15048 13492 15076
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 14977 5687 15011
rect 5629 14971 5687 14977
rect 5721 15011 5779 15017
rect 5721 14977 5733 15011
rect 5767 15008 5779 15011
rect 6178 15008 6184 15020
rect 5767 14980 6184 15008
rect 5767 14977 5779 14980
rect 5721 14971 5779 14977
rect 4488 14912 4752 14940
rect 4488 14900 4494 14912
rect 3200 14844 3648 14872
rect 3200 14832 3206 14844
rect 4522 14832 4528 14884
rect 4580 14872 4586 14884
rect 5261 14875 5319 14881
rect 5261 14872 5273 14875
rect 4580 14844 5273 14872
rect 4580 14832 4586 14844
rect 5261 14841 5273 14844
rect 5307 14841 5319 14875
rect 5261 14835 5319 14841
rect 3513 14807 3571 14813
rect 3513 14773 3525 14807
rect 3559 14804 3571 14807
rect 3970 14804 3976 14816
rect 3559 14776 3976 14804
rect 3559 14773 3571 14776
rect 3513 14767 3571 14773
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 4065 14807 4123 14813
rect 4065 14773 4077 14807
rect 4111 14804 4123 14807
rect 5350 14804 5356 14816
rect 4111 14776 5356 14804
rect 4111 14773 4123 14776
rect 4065 14767 4123 14773
rect 5350 14764 5356 14776
rect 5408 14804 5414 14816
rect 5644 14804 5672 14971
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 15008 9735 15011
rect 9766 15008 9772 15020
rect 9723 14980 9772 15008
rect 9723 14977 9735 14980
rect 9677 14971 9735 14977
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 10042 14968 10048 15020
rect 10100 15008 10106 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 10100 14980 10517 15008
rect 10100 14968 10106 14980
rect 10505 14977 10517 14980
rect 10551 14977 10563 15011
rect 10778 15008 10784 15020
rect 10739 14980 10784 15008
rect 10505 14971 10563 14977
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 12621 15011 12679 15017
rect 12621 14977 12633 15011
rect 12667 15008 12679 15011
rect 12710 15008 12716 15020
rect 12667 14980 12716 15008
rect 12667 14977 12679 14980
rect 12621 14971 12679 14977
rect 6638 14900 6644 14952
rect 6696 14940 6702 14952
rect 7374 14940 7380 14952
rect 6696 14912 7380 14940
rect 6696 14900 6702 14912
rect 7374 14900 7380 14912
rect 7432 14940 7438 14952
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 7432 14912 7481 14940
rect 7432 14900 7438 14912
rect 7469 14909 7481 14912
rect 7515 14909 7527 14943
rect 12360 14940 12388 14971
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 12820 15017 12848 15048
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 14977 12863 15011
rect 12805 14971 12863 14977
rect 13081 15011 13139 15017
rect 13081 14977 13093 15011
rect 13127 15008 13139 15011
rect 13262 15008 13268 15020
rect 13127 14980 13268 15008
rect 13127 14977 13139 14980
rect 13081 14971 13139 14977
rect 13096 14940 13124 14971
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 13464 15017 13492 15048
rect 13538 15036 13544 15088
rect 13596 15076 13602 15088
rect 16132 15076 16160 15104
rect 18782 15076 18788 15088
rect 13596 15048 13952 15076
rect 13596 15036 13602 15048
rect 13924 15017 13952 15048
rect 14476 15048 16160 15076
rect 18743 15048 18788 15076
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 14977 13507 15011
rect 13449 14971 13507 14977
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 14977 13783 15011
rect 13725 14971 13783 14977
rect 13909 15011 13967 15017
rect 13909 14977 13921 15011
rect 13955 14977 13967 15011
rect 14274 15008 14280 15020
rect 14235 14980 14280 15008
rect 13909 14971 13967 14977
rect 12360 14912 13124 14940
rect 7469 14903 7527 14909
rect 12342 14832 12348 14884
rect 12400 14872 12406 14884
rect 12437 14875 12495 14881
rect 12437 14872 12449 14875
rect 12400 14844 12449 14872
rect 12400 14832 12406 14844
rect 12437 14841 12449 14844
rect 12483 14841 12495 14875
rect 12437 14835 12495 14841
rect 12526 14832 12532 14884
rect 12584 14872 12590 14884
rect 13372 14872 13400 14971
rect 13740 14940 13768 14971
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 14476 15017 14504 15048
rect 18782 15036 18788 15048
rect 18840 15036 18846 15088
rect 19337 15079 19395 15085
rect 19337 15045 19349 15079
rect 19383 15076 19395 15079
rect 19518 15076 19524 15088
rect 19383 15048 19524 15076
rect 19383 15045 19395 15048
rect 19337 15039 19395 15045
rect 19518 15036 19524 15048
rect 19576 15076 19582 15088
rect 19576 15048 20576 15076
rect 19576 15036 19582 15048
rect 14461 15011 14519 15017
rect 14461 14977 14473 15011
rect 14507 14977 14519 15011
rect 14461 14971 14519 14977
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 14829 15011 14887 15017
rect 14608 14980 14653 15008
rect 14608 14968 14614 14980
rect 14829 14977 14841 15011
rect 14875 14977 14887 15011
rect 15010 15008 15016 15020
rect 14971 14980 15016 15008
rect 14829 14971 14887 14977
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 13740 14912 14657 14940
rect 14645 14909 14657 14912
rect 14691 14909 14703 14943
rect 14645 14903 14703 14909
rect 14090 14872 14096 14884
rect 12584 14844 12629 14872
rect 13372 14844 14096 14872
rect 12584 14832 12590 14844
rect 14090 14832 14096 14844
rect 14148 14832 14154 14884
rect 14844 14872 14872 14971
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 15197 15012 15255 15017
rect 15120 15011 15255 15012
rect 15120 14984 15209 15011
rect 14918 14900 14924 14952
rect 14976 14940 14982 14952
rect 15120 14940 15148 14984
rect 15197 14977 15209 14984
rect 15243 14977 15255 15011
rect 15562 15008 15568 15020
rect 15523 14980 15568 15008
rect 15197 14971 15255 14977
rect 15562 14968 15568 14980
rect 15620 14968 15626 15020
rect 16022 15008 16028 15020
rect 15983 14980 16028 15008
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 16132 14980 16712 15008
rect 14976 14912 15148 14940
rect 14976 14900 14982 14912
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 15841 14943 15899 14949
rect 15841 14940 15853 14943
rect 15344 14912 15853 14940
rect 15344 14900 15350 14912
rect 15841 14909 15853 14912
rect 15887 14940 15899 14943
rect 16132 14940 16160 14980
rect 15887 14912 16160 14940
rect 16301 14943 16359 14949
rect 15887 14909 15899 14912
rect 15841 14903 15899 14909
rect 16301 14909 16313 14943
rect 16347 14940 16359 14943
rect 16684 14940 16712 14980
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16816 14980 16865 15008
rect 16816 14968 16822 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 18966 15008 18972 15020
rect 18927 14980 18972 15008
rect 16853 14971 16911 14977
rect 18966 14968 18972 14980
rect 19024 14968 19030 15020
rect 19429 15011 19487 15017
rect 19429 15008 19441 15011
rect 19168 14980 19441 15008
rect 17218 14940 17224 14952
rect 16347 14912 16620 14940
rect 16684 14912 17224 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 16482 14872 16488 14884
rect 14844 14844 16488 14872
rect 16482 14832 16488 14844
rect 16540 14832 16546 14884
rect 16592 14872 16620 14912
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 17586 14872 17592 14884
rect 16592 14844 17592 14872
rect 17586 14832 17592 14844
rect 17644 14832 17650 14884
rect 19168 14881 19196 14980
rect 19429 14977 19441 14980
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 19794 14968 19800 15020
rect 19852 15008 19858 15020
rect 20548 15017 20576 15048
rect 20916 15048 21220 15076
rect 20714 15017 20720 15020
rect 19889 15011 19947 15017
rect 19889 15008 19901 15011
rect 19852 14980 19901 15008
rect 19852 14968 19858 14980
rect 19889 14977 19901 14980
rect 19935 14977 19947 15011
rect 20257 15011 20315 15017
rect 20257 15008 20269 15011
rect 19889 14971 19947 14977
rect 19996 14980 20269 15008
rect 19153 14875 19211 14881
rect 19153 14841 19165 14875
rect 19199 14841 19211 14875
rect 19153 14835 19211 14841
rect 19613 14875 19671 14881
rect 19613 14841 19625 14875
rect 19659 14872 19671 14875
rect 19702 14872 19708 14884
rect 19659 14844 19708 14872
rect 19659 14841 19671 14844
rect 19613 14835 19671 14841
rect 19702 14832 19708 14844
rect 19760 14832 19766 14884
rect 5813 14807 5871 14813
rect 5813 14804 5825 14807
rect 5408 14776 5825 14804
rect 5408 14764 5414 14776
rect 5813 14773 5825 14776
rect 5859 14773 5871 14807
rect 9214 14804 9220 14816
rect 9175 14776 9220 14804
rect 5813 14767 5871 14773
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 9861 14807 9919 14813
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 9950 14804 9956 14816
rect 9907 14776 9956 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 12158 14764 12164 14816
rect 12216 14804 12222 14816
rect 12802 14804 12808 14816
rect 12216 14776 12808 14804
rect 12216 14764 12222 14776
rect 12802 14764 12808 14776
rect 12860 14804 12866 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12860 14776 12909 14804
rect 12860 14764 12866 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 12897 14767 12955 14773
rect 13173 14807 13231 14813
rect 13173 14773 13185 14807
rect 13219 14804 13231 14807
rect 13262 14804 13268 14816
rect 13219 14776 13268 14804
rect 13219 14773 13231 14776
rect 13173 14767 13231 14773
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13354 14764 13360 14816
rect 13412 14804 13418 14816
rect 13541 14807 13599 14813
rect 13541 14804 13553 14807
rect 13412 14776 13553 14804
rect 13412 14764 13418 14776
rect 13541 14773 13553 14776
rect 13587 14773 13599 14807
rect 13541 14767 13599 14773
rect 14826 14764 14832 14816
rect 14884 14804 14890 14816
rect 16206 14804 16212 14816
rect 14884 14776 16212 14804
rect 14884 14764 14890 14776
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 19996 14804 20024 14980
rect 20257 14977 20269 14980
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 20533 15011 20591 15017
rect 20533 14977 20545 15011
rect 20579 14977 20591 15011
rect 20533 14971 20591 14977
rect 20677 15011 20720 15017
rect 20677 14977 20689 15011
rect 20772 15008 20778 15020
rect 20916 15008 20944 15048
rect 21082 15008 21088 15020
rect 20772 14980 20944 15008
rect 21043 14980 21088 15008
rect 20677 14971 20720 14977
rect 20456 14940 20484 14971
rect 20714 14968 20720 14971
rect 20772 14968 20778 14980
rect 21082 14968 21088 14980
rect 21140 14968 21146 15020
rect 21192 15008 21220 15048
rect 21453 15011 21511 15017
rect 21192 14980 21404 15008
rect 21376 14940 21404 14980
rect 21453 14977 21465 15011
rect 21499 15008 21511 15011
rect 21821 15011 21879 15017
rect 21821 15008 21833 15011
rect 21499 14980 21833 15008
rect 21499 14977 21511 14980
rect 21453 14971 21511 14977
rect 21821 14977 21833 14980
rect 21867 14977 21879 15011
rect 21821 14971 21879 14977
rect 21910 14968 21916 15020
rect 21968 15017 21974 15020
rect 22066 15017 22094 15116
rect 22741 15113 22753 15147
rect 22787 15144 22799 15147
rect 23382 15144 23388 15156
rect 22787 15116 23388 15144
rect 22787 15113 22799 15116
rect 22741 15107 22799 15113
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 24394 15144 24400 15156
rect 24320 15116 24400 15144
rect 24320 15076 24348 15116
rect 24394 15104 24400 15116
rect 24452 15104 24458 15156
rect 26326 15144 26332 15156
rect 26239 15116 26332 15144
rect 26326 15104 26332 15116
rect 26384 15144 26390 15156
rect 27522 15144 27528 15156
rect 26384 15116 27528 15144
rect 26384 15104 26390 15116
rect 27522 15104 27528 15116
rect 27580 15104 27586 15156
rect 24320 15048 25084 15076
rect 22278 15017 22284 15020
rect 21968 15011 22017 15017
rect 21968 14977 21971 15011
rect 22005 14977 22017 15011
rect 22066 15011 22152 15017
rect 22066 14980 22106 15011
rect 21968 14971 22017 14977
rect 22094 14977 22106 14980
rect 22140 14977 22152 15011
rect 22094 14971 22152 14977
rect 22241 15011 22284 15017
rect 22241 14977 22253 15011
rect 22241 14971 22284 14977
rect 21968 14968 21974 14971
rect 22256 14940 22284 14971
rect 22336 14968 22342 15020
rect 22554 15008 22560 15020
rect 22467 14980 22560 15008
rect 22554 14968 22560 14980
rect 22612 15008 22618 15020
rect 23566 15008 23572 15020
rect 22612 14980 23572 15008
rect 22612 14968 22618 14980
rect 23566 14968 23572 14980
rect 23624 14968 23630 15020
rect 24302 15008 24308 15020
rect 24263 14980 24308 15008
rect 24302 14968 24308 14980
rect 24360 15008 24366 15020
rect 25056 15017 25084 15048
rect 24581 15011 24639 15017
rect 24581 15008 24593 15011
rect 24360 14980 24593 15008
rect 24360 14968 24366 14980
rect 24581 14977 24593 14980
rect 24627 14977 24639 15011
rect 24581 14971 24639 14977
rect 25041 15011 25099 15017
rect 25041 14977 25053 15011
rect 25087 14977 25099 15011
rect 25041 14971 25099 14977
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 26513 15011 26571 15017
rect 26513 14977 26525 15011
rect 26559 15008 26571 15011
rect 26602 15008 26608 15020
rect 26559 14980 26608 15008
rect 26559 14977 26571 14980
rect 26513 14971 26571 14977
rect 20456 14912 21312 14940
rect 21376 14912 22284 14940
rect 20806 14872 20812 14884
rect 20767 14844 20812 14872
rect 20806 14832 20812 14844
rect 20864 14832 20870 14884
rect 21284 14872 21312 14912
rect 23474 14900 23480 14952
rect 23532 14940 23538 14952
rect 26160 14940 26188 14971
rect 26602 14968 26608 14980
rect 26660 14968 26666 15020
rect 23532 14912 26188 14940
rect 23532 14900 23538 14912
rect 22278 14872 22284 14884
rect 21284 14844 22284 14872
rect 22278 14832 22284 14844
rect 22336 14832 22342 14884
rect 22373 14875 22431 14881
rect 22373 14841 22385 14875
rect 22419 14872 22431 14875
rect 22830 14872 22836 14884
rect 22419 14844 22836 14872
rect 22419 14841 22431 14844
rect 22373 14835 22431 14841
rect 22830 14832 22836 14844
rect 22888 14832 22894 14884
rect 24486 14832 24492 14884
rect 24544 14872 24550 14884
rect 24857 14875 24915 14881
rect 24857 14872 24869 14875
rect 24544 14844 24869 14872
rect 24544 14832 24550 14844
rect 24857 14841 24869 14844
rect 24903 14841 24915 14875
rect 24857 14835 24915 14841
rect 21174 14804 21180 14816
rect 16448 14776 21180 14804
rect 16448 14764 16454 14776
rect 21174 14764 21180 14776
rect 21232 14764 21238 14816
rect 21269 14807 21327 14813
rect 21269 14773 21281 14807
rect 21315 14804 21327 14807
rect 21358 14804 21364 14816
rect 21315 14776 21364 14804
rect 21315 14773 21327 14776
rect 21269 14767 21327 14773
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 23934 14764 23940 14816
rect 23992 14804 23998 14816
rect 24765 14807 24823 14813
rect 24765 14804 24777 14807
rect 23992 14776 24777 14804
rect 23992 14764 23998 14776
rect 24765 14773 24777 14776
rect 24811 14804 24823 14807
rect 25222 14804 25228 14816
rect 24811 14776 25228 14804
rect 24811 14773 24823 14776
rect 24765 14767 24823 14773
rect 25222 14764 25228 14776
rect 25280 14764 25286 14816
rect 26697 14807 26755 14813
rect 26697 14773 26709 14807
rect 26743 14804 26755 14807
rect 26786 14804 26792 14816
rect 26743 14776 26792 14804
rect 26743 14773 26755 14776
rect 26697 14767 26755 14773
rect 26786 14764 26792 14776
rect 26844 14764 26850 14816
rect 1104 14714 29532 14736
rect 1104 14662 5688 14714
rect 5740 14662 5752 14714
rect 5804 14662 5816 14714
rect 5868 14662 5880 14714
rect 5932 14662 5944 14714
rect 5996 14662 15163 14714
rect 15215 14662 15227 14714
rect 15279 14662 15291 14714
rect 15343 14662 15355 14714
rect 15407 14662 15419 14714
rect 15471 14662 24639 14714
rect 24691 14662 24703 14714
rect 24755 14662 24767 14714
rect 24819 14662 24831 14714
rect 24883 14662 24895 14714
rect 24947 14662 29532 14714
rect 1104 14640 29532 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 3234 14600 3240 14612
rect 3195 14572 3240 14600
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 3786 14600 3792 14612
rect 3747 14572 3792 14600
rect 3786 14560 3792 14572
rect 3844 14560 3850 14612
rect 12986 14600 12992 14612
rect 12947 14572 12992 14600
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 13228 14572 13461 14600
rect 13228 14560 13234 14572
rect 13449 14569 13461 14572
rect 13495 14569 13507 14603
rect 13449 14563 13507 14569
rect 14090 14560 14096 14612
rect 14148 14600 14154 14612
rect 14185 14603 14243 14609
rect 14185 14600 14197 14603
rect 14148 14572 14197 14600
rect 14148 14560 14154 14572
rect 14185 14569 14197 14572
rect 14231 14569 14243 14603
rect 14185 14563 14243 14569
rect 14553 14603 14611 14609
rect 14553 14569 14565 14603
rect 14599 14600 14611 14603
rect 15010 14600 15016 14612
rect 14599 14572 15016 14600
rect 14599 14569 14611 14572
rect 14553 14563 14611 14569
rect 15010 14560 15016 14572
rect 15068 14560 15074 14612
rect 15562 14600 15568 14612
rect 15523 14572 15568 14600
rect 15562 14560 15568 14572
rect 15620 14560 15626 14612
rect 16758 14600 16764 14612
rect 16719 14572 16764 14600
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 19061 14603 19119 14609
rect 19061 14569 19073 14603
rect 19107 14600 19119 14603
rect 19429 14603 19487 14609
rect 19429 14600 19441 14603
rect 19107 14572 19441 14600
rect 19107 14569 19119 14572
rect 19061 14563 19119 14569
rect 19429 14569 19441 14572
rect 19475 14600 19487 14603
rect 19610 14600 19616 14612
rect 19475 14572 19616 14600
rect 19475 14569 19487 14572
rect 19429 14563 19487 14569
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 20349 14603 20407 14609
rect 20349 14569 20361 14603
rect 20395 14600 20407 14603
rect 20714 14600 20720 14612
rect 20395 14572 20720 14600
rect 20395 14569 20407 14572
rect 20349 14563 20407 14569
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 22278 14560 22284 14612
rect 22336 14600 22342 14612
rect 25774 14600 25780 14612
rect 22336 14572 25780 14600
rect 22336 14560 22342 14572
rect 25774 14560 25780 14572
rect 25832 14560 25838 14612
rect 9766 14424 9772 14476
rect 9824 14464 9830 14476
rect 11701 14467 11759 14473
rect 11701 14464 11713 14467
rect 9824 14436 11713 14464
rect 9824 14424 9830 14436
rect 11701 14433 11713 14436
rect 11747 14433 11759 14467
rect 12250 14464 12256 14476
rect 11701 14427 11759 14433
rect 11900 14436 12256 14464
rect 2038 14396 2044 14408
rect 1999 14368 2044 14396
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 3142 14396 3148 14408
rect 3103 14368 3148 14396
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4246 14396 4252 14408
rect 4019 14368 4252 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4246 14356 4252 14368
rect 4304 14356 4310 14408
rect 5074 14356 5080 14408
rect 5132 14396 5138 14408
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 5132 14368 5641 14396
rect 5132 14356 5138 14368
rect 5629 14365 5641 14368
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 5905 14399 5963 14405
rect 5905 14365 5917 14399
rect 5951 14396 5963 14399
rect 8205 14399 8263 14405
rect 8205 14396 8217 14399
rect 5951 14368 8217 14396
rect 5951 14365 5963 14368
rect 5905 14359 5963 14365
rect 8205 14365 8217 14368
rect 8251 14365 8263 14399
rect 8205 14359 8263 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14365 8355 14399
rect 8478 14396 8484 14408
rect 8439 14368 8484 14396
rect 8297 14359 8355 14365
rect 4338 14288 4344 14340
rect 4396 14328 4402 14340
rect 5920 14328 5948 14359
rect 4396 14300 5948 14328
rect 8312 14328 8340 14359
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 9950 14396 9956 14408
rect 9911 14368 9956 14396
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 11330 14396 11336 14408
rect 11291 14368 11336 14396
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 11900 14405 11928 14436
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 12529 14467 12587 14473
rect 12529 14433 12541 14467
rect 12575 14464 12587 14467
rect 13004 14464 13032 14560
rect 13262 14492 13268 14544
rect 13320 14532 13326 14544
rect 14458 14532 14464 14544
rect 13320 14504 14464 14532
rect 13320 14492 13326 14504
rect 14458 14492 14464 14504
rect 14516 14492 14522 14544
rect 16390 14532 16396 14544
rect 15212 14504 16396 14532
rect 12575 14436 13032 14464
rect 12575 14433 12587 14436
rect 12529 14427 12587 14433
rect 13998 14424 14004 14476
rect 14056 14464 14062 14476
rect 15212 14464 15240 14504
rect 16390 14492 16396 14504
rect 16448 14492 16454 14544
rect 16945 14535 17003 14541
rect 16945 14501 16957 14535
rect 16991 14501 17003 14535
rect 16945 14495 17003 14501
rect 15562 14464 15568 14476
rect 14056 14436 15240 14464
rect 15304 14436 15568 14464
rect 14056 14424 14062 14436
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 12710 14396 12716 14408
rect 12115 14368 12572 14396
rect 12671 14368 12716 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 8846 14328 8852 14340
rect 8312 14300 8852 14328
rect 4396 14288 4402 14300
rect 8846 14288 8852 14300
rect 8904 14288 8910 14340
rect 9122 14288 9128 14340
rect 9180 14328 9186 14340
rect 11624 14328 11652 14359
rect 12345 14331 12403 14337
rect 12345 14328 12357 14331
rect 9180 14300 10272 14328
rect 11624 14300 12357 14328
rect 9180 14288 9186 14300
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 5721 14263 5779 14269
rect 5721 14260 5733 14263
rect 5684 14232 5733 14260
rect 5684 14220 5690 14232
rect 5721 14229 5733 14232
rect 5767 14229 5779 14263
rect 10134 14260 10140 14272
rect 10095 14232 10140 14260
rect 5721 14223 5779 14229
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 10244 14260 10272 14300
rect 12345 14297 12357 14300
rect 12391 14297 12403 14331
rect 12544 14328 12572 14368
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 12802 14356 12808 14408
rect 12860 14396 12866 14408
rect 13081 14399 13139 14405
rect 12860 14368 12905 14396
rect 12860 14356 12866 14368
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13541 14399 13599 14405
rect 13541 14396 13553 14399
rect 13127 14368 13553 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 13541 14365 13553 14368
rect 13587 14396 13599 14399
rect 14366 14396 14372 14408
rect 13587 14368 14372 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 14366 14356 14372 14368
rect 14424 14356 14430 14408
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14396 14611 14399
rect 14642 14396 14648 14408
rect 14599 14368 14648 14396
rect 14599 14365 14611 14368
rect 14553 14359 14611 14365
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 15304 14405 15332 14436
rect 15562 14424 15568 14436
rect 15620 14424 15626 14476
rect 16960 14464 16988 14495
rect 22186 14492 22192 14544
rect 22244 14532 22250 14544
rect 23750 14532 23756 14544
rect 22244 14504 23756 14532
rect 22244 14492 22250 14504
rect 23750 14492 23756 14504
rect 23808 14492 23814 14544
rect 23842 14492 23848 14544
rect 23900 14532 23906 14544
rect 24121 14535 24179 14541
rect 24121 14532 24133 14535
rect 23900 14504 24133 14532
rect 23900 14492 23906 14504
rect 24121 14501 24133 14504
rect 24167 14501 24179 14535
rect 24121 14495 24179 14501
rect 24673 14535 24731 14541
rect 24673 14501 24685 14535
rect 24719 14532 24731 14535
rect 25038 14532 25044 14544
rect 24719 14504 25044 14532
rect 24719 14501 24731 14504
rect 24673 14495 24731 14501
rect 25038 14492 25044 14504
rect 25096 14492 25102 14544
rect 25317 14535 25375 14541
rect 25317 14501 25329 14535
rect 25363 14532 25375 14535
rect 25363 14504 25636 14532
rect 25363 14501 25375 14504
rect 25317 14495 25375 14501
rect 19429 14467 19487 14473
rect 19429 14464 19441 14467
rect 15764 14436 16988 14464
rect 17420 14436 19441 14464
rect 15289 14399 15347 14405
rect 15289 14365 15301 14399
rect 15335 14365 15347 14399
rect 15289 14359 15347 14365
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14396 15531 14399
rect 15654 14396 15660 14408
rect 15519 14368 15660 14396
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 15764 14405 15792 14436
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 15838 14356 15844 14408
rect 15896 14396 15902 14408
rect 15979 14399 16037 14405
rect 15979 14396 15991 14399
rect 15896 14368 15991 14396
rect 15896 14356 15902 14368
rect 15979 14365 15991 14368
rect 16025 14365 16037 14399
rect 16298 14396 16304 14408
rect 16259 14368 16304 14396
rect 15979 14359 16037 14365
rect 16298 14356 16304 14368
rect 16356 14396 16362 14408
rect 16393 14399 16451 14405
rect 16393 14396 16405 14399
rect 16356 14368 16405 14396
rect 16356 14356 16362 14368
rect 16393 14365 16405 14368
rect 16439 14365 16451 14399
rect 16393 14359 16451 14365
rect 16482 14356 16488 14408
rect 16540 14396 16546 14408
rect 17420 14405 17448 14436
rect 19429 14433 19441 14436
rect 19475 14433 19487 14467
rect 24486 14464 24492 14476
rect 19429 14427 19487 14433
rect 23584 14436 24492 14464
rect 23584 14408 23612 14436
rect 24486 14424 24492 14436
rect 24544 14424 24550 14476
rect 25056 14464 25084 14492
rect 25501 14467 25559 14473
rect 25501 14464 25513 14467
rect 25056 14436 25513 14464
rect 25501 14433 25513 14436
rect 25547 14433 25559 14467
rect 25608 14464 25636 14504
rect 25777 14467 25835 14473
rect 25777 14464 25789 14467
rect 25608 14436 25789 14464
rect 25501 14427 25559 14433
rect 25777 14433 25789 14436
rect 25823 14433 25835 14467
rect 25777 14427 25835 14433
rect 17405 14399 17463 14405
rect 17405 14396 17417 14399
rect 16540 14368 17417 14396
rect 16540 14356 16546 14368
rect 17405 14365 17417 14368
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 17678 14356 17684 14408
rect 17736 14396 17742 14408
rect 17865 14399 17923 14405
rect 17865 14396 17877 14399
rect 17736 14368 17877 14396
rect 17736 14356 17742 14368
rect 17865 14365 17877 14368
rect 17911 14396 17923 14399
rect 17954 14396 17960 14408
rect 17911 14368 17960 14396
rect 17911 14365 17923 14368
rect 17865 14359 17923 14365
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 19518 14356 19524 14408
rect 19576 14396 19582 14408
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 19576 14368 19809 14396
rect 19576 14356 19582 14368
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14365 20223 14399
rect 21358 14396 21364 14408
rect 21319 14368 21364 14396
rect 20165 14359 20223 14365
rect 12894 14328 12900 14340
rect 12544 14300 12900 14328
rect 12345 14291 12403 14297
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 13265 14331 13323 14337
rect 13265 14297 13277 14331
rect 13311 14328 13323 14331
rect 13446 14328 13452 14340
rect 13311 14300 13452 14328
rect 13311 14297 13323 14300
rect 13265 14291 13323 14297
rect 13446 14288 13452 14300
rect 13504 14288 13510 14340
rect 15105 14331 15163 14337
rect 15105 14297 15117 14331
rect 15151 14328 15163 14331
rect 15562 14328 15568 14340
rect 15151 14300 15568 14328
rect 15151 14297 15163 14300
rect 15105 14291 15163 14297
rect 15562 14288 15568 14300
rect 15620 14288 15626 14340
rect 16132 14300 16436 14328
rect 13354 14260 13360 14272
rect 10244 14232 13360 14260
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 13464 14260 13492 14288
rect 16132 14269 16160 14300
rect 16408 14272 16436 14300
rect 16666 14288 16672 14340
rect 16724 14328 16730 14340
rect 16770 14331 16828 14337
rect 16770 14328 16782 14331
rect 16724 14300 16782 14328
rect 16724 14288 16730 14300
rect 16770 14297 16782 14300
rect 16816 14297 16828 14331
rect 16770 14291 16828 14297
rect 17034 14288 17040 14340
rect 17092 14328 17098 14340
rect 17221 14331 17279 14337
rect 17221 14328 17233 14331
rect 17092 14300 17233 14328
rect 17092 14288 17098 14300
rect 17221 14297 17233 14300
rect 17267 14297 17279 14331
rect 17586 14328 17592 14340
rect 17499 14300 17592 14328
rect 17221 14291 17279 14297
rect 17586 14288 17592 14300
rect 17644 14328 17650 14340
rect 19061 14331 19119 14337
rect 19061 14328 19073 14331
rect 17644 14300 19073 14328
rect 17644 14288 17650 14300
rect 19061 14297 19073 14300
rect 19107 14297 19119 14331
rect 20180 14328 20208 14359
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14396 23259 14399
rect 23290 14396 23296 14408
rect 23247 14368 23296 14396
rect 23247 14365 23259 14368
rect 23201 14359 23259 14365
rect 23290 14356 23296 14368
rect 23348 14356 23354 14408
rect 23566 14396 23572 14408
rect 23479 14368 23572 14396
rect 23566 14356 23572 14368
rect 23624 14356 23630 14408
rect 23845 14399 23903 14405
rect 23845 14396 23857 14399
rect 23676 14368 23857 14396
rect 20254 14328 20260 14340
rect 19061 14291 19119 14297
rect 19628 14300 20260 14328
rect 16117 14263 16175 14269
rect 16117 14260 16129 14263
rect 13464 14232 16129 14260
rect 16117 14229 16129 14232
rect 16163 14229 16175 14263
rect 16117 14223 16175 14229
rect 16206 14220 16212 14272
rect 16264 14260 16270 14272
rect 16264 14232 16309 14260
rect 16264 14220 16270 14232
rect 16390 14220 16396 14272
rect 16448 14220 16454 14272
rect 17494 14220 17500 14272
rect 17552 14260 17558 14272
rect 19628 14269 19656 14300
rect 20254 14288 20260 14300
rect 20312 14288 20318 14340
rect 23676 14328 23704 14368
rect 23845 14365 23857 14368
rect 23891 14365 23903 14399
rect 23845 14359 23903 14365
rect 23934 14356 23940 14408
rect 23992 14405 23998 14408
rect 23992 14396 24000 14405
rect 24504 14396 24532 14424
rect 25222 14405 25228 14408
rect 24765 14399 24823 14405
rect 23992 14368 24037 14396
rect 24504 14392 24716 14396
rect 24765 14392 24777 14399
rect 24504 14368 24777 14392
rect 23992 14359 24000 14368
rect 24688 14365 24777 14368
rect 24811 14365 24823 14399
rect 24688 14364 24823 14365
rect 24765 14359 24823 14364
rect 25185 14399 25228 14405
rect 25185 14365 25197 14399
rect 25185 14359 25228 14365
rect 23992 14356 23998 14359
rect 25222 14356 25228 14359
rect 25280 14356 25286 14408
rect 27522 14356 27528 14408
rect 27580 14396 27586 14408
rect 27985 14399 28043 14405
rect 27985 14396 27997 14399
rect 27580 14368 27997 14396
rect 27580 14356 27586 14368
rect 27985 14365 27997 14368
rect 28031 14365 28043 14399
rect 28353 14399 28411 14405
rect 28353 14396 28365 14399
rect 27985 14359 28043 14365
rect 28184 14368 28365 14396
rect 23032 14300 23704 14328
rect 17773 14263 17831 14269
rect 17773 14260 17785 14263
rect 17552 14232 17785 14260
rect 17552 14220 17558 14232
rect 17773 14229 17785 14232
rect 17819 14229 17831 14263
rect 17773 14223 17831 14229
rect 19613 14263 19671 14269
rect 19613 14229 19625 14263
rect 19659 14229 19671 14263
rect 21542 14260 21548 14272
rect 21503 14232 21548 14260
rect 19613 14223 19671 14229
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 22646 14220 22652 14272
rect 22704 14260 22710 14272
rect 23032 14269 23060 14300
rect 23750 14288 23756 14340
rect 23808 14328 23814 14340
rect 24486 14328 24492 14340
rect 23808 14300 23853 14328
rect 24447 14300 24492 14328
rect 23808 14288 23814 14300
rect 24486 14288 24492 14300
rect 24544 14288 24550 14340
rect 24946 14328 24952 14340
rect 24907 14300 24952 14328
rect 24946 14288 24952 14300
rect 25004 14288 25010 14340
rect 25041 14331 25099 14337
rect 25041 14297 25053 14331
rect 25087 14297 25099 14331
rect 25041 14291 25099 14297
rect 23017 14263 23075 14269
rect 23017 14260 23029 14263
rect 22704 14232 23029 14260
rect 22704 14220 22710 14232
rect 23017 14229 23029 14232
rect 23063 14229 23075 14263
rect 23017 14223 23075 14229
rect 23385 14263 23443 14269
rect 23385 14229 23397 14263
rect 23431 14260 23443 14263
rect 24394 14260 24400 14272
rect 23431 14232 24400 14260
rect 23431 14229 23443 14232
rect 23385 14223 23443 14229
rect 24394 14220 24400 14232
rect 24452 14220 24458 14272
rect 25056 14260 25084 14291
rect 26786 14288 26792 14340
rect 26844 14288 26850 14340
rect 27249 14263 27307 14269
rect 27249 14260 27261 14263
rect 25056 14232 27261 14260
rect 27249 14229 27261 14232
rect 27295 14260 27307 14263
rect 27522 14260 27528 14272
rect 27295 14232 27528 14260
rect 27295 14229 27307 14232
rect 27249 14223 27307 14229
rect 27522 14220 27528 14232
rect 27580 14220 27586 14272
rect 28184 14269 28212 14368
rect 28353 14365 28365 14368
rect 28399 14365 28411 14399
rect 28353 14359 28411 14365
rect 28169 14263 28227 14269
rect 28169 14229 28181 14263
rect 28215 14229 28227 14263
rect 28169 14223 28227 14229
rect 28537 14263 28595 14269
rect 28537 14229 28549 14263
rect 28583 14260 28595 14263
rect 28626 14260 28632 14272
rect 28583 14232 28632 14260
rect 28583 14229 28595 14232
rect 28537 14223 28595 14229
rect 28626 14220 28632 14232
rect 28684 14220 28690 14272
rect 1104 14170 29532 14192
rect 1104 14118 10425 14170
rect 10477 14118 10489 14170
rect 10541 14118 10553 14170
rect 10605 14118 10617 14170
rect 10669 14118 10681 14170
rect 10733 14118 19901 14170
rect 19953 14118 19965 14170
rect 20017 14118 20029 14170
rect 20081 14118 20093 14170
rect 20145 14118 20157 14170
rect 20209 14118 29532 14170
rect 1104 14096 29532 14118
rect 3329 14059 3387 14065
rect 3329 14025 3341 14059
rect 3375 14056 3387 14059
rect 3418 14056 3424 14068
rect 3375 14028 3424 14056
rect 3375 14025 3387 14028
rect 3329 14019 3387 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 4890 14056 4896 14068
rect 3896 14028 4896 14056
rect 3896 13997 3924 14028
rect 4890 14016 4896 14028
rect 4948 14016 4954 14068
rect 5074 14056 5080 14068
rect 5035 14028 5080 14056
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 6181 14059 6239 14065
rect 6181 14025 6193 14059
rect 6227 14025 6239 14059
rect 6181 14019 6239 14025
rect 8021 14059 8079 14065
rect 8021 14025 8033 14059
rect 8067 14056 8079 14059
rect 8478 14056 8484 14068
rect 8067 14028 8484 14056
rect 8067 14025 8079 14028
rect 8021 14019 8079 14025
rect 3881 13991 3939 13997
rect 3881 13957 3893 13991
rect 3927 13957 3939 13991
rect 3881 13951 3939 13957
rect 4430 13948 4436 14000
rect 4488 13948 4494 14000
rect 4706 13988 4712 14000
rect 4632 13960 4712 13988
rect 4434 13945 4492 13948
rect 2866 13880 2872 13932
rect 2924 13920 2930 13932
rect 3145 13923 3203 13929
rect 3145 13920 3157 13923
rect 2924 13892 3157 13920
rect 2924 13880 2930 13892
rect 3145 13889 3157 13892
rect 3191 13889 3203 13923
rect 3694 13920 3700 13932
rect 3655 13892 3700 13920
rect 3145 13883 3203 13889
rect 3694 13880 3700 13892
rect 3752 13880 3758 13932
rect 4154 13920 4160 13932
rect 4115 13892 4160 13920
rect 4154 13880 4160 13892
rect 4212 13880 4218 13932
rect 4338 13920 4344 13932
rect 4299 13892 4344 13920
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 4434 13911 4446 13945
rect 4480 13911 4492 13945
rect 4434 13905 4492 13911
rect 4542 13923 4600 13929
rect 4542 13889 4554 13923
rect 4588 13920 4600 13923
rect 4632 13920 4660 13960
rect 4706 13948 4712 13960
rect 4764 13988 4770 14000
rect 5092 13988 5120 14016
rect 4764 13960 5120 13988
rect 4764 13948 4770 13960
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 5813 13991 5871 13997
rect 5813 13988 5825 13991
rect 5592 13960 5825 13988
rect 5592 13948 5598 13960
rect 5813 13957 5825 13960
rect 5859 13957 5871 13991
rect 6196 13988 6224 14019
rect 8478 14016 8484 14028
rect 8536 14056 8542 14068
rect 9122 14056 9128 14068
rect 8536 14028 8616 14056
rect 8536 14016 8542 14028
rect 8588 13997 8616 14028
rect 8772 14028 9128 14056
rect 8772 13997 8800 14028
rect 9122 14016 9128 14028
rect 9180 14056 9186 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 9180 14028 11345 14056
rect 9180 14016 9186 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11333 14019 11391 14025
rect 12529 14059 12587 14065
rect 12529 14025 12541 14059
rect 12575 14056 12587 14059
rect 12710 14056 12716 14068
rect 12575 14028 12716 14056
rect 12575 14025 12587 14028
rect 12529 14019 12587 14025
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 13081 14059 13139 14065
rect 13081 14025 13093 14059
rect 13127 14025 13139 14059
rect 13081 14019 13139 14025
rect 13173 14059 13231 14065
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 14366 14056 14372 14068
rect 13219 14028 14372 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 6886 13991 6944 13997
rect 6886 13988 6898 13991
rect 6196 13960 6898 13988
rect 5813 13951 5871 13957
rect 6886 13957 6898 13960
rect 6932 13957 6944 13991
rect 6886 13951 6944 13957
rect 8573 13991 8631 13997
rect 8573 13957 8585 13991
rect 8619 13957 8631 13991
rect 8573 13951 8631 13957
rect 8757 13991 8815 13997
rect 8757 13957 8769 13991
rect 8803 13957 8815 13991
rect 9674 13988 9680 14000
rect 8757 13951 8815 13957
rect 9140 13960 9680 13988
rect 4798 13920 4804 13932
rect 4588 13892 4660 13920
rect 4759 13892 4804 13920
rect 4588 13889 4600 13892
rect 4542 13883 4600 13889
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13920 4951 13923
rect 4982 13920 4988 13932
rect 4939 13892 4988 13920
rect 4939 13889 4951 13892
rect 4893 13883 4951 13889
rect 4982 13880 4988 13892
rect 5040 13880 5046 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5500 13892 5733 13920
rect 5500 13880 5506 13892
rect 5721 13889 5733 13892
rect 5767 13889 5779 13923
rect 8386 13920 8392 13932
rect 8347 13892 8392 13920
rect 5721 13883 5779 13889
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 8846 13920 8852 13932
rect 8807 13892 8852 13920
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9140 13929 9168 13960
rect 9674 13948 9680 13960
rect 9732 13948 9738 14000
rect 10134 13948 10140 14000
rect 10192 13948 10198 14000
rect 12342 13988 12348 14000
rect 12176 13960 12348 13988
rect 9125 13923 9183 13929
rect 9125 13889 9137 13923
rect 9171 13889 9183 13923
rect 11057 13923 11115 13929
rect 11057 13920 11069 13923
rect 9125 13883 9183 13889
rect 10888 13892 11069 13920
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13852 4123 13855
rect 4246 13852 4252 13864
rect 4111 13824 4252 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 4246 13812 4252 13824
rect 4304 13852 4310 13864
rect 5626 13852 5632 13864
rect 4304 13824 4936 13852
rect 5587 13824 5632 13852
rect 4304 13812 4310 13824
rect 4908 13796 4936 13824
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 6638 13852 6644 13864
rect 6599 13824 6644 13852
rect 6638 13812 6644 13824
rect 6696 13812 6702 13864
rect 9401 13855 9459 13861
rect 9401 13821 9413 13855
rect 9447 13852 9459 13855
rect 9766 13852 9772 13864
rect 9447 13824 9772 13852
rect 9447 13821 9459 13824
rect 9401 13815 9459 13821
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 10888 13861 10916 13892
rect 11057 13889 11069 13892
rect 11103 13889 11115 13923
rect 11057 13883 11115 13889
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12176 13929 12204 13960
rect 12342 13948 12348 13960
rect 12400 13948 12406 14000
rect 13096 13988 13124 14019
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 14844 14028 15485 14056
rect 14844 13997 14872 14028
rect 15473 14025 15485 14028
rect 15519 14056 15531 14059
rect 15746 14056 15752 14068
rect 15519 14028 15752 14056
rect 15519 14025 15531 14028
rect 15473 14019 15531 14025
rect 15746 14016 15752 14028
rect 15804 14016 15810 14068
rect 15841 14059 15899 14065
rect 15841 14025 15853 14059
rect 15887 14056 15899 14059
rect 15930 14056 15936 14068
rect 15887 14028 15936 14056
rect 15887 14025 15899 14028
rect 15841 14019 15899 14025
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16669 14059 16727 14065
rect 16669 14025 16681 14059
rect 16715 14025 16727 14059
rect 16669 14019 16727 14025
rect 14645 13991 14703 13997
rect 14645 13988 14657 13991
rect 13096 13960 14657 13988
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 12032 13892 12081 13920
rect 12032 13880 12038 13892
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12492 13892 13001 13920
rect 12492 13880 12498 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 10873 13855 10931 13861
rect 10873 13821 10885 13855
rect 10919 13821 10931 13855
rect 10873 13815 10931 13821
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 11330 13852 11336 13864
rect 11195 13824 11336 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 11330 13812 11336 13824
rect 11388 13852 11394 13864
rect 11698 13852 11704 13864
rect 11388 13824 11704 13852
rect 11388 13812 11394 13824
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 12345 13855 12403 13861
rect 12345 13821 12357 13855
rect 12391 13852 12403 13855
rect 13096 13852 13124 13960
rect 14645 13957 14657 13960
rect 14691 13957 14703 13991
rect 14645 13951 14703 13957
rect 14829 13991 14887 13997
rect 14829 13957 14841 13991
rect 14875 13957 14887 13991
rect 15010 13988 15016 14000
rect 14971 13960 15016 13988
rect 14829 13951 14887 13957
rect 15010 13948 15016 13960
rect 15068 13948 15074 14000
rect 16298 13988 16304 14000
rect 16259 13960 16304 13988
rect 16298 13948 16304 13960
rect 16356 13948 16362 14000
rect 16390 13948 16396 14000
rect 16448 13988 16454 14000
rect 16684 13988 16712 14019
rect 17218 14016 17224 14068
rect 17276 14056 17282 14068
rect 19518 14056 19524 14068
rect 17276 14028 19524 14056
rect 17276 14016 17282 14028
rect 19518 14016 19524 14028
rect 19576 14016 19582 14068
rect 20714 14016 20720 14068
rect 20772 14016 20778 14068
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 21269 14059 21327 14065
rect 21269 14056 21281 14059
rect 21232 14028 21281 14056
rect 21232 14016 21238 14028
rect 21269 14025 21281 14028
rect 21315 14025 21327 14059
rect 22370 14056 22376 14068
rect 21269 14019 21327 14025
rect 22066 14028 22376 14056
rect 16448 13960 16712 13988
rect 16448 13948 16454 13960
rect 16942 13948 16948 14000
rect 17000 13988 17006 14000
rect 17313 13991 17371 13997
rect 17313 13988 17325 13991
rect 17000 13960 17325 13988
rect 17000 13948 17006 13960
rect 17313 13957 17325 13960
rect 17359 13957 17371 13991
rect 17313 13951 17371 13957
rect 18690 13948 18696 14000
rect 18748 13948 18754 14000
rect 20732 13988 20760 14016
rect 20635 13960 20760 13988
rect 20809 13991 20867 13997
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 13998 13920 14004 13932
rect 13403 13892 14004 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 14093 13923 14151 13929
rect 14093 13889 14105 13923
rect 14139 13889 14151 13923
rect 14093 13883 14151 13889
rect 12391 13824 13124 13852
rect 12391 13821 12403 13824
rect 12345 13815 12403 13821
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 14108 13852 14136 13883
rect 14734 13880 14740 13932
rect 14792 13920 14798 13932
rect 15105 13923 15163 13929
rect 15105 13920 15117 13923
rect 14792 13892 15117 13920
rect 14792 13880 14798 13892
rect 15105 13889 15117 13892
rect 15151 13889 15163 13923
rect 15105 13883 15163 13889
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13920 15623 13923
rect 15654 13920 15660 13932
rect 15611 13892 15660 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 15930 13920 15936 13932
rect 15891 13892 15936 13920
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 16132 13852 16160 13883
rect 16758 13880 16764 13932
rect 16816 13920 16822 13932
rect 16853 13923 16911 13929
rect 16853 13920 16865 13923
rect 16816 13892 16865 13920
rect 16816 13880 16822 13892
rect 16853 13889 16865 13892
rect 16899 13889 16911 13923
rect 17034 13920 17040 13932
rect 16995 13892 17040 13920
rect 16853 13883 16911 13889
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 17218 13920 17224 13932
rect 17179 13892 17224 13920
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 17494 13929 17500 13932
rect 17457 13923 17500 13929
rect 17457 13889 17469 13923
rect 17457 13883 17500 13889
rect 17494 13880 17500 13883
rect 17552 13880 17558 13932
rect 17770 13920 17776 13932
rect 17731 13892 17776 13920
rect 17770 13880 17776 13892
rect 17828 13880 17834 13932
rect 20073 13923 20131 13929
rect 20073 13889 20085 13923
rect 20119 13920 20131 13923
rect 20254 13920 20260 13932
rect 20119 13892 20260 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 20635 13929 20663 13960
rect 20809 13957 20821 13991
rect 20855 13988 20867 13991
rect 22066 13988 22094 14028
rect 22370 14016 22376 14028
rect 22428 14056 22434 14068
rect 23750 14056 23756 14068
rect 22428 14028 23756 14056
rect 22428 14016 22434 14028
rect 23750 14016 23756 14028
rect 23808 14016 23814 14068
rect 24213 14059 24271 14065
rect 24213 14025 24225 14059
rect 24259 14025 24271 14059
rect 24213 14019 24271 14025
rect 24228 13988 24256 14019
rect 24946 14016 24952 14068
rect 25004 14056 25010 14068
rect 25774 14056 25780 14068
rect 25004 14028 25780 14056
rect 25004 14016 25010 14028
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 26602 14056 26608 14068
rect 26563 14028 26608 14056
rect 26602 14016 26608 14028
rect 26660 14016 26666 14068
rect 27430 14016 27436 14068
rect 27488 14056 27494 14068
rect 29086 14056 29092 14068
rect 27488 14028 29092 14056
rect 27488 14016 27494 14028
rect 29086 14016 29092 14028
rect 29144 14016 29150 14068
rect 27614 13988 27620 14000
rect 20855 13960 22094 13988
rect 23414 13960 24256 13988
rect 27575 13960 27620 13988
rect 20855 13957 20867 13960
rect 20809 13951 20867 13957
rect 27614 13948 27620 13960
rect 27672 13948 27678 14000
rect 28626 13948 28632 14000
rect 28684 13948 28690 14000
rect 20620 13923 20678 13929
rect 20620 13889 20632 13923
rect 20666 13889 20678 13923
rect 20620 13883 20678 13889
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 20993 13923 21051 13929
rect 20772 13892 20817 13920
rect 20772 13880 20778 13892
rect 20993 13889 21005 13923
rect 21039 13920 21051 13923
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 21039 13892 21097 13920
rect 21039 13889 21051 13892
rect 20993 13883 21051 13889
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 24394 13920 24400 13932
rect 24355 13892 24400 13920
rect 21085 13883 21143 13889
rect 16390 13852 16396 13864
rect 13688 13824 14136 13852
rect 14200 13824 16396 13852
rect 13688 13812 13694 13824
rect 4890 13744 4896 13796
rect 4948 13744 4954 13796
rect 5644 13784 5672 13812
rect 6086 13784 6092 13796
rect 5644 13756 6092 13784
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 12802 13784 12808 13796
rect 12763 13756 12808 13784
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 5258 13716 5264 13728
rect 3936 13688 5264 13716
rect 3936 13676 3942 13688
rect 5258 13676 5264 13688
rect 5316 13676 5322 13728
rect 9030 13716 9036 13728
rect 8991 13688 9036 13716
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 11333 13719 11391 13725
rect 11333 13685 11345 13719
rect 11379 13716 11391 13719
rect 14200 13716 14228 13824
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17604 13824 18061 13852
rect 15010 13744 15016 13796
rect 15068 13784 15074 13796
rect 15289 13787 15347 13793
rect 15289 13784 15301 13787
rect 15068 13756 15301 13784
rect 15068 13744 15074 13756
rect 15289 13753 15301 13756
rect 15335 13784 15347 13787
rect 16482 13784 16488 13796
rect 15335 13756 16488 13784
rect 15335 13753 15347 13756
rect 15289 13747 15347 13753
rect 16482 13744 16488 13756
rect 16540 13744 16546 13796
rect 17604 13793 17632 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 20165 13855 20223 13861
rect 20165 13821 20177 13855
rect 20211 13852 20223 13855
rect 21008 13852 21036 13883
rect 24394 13880 24400 13892
rect 24452 13880 24458 13932
rect 26326 13880 26332 13932
rect 26384 13920 26390 13932
rect 26421 13923 26479 13929
rect 26421 13920 26433 13923
rect 26384 13892 26433 13920
rect 26384 13880 26390 13892
rect 26421 13889 26433 13892
rect 26467 13889 26479 13923
rect 26421 13883 26479 13889
rect 21361 13855 21419 13861
rect 21361 13852 21373 13855
rect 20211 13824 21036 13852
rect 21100 13824 21373 13852
rect 20211 13821 20223 13824
rect 20165 13815 20223 13821
rect 17589 13787 17647 13793
rect 17589 13753 17601 13787
rect 17635 13753 17647 13787
rect 17589 13747 17647 13753
rect 20714 13744 20720 13796
rect 20772 13784 20778 13796
rect 21100 13784 21128 13824
rect 21361 13821 21373 13824
rect 21407 13852 21419 13855
rect 22278 13852 22284 13864
rect 21407 13824 22284 13852
rect 21407 13821 21419 13824
rect 21361 13815 21419 13821
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 22373 13855 22431 13861
rect 22373 13821 22385 13855
rect 22419 13852 22431 13855
rect 22646 13852 22652 13864
rect 22419 13824 22652 13852
rect 22419 13821 22431 13824
rect 22373 13815 22431 13821
rect 22646 13812 22652 13824
rect 22704 13812 22710 13864
rect 23842 13852 23848 13864
rect 23803 13824 23848 13852
rect 23842 13812 23848 13824
rect 23900 13812 23906 13864
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13852 24179 13855
rect 25038 13852 25044 13864
rect 24167 13824 25044 13852
rect 24167 13821 24179 13824
rect 24121 13815 24179 13821
rect 25038 13812 25044 13824
rect 25096 13852 25102 13864
rect 27341 13855 27399 13861
rect 27341 13852 27353 13855
rect 25096 13824 27353 13852
rect 25096 13812 25102 13824
rect 27341 13821 27353 13824
rect 27387 13821 27399 13855
rect 27341 13815 27399 13821
rect 20772 13756 21128 13784
rect 20772 13744 20778 13756
rect 11379 13688 14228 13716
rect 14277 13719 14335 13725
rect 11379 13685 11391 13688
rect 11333 13679 11391 13685
rect 14277 13685 14289 13719
rect 14323 13716 14335 13719
rect 14458 13716 14464 13728
rect 14323 13688 14464 13716
rect 14323 13685 14335 13688
rect 14277 13679 14335 13685
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 20441 13719 20499 13725
rect 20441 13685 20453 13719
rect 20487 13716 20499 13719
rect 20806 13716 20812 13728
rect 20487 13688 20812 13716
rect 20487 13685 20499 13688
rect 20441 13679 20499 13685
rect 20806 13676 20812 13688
rect 20864 13676 20870 13728
rect 1104 13626 29532 13648
rect 1104 13574 5688 13626
rect 5740 13574 5752 13626
rect 5804 13574 5816 13626
rect 5868 13574 5880 13626
rect 5932 13574 5944 13626
rect 5996 13574 15163 13626
rect 15215 13574 15227 13626
rect 15279 13574 15291 13626
rect 15343 13574 15355 13626
rect 15407 13574 15419 13626
rect 15471 13574 24639 13626
rect 24691 13574 24703 13626
rect 24755 13574 24767 13626
rect 24819 13574 24831 13626
rect 24883 13574 24895 13626
rect 24947 13574 29532 13626
rect 1104 13552 29532 13574
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 5040 13484 8708 13512
rect 5040 13472 5046 13484
rect 3418 13404 3424 13456
rect 3476 13444 3482 13456
rect 5258 13444 5264 13456
rect 3476 13416 5264 13444
rect 3476 13404 3482 13416
rect 5258 13404 5264 13416
rect 5316 13404 5322 13456
rect 5445 13447 5503 13453
rect 5445 13413 5457 13447
rect 5491 13444 5503 13447
rect 5534 13444 5540 13456
rect 5491 13416 5540 13444
rect 5491 13413 5503 13416
rect 5445 13407 5503 13413
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 8021 13447 8079 13453
rect 8021 13413 8033 13447
rect 8067 13444 8079 13447
rect 8386 13444 8392 13456
rect 8067 13416 8392 13444
rect 8067 13413 8079 13416
rect 8021 13407 8079 13413
rect 8386 13404 8392 13416
rect 8444 13404 8450 13456
rect 4154 13376 4160 13388
rect 3344 13348 4160 13376
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 3344 13317 3372 13348
rect 4154 13336 4160 13348
rect 4212 13336 4218 13388
rect 4617 13379 4675 13385
rect 4617 13345 4629 13379
rect 4663 13376 4675 13379
rect 5997 13379 6055 13385
rect 4663 13348 5212 13376
rect 4663 13345 4675 13348
rect 4617 13339 4675 13345
rect 2869 13311 2927 13317
rect 2869 13308 2881 13311
rect 2832 13280 2881 13308
rect 2832 13268 2838 13280
rect 2869 13277 2881 13280
rect 2915 13277 2927 13311
rect 2869 13271 2927 13277
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13277 3203 13311
rect 3145 13271 3203 13277
rect 3329 13311 3387 13317
rect 3329 13277 3341 13311
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 3605 13311 3663 13317
rect 3605 13277 3617 13311
rect 3651 13308 3663 13311
rect 4338 13308 4344 13320
rect 3651 13280 4344 13308
rect 3651 13277 3663 13280
rect 3605 13271 3663 13277
rect 2406 13200 2412 13252
rect 2464 13240 2470 13252
rect 2602 13243 2660 13249
rect 2602 13240 2614 13243
rect 2464 13212 2614 13240
rect 2464 13200 2470 13212
rect 2602 13209 2614 13212
rect 2648 13209 2660 13243
rect 2961 13243 3019 13249
rect 2961 13240 2973 13243
rect 2602 13203 2660 13209
rect 2746 13212 2973 13240
rect 2746 13184 2774 13212
rect 2961 13209 2973 13212
rect 3007 13209 3019 13243
rect 3160 13240 3188 13271
rect 3620 13240 3648 13271
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 4706 13308 4712 13320
rect 4667 13280 4712 13308
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 4798 13268 4804 13320
rect 4856 13308 4862 13320
rect 5097 13311 5155 13317
rect 4856 13280 4901 13308
rect 4856 13268 4862 13280
rect 5097 13277 5109 13311
rect 5143 13277 5155 13311
rect 5184 13308 5212 13348
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6086 13376 6092 13388
rect 6043 13348 6092 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 8680 13385 8708 13484
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8904 13484 9045 13512
rect 8904 13472 8910 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 9033 13475 9091 13481
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11848 13484 12081 13512
rect 11848 13472 11854 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 12253 13515 12311 13521
rect 12253 13481 12265 13515
rect 12299 13512 12311 13515
rect 12434 13512 12440 13524
rect 12299 13484 12440 13512
rect 12299 13481 12311 13484
rect 12253 13475 12311 13481
rect 12084 13444 12112 13475
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 16390 13472 16396 13524
rect 16448 13512 16454 13524
rect 18690 13512 18696 13524
rect 16448 13484 17724 13512
rect 18651 13484 18696 13512
rect 16448 13472 16454 13484
rect 14458 13444 14464 13456
rect 12084 13416 14464 13444
rect 14458 13404 14464 13416
rect 14516 13404 14522 13456
rect 17126 13404 17132 13456
rect 17184 13444 17190 13456
rect 17313 13447 17371 13453
rect 17313 13444 17325 13447
rect 17184 13416 17325 13444
rect 17184 13404 17190 13416
rect 17313 13413 17325 13416
rect 17359 13413 17371 13447
rect 17313 13407 17371 13413
rect 8665 13379 8723 13385
rect 8665 13345 8677 13379
rect 8711 13345 8723 13379
rect 8665 13339 8723 13345
rect 15654 13336 15660 13388
rect 15712 13336 15718 13388
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 16761 13379 16819 13385
rect 16761 13376 16773 13379
rect 16632 13348 16773 13376
rect 16632 13336 16638 13348
rect 16761 13345 16773 13348
rect 16807 13345 16819 13379
rect 16761 13339 16819 13345
rect 16853 13379 16911 13385
rect 16853 13345 16865 13379
rect 16899 13376 16911 13379
rect 17494 13376 17500 13388
rect 16899 13348 17500 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 5534 13308 5540 13320
rect 5184 13280 5540 13308
rect 5097 13271 5155 13277
rect 3160 13212 3648 13240
rect 4724 13240 4752 13268
rect 5009 13243 5067 13249
rect 5009 13240 5021 13243
rect 4724 13212 5021 13240
rect 2961 13203 3019 13209
rect 5009 13209 5021 13212
rect 5055 13209 5067 13243
rect 5009 13203 5067 13209
rect 5112 13184 5140 13271
rect 5534 13268 5540 13280
rect 5592 13308 5598 13320
rect 6638 13308 6644 13320
rect 5592 13280 6132 13308
rect 6599 13280 6644 13308
rect 5592 13268 5598 13280
rect 5258 13200 5264 13252
rect 5316 13240 5322 13252
rect 6104 13249 6132 13280
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 8386 13308 8392 13320
rect 8347 13280 8392 13308
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13308 8631 13311
rect 9030 13308 9036 13320
rect 8619 13280 9036 13308
rect 8619 13277 8631 13280
rect 8573 13271 8631 13277
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13308 9183 13311
rect 11882 13308 11888 13320
rect 9171 13280 9352 13308
rect 11843 13280 11888 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 5353 13243 5411 13249
rect 5353 13240 5365 13243
rect 5316 13212 5365 13240
rect 5316 13200 5322 13212
rect 5353 13209 5365 13212
rect 5399 13209 5411 13243
rect 5353 13203 5411 13209
rect 6089 13243 6147 13249
rect 6089 13209 6101 13243
rect 6135 13209 6147 13243
rect 6886 13243 6944 13249
rect 6886 13240 6898 13243
rect 6089 13203 6147 13209
rect 6564 13212 6898 13240
rect 1489 13175 1547 13181
rect 1489 13141 1501 13175
rect 1535 13172 1547 13175
rect 1762 13172 1768 13184
rect 1535 13144 1768 13172
rect 1535 13141 1547 13144
rect 1489 13135 1547 13141
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 2682 13132 2688 13184
rect 2740 13144 2774 13184
rect 3513 13175 3571 13181
rect 2740 13132 2746 13144
rect 3513 13141 3525 13175
rect 3559 13172 3571 13175
rect 3694 13172 3700 13184
rect 3559 13144 3700 13172
rect 3559 13141 3571 13144
rect 3513 13135 3571 13141
rect 3694 13132 3700 13144
rect 3752 13172 3758 13184
rect 4706 13172 4712 13184
rect 3752 13144 4712 13172
rect 3752 13132 3758 13144
rect 4706 13132 4712 13144
rect 4764 13172 4770 13184
rect 4893 13175 4951 13181
rect 4893 13172 4905 13175
rect 4764 13144 4905 13172
rect 4764 13132 4770 13144
rect 4893 13141 4905 13144
rect 4939 13141 4951 13175
rect 4893 13135 4951 13141
rect 5094 13132 5100 13184
rect 5152 13132 5158 13184
rect 6178 13132 6184 13184
rect 6236 13172 6242 13184
rect 6564 13181 6592 13212
rect 6886 13209 6898 13212
rect 6932 13209 6944 13243
rect 6886 13203 6944 13209
rect 9324 13184 9352 13280
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 11974 13268 11980 13320
rect 12032 13308 12038 13320
rect 12032 13280 12077 13308
rect 12032 13268 12038 13280
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 13633 13311 13691 13317
rect 13633 13308 13645 13311
rect 13504 13280 13645 13308
rect 13504 13268 13510 13280
rect 13633 13277 13645 13280
rect 13679 13277 13691 13311
rect 15562 13308 15568 13320
rect 15523 13280 15568 13308
rect 13633 13271 13691 13277
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 15672 13308 15700 13336
rect 17057 13311 17115 13317
rect 17057 13308 17069 13311
rect 15672 13280 17069 13308
rect 17057 13277 17069 13280
rect 17103 13277 17115 13311
rect 17057 13271 17115 13277
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13308 17371 13311
rect 17589 13311 17647 13317
rect 17589 13308 17601 13311
rect 17359 13280 17601 13308
rect 17359 13277 17371 13280
rect 17313 13271 17371 13277
rect 17589 13277 17601 13280
rect 17635 13277 17647 13311
rect 17696 13308 17724 13484
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 22278 13512 22284 13524
rect 22239 13484 22284 13512
rect 22278 13472 22284 13484
rect 22336 13472 22342 13524
rect 23109 13515 23167 13521
rect 23109 13481 23121 13515
rect 23155 13512 23167 13515
rect 23842 13512 23848 13524
rect 23155 13484 23848 13512
rect 23155 13481 23167 13484
rect 23109 13475 23167 13481
rect 23842 13472 23848 13484
rect 23900 13512 23906 13524
rect 24486 13512 24492 13524
rect 23900 13484 24492 13512
rect 23900 13472 23906 13484
rect 24486 13472 24492 13484
rect 24544 13472 24550 13524
rect 25222 13444 25228 13456
rect 23860 13416 25228 13444
rect 20530 13376 20536 13388
rect 20491 13348 20536 13376
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 20806 13376 20812 13388
rect 20767 13348 20812 13376
rect 20806 13336 20812 13348
rect 20864 13336 20870 13388
rect 17773 13311 17831 13317
rect 17773 13308 17785 13311
rect 17696 13280 17785 13308
rect 17589 13271 17647 13277
rect 17773 13277 17785 13280
rect 17819 13277 17831 13311
rect 17954 13308 17960 13320
rect 17915 13280 17960 13308
rect 17773 13271 17831 13277
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 18049 13311 18107 13317
rect 18049 13277 18061 13311
rect 18095 13277 18107 13311
rect 18509 13311 18567 13317
rect 18509 13308 18521 13311
rect 18049 13271 18107 13277
rect 18248 13280 18521 13308
rect 15654 13200 15660 13252
rect 15712 13240 15718 13252
rect 15712 13212 17080 13240
rect 15712 13200 15718 13212
rect 6549 13175 6607 13181
rect 6236 13144 6281 13172
rect 6236 13132 6242 13144
rect 6549 13141 6561 13175
rect 6595 13141 6607 13175
rect 9306 13172 9312 13184
rect 9267 13144 9312 13172
rect 6549 13135 6607 13141
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 13814 13172 13820 13184
rect 13775 13144 13820 13172
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 15010 13132 15016 13184
rect 15068 13172 15074 13184
rect 15381 13175 15439 13181
rect 15381 13172 15393 13175
rect 15068 13144 15393 13172
rect 15068 13132 15074 13144
rect 15381 13141 15393 13144
rect 15427 13141 15439 13175
rect 16942 13172 16948 13184
rect 16903 13144 16948 13172
rect 15381 13135 15439 13141
rect 16942 13132 16948 13144
rect 17000 13132 17006 13184
rect 17052 13172 17080 13212
rect 18064 13172 18092 13271
rect 18248 13181 18276 13280
rect 18509 13277 18521 13280
rect 18555 13277 18567 13311
rect 23474 13308 23480 13320
rect 23435 13280 23480 13308
rect 18509 13271 18567 13277
rect 23474 13268 23480 13280
rect 23532 13268 23538 13320
rect 23566 13268 23572 13320
rect 23624 13308 23630 13320
rect 23750 13308 23756 13320
rect 23624 13280 23669 13308
rect 23711 13280 23756 13308
rect 23624 13268 23630 13280
rect 23750 13268 23756 13280
rect 23808 13268 23814 13320
rect 21542 13200 21548 13252
rect 21600 13200 21606 13252
rect 23017 13243 23075 13249
rect 23017 13240 23029 13243
rect 22756 13212 23029 13240
rect 22756 13184 22784 13212
rect 23017 13209 23029 13212
rect 23063 13209 23075 13243
rect 23017 13203 23075 13209
rect 17052 13144 18092 13172
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13141 18291 13175
rect 22738 13172 22744 13184
rect 22699 13144 22744 13172
rect 18233 13135 18291 13141
rect 22738 13132 22744 13144
rect 22796 13132 22802 13184
rect 23290 13172 23296 13184
rect 23251 13144 23296 13172
rect 23290 13132 23296 13144
rect 23348 13132 23354 13184
rect 23584 13172 23612 13268
rect 23860 13249 23888 13416
rect 25222 13404 25228 13416
rect 25280 13404 25286 13456
rect 25317 13447 25375 13453
rect 25317 13413 25329 13447
rect 25363 13444 25375 13447
rect 25363 13416 25636 13444
rect 25363 13413 25375 13416
rect 25317 13407 25375 13413
rect 23957 13348 24900 13376
rect 23957 13320 23985 13348
rect 23934 13268 23940 13320
rect 23992 13317 23998 13320
rect 23992 13308 24000 13317
rect 24765 13311 24823 13317
rect 23992 13280 24037 13308
rect 23992 13271 24000 13280
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 24872 13308 24900 13348
rect 25038 13336 25044 13388
rect 25096 13376 25102 13388
rect 25501 13379 25559 13385
rect 25501 13376 25513 13379
rect 25096 13348 25513 13376
rect 25096 13336 25102 13348
rect 25501 13345 25513 13348
rect 25547 13345 25559 13379
rect 25608 13376 25636 13416
rect 25777 13379 25835 13385
rect 25777 13376 25789 13379
rect 25608 13348 25789 13376
rect 25501 13339 25559 13345
rect 25777 13345 25789 13348
rect 25823 13345 25835 13379
rect 25777 13339 25835 13345
rect 25138 13311 25196 13317
rect 25138 13308 25150 13311
rect 24872 13280 25150 13308
rect 24765 13271 24823 13277
rect 25138 13277 25150 13280
rect 25184 13277 25196 13311
rect 25138 13271 25196 13277
rect 23992 13268 23998 13271
rect 23845 13243 23903 13249
rect 23845 13209 23857 13243
rect 23891 13209 23903 13243
rect 24780 13240 24808 13271
rect 24946 13240 24952 13252
rect 23845 13203 23903 13209
rect 24044 13212 24808 13240
rect 24907 13212 24952 13240
rect 24044 13172 24072 13212
rect 24946 13200 24952 13212
rect 25004 13200 25010 13252
rect 25041 13243 25099 13249
rect 25041 13209 25053 13243
rect 25087 13209 25099 13243
rect 25041 13203 25099 13209
rect 23584 13144 24072 13172
rect 24138 13175 24196 13181
rect 24138 13141 24150 13175
rect 24184 13172 24196 13175
rect 24394 13172 24400 13184
rect 24184 13144 24400 13172
rect 24184 13141 24196 13144
rect 24138 13135 24196 13141
rect 24394 13132 24400 13144
rect 24452 13132 24458 13184
rect 25056 13172 25084 13203
rect 26510 13200 26516 13252
rect 26568 13200 26574 13252
rect 27154 13172 27160 13184
rect 25056 13144 27160 13172
rect 27154 13132 27160 13144
rect 27212 13172 27218 13184
rect 27249 13175 27307 13181
rect 27249 13172 27261 13175
rect 27212 13144 27261 13172
rect 27212 13132 27218 13144
rect 27249 13141 27261 13144
rect 27295 13141 27307 13175
rect 27249 13135 27307 13141
rect 1104 13082 29532 13104
rect 1104 13030 10425 13082
rect 10477 13030 10489 13082
rect 10541 13030 10553 13082
rect 10605 13030 10617 13082
rect 10669 13030 10681 13082
rect 10733 13030 19901 13082
rect 19953 13030 19965 13082
rect 20017 13030 20029 13082
rect 20081 13030 20093 13082
rect 20145 13030 20157 13082
rect 20209 13030 29532 13082
rect 1104 13008 29532 13030
rect 2866 12928 2872 12980
rect 2924 12968 2930 12980
rect 2961 12971 3019 12977
rect 2961 12968 2973 12971
rect 2924 12940 2973 12968
rect 2924 12928 2930 12940
rect 2961 12937 2973 12940
rect 3007 12968 3019 12971
rect 3418 12968 3424 12980
rect 3007 12940 3424 12968
rect 3007 12937 3019 12940
rect 2961 12931 3019 12937
rect 3418 12928 3424 12940
rect 3476 12968 3482 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3476 12940 3525 12968
rect 3476 12928 3482 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 3513 12931 3571 12937
rect 3973 12971 4031 12977
rect 3973 12937 3985 12971
rect 4019 12968 4031 12971
rect 4062 12968 4068 12980
rect 4019 12940 4068 12968
rect 4019 12937 4031 12940
rect 3973 12931 4031 12937
rect 2406 12900 2412 12912
rect 2367 12872 2412 12900
rect 2406 12860 2412 12872
rect 2464 12860 2470 12912
rect 2593 12903 2651 12909
rect 2593 12869 2605 12903
rect 2639 12900 2651 12903
rect 2682 12900 2688 12912
rect 2639 12872 2688 12900
rect 2639 12869 2651 12872
rect 2593 12863 2651 12869
rect 2682 12860 2688 12872
rect 2740 12860 2746 12912
rect 3988 12900 4016 12931
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4430 12968 4436 12980
rect 4203 12940 4436 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4430 12928 4436 12940
rect 4488 12968 4494 12980
rect 4798 12968 4804 12980
rect 4488 12940 4804 12968
rect 4488 12928 4494 12940
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 4982 12968 4988 12980
rect 4943 12940 4988 12968
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 5442 12968 5448 12980
rect 5403 12940 5448 12968
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 12253 12971 12311 12977
rect 12253 12968 12265 12971
rect 9876 12940 12265 12968
rect 3160 12872 4016 12900
rect 1762 12792 1768 12844
rect 1820 12832 1826 12844
rect 3160 12841 3188 12872
rect 5074 12860 5080 12912
rect 5132 12900 5138 12912
rect 5132 12872 5488 12900
rect 5132 12860 5138 12872
rect 2823 12835 2881 12841
rect 2823 12832 2835 12835
rect 1820 12804 2835 12832
rect 1820 12792 1826 12804
rect 2823 12801 2835 12804
rect 2869 12801 2881 12835
rect 2823 12795 2881 12801
rect 3145 12835 3203 12841
rect 3145 12801 3157 12835
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 4155 12835 4213 12841
rect 4155 12832 4167 12835
rect 3743 12804 4167 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 4155 12801 4167 12804
rect 4201 12832 4213 12835
rect 4801 12835 4859 12841
rect 4801 12832 4813 12835
rect 4201 12804 4813 12832
rect 4201 12801 4213 12804
rect 4155 12795 4213 12801
rect 4801 12801 4813 12804
rect 4847 12801 4859 12835
rect 4801 12795 4859 12801
rect 4890 12792 4896 12844
rect 4948 12832 4954 12844
rect 4948 12804 4993 12832
rect 4948 12792 4954 12804
rect 5166 12792 5172 12844
rect 5224 12832 5230 12844
rect 5350 12832 5356 12844
rect 5224 12804 5356 12832
rect 5224 12792 5230 12804
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 5460 12832 5488 12872
rect 6549 12835 6607 12841
rect 5460 12804 5580 12832
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 4522 12764 4528 12776
rect 3099 12736 4528 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 4617 12767 4675 12773
rect 4617 12733 4629 12767
rect 4663 12764 4675 12767
rect 5442 12764 5448 12776
rect 4663 12736 5448 12764
rect 4663 12733 4675 12736
rect 4617 12727 4675 12733
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5552 12773 5580 12804
rect 6549 12801 6561 12835
rect 6595 12832 6607 12835
rect 6914 12832 6920 12844
rect 6595 12804 6920 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 9876 12841 9904 12940
rect 12253 12937 12265 12940
rect 12299 12968 12311 12971
rect 13538 12968 13544 12980
rect 12299 12940 13544 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 10870 12860 10876 12912
rect 10928 12900 10934 12912
rect 12161 12903 12219 12909
rect 12161 12900 12173 12903
rect 10928 12872 12173 12900
rect 10928 12860 10934 12872
rect 12161 12869 12173 12872
rect 12207 12869 12219 12903
rect 12161 12863 12219 12869
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9732 12804 9873 12832
rect 9732 12792 9738 12804
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 9950 12792 9956 12844
rect 10008 12832 10014 12844
rect 10117 12835 10175 12841
rect 10117 12832 10129 12835
rect 10008 12804 10129 12832
rect 10008 12792 10014 12804
rect 10117 12801 10129 12804
rect 10163 12801 10175 12835
rect 10117 12795 10175 12801
rect 11609 12835 11667 12841
rect 11609 12801 11621 12835
rect 11655 12801 11667 12835
rect 11790 12832 11796 12844
rect 11751 12804 11796 12832
rect 11609 12795 11667 12801
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 11624 12764 11652 12795
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 12406 12832 12434 12940
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 14277 12971 14335 12977
rect 14277 12937 14289 12971
rect 14323 12968 14335 12971
rect 14366 12968 14372 12980
rect 14323 12940 14372 12968
rect 14323 12937 14335 12940
rect 14277 12931 14335 12937
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 16040 12940 16681 12968
rect 12802 12900 12808 12912
rect 12763 12872 12808 12900
rect 12802 12860 12808 12872
rect 12860 12860 12866 12912
rect 13814 12860 13820 12912
rect 13872 12860 13878 12912
rect 16040 12886 16068 12940
rect 16669 12937 16681 12940
rect 16715 12937 16727 12971
rect 23017 12971 23075 12977
rect 23017 12968 23029 12971
rect 16669 12931 16727 12937
rect 18524 12940 23029 12968
rect 16485 12903 16543 12909
rect 16485 12869 16497 12903
rect 16531 12900 16543 12903
rect 16758 12900 16764 12912
rect 16531 12872 16764 12900
rect 16531 12869 16543 12872
rect 16485 12863 16543 12869
rect 16758 12860 16764 12872
rect 16816 12860 16822 12912
rect 12529 12835 12587 12841
rect 12529 12832 12541 12835
rect 12406 12804 12541 12832
rect 12529 12801 12541 12804
rect 12575 12801 12587 12835
rect 15010 12832 15016 12844
rect 14971 12804 15016 12832
rect 12529 12795 12587 12801
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 18524 12841 18552 12940
rect 23017 12937 23029 12940
rect 23063 12937 23075 12971
rect 25038 12968 25044 12980
rect 23017 12931 23075 12937
rect 24228 12940 25044 12968
rect 20530 12900 20536 12912
rect 19628 12872 20536 12900
rect 19628 12841 19656 12872
rect 20530 12860 20536 12872
rect 20588 12860 20594 12912
rect 24228 12900 24256 12940
rect 25038 12928 25044 12940
rect 25096 12928 25102 12980
rect 25222 12928 25228 12980
rect 25280 12968 25286 12980
rect 25869 12971 25927 12977
rect 25869 12968 25881 12971
rect 25280 12940 25881 12968
rect 25280 12928 25286 12940
rect 25869 12937 25881 12940
rect 25915 12937 25927 12971
rect 26510 12968 26516 12980
rect 26471 12940 26516 12968
rect 25869 12931 25927 12937
rect 24394 12900 24400 12912
rect 24136 12872 24256 12900
rect 24355 12872 24400 12900
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16724 12804 16865 12832
rect 16724 12792 16730 12804
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 18509 12835 18567 12841
rect 18509 12801 18521 12835
rect 18555 12801 18567 12835
rect 18509 12795 18567 12801
rect 19613 12835 19671 12841
rect 19613 12801 19625 12835
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 19880 12835 19938 12841
rect 19880 12801 19892 12835
rect 19926 12832 19938 12835
rect 20438 12832 20444 12844
rect 19926 12804 20444 12832
rect 19926 12801 19938 12804
rect 19880 12795 19938 12801
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 22370 12832 22376 12844
rect 22331 12804 22376 12832
rect 22370 12792 22376 12804
rect 22428 12792 22434 12844
rect 24136 12841 24164 12872
rect 24394 12860 24400 12872
rect 24452 12860 24458 12912
rect 25406 12860 25412 12912
rect 25464 12860 25470 12912
rect 25884 12900 25912 12931
rect 26510 12928 26516 12940
rect 26568 12928 26574 12980
rect 27062 12900 27068 12912
rect 25884 12872 27068 12900
rect 27062 12860 27068 12872
rect 27120 12860 27126 12912
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 26053 12835 26111 12841
rect 26053 12801 26065 12835
rect 26099 12801 26111 12835
rect 26329 12835 26387 12841
rect 26329 12832 26341 12835
rect 26053 12795 26111 12801
rect 26252 12804 26341 12832
rect 12066 12764 12072 12776
rect 5537 12727 5595 12733
rect 11256 12736 12072 12764
rect 2774 12656 2780 12708
rect 2832 12696 2838 12708
rect 6365 12699 6423 12705
rect 6365 12696 6377 12699
rect 2832 12668 6377 12696
rect 2832 12656 2838 12668
rect 6365 12665 6377 12668
rect 6411 12696 6423 12699
rect 6638 12696 6644 12708
rect 6411 12668 6644 12696
rect 6411 12665 6423 12668
rect 6365 12659 6423 12665
rect 6638 12656 6644 12668
rect 6696 12656 6702 12708
rect 11256 12705 11284 12736
rect 12066 12724 12072 12736
rect 12124 12724 12130 12776
rect 13538 12724 13544 12776
rect 13596 12764 13602 12776
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 13596 12736 14657 12764
rect 13596 12724 13602 12736
rect 14645 12733 14657 12736
rect 14691 12733 14703 12767
rect 23216 12764 23244 12795
rect 23290 12764 23296 12776
rect 23203 12736 23296 12764
rect 14645 12727 14703 12733
rect 23290 12724 23296 12736
rect 23348 12764 23354 12776
rect 24486 12764 24492 12776
rect 23348 12736 24492 12764
rect 23348 12724 23354 12736
rect 24486 12724 24492 12736
rect 24544 12764 24550 12776
rect 26068 12764 26096 12795
rect 24544 12736 26096 12764
rect 24544 12724 24550 12736
rect 11241 12699 11299 12705
rect 11241 12665 11253 12699
rect 11287 12665 11299 12699
rect 11241 12659 11299 12665
rect 11885 12699 11943 12705
rect 11885 12665 11897 12699
rect 11931 12696 11943 12699
rect 12526 12696 12532 12708
rect 11931 12668 12532 12696
rect 11931 12665 11943 12668
rect 11885 12659 11943 12665
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 26252 12705 26280 12804
rect 26329 12801 26341 12804
rect 26375 12801 26387 12835
rect 26329 12795 26387 12801
rect 26237 12699 26295 12705
rect 26237 12665 26249 12699
rect 26283 12665 26295 12699
rect 26237 12659 26295 12665
rect 4525 12631 4583 12637
rect 4525 12597 4537 12631
rect 4571 12628 4583 12631
rect 5534 12628 5540 12640
rect 4571 12600 5540 12628
rect 4571 12597 4583 12600
rect 4525 12591 4583 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 9306 12588 9312 12640
rect 9364 12628 9370 12640
rect 13354 12628 13360 12640
rect 9364 12600 13360 12628
rect 9364 12588 9370 12600
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 18230 12588 18236 12640
rect 18288 12628 18294 12640
rect 18325 12631 18383 12637
rect 18325 12628 18337 12631
rect 18288 12600 18337 12628
rect 18288 12588 18294 12600
rect 18325 12597 18337 12600
rect 18371 12597 18383 12631
rect 18325 12591 18383 12597
rect 19242 12588 19248 12640
rect 19300 12628 19306 12640
rect 20714 12628 20720 12640
rect 19300 12600 20720 12628
rect 19300 12588 19306 12600
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 20993 12631 21051 12637
rect 20993 12597 21005 12631
rect 21039 12628 21051 12631
rect 21174 12628 21180 12640
rect 21039 12600 21180 12628
rect 21039 12597 21051 12600
rect 20993 12591 21051 12597
rect 21174 12588 21180 12600
rect 21232 12588 21238 12640
rect 22462 12628 22468 12640
rect 22423 12600 22468 12628
rect 22462 12588 22468 12600
rect 22520 12588 22526 12640
rect 1104 12538 29532 12560
rect 1104 12486 5688 12538
rect 5740 12486 5752 12538
rect 5804 12486 5816 12538
rect 5868 12486 5880 12538
rect 5932 12486 5944 12538
rect 5996 12486 15163 12538
rect 15215 12486 15227 12538
rect 15279 12486 15291 12538
rect 15343 12486 15355 12538
rect 15407 12486 15419 12538
rect 15471 12486 24639 12538
rect 24691 12486 24703 12538
rect 24755 12486 24767 12538
rect 24819 12486 24831 12538
rect 24883 12486 24895 12538
rect 24947 12486 29532 12538
rect 1104 12464 29532 12486
rect 4430 12384 4436 12436
rect 4488 12424 4494 12436
rect 5074 12424 5080 12436
rect 4488 12396 5080 12424
rect 4488 12384 4494 12396
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 14274 12424 14280 12436
rect 6196 12396 14136 12424
rect 14235 12396 14280 12424
rect 2961 12359 3019 12365
rect 2961 12325 2973 12359
rect 3007 12356 3019 12359
rect 4982 12356 4988 12368
rect 3007 12328 4988 12356
rect 3007 12325 3019 12328
rect 2961 12319 3019 12325
rect 4982 12316 4988 12328
rect 5040 12316 5046 12368
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 4798 12288 4804 12300
rect 4479 12260 4804 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 5092 12288 5120 12384
rect 5353 12291 5411 12297
rect 5353 12288 5365 12291
rect 5092 12260 5365 12288
rect 5353 12257 5365 12260
rect 5399 12257 5411 12291
rect 5534 12288 5540 12300
rect 5495 12260 5540 12288
rect 5353 12251 5411 12257
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 1581 12223 1639 12229
rect 1581 12189 1593 12223
rect 1627 12220 1639 12223
rect 2774 12220 2780 12232
rect 1627 12192 2780 12220
rect 1627 12189 1639 12192
rect 1581 12183 1639 12189
rect 2774 12180 2780 12192
rect 2832 12180 2838 12232
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12220 4307 12223
rect 4522 12220 4528 12232
rect 4295 12192 4528 12220
rect 4295 12189 4307 12192
rect 4249 12183 4307 12189
rect 4522 12180 4528 12192
rect 4580 12180 4586 12232
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12220 5687 12223
rect 6086 12220 6092 12232
rect 5675 12192 6092 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 1848 12155 1906 12161
rect 1848 12121 1860 12155
rect 1894 12152 1906 12155
rect 1894 12124 3832 12152
rect 1894 12121 1906 12124
rect 1848 12115 1906 12121
rect 3804 12093 3832 12124
rect 4062 12112 4068 12164
rect 4120 12152 4126 12164
rect 4120 12124 4476 12152
rect 4120 12112 4126 12124
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12053 3847 12087
rect 3789 12047 3847 12053
rect 3878 12044 3884 12096
rect 3936 12084 3942 12096
rect 4157 12087 4215 12093
rect 4157 12084 4169 12087
rect 3936 12056 4169 12084
rect 3936 12044 3942 12056
rect 4157 12053 4169 12056
rect 4203 12053 4215 12087
rect 4448 12084 4476 12124
rect 5534 12112 5540 12164
rect 5592 12152 5598 12164
rect 5644 12152 5672 12183
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 6196 12152 6224 12396
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 8938 12356 8944 12368
rect 8352 12328 8944 12356
rect 8352 12316 8358 12328
rect 8938 12316 8944 12328
rect 8996 12356 9002 12368
rect 9582 12356 9588 12368
rect 8996 12328 9588 12356
rect 8996 12316 9002 12328
rect 9582 12316 9588 12328
rect 9640 12316 9646 12368
rect 9769 12359 9827 12365
rect 9769 12325 9781 12359
rect 9815 12356 9827 12359
rect 9950 12356 9956 12368
rect 9815 12328 9956 12356
rect 9815 12325 9827 12328
rect 9769 12319 9827 12325
rect 9950 12316 9956 12328
rect 10008 12316 10014 12368
rect 10778 12356 10784 12368
rect 10739 12328 10784 12356
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 11572 12328 12296 12356
rect 11572 12316 11578 12328
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 9677 12291 9735 12297
rect 9677 12288 9689 12291
rect 8536 12260 9689 12288
rect 8536 12248 8542 12260
rect 9677 12257 9689 12260
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12288 10287 12291
rect 10318 12288 10324 12300
rect 10275 12260 10324 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 6362 12180 6368 12232
rect 6420 12220 6426 12232
rect 6638 12220 6644 12232
rect 6420 12192 6644 12220
rect 6420 12180 6426 12192
rect 6638 12180 6644 12192
rect 6696 12220 6702 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 6696 12192 7297 12220
rect 6696 12180 6702 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 9585 12223 9643 12229
rect 9585 12220 9597 12223
rect 8444 12192 9597 12220
rect 8444 12180 8450 12192
rect 9585 12189 9597 12192
rect 9631 12189 9643 12223
rect 9585 12183 9643 12189
rect 5592 12124 5672 12152
rect 5736 12124 6224 12152
rect 7552 12155 7610 12161
rect 5592 12112 5598 12124
rect 5736 12084 5764 12124
rect 7552 12121 7564 12155
rect 7598 12152 7610 12155
rect 7650 12152 7656 12164
rect 7598 12124 7656 12152
rect 7598 12121 7610 12124
rect 7552 12115 7610 12121
rect 7650 12112 7656 12124
rect 7708 12112 7714 12164
rect 5994 12084 6000 12096
rect 4448 12056 5764 12084
rect 5955 12056 6000 12084
rect 4157 12047 4215 12053
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 8665 12087 8723 12093
rect 8665 12053 8677 12087
rect 8711 12084 8723 12087
rect 8754 12084 8760 12096
rect 8711 12056 8760 12084
rect 8711 12053 8723 12056
rect 8665 12047 8723 12053
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8904 12056 8953 12084
rect 8904 12044 8910 12056
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 9692 12084 9720 12251
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 11882 12288 11888 12300
rect 10428 12260 11888 12288
rect 10137 12223 10195 12229
rect 10137 12189 10149 12223
rect 10183 12220 10195 12223
rect 10428 12220 10456 12260
rect 11882 12248 11888 12260
rect 11940 12288 11946 12300
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 11940 12260 12173 12288
rect 11940 12248 11946 12260
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 10183 12192 10456 12220
rect 10505 12223 10563 12229
rect 10183 12189 10195 12192
rect 10137 12183 10195 12189
rect 10505 12189 10517 12223
rect 10551 12189 10563 12223
rect 10505 12183 10563 12189
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12220 10747 12223
rect 10778 12220 10784 12232
rect 10735 12192 10784 12220
rect 10735 12189 10747 12192
rect 10689 12183 10747 12189
rect 10520 12152 10548 12183
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 11790 12220 11796 12232
rect 11664 12192 11796 12220
rect 11664 12180 11670 12192
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 12066 12220 12072 12232
rect 12027 12192 12072 12220
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 12268 12220 12296 12328
rect 12894 12316 12900 12368
rect 12952 12356 12958 12368
rect 13725 12359 13783 12365
rect 13725 12356 13737 12359
rect 12952 12328 13737 12356
rect 12952 12316 12958 12328
rect 13725 12325 13737 12328
rect 13771 12325 13783 12359
rect 14108 12356 14136 12396
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 14458 12384 14464 12436
rect 14516 12424 14522 12436
rect 14826 12424 14832 12436
rect 14516 12396 14832 12424
rect 14516 12384 14522 12396
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 15749 12427 15807 12433
rect 15749 12393 15761 12427
rect 15795 12424 15807 12427
rect 16666 12424 16672 12436
rect 15795 12396 16672 12424
rect 15795 12393 15807 12396
rect 15749 12387 15807 12393
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 19242 12424 19248 12436
rect 16776 12396 19248 12424
rect 16776 12356 16804 12396
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 22370 12424 22376 12436
rect 22331 12396 22376 12424
rect 22370 12384 22376 12396
rect 22428 12384 22434 12436
rect 25317 12427 25375 12433
rect 25317 12393 25329 12427
rect 25363 12424 25375 12427
rect 25406 12424 25412 12436
rect 25363 12396 25412 12424
rect 25363 12393 25375 12396
rect 25317 12387 25375 12393
rect 25406 12384 25412 12396
rect 25464 12384 25470 12436
rect 22738 12356 22744 12368
rect 14108 12328 16804 12356
rect 19904 12328 22744 12356
rect 13725 12319 13783 12325
rect 14737 12291 14795 12297
rect 13464 12260 14688 12288
rect 12345 12223 12403 12229
rect 12345 12220 12357 12223
rect 12268 12192 12357 12220
rect 12345 12189 12357 12192
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 12618 12180 12624 12232
rect 12676 12220 12682 12232
rect 13464 12229 13492 12260
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 12676 12192 13461 12220
rect 12676 12180 12682 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 13909 12223 13967 12229
rect 13909 12220 13921 12223
rect 13872 12192 13921 12220
rect 13872 12180 13878 12192
rect 13909 12189 13921 12192
rect 13955 12220 13967 12223
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13955 12192 14105 12220
rect 13955 12189 13967 12192
rect 13909 12183 13967 12189
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14458 12220 14464 12232
rect 14419 12192 14464 12220
rect 14093 12183 14151 12189
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12189 14611 12223
rect 14660 12220 14688 12260
rect 14737 12257 14749 12291
rect 14783 12288 14795 12291
rect 15470 12288 15476 12300
rect 14783 12260 15476 12288
rect 14783 12257 14795 12260
rect 14737 12251 14795 12257
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 17126 12288 17132 12300
rect 17087 12260 17132 12288
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19613 12291 19671 12297
rect 19613 12288 19625 12291
rect 19392 12260 19625 12288
rect 19392 12248 19398 12260
rect 19613 12257 19625 12260
rect 19659 12288 19671 12291
rect 19904 12288 19932 12328
rect 22738 12316 22744 12328
rect 22796 12316 22802 12368
rect 20438 12288 20444 12300
rect 19659 12260 19932 12288
rect 20399 12260 20444 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 15565 12223 15623 12229
rect 15565 12220 15577 12223
rect 14660 12192 15577 12220
rect 14553 12183 14611 12189
rect 15565 12189 15577 12192
rect 15611 12220 15623 12223
rect 15654 12220 15660 12232
rect 15611 12192 15660 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 10965 12155 11023 12161
rect 10965 12152 10977 12155
rect 10520 12124 10977 12152
rect 10965 12121 10977 12124
rect 11011 12152 11023 12155
rect 11054 12152 11060 12164
rect 11011 12124 11060 12152
rect 11011 12121 11023 12124
rect 10965 12115 11023 12121
rect 11054 12112 11060 12124
rect 11112 12112 11118 12164
rect 11149 12155 11207 12161
rect 11149 12121 11161 12155
rect 11195 12152 11207 12155
rect 12437 12155 12495 12161
rect 11195 12124 12112 12152
rect 11195 12121 11207 12124
rect 11149 12115 11207 12121
rect 12084 12096 12112 12124
rect 12437 12121 12449 12155
rect 12483 12152 12495 12155
rect 13722 12152 13728 12164
rect 12483 12124 13728 12152
rect 12483 12121 12495 12124
rect 12437 12115 12495 12121
rect 13722 12112 13728 12124
rect 13780 12152 13786 12164
rect 14568 12152 14596 12183
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 16390 12180 16396 12232
rect 16448 12220 16454 12232
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 16448 12192 16681 12220
rect 16448 12180 16454 12192
rect 16669 12189 16681 12192
rect 16715 12189 16727 12223
rect 16669 12183 16727 12189
rect 16758 12180 16764 12232
rect 16816 12220 16822 12232
rect 16853 12223 16911 12229
rect 16853 12220 16865 12223
rect 16816 12192 16865 12220
rect 16816 12180 16822 12192
rect 16853 12189 16865 12192
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 18230 12180 18236 12232
rect 18288 12180 18294 12232
rect 19061 12223 19119 12229
rect 19061 12189 19073 12223
rect 19107 12220 19119 12223
rect 19150 12220 19156 12232
rect 19107 12192 19156 12220
rect 19107 12189 19119 12192
rect 19061 12183 19119 12189
rect 19150 12180 19156 12192
rect 19208 12220 19214 12232
rect 19904 12229 19932 12260
rect 20438 12248 20444 12260
rect 20496 12248 20502 12300
rect 21266 12288 21272 12300
rect 20548 12260 21272 12288
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 19208 12192 19257 12220
rect 19208 12180 19214 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12189 19947 12223
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 19889 12183 19947 12189
rect 19996 12192 20085 12220
rect 13780 12124 14596 12152
rect 13780 12112 13786 12124
rect 14642 12112 14648 12164
rect 14700 12152 14706 12164
rect 14829 12155 14887 12161
rect 14829 12152 14841 12155
rect 14700 12124 14841 12152
rect 14700 12112 14706 12124
rect 14829 12121 14841 12124
rect 14875 12121 14887 12155
rect 14829 12115 14887 12121
rect 14921 12155 14979 12161
rect 14921 12121 14933 12155
rect 14967 12152 14979 12155
rect 15286 12152 15292 12164
rect 14967 12124 15292 12152
rect 14967 12121 14979 12124
rect 14921 12115 14979 12121
rect 15286 12112 15292 12124
rect 15344 12112 15350 12164
rect 18969 12155 19027 12161
rect 15396 12124 16712 12152
rect 11330 12084 11336 12096
rect 9692 12056 11336 12084
rect 8941 12047 8999 12053
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 11974 12084 11980 12096
rect 11848 12056 11980 12084
rect 11848 12044 11854 12056
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12066 12044 12072 12096
rect 12124 12044 12130 12096
rect 13538 12044 13544 12096
rect 13596 12084 13602 12096
rect 13633 12087 13691 12093
rect 13633 12084 13645 12087
rect 13596 12056 13645 12084
rect 13596 12044 13602 12056
rect 13633 12053 13645 12056
rect 13679 12053 13691 12087
rect 13633 12047 13691 12053
rect 14093 12087 14151 12093
rect 14093 12053 14105 12087
rect 14139 12084 14151 12087
rect 15396 12084 15424 12124
rect 16574 12084 16580 12096
rect 14139 12056 15424 12084
rect 16535 12056 16580 12084
rect 14139 12053 14151 12056
rect 14093 12047 14151 12053
rect 16574 12044 16580 12056
rect 16632 12044 16638 12096
rect 16684 12084 16712 12124
rect 18969 12121 18981 12155
rect 19015 12152 19027 12155
rect 19518 12152 19524 12164
rect 19015 12124 19524 12152
rect 19015 12121 19027 12124
rect 18969 12115 19027 12121
rect 19518 12112 19524 12124
rect 19576 12112 19582 12164
rect 19702 12152 19708 12164
rect 19663 12124 19708 12152
rect 19702 12112 19708 12124
rect 19760 12112 19766 12164
rect 19996 12152 20024 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 20349 12223 20407 12229
rect 20349 12220 20361 12223
rect 20312 12192 20361 12220
rect 20312 12180 20318 12192
rect 20349 12189 20361 12192
rect 20395 12189 20407 12223
rect 20349 12183 20407 12189
rect 20548 12152 20576 12260
rect 21266 12248 21272 12260
rect 21324 12288 21330 12300
rect 21821 12291 21879 12297
rect 21324 12260 21404 12288
rect 21324 12248 21330 12260
rect 20625 12223 20683 12229
rect 20625 12189 20637 12223
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 19996 12124 20576 12152
rect 20640 12152 20668 12183
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 20809 12223 20867 12229
rect 20809 12220 20821 12223
rect 20772 12192 20821 12220
rect 20772 12180 20778 12192
rect 20809 12189 20821 12192
rect 20855 12220 20867 12223
rect 21085 12223 21143 12229
rect 21085 12220 21097 12223
rect 20855 12192 21097 12220
rect 20855 12189 20867 12192
rect 20809 12183 20867 12189
rect 21085 12189 21097 12192
rect 21131 12189 21143 12223
rect 21085 12183 21143 12189
rect 21174 12180 21180 12232
rect 21232 12220 21238 12232
rect 21376 12229 21404 12260
rect 21821 12257 21833 12291
rect 21867 12288 21879 12291
rect 23753 12291 23811 12297
rect 21867 12260 22600 12288
rect 21867 12257 21879 12260
rect 21821 12251 21879 12257
rect 21361 12223 21419 12229
rect 21232 12192 21277 12220
rect 21232 12180 21238 12192
rect 21361 12189 21373 12223
rect 21407 12189 21419 12223
rect 21634 12220 21640 12232
rect 21595 12192 21640 12220
rect 21361 12183 21419 12189
rect 21634 12180 21640 12192
rect 21692 12180 21698 12232
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12220 22155 12223
rect 22186 12220 22192 12232
rect 22143 12192 22192 12220
rect 22143 12189 22155 12192
rect 22097 12183 22155 12189
rect 21450 12152 21456 12164
rect 20640 12124 21456 12152
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 16684 12056 18613 12084
rect 18601 12053 18613 12056
rect 18647 12053 18659 12087
rect 18601 12047 18659 12053
rect 19429 12087 19487 12093
rect 19429 12053 19441 12087
rect 19475 12084 19487 12087
rect 19996 12084 20024 12124
rect 21450 12112 21456 12124
rect 21508 12152 21514 12164
rect 21928 12152 21956 12183
rect 22186 12180 22192 12192
rect 22244 12220 22250 12232
rect 22462 12220 22468 12232
rect 22244 12192 22468 12220
rect 22244 12180 22250 12192
rect 22462 12180 22468 12192
rect 22520 12180 22526 12232
rect 22572 12220 22600 12260
rect 23753 12257 23765 12291
rect 23799 12288 23811 12291
rect 25038 12288 25044 12300
rect 23799 12260 25044 12288
rect 23799 12257 23811 12260
rect 23753 12251 23811 12257
rect 25038 12248 25044 12260
rect 25096 12248 25102 12300
rect 23486 12223 23544 12229
rect 23486 12220 23498 12223
rect 22572 12192 23498 12220
rect 23486 12189 23498 12192
rect 23532 12189 23544 12223
rect 23486 12183 23544 12189
rect 24486 12180 24492 12232
rect 24544 12220 24550 12232
rect 24857 12223 24915 12229
rect 24857 12220 24869 12223
rect 24544 12192 24869 12220
rect 24544 12180 24550 12192
rect 24857 12189 24869 12192
rect 24903 12189 24915 12223
rect 25133 12223 25191 12229
rect 25133 12220 25145 12223
rect 24857 12183 24915 12189
rect 25056 12192 25145 12220
rect 21508 12124 21956 12152
rect 21508 12112 21514 12124
rect 25056 12093 25084 12192
rect 25133 12189 25145 12192
rect 25179 12189 25191 12223
rect 25133 12183 25191 12189
rect 19475 12056 20024 12084
rect 25041 12087 25099 12093
rect 19475 12053 19487 12056
rect 19429 12047 19487 12053
rect 25041 12053 25053 12087
rect 25087 12053 25099 12087
rect 25041 12047 25099 12053
rect 1104 11994 29532 12016
rect 1104 11942 10425 11994
rect 10477 11942 10489 11994
rect 10541 11942 10553 11994
rect 10605 11942 10617 11994
rect 10669 11942 10681 11994
rect 10733 11942 19901 11994
rect 19953 11942 19965 11994
rect 20017 11942 20029 11994
rect 20081 11942 20093 11994
rect 20145 11942 20157 11994
rect 20209 11942 29532 11994
rect 1104 11920 29532 11942
rect 3786 11880 3792 11892
rect 3747 11852 3792 11880
rect 3786 11840 3792 11852
rect 3844 11840 3850 11892
rect 4065 11883 4123 11889
rect 4065 11849 4077 11883
rect 4111 11849 4123 11883
rect 4065 11843 4123 11849
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 5166 11880 5172 11892
rect 4479 11852 5172 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 3418 11812 3424 11824
rect 3379 11784 3424 11812
rect 3418 11772 3424 11784
rect 3476 11772 3482 11824
rect 3878 11812 3884 11824
rect 3620 11784 3884 11812
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 3620 11744 3648 11784
rect 3878 11772 3884 11784
rect 3936 11772 3942 11824
rect 3283 11716 3648 11744
rect 3677 11747 3735 11753
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 3677 11713 3689 11747
rect 3723 11744 3735 11747
rect 4080 11744 4108 11843
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 7558 11880 7564 11892
rect 5736 11852 7564 11880
rect 3723 11716 4108 11744
rect 3723 11713 3735 11716
rect 3677 11707 3735 11713
rect 4430 11704 4436 11756
rect 4488 11744 4494 11756
rect 4488 11716 4752 11744
rect 4488 11704 4494 11716
rect 4724 11688 4752 11716
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 4948 11716 5181 11744
rect 4948 11704 4954 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5442 11744 5448 11756
rect 5403 11716 5448 11744
rect 5169 11707 5227 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 5736 11753 5764 11852
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 7745 11883 7803 11889
rect 7745 11849 7757 11883
rect 7791 11849 7803 11883
rect 8386 11880 8392 11892
rect 8347 11852 8392 11880
rect 7745 11843 7803 11849
rect 5818 11815 5876 11821
rect 5818 11781 5830 11815
rect 5864 11812 5876 11815
rect 5994 11812 6000 11824
rect 5864 11784 6000 11812
rect 5864 11781 5876 11784
rect 5818 11775 5876 11781
rect 5994 11772 6000 11784
rect 6052 11772 6058 11824
rect 7760 11812 7788 11843
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 10873 11883 10931 11889
rect 10873 11880 10885 11883
rect 10836 11852 10885 11880
rect 10836 11840 10842 11852
rect 10873 11849 10885 11852
rect 10919 11849 10931 11883
rect 10873 11843 10931 11849
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 13078 11880 13084 11892
rect 11388 11852 13084 11880
rect 11388 11840 11394 11852
rect 8113 11815 8171 11821
rect 7760 11784 8064 11812
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 3878 11676 3884 11688
rect 3839 11648 3884 11676
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11676 4031 11679
rect 4522 11676 4528 11688
rect 4019 11648 4528 11676
rect 4019 11645 4031 11648
rect 3973 11639 4031 11645
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 4706 11676 4712 11688
rect 4667 11648 4712 11676
rect 4706 11636 4712 11648
rect 4764 11636 4770 11688
rect 5552 11676 5580 11707
rect 5902 11704 5908 11756
rect 5960 11753 5966 11756
rect 5960 11744 5968 11753
rect 6086 11744 6092 11756
rect 5960 11716 6092 11744
rect 5960 11707 5968 11716
rect 5960 11704 5966 11707
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 6362 11744 6368 11756
rect 6323 11716 6368 11744
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 6621 11747 6679 11753
rect 6621 11744 6633 11747
rect 6472 11716 6633 11744
rect 6270 11676 6276 11688
rect 5092 11648 6276 11676
rect 4246 11568 4252 11620
rect 4304 11608 4310 11620
rect 4985 11611 5043 11617
rect 4985 11608 4997 11611
rect 4304 11580 4997 11608
rect 4304 11568 4310 11580
rect 4985 11577 4997 11580
rect 5031 11577 5043 11611
rect 4985 11571 5043 11577
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 5092 11540 5120 11648
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 6472 11676 6500 11716
rect 6621 11713 6633 11716
rect 6667 11713 6679 11747
rect 6621 11707 6679 11713
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 8036 11744 8064 11784
rect 8113 11781 8125 11815
rect 8159 11812 8171 11815
rect 9769 11815 9827 11821
rect 9769 11812 9781 11815
rect 8159 11784 9781 11812
rect 8159 11781 8171 11784
rect 8113 11775 8171 11781
rect 9769 11781 9781 11784
rect 9815 11812 9827 11815
rect 9858 11812 9864 11824
rect 9815 11784 9864 11812
rect 9815 11781 9827 11784
rect 9769 11775 9827 11781
rect 9858 11772 9864 11784
rect 9916 11812 9922 11824
rect 10505 11815 10563 11821
rect 10505 11812 10517 11815
rect 9916 11784 10517 11812
rect 9916 11772 9922 11784
rect 10505 11781 10517 11784
rect 10551 11812 10563 11815
rect 11057 11815 11115 11821
rect 11057 11812 11069 11815
rect 10551 11784 11069 11812
rect 10551 11781 10563 11784
rect 10505 11775 10563 11781
rect 11057 11781 11069 11784
rect 11103 11781 11115 11815
rect 11057 11775 11115 11781
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 6972 11716 7972 11744
rect 8036 11716 8309 11744
rect 6972 11704 6978 11716
rect 6380 11648 6500 11676
rect 5353 11611 5411 11617
rect 5353 11577 5365 11611
rect 5399 11577 5411 11611
rect 5353 11571 5411 11577
rect 6089 11611 6147 11617
rect 6089 11577 6101 11611
rect 6135 11608 6147 11611
rect 6178 11608 6184 11620
rect 6135 11580 6184 11608
rect 6135 11577 6147 11580
rect 6089 11571 6147 11577
rect 4028 11512 5120 11540
rect 5368 11540 5396 11571
rect 6178 11568 6184 11580
rect 6236 11568 6242 11620
rect 6380 11540 6408 11648
rect 7944 11620 7972 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8754 11744 8760 11756
rect 8715 11716 8760 11744
rect 8297 11707 8355 11713
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 8938 11744 8944 11756
rect 8899 11716 8944 11744
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 9122 11744 9128 11756
rect 9083 11716 9128 11744
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11713 9275 11747
rect 9950 11744 9956 11756
rect 9911 11716 9956 11744
rect 9217 11707 9275 11713
rect 7926 11608 7932 11620
rect 7887 11580 7932 11608
rect 7926 11568 7932 11580
rect 7984 11568 7990 11620
rect 6730 11540 6736 11552
rect 5368 11512 6736 11540
rect 4028 11500 4034 11512
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 8202 11500 8208 11552
rect 8260 11540 8266 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 8260 11512 8585 11540
rect 8260 11500 8266 11512
rect 8573 11509 8585 11512
rect 8619 11509 8631 11543
rect 8772 11540 8800 11704
rect 8941 11543 8999 11549
rect 8941 11540 8953 11543
rect 8772 11512 8953 11540
rect 8573 11503 8631 11509
rect 8941 11509 8953 11512
rect 8987 11509 8999 11543
rect 9232 11540 9260 11707
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 10134 11744 10140 11756
rect 10095 11716 10140 11744
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10318 11744 10324 11756
rect 10279 11716 10324 11744
rect 10318 11704 10324 11716
rect 10376 11744 10382 11756
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 10376 11716 10793 11744
rect 10376 11704 10382 11716
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 11882 11744 11888 11756
rect 11843 11716 11888 11744
rect 10781 11707 10839 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 11992 11753 12020 11852
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 15286 11880 15292 11892
rect 15247 11852 15292 11880
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 15473 11883 15531 11889
rect 15473 11849 15485 11883
rect 15519 11880 15531 11883
rect 15838 11880 15844 11892
rect 15519 11852 15844 11880
rect 15519 11849 15531 11852
rect 15473 11843 15531 11849
rect 15838 11840 15844 11852
rect 15896 11840 15902 11892
rect 16942 11840 16948 11892
rect 17000 11880 17006 11892
rect 17037 11883 17095 11889
rect 17037 11880 17049 11883
rect 17000 11852 17049 11880
rect 17000 11840 17006 11852
rect 17037 11849 17049 11852
rect 17083 11849 17095 11883
rect 19794 11880 19800 11892
rect 19707 11852 19800 11880
rect 17037 11843 17095 11849
rect 19794 11840 19800 11852
rect 19852 11880 19858 11892
rect 21450 11880 21456 11892
rect 19852 11852 20944 11880
rect 21411 11852 21456 11880
rect 19852 11840 19858 11852
rect 13725 11815 13783 11821
rect 13725 11781 13737 11815
rect 13771 11812 13783 11815
rect 16574 11812 16580 11824
rect 13771 11784 16580 11812
rect 13771 11781 13783 11784
rect 13725 11775 13783 11781
rect 16574 11772 16580 11784
rect 16632 11812 16638 11824
rect 16632 11784 16896 11812
rect 16632 11772 16638 11784
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11713 12035 11747
rect 12158 11744 12164 11756
rect 12119 11716 12164 11744
rect 11977 11707 12035 11713
rect 12158 11704 12164 11716
rect 12216 11704 12222 11756
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 11514 11676 11520 11688
rect 9416 11648 11520 11676
rect 9416 11617 9444 11648
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 12452 11676 12480 11707
rect 11848 11648 12480 11676
rect 13556 11676 13584 11707
rect 13722 11676 13728 11688
rect 13556 11648 13728 11676
rect 11848 11636 11854 11648
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 15396 11676 15424 11707
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 16868 11753 16896 11784
rect 15657 11747 15715 11753
rect 15657 11744 15669 11747
rect 15620 11716 15669 11744
rect 15620 11704 15626 11716
rect 15657 11713 15669 11716
rect 15703 11713 15715 11747
rect 15657 11707 15715 11713
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 18684 11747 18742 11753
rect 18684 11713 18696 11747
rect 18730 11744 18742 11747
rect 19242 11744 19248 11756
rect 18730 11716 19248 11744
rect 18730 11713 18742 11716
rect 18684 11707 18742 11713
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 20451 11753 20479 11852
rect 20533 11815 20591 11821
rect 20533 11781 20545 11815
rect 20579 11812 20591 11815
rect 20714 11812 20720 11824
rect 20579 11784 20720 11812
rect 20579 11781 20591 11784
rect 20533 11775 20591 11781
rect 20714 11772 20720 11784
rect 20772 11772 20778 11824
rect 20916 11821 20944 11852
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 21634 11840 21640 11892
rect 21692 11880 21698 11892
rect 22005 11883 22063 11889
rect 22005 11880 22017 11883
rect 21692 11852 22017 11880
rect 21692 11840 21698 11852
rect 22005 11849 22017 11852
rect 22051 11849 22063 11883
rect 22833 11883 22891 11889
rect 22833 11880 22845 11883
rect 22005 11843 22063 11849
rect 22112 11852 22845 11880
rect 20901 11815 20959 11821
rect 20901 11781 20913 11815
rect 20947 11781 20959 11815
rect 20901 11775 20959 11781
rect 21085 11815 21143 11821
rect 21085 11781 21097 11815
rect 21131 11812 21143 11815
rect 21174 11812 21180 11824
rect 21131 11784 21180 11812
rect 21131 11781 21143 11784
rect 21085 11775 21143 11781
rect 21174 11772 21180 11784
rect 21232 11772 21238 11824
rect 21468 11812 21496 11840
rect 22112 11812 22140 11852
rect 22833 11849 22845 11852
rect 22879 11849 22891 11883
rect 22833 11843 22891 11849
rect 22649 11815 22707 11821
rect 22649 11812 22661 11815
rect 21468 11784 22140 11812
rect 22204 11784 22661 11812
rect 22204 11756 22232 11784
rect 22649 11781 22661 11784
rect 22695 11781 22707 11815
rect 22649 11775 22707 11781
rect 20436 11747 20494 11753
rect 20436 11713 20448 11747
rect 20482 11713 20494 11747
rect 20436 11707 20494 11713
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11744 20683 11747
rect 20809 11747 20867 11753
rect 20671 11716 20760 11744
rect 20671 11713 20683 11716
rect 20625 11707 20683 11713
rect 20732 11688 20760 11716
rect 20809 11713 20821 11747
rect 20855 11713 20867 11747
rect 21545 11747 21603 11753
rect 21545 11744 21557 11747
rect 20809 11707 20867 11713
rect 21008 11716 21557 11744
rect 15838 11676 15844 11688
rect 15396 11648 15844 11676
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 18417 11679 18475 11685
rect 18417 11645 18429 11679
rect 18463 11645 18475 11679
rect 18417 11639 18475 11645
rect 9401 11611 9459 11617
rect 9401 11577 9413 11611
rect 9447 11577 9459 11611
rect 9401 11571 9459 11577
rect 10689 11611 10747 11617
rect 10689 11577 10701 11611
rect 10735 11608 10747 11611
rect 10778 11608 10784 11620
rect 10735 11580 10784 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 10778 11568 10784 11580
rect 10836 11568 10842 11620
rect 10962 11568 10968 11620
rect 11020 11608 11026 11620
rect 12250 11608 12256 11620
rect 11020 11580 11836 11608
rect 12211 11580 12256 11608
rect 11020 11568 11026 11580
rect 9677 11543 9735 11549
rect 9677 11540 9689 11543
rect 9232 11512 9689 11540
rect 8941 11503 8999 11509
rect 9677 11509 9689 11512
rect 9723 11540 9735 11543
rect 9858 11540 9864 11552
rect 9723 11512 9864 11540
rect 9723 11509 9735 11512
rect 9677 11503 9735 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 11146 11500 11152 11552
rect 11204 11540 11210 11552
rect 11606 11540 11612 11552
rect 11204 11512 11612 11540
rect 11204 11500 11210 11512
rect 11606 11500 11612 11512
rect 11664 11540 11670 11552
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 11664 11512 11713 11540
rect 11664 11500 11670 11512
rect 11701 11509 11713 11512
rect 11747 11509 11759 11543
rect 11808 11540 11836 11580
rect 12250 11568 12256 11580
rect 12308 11568 12314 11620
rect 13357 11611 13415 11617
rect 13357 11608 13369 11611
rect 12406 11580 13369 11608
rect 12406 11540 12434 11580
rect 13357 11577 13369 11580
rect 13403 11577 13415 11611
rect 13357 11571 13415 11577
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 15746 11608 15752 11620
rect 15344 11580 15752 11608
rect 15344 11568 15350 11580
rect 15746 11568 15752 11580
rect 15804 11568 15810 11620
rect 12526 11540 12532 11552
rect 11808 11512 12434 11540
rect 12487 11512 12532 11540
rect 11701 11503 11759 11509
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 18432 11540 18460 11639
rect 20714 11636 20720 11688
rect 20772 11636 20778 11688
rect 20824 11620 20852 11707
rect 20254 11608 20260 11620
rect 20215 11580 20260 11608
rect 20254 11568 20260 11580
rect 20312 11568 20318 11620
rect 20806 11568 20812 11620
rect 20864 11568 20870 11620
rect 19334 11540 19340 11552
rect 18432 11512 19340 11540
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 19610 11500 19616 11552
rect 19668 11540 19674 11552
rect 21008 11540 21036 11716
rect 21545 11713 21557 11716
rect 21591 11713 21603 11747
rect 22186 11744 22192 11756
rect 22147 11716 22192 11744
rect 21545 11707 21603 11713
rect 22186 11704 22192 11716
rect 22244 11704 22250 11756
rect 22278 11704 22284 11756
rect 22336 11744 22342 11756
rect 22554 11744 22560 11756
rect 22336 11716 22381 11744
rect 22515 11716 22560 11744
rect 22336 11704 22342 11716
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 27246 11753 27252 11756
rect 27240 11707 27252 11753
rect 27304 11744 27310 11756
rect 27304 11716 27340 11744
rect 27246 11704 27252 11707
rect 27304 11704 27310 11716
rect 22465 11679 22523 11685
rect 22465 11676 22477 11679
rect 21192 11648 22477 11676
rect 21192 11552 21220 11648
rect 22465 11645 22477 11648
rect 22511 11645 22523 11679
rect 22465 11639 22523 11645
rect 25038 11636 25044 11688
rect 25096 11676 25102 11688
rect 26973 11679 27031 11685
rect 26973 11676 26985 11679
rect 25096 11648 26985 11676
rect 25096 11636 25102 11648
rect 26973 11645 26985 11648
rect 27019 11645 27031 11679
rect 26973 11639 27031 11645
rect 22278 11568 22284 11620
rect 22336 11608 22342 11620
rect 22336 11580 22876 11608
rect 22336 11568 22342 11580
rect 21174 11540 21180 11552
rect 19668 11512 21036 11540
rect 21135 11512 21180 11540
rect 19668 11500 19674 11512
rect 21174 11500 21180 11512
rect 21232 11500 21238 11552
rect 22848 11549 22876 11580
rect 22833 11543 22891 11549
rect 22833 11509 22845 11543
rect 22879 11509 22891 11543
rect 23014 11540 23020 11552
rect 22975 11512 23020 11540
rect 22833 11503 22891 11509
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 28350 11540 28356 11552
rect 28311 11512 28356 11540
rect 28350 11500 28356 11512
rect 28408 11500 28414 11552
rect 1104 11450 29532 11472
rect 1104 11398 5688 11450
rect 5740 11398 5752 11450
rect 5804 11398 5816 11450
rect 5868 11398 5880 11450
rect 5932 11398 5944 11450
rect 5996 11398 15163 11450
rect 15215 11398 15227 11450
rect 15279 11398 15291 11450
rect 15343 11398 15355 11450
rect 15407 11398 15419 11450
rect 15471 11398 24639 11450
rect 24691 11398 24703 11450
rect 24755 11398 24767 11450
rect 24819 11398 24831 11450
rect 24883 11398 24895 11450
rect 24947 11398 29532 11450
rect 1104 11376 29532 11398
rect 3786 11296 3792 11348
rect 3844 11336 3850 11348
rect 3844 11308 6684 11336
rect 3844 11296 3850 11308
rect 1946 11268 1952 11280
rect 1907 11240 1952 11268
rect 1946 11228 1952 11240
rect 2004 11228 2010 11280
rect 5721 11271 5779 11277
rect 5721 11237 5733 11271
rect 5767 11237 5779 11271
rect 5721 11231 5779 11237
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4706 11200 4712 11212
rect 4212 11172 4712 11200
rect 4212 11160 4218 11172
rect 4706 11160 4712 11172
rect 4764 11200 4770 11212
rect 5077 11203 5135 11209
rect 5077 11200 5089 11203
rect 4764 11172 5089 11200
rect 4764 11160 4770 11172
rect 5077 11169 5089 11172
rect 5123 11169 5135 11203
rect 5736 11200 5764 11231
rect 6086 11228 6092 11280
rect 6144 11268 6150 11280
rect 6365 11271 6423 11277
rect 6365 11268 6377 11271
rect 6144 11240 6377 11268
rect 6144 11228 6150 11240
rect 6365 11237 6377 11240
rect 6411 11237 6423 11271
rect 6656 11268 6684 11308
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 6788 11308 6929 11336
rect 6788 11296 6794 11308
rect 6917 11305 6929 11308
rect 6963 11305 6975 11339
rect 6917 11299 6975 11305
rect 8938 11296 8944 11348
rect 8996 11336 9002 11348
rect 9033 11339 9091 11345
rect 9033 11336 9045 11339
rect 8996 11308 9045 11336
rect 8996 11296 9002 11308
rect 9033 11305 9045 11308
rect 9079 11305 9091 11339
rect 9033 11299 9091 11305
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 9180 11308 9229 11336
rect 9180 11296 9186 11308
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 9217 11299 9275 11305
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 11330 11336 11336 11348
rect 10192 11308 11336 11336
rect 10192 11296 10198 11308
rect 11330 11296 11336 11308
rect 11388 11336 11394 11348
rect 11606 11336 11612 11348
rect 11388 11308 11612 11336
rect 11388 11296 11394 11308
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 11977 11339 12035 11345
rect 11977 11305 11989 11339
rect 12023 11336 12035 11339
rect 12158 11336 12164 11348
rect 12023 11308 12164 11336
rect 12023 11305 12035 11308
rect 11977 11299 12035 11305
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 13909 11339 13967 11345
rect 13909 11336 13921 11339
rect 13780 11308 13921 11336
rect 13780 11296 13786 11308
rect 13909 11305 13921 11308
rect 13955 11305 13967 11339
rect 14642 11336 14648 11348
rect 14603 11308 14648 11336
rect 13909 11299 13967 11305
rect 7006 11268 7012 11280
rect 6656 11240 7012 11268
rect 6365 11231 6423 11237
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 7650 11268 7656 11280
rect 7611 11240 7656 11268
rect 7650 11228 7656 11240
rect 7708 11228 7714 11280
rect 10962 11268 10968 11280
rect 7760 11240 10968 11268
rect 7760 11200 7788 11240
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 11348 11240 12434 11268
rect 9214 11200 9220 11212
rect 5736 11172 6132 11200
rect 5077 11163 5135 11169
rect 2222 11132 2228 11144
rect 2135 11104 2228 11132
rect 2222 11092 2228 11104
rect 2280 11132 2286 11144
rect 4246 11132 4252 11144
rect 2280 11104 4252 11132
rect 2280 11092 2286 11104
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11132 5411 11135
rect 5534 11132 5540 11144
rect 5399 11104 5540 11132
rect 5399 11101 5411 11104
rect 5353 11095 5411 11101
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 5810 11132 5816 11144
rect 5771 11104 5816 11132
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 6104 11141 6132 11172
rect 7392 11172 7788 11200
rect 8036 11172 9220 11200
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 6178 11092 6184 11144
rect 6236 11141 6242 11144
rect 7392 11141 7420 11172
rect 6236 11132 6244 11141
rect 7009 11135 7067 11141
rect 6236 11104 6281 11132
rect 6236 11095 6244 11104
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7055 11104 7389 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 6236 11092 6242 11095
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 8036 11141 8064 11172
rect 9214 11160 9220 11172
rect 9272 11200 9278 11212
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 9272 11172 9321 11200
rect 9272 11160 9278 11172
rect 9309 11169 9321 11172
rect 9355 11169 9367 11203
rect 9953 11203 10011 11209
rect 9953 11200 9965 11203
rect 9309 11163 9367 11169
rect 9416 11172 9965 11200
rect 7895 11135 7953 11141
rect 7895 11132 7907 11135
rect 7524 11104 7907 11132
rect 7524 11092 7530 11104
rect 7895 11101 7907 11104
rect 7941 11101 7953 11135
rect 7895 11095 7953 11101
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8110 11092 8116 11144
rect 8168 11132 8174 11144
rect 8294 11132 8300 11144
rect 8168 11104 8213 11132
rect 8255 11104 8300 11132
rect 8168 11092 8174 11104
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 9416 11141 9444 11172
rect 9953 11169 9965 11172
rect 9999 11200 10011 11203
rect 10134 11200 10140 11212
rect 9999 11172 10140 11200
rect 9999 11169 10011 11172
rect 9953 11163 10011 11169
rect 10134 11160 10140 11172
rect 10192 11200 10198 11212
rect 10192 11172 11284 11200
rect 10192 11160 10198 11172
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11132 8539 11135
rect 9401 11135 9459 11141
rect 9401 11132 9413 11135
rect 8527 11104 9413 11132
rect 8527 11101 8539 11104
rect 8481 11095 8539 11101
rect 9401 11101 9413 11104
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9539 11104 9781 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 10318 11132 10324 11144
rect 10279 11104 10324 11132
rect 9769 11095 9827 11101
rect 5997 11067 6055 11073
rect 5997 11033 6009 11067
rect 6043 11033 6055 11067
rect 5997 11027 6055 11033
rect 8665 11067 8723 11073
rect 8665 11033 8677 11067
rect 8711 11064 8723 11067
rect 9030 11064 9036 11076
rect 8711 11036 9036 11064
rect 8711 11033 8723 11036
rect 8665 11027 8723 11033
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 1765 10999 1823 11005
rect 1765 10996 1777 10999
rect 1544 10968 1777 10996
rect 1544 10956 1550 10968
rect 1765 10965 1777 10968
rect 1811 10965 1823 10999
rect 5258 10996 5264 11008
rect 5219 10968 5264 10996
rect 1765 10959 1823 10965
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 6012 10996 6040 11027
rect 9030 11024 9036 11036
rect 9088 11064 9094 11076
rect 9508 11064 9536 11095
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 10686 11132 10692 11144
rect 10647 11104 10692 11132
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11132 11115 11135
rect 11146 11132 11152 11144
rect 11103 11104 11152 11132
rect 11103 11101 11115 11104
rect 11057 11095 11115 11101
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11256 11141 11284 11172
rect 11348 11141 11376 11240
rect 11698 11200 11704 11212
rect 11659 11172 11704 11200
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 11790 11160 11796 11212
rect 11848 11200 11854 11212
rect 12406 11200 12434 11240
rect 12526 11200 12532 11212
rect 11848 11172 11893 11200
rect 12406 11172 12532 11200
rect 11848 11160 11854 11172
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 13924 11200 13952 11299
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 15013 11339 15071 11345
rect 15013 11336 15025 11339
rect 14792 11308 15025 11336
rect 14792 11296 14798 11308
rect 15013 11305 15025 11308
rect 15059 11305 15071 11339
rect 15013 11299 15071 11305
rect 15381 11339 15439 11345
rect 15381 11305 15393 11339
rect 15427 11305 15439 11339
rect 15562 11336 15568 11348
rect 15523 11308 15568 11336
rect 15381 11299 15439 11305
rect 14660 11268 14688 11296
rect 15396 11268 15424 11299
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 16485 11339 16543 11345
rect 16485 11305 16497 11339
rect 16531 11336 16543 11339
rect 18138 11336 18144 11348
rect 16531 11308 18144 11336
rect 16531 11305 16543 11308
rect 16485 11299 16543 11305
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 19242 11296 19248 11348
rect 19300 11336 19306 11348
rect 19337 11339 19395 11345
rect 19337 11336 19349 11339
rect 19300 11308 19349 11336
rect 19300 11296 19306 11308
rect 19337 11305 19349 11308
rect 19383 11305 19395 11339
rect 19337 11299 19395 11305
rect 19518 11296 19524 11348
rect 19576 11336 19582 11348
rect 19797 11339 19855 11345
rect 19797 11336 19809 11339
rect 19576 11308 19809 11336
rect 19576 11296 19582 11308
rect 19797 11305 19809 11308
rect 19843 11305 19855 11339
rect 20806 11336 20812 11348
rect 19797 11299 19855 11305
rect 20364 11308 20812 11336
rect 14660 11240 15424 11268
rect 15378 11200 15384 11212
rect 13924 11172 15384 11200
rect 15378 11160 15384 11172
rect 15436 11200 15442 11212
rect 15436 11172 15976 11200
rect 15436 11160 15442 11172
rect 11241 11135 11299 11141
rect 11241 11101 11253 11135
rect 11287 11101 11299 11135
rect 11241 11095 11299 11101
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11101 11391 11135
rect 11514 11132 11520 11144
rect 11475 11104 11520 11132
rect 11333 11095 11391 11101
rect 9088 11036 9536 11064
rect 9585 11067 9643 11073
rect 9088 11024 9094 11036
rect 9585 11033 9597 11067
rect 9631 11064 9643 11067
rect 10226 11064 10232 11076
rect 9631 11036 10232 11064
rect 9631 11033 9643 11036
rect 9585 11027 9643 11033
rect 10226 11024 10232 11036
rect 10284 11024 10290 11076
rect 10413 11067 10471 11073
rect 10413 11033 10425 11067
rect 10459 11064 10471 11067
rect 10962 11064 10968 11076
rect 10459 11036 10968 11064
rect 10459 11033 10471 11036
rect 10413 11027 10471 11033
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 11256 11064 11284 11095
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11606 11092 11612 11144
rect 11664 11132 11670 11144
rect 11664 11104 11709 11132
rect 11664 11092 11670 11104
rect 12250 11092 12256 11144
rect 12308 11132 12314 11144
rect 13366 11135 13424 11141
rect 13366 11132 13378 11135
rect 12308 11104 13378 11132
rect 12308 11092 12314 11104
rect 13366 11101 13378 11104
rect 13412 11101 13424 11135
rect 13366 11095 13424 11101
rect 13538 11092 13544 11144
rect 13596 11132 13602 11144
rect 13725 11135 13783 11141
rect 13725 11132 13737 11135
rect 13596 11104 13737 11132
rect 13596 11092 13602 11104
rect 13725 11101 13737 11104
rect 13771 11132 13783 11135
rect 13906 11132 13912 11144
rect 13771 11104 13912 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 13906 11092 13912 11104
rect 13964 11132 13970 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13964 11104 14105 11132
rect 13964 11092 13970 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11132 14427 11135
rect 14642 11132 14648 11144
rect 14415 11104 14648 11132
rect 14415 11101 14427 11104
rect 14369 11095 14427 11101
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 14829 11135 14887 11141
rect 14829 11101 14841 11135
rect 14875 11101 14887 11135
rect 15746 11132 15752 11144
rect 15707 11104 15752 11132
rect 14829 11095 14887 11101
rect 11790 11064 11796 11076
rect 11256 11036 11796 11064
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 14844 11064 14872 11095
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 15948 11141 15976 11172
rect 19794 11160 19800 11212
rect 19852 11200 19858 11212
rect 19889 11203 19947 11209
rect 19889 11200 19901 11203
rect 19852 11172 19901 11200
rect 19852 11160 19858 11172
rect 19889 11169 19901 11172
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11132 16175 11135
rect 16301 11135 16359 11141
rect 16301 11132 16313 11135
rect 16163 11104 16313 11132
rect 16163 11101 16175 11104
rect 16117 11095 16175 11101
rect 16301 11101 16313 11104
rect 16347 11101 16359 11135
rect 16301 11095 16359 11101
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 18141 11135 18199 11141
rect 18141 11132 18153 11135
rect 16724 11104 18153 11132
rect 16724 11092 16730 11104
rect 18141 11101 18153 11104
rect 18187 11132 18199 11135
rect 19334 11132 19340 11144
rect 18187 11104 19340 11132
rect 18187 11101 18199 11104
rect 18141 11095 18199 11101
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 15197 11067 15255 11073
rect 15197 11064 15209 11067
rect 14844 11036 15209 11064
rect 15197 11033 15209 11036
rect 15243 11064 15255 11067
rect 15562 11064 15568 11076
rect 15243 11036 15568 11064
rect 15243 11033 15255 11036
rect 15197 11027 15255 11033
rect 15562 11024 15568 11036
rect 15620 11064 15626 11076
rect 15838 11064 15844 11076
rect 15620 11036 15844 11064
rect 15620 11024 15626 11036
rect 15838 11024 15844 11036
rect 15896 11064 15902 11076
rect 17896 11067 17954 11073
rect 15896 11036 16804 11064
rect 15896 11024 15902 11036
rect 6270 10996 6276 11008
rect 6012 10968 6276 10996
rect 6270 10956 6276 10968
rect 6328 10996 6334 11008
rect 7190 10996 7196 11008
rect 6328 10968 7196 10996
rect 6328 10956 6334 10968
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 10781 10999 10839 11005
rect 10781 10965 10793 10999
rect 10827 10996 10839 10999
rect 10870 10996 10876 11008
rect 10827 10968 10876 10996
rect 10827 10965 10839 10968
rect 10781 10959 10839 10965
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 12253 10999 12311 11005
rect 12253 10996 12265 10999
rect 11940 10968 12265 10996
rect 11940 10956 11946 10968
rect 12253 10965 12265 10968
rect 12299 10965 12311 10999
rect 12253 10959 12311 10965
rect 14553 10999 14611 11005
rect 14553 10965 14565 10999
rect 14599 10996 14611 10999
rect 15102 10996 15108 11008
rect 14599 10968 15108 10996
rect 14599 10965 14611 10968
rect 14553 10959 14611 10965
rect 15102 10956 15108 10968
rect 15160 10956 15166 11008
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 16776 11005 16804 11036
rect 17896 11033 17908 11067
rect 17942 11064 17954 11067
rect 18046 11064 18052 11076
rect 17942 11036 18052 11064
rect 17942 11033 17954 11036
rect 17896 11027 17954 11033
rect 18046 11024 18052 11036
rect 18104 11024 18110 11076
rect 19536 11064 19564 11095
rect 19610 11092 19616 11144
rect 19668 11132 19674 11144
rect 19904 11132 19932 11163
rect 20257 11135 20315 11141
rect 20257 11132 20269 11135
rect 19668 11104 19713 11132
rect 19904 11104 20269 11132
rect 19668 11092 19674 11104
rect 20257 11101 20269 11104
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 20165 11067 20223 11073
rect 20165 11064 20177 11067
rect 19536 11036 20177 11064
rect 20165 11033 20177 11036
rect 20211 11064 20223 11067
rect 20364 11064 20392 11308
rect 20806 11296 20812 11308
rect 20864 11336 20870 11348
rect 20901 11339 20959 11345
rect 20901 11336 20913 11339
rect 20864 11308 20913 11336
rect 20864 11296 20870 11308
rect 20901 11305 20913 11308
rect 20947 11305 20959 11339
rect 20901 11299 20959 11305
rect 22278 11296 22284 11348
rect 22336 11336 22342 11348
rect 22373 11339 22431 11345
rect 22373 11336 22385 11339
rect 22336 11308 22385 11336
rect 22336 11296 22342 11308
rect 22373 11305 22385 11308
rect 22419 11305 22431 11339
rect 27246 11336 27252 11348
rect 27207 11308 27252 11336
rect 22373 11299 22431 11305
rect 27246 11296 27252 11308
rect 27304 11296 27310 11348
rect 27157 11271 27215 11277
rect 27157 11237 27169 11271
rect 27203 11237 27215 11271
rect 27157 11231 27215 11237
rect 21085 11203 21143 11209
rect 21085 11169 21097 11203
rect 21131 11200 21143 11203
rect 21266 11200 21272 11212
rect 21131 11172 21272 11200
rect 21131 11169 21143 11172
rect 21085 11163 21143 11169
rect 21266 11160 21272 11172
rect 21324 11200 21330 11212
rect 21324 11172 23060 11200
rect 21324 11160 21330 11172
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 20990 11132 20996 11144
rect 20772 11104 20996 11132
rect 20772 11092 20778 11104
rect 20990 11092 20996 11104
rect 21048 11132 21054 11144
rect 21177 11135 21235 11141
rect 21177 11132 21189 11135
rect 21048 11104 21189 11132
rect 21048 11092 21054 11104
rect 21177 11101 21189 11104
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 21358 11092 21364 11144
rect 21416 11132 21422 11144
rect 23032 11141 23060 11172
rect 22281 11135 22339 11141
rect 22281 11132 22293 11135
rect 21416 11104 22293 11132
rect 21416 11092 21422 11104
rect 22281 11101 22293 11104
rect 22327 11101 22339 11135
rect 22281 11095 22339 11101
rect 23017 11135 23075 11141
rect 23017 11101 23029 11135
rect 23063 11132 23075 11135
rect 23106 11132 23112 11144
rect 23063 11104 23112 11132
rect 23063 11101 23075 11104
rect 23017 11095 23075 11101
rect 23106 11092 23112 11104
rect 23164 11092 23170 11144
rect 23842 11132 23848 11144
rect 23803 11104 23848 11132
rect 23842 11092 23848 11104
rect 23900 11092 23906 11144
rect 24026 11132 24032 11144
rect 23987 11104 24032 11132
rect 24026 11092 24032 11104
rect 24084 11092 24090 11144
rect 24397 11135 24455 11141
rect 24397 11101 24409 11135
rect 24443 11132 24455 11135
rect 25038 11132 25044 11144
rect 24443 11104 25044 11132
rect 24443 11101 24455 11104
rect 24397 11095 24455 11101
rect 20211 11036 20392 11064
rect 20901 11067 20959 11073
rect 20211 11033 20223 11036
rect 20165 11027 20223 11033
rect 20901 11033 20913 11067
rect 20947 11064 20959 11067
rect 21450 11064 21456 11076
rect 20947 11036 21456 11064
rect 20947 11033 20959 11036
rect 20901 11027 20959 11033
rect 21450 11024 21456 11036
rect 21508 11064 21514 11076
rect 22370 11064 22376 11076
rect 21508 11036 22376 11064
rect 21508 11024 21514 11036
rect 22370 11024 22376 11036
rect 22428 11024 22434 11076
rect 23661 11067 23719 11073
rect 23661 11033 23673 11067
rect 23707 11064 23719 11067
rect 24412 11064 24440 11095
rect 25038 11092 25044 11104
rect 25096 11092 25102 11144
rect 26970 11132 26976 11144
rect 26931 11104 26976 11132
rect 26970 11092 26976 11104
rect 27028 11092 27034 11144
rect 27172 11132 27200 11231
rect 27893 11203 27951 11209
rect 27893 11169 27905 11203
rect 27939 11200 27951 11203
rect 28442 11200 28448 11212
rect 27939 11172 28448 11200
rect 27939 11169 27951 11172
rect 27893 11163 27951 11169
rect 28442 11160 28448 11172
rect 28500 11160 28506 11212
rect 27617 11135 27675 11141
rect 27617 11132 27629 11135
rect 27172 11104 27629 11132
rect 27617 11101 27629 11104
rect 27663 11101 27675 11135
rect 27617 11095 27675 11101
rect 23707 11036 24440 11064
rect 23707 11033 23719 11036
rect 23661 11027 23719 11033
rect 24486 11024 24492 11076
rect 24544 11064 24550 11076
rect 24642 11067 24700 11073
rect 24642 11064 24654 11067
rect 24544 11036 24654 11064
rect 24544 11024 24550 11036
rect 24642 11033 24654 11036
rect 24688 11033 24700 11067
rect 26050 11064 26056 11076
rect 26011 11036 26056 11064
rect 24642 11027 24700 11033
rect 26050 11024 26056 11036
rect 26108 11024 26114 11076
rect 26237 11067 26295 11073
rect 26237 11033 26249 11067
rect 26283 11064 26295 11067
rect 26418 11064 26424 11076
rect 26283 11036 26317 11064
rect 26379 11036 26424 11064
rect 26283 11033 26295 11036
rect 26237 11027 26295 11033
rect 15381 10999 15439 11005
rect 15381 10996 15393 10999
rect 15344 10968 15393 10996
rect 15344 10956 15350 10968
rect 15381 10965 15393 10968
rect 15427 10965 15439 10999
rect 15381 10959 15439 10965
rect 16761 10999 16819 11005
rect 16761 10965 16773 10999
rect 16807 10965 16819 10999
rect 21358 10996 21364 11008
rect 21319 10968 21364 10996
rect 16761 10959 16819 10965
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 22738 10956 22744 11008
rect 22796 10996 22802 11008
rect 22925 10999 22983 11005
rect 22925 10996 22937 10999
rect 22796 10968 22937 10996
rect 22796 10956 22802 10968
rect 22925 10965 22937 10968
rect 22971 10965 22983 10999
rect 22925 10959 22983 10965
rect 24213 10999 24271 11005
rect 24213 10965 24225 10999
rect 24259 10996 24271 10999
rect 24762 10996 24768 11008
rect 24259 10968 24768 10996
rect 24259 10965 24271 10968
rect 24213 10959 24271 10965
rect 24762 10956 24768 10968
rect 24820 10956 24826 11008
rect 25777 10999 25835 11005
rect 25777 10965 25789 10999
rect 25823 10996 25835 10999
rect 26252 10996 26280 11027
rect 26418 11024 26424 11036
rect 26476 11024 26482 11076
rect 27632 11064 27660 11095
rect 27982 11092 27988 11144
rect 28040 11132 28046 11144
rect 28077 11135 28135 11141
rect 28077 11132 28089 11135
rect 28040 11104 28089 11132
rect 28040 11092 28046 11104
rect 28077 11101 28089 11104
rect 28123 11101 28135 11135
rect 28077 11095 28135 11101
rect 28261 11135 28319 11141
rect 28261 11101 28273 11135
rect 28307 11101 28319 11135
rect 28261 11095 28319 11101
rect 28276 11064 28304 11095
rect 27632 11036 28304 11064
rect 26326 10996 26332 11008
rect 25823 10968 26332 10996
rect 25823 10965 25835 10968
rect 25777 10959 25835 10965
rect 26326 10956 26332 10968
rect 26384 10956 26390 11008
rect 27706 10956 27712 11008
rect 27764 10996 27770 11008
rect 27764 10968 27809 10996
rect 27764 10956 27770 10968
rect 27890 10956 27896 11008
rect 27948 10996 27954 11008
rect 28445 10999 28503 11005
rect 28445 10996 28457 10999
rect 27948 10968 28457 10996
rect 27948 10956 27954 10968
rect 28445 10965 28457 10968
rect 28491 10965 28503 10999
rect 28445 10959 28503 10965
rect 1104 10906 29532 10928
rect 1104 10854 10425 10906
rect 10477 10854 10489 10906
rect 10541 10854 10553 10906
rect 10605 10854 10617 10906
rect 10669 10854 10681 10906
rect 10733 10854 19901 10906
rect 19953 10854 19965 10906
rect 20017 10854 20029 10906
rect 20081 10854 20093 10906
rect 20145 10854 20157 10906
rect 20209 10854 29532 10906
rect 1104 10832 29532 10854
rect 4154 10792 4160 10804
rect 4115 10764 4160 10792
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 5460 10764 6561 10792
rect 5460 10733 5488 10764
rect 6549 10761 6561 10764
rect 6595 10792 6607 10795
rect 7466 10792 7472 10804
rect 6595 10764 7472 10792
rect 6595 10761 6607 10764
rect 6549 10755 6607 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7561 10795 7619 10801
rect 7561 10761 7573 10795
rect 7607 10792 7619 10795
rect 8294 10792 8300 10804
rect 7607 10764 8300 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 9033 10795 9091 10801
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9674 10792 9680 10804
rect 9079 10764 9680 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 9674 10752 9680 10764
rect 9732 10792 9738 10804
rect 10042 10792 10048 10804
rect 9732 10764 10048 10792
rect 9732 10752 9738 10764
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 10376 10764 10517 10792
rect 10376 10752 10382 10764
rect 10505 10761 10517 10764
rect 10551 10761 10563 10795
rect 10505 10755 10563 10761
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11149 10795 11207 10801
rect 11149 10792 11161 10795
rect 11112 10764 11161 10792
rect 11112 10752 11118 10764
rect 11149 10761 11161 10764
rect 11195 10761 11207 10795
rect 11149 10755 11207 10761
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 12069 10795 12127 10801
rect 12069 10792 12081 10795
rect 11664 10764 12081 10792
rect 11664 10752 11670 10764
rect 12069 10761 12081 10764
rect 12115 10761 12127 10795
rect 13078 10792 13084 10804
rect 13039 10764 13084 10792
rect 12069 10755 12127 10761
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 14642 10752 14648 10804
rect 14700 10792 14706 10804
rect 14737 10795 14795 10801
rect 14737 10792 14749 10795
rect 14700 10764 14749 10792
rect 14700 10752 14706 10764
rect 14737 10761 14749 10764
rect 14783 10761 14795 10795
rect 14737 10755 14795 10761
rect 15105 10795 15163 10801
rect 15105 10761 15117 10795
rect 15151 10792 15163 10795
rect 15286 10792 15292 10804
rect 15151 10764 15292 10792
rect 15151 10761 15163 10764
rect 15105 10755 15163 10761
rect 15286 10752 15292 10764
rect 15344 10792 15350 10804
rect 16482 10792 16488 10804
rect 15344 10764 16488 10792
rect 15344 10752 15350 10764
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 17310 10792 17316 10804
rect 17000 10764 17316 10792
rect 17000 10752 17006 10764
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17957 10795 18015 10801
rect 17957 10761 17969 10795
rect 18003 10792 18015 10795
rect 18046 10792 18052 10804
rect 18003 10764 18052 10792
rect 18003 10761 18015 10764
rect 17957 10755 18015 10761
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 18156 10764 23060 10792
rect 5445 10727 5503 10733
rect 5445 10693 5457 10727
rect 5491 10693 5503 10727
rect 5445 10687 5503 10693
rect 5629 10727 5687 10733
rect 5629 10693 5641 10727
rect 5675 10724 5687 10727
rect 5810 10724 5816 10736
rect 5675 10696 5816 10724
rect 5675 10693 5687 10696
rect 5629 10687 5687 10693
rect 5810 10684 5816 10696
rect 5868 10684 5874 10736
rect 7377 10727 7435 10733
rect 7377 10693 7389 10727
rect 7423 10724 7435 10727
rect 8386 10724 8392 10736
rect 7423 10696 8392 10724
rect 7423 10693 7435 10696
rect 7377 10687 7435 10693
rect 8386 10684 8392 10696
rect 8444 10684 8450 10736
rect 9950 10724 9956 10736
rect 9600 10696 9956 10724
rect 1486 10656 1492 10668
rect 1447 10628 1492 10656
rect 1486 10616 1492 10628
rect 1544 10616 1550 10668
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 2021 10659 2079 10665
rect 2021 10656 2033 10659
rect 1912 10628 2033 10656
rect 1912 10616 1918 10628
rect 2021 10625 2033 10628
rect 2067 10625 2079 10659
rect 2021 10619 2079 10625
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3200 10628 3985 10656
rect 3200 10616 3206 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 5258 10656 5264 10668
rect 5219 10628 5264 10656
rect 3973 10619 4031 10625
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5592 10628 6377 10656
rect 5592 10616 5598 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1728 10560 1777 10588
rect 1728 10548 1734 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 6380 10520 6408 10619
rect 7742 10616 7748 10668
rect 7800 10656 7806 10668
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 7800 10628 7941 10656
rect 7800 10616 7806 10628
rect 7929 10625 7941 10628
rect 7975 10625 7987 10659
rect 8202 10656 8208 10668
rect 8115 10628 8208 10656
rect 7929 10619 7987 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 9600 10665 9628 10696
rect 9950 10684 9956 10696
rect 10008 10684 10014 10736
rect 10134 10724 10140 10736
rect 10095 10696 10140 10724
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 10226 10684 10232 10736
rect 10284 10724 10290 10736
rect 10597 10727 10655 10733
rect 10597 10724 10609 10727
rect 10284 10696 10609 10724
rect 10284 10684 10290 10696
rect 10597 10693 10609 10696
rect 10643 10693 10655 10727
rect 18156 10724 18184 10764
rect 19334 10724 19340 10736
rect 10597 10687 10655 10693
rect 11348 10696 12020 10724
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10588 7895 10591
rect 8110 10588 8116 10600
rect 7883 10560 8116 10588
rect 7883 10557 7895 10560
rect 7837 10551 7895 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8220 10520 8248 10616
rect 6380 10492 8248 10520
rect 1673 10455 1731 10461
rect 1673 10421 1685 10455
rect 1719 10452 1731 10455
rect 2130 10452 2136 10464
rect 1719 10424 2136 10452
rect 1719 10421 1731 10424
rect 1673 10415 1731 10421
rect 2130 10412 2136 10424
rect 2188 10412 2194 10464
rect 3145 10455 3203 10461
rect 3145 10421 3157 10455
rect 3191 10452 3203 10455
rect 3234 10452 3240 10464
rect 3191 10424 3240 10452
rect 3191 10421 3203 10424
rect 3145 10415 3203 10421
rect 3234 10412 3240 10424
rect 3292 10452 3298 10464
rect 4062 10452 4068 10464
rect 3292 10424 4068 10452
rect 3292 10412 3298 10424
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 7377 10455 7435 10461
rect 7377 10421 7389 10455
rect 7423 10452 7435 10455
rect 7745 10455 7803 10461
rect 7745 10452 7757 10455
rect 7423 10424 7757 10452
rect 7423 10421 7435 10424
rect 7377 10415 7435 10421
rect 7745 10421 7757 10424
rect 7791 10421 7803 10455
rect 8110 10452 8116 10464
rect 8071 10424 8116 10452
rect 7745 10415 7803 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 9214 10452 9220 10464
rect 9175 10424 9220 10452
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 9416 10452 9444 10619
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 9861 10659 9919 10665
rect 9732 10628 9777 10656
rect 9732 10616 9738 10628
rect 9861 10625 9873 10659
rect 9907 10656 9919 10659
rect 10042 10656 10048 10668
rect 9907 10628 10048 10656
rect 9907 10625 9919 10628
rect 9861 10619 9919 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 10393 10659 10451 10665
rect 10393 10625 10405 10659
rect 10439 10656 10451 10659
rect 10502 10656 10508 10668
rect 10439 10628 10508 10656
rect 10439 10625 10451 10628
rect 10393 10619 10451 10625
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 10612 10588 10640 10687
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10654 10747 10659
rect 10870 10656 10876 10668
rect 10796 10654 10876 10656
rect 10735 10628 10876 10654
rect 10735 10626 10824 10628
rect 10735 10625 10747 10626
rect 10689 10619 10747 10625
rect 10870 10616 10876 10628
rect 10928 10656 10934 10668
rect 11348 10665 11376 10696
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 10928 10628 11345 10656
rect 10928 10616 10934 10628
rect 11333 10625 11345 10628
rect 11379 10625 11391 10659
rect 11698 10656 11704 10668
rect 11659 10628 11704 10656
rect 11333 10619 11391 10625
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 11882 10656 11888 10668
rect 11843 10628 11888 10656
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 11992 10665 12020 10696
rect 12406 10696 18184 10724
rect 19295 10696 19340 10724
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 12161 10659 12219 10665
rect 12161 10656 12173 10659
rect 12124 10628 12173 10656
rect 12124 10616 12130 10628
rect 12161 10625 12173 10628
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 10962 10588 10968 10600
rect 10612 10560 10824 10588
rect 10923 10560 10968 10588
rect 9493 10523 9551 10529
rect 9493 10489 9505 10523
rect 9539 10520 9551 10523
rect 10410 10520 10416 10532
rect 9539 10492 10416 10520
rect 9539 10489 9551 10492
rect 9493 10483 9551 10489
rect 10410 10480 10416 10492
rect 10468 10480 10474 10532
rect 10686 10452 10692 10464
rect 9416 10424 10692 10452
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 10796 10461 10824 10560
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 12406 10588 12434 10696
rect 19334 10684 19340 10696
rect 19392 10684 19398 10736
rect 19521 10727 19579 10733
rect 19521 10693 19533 10727
rect 19567 10724 19579 10727
rect 19702 10724 19708 10736
rect 19567 10696 19708 10724
rect 19567 10693 19579 10696
rect 19521 10687 19579 10693
rect 19702 10684 19708 10696
rect 19760 10684 19766 10736
rect 13265 10659 13323 10665
rect 13265 10625 13277 10659
rect 13311 10656 13323 10659
rect 13722 10656 13728 10668
rect 13311 10628 13728 10656
rect 13311 10625 13323 10628
rect 13265 10619 13323 10625
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 14826 10656 14832 10668
rect 14787 10628 14832 10656
rect 14826 10616 14832 10628
rect 14884 10656 14890 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 14884 10628 14933 10656
rect 14884 10616 14890 10628
rect 14921 10625 14933 10628
rect 14967 10625 14979 10659
rect 15194 10656 15200 10668
rect 15107 10628 15200 10656
rect 14921 10619 14979 10625
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 15378 10656 15384 10668
rect 15339 10628 15384 10656
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 15657 10659 15715 10665
rect 15657 10656 15669 10659
rect 15611 10628 15669 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 15657 10625 15669 10628
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 17589 10659 17647 10665
rect 17589 10625 17601 10659
rect 17635 10625 17647 10659
rect 18138 10656 18144 10668
rect 18099 10628 18144 10656
rect 17589 10619 17647 10625
rect 11112 10560 12434 10588
rect 15212 10588 15240 10616
rect 17310 10588 17316 10600
rect 15212 10560 15700 10588
rect 17271 10560 17316 10588
rect 11112 10548 11118 10560
rect 15672 10532 15700 10560
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 17497 10591 17555 10597
rect 17497 10557 17509 10591
rect 17543 10557 17555 10591
rect 17604 10588 17632 10619
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 18233 10659 18291 10665
rect 18233 10625 18245 10659
rect 18279 10656 18291 10659
rect 18322 10656 18328 10668
rect 18279 10628 18328 10656
rect 18279 10625 18291 10628
rect 18233 10619 18291 10625
rect 18322 10616 18328 10628
rect 18380 10656 18386 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18380 10628 18613 10656
rect 18380 10616 18386 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 18414 10588 18420 10600
rect 17604 10560 18420 10588
rect 17497 10551 17555 10557
rect 10870 10480 10876 10532
rect 10928 10520 10934 10532
rect 11609 10523 11667 10529
rect 11609 10520 11621 10523
rect 10928 10492 11621 10520
rect 10928 10480 10934 10492
rect 11609 10489 11621 10492
rect 11655 10489 11667 10523
rect 11609 10483 11667 10489
rect 15654 10480 15660 10532
rect 15712 10480 15718 10532
rect 17402 10480 17408 10532
rect 17460 10520 17466 10532
rect 17512 10520 17540 10551
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 19352 10588 19380 10684
rect 20438 10616 20444 10668
rect 20496 10656 20502 10668
rect 21085 10659 21143 10665
rect 21085 10656 21097 10659
rect 20496 10628 21097 10656
rect 20496 10616 20502 10628
rect 21085 10625 21097 10628
rect 21131 10625 21143 10659
rect 21085 10619 21143 10625
rect 21174 10616 21180 10668
rect 21232 10656 21238 10668
rect 21269 10659 21327 10665
rect 21269 10656 21281 10659
rect 21232 10628 21281 10656
rect 21232 10616 21238 10628
rect 21269 10625 21281 10628
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 21361 10659 21419 10665
rect 21361 10625 21373 10659
rect 21407 10656 21419 10659
rect 21450 10656 21456 10668
rect 21407 10628 21456 10656
rect 21407 10625 21419 10628
rect 21361 10619 21419 10625
rect 21450 10616 21456 10628
rect 21508 10616 21514 10668
rect 22370 10616 22376 10668
rect 22428 10656 22434 10668
rect 22537 10659 22595 10665
rect 22537 10656 22549 10659
rect 22428 10628 22549 10656
rect 22428 10616 22434 10628
rect 22537 10625 22549 10628
rect 22583 10625 22595 10659
rect 23032 10656 23060 10764
rect 23106 10752 23112 10804
rect 23164 10792 23170 10804
rect 23661 10795 23719 10801
rect 23661 10792 23673 10795
rect 23164 10764 23673 10792
rect 23164 10752 23170 10764
rect 23661 10761 23673 10764
rect 23707 10761 23719 10795
rect 23661 10755 23719 10761
rect 24305 10795 24363 10801
rect 24305 10761 24317 10795
rect 24351 10792 24363 10795
rect 24486 10792 24492 10804
rect 24351 10764 24492 10792
rect 24351 10761 24363 10764
rect 24305 10755 24363 10761
rect 24486 10752 24492 10764
rect 24544 10752 24550 10804
rect 24762 10792 24768 10804
rect 24723 10764 24768 10792
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 25133 10795 25191 10801
rect 25133 10761 25145 10795
rect 25179 10761 25191 10795
rect 27706 10792 27712 10804
rect 27667 10764 27712 10792
rect 25133 10755 25191 10761
rect 24673 10727 24731 10733
rect 24673 10724 24685 10727
rect 24504 10696 24685 10724
rect 24504 10668 24532 10696
rect 24673 10693 24685 10696
rect 24719 10724 24731 10727
rect 25148 10724 25176 10755
rect 27706 10752 27712 10764
rect 27764 10752 27770 10804
rect 26329 10727 26387 10733
rect 26329 10724 26341 10727
rect 24719 10696 25176 10724
rect 26252 10696 26341 10724
rect 24719 10693 24731 10696
rect 24673 10687 24731 10693
rect 23032 10628 23336 10656
rect 22537 10619 22595 10625
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 19352 10560 22293 10588
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 21177 10523 21235 10529
rect 17460 10492 18460 10520
rect 17460 10480 17466 10492
rect 10781 10455 10839 10461
rect 10781 10421 10793 10455
rect 10827 10421 10839 10455
rect 10781 10415 10839 10421
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 18432 10461 18460 10492
rect 21177 10489 21189 10523
rect 21223 10520 21235 10523
rect 21266 10520 21272 10532
rect 21223 10492 21272 10520
rect 21223 10489 21235 10492
rect 21177 10483 21235 10489
rect 21266 10480 21272 10492
rect 21324 10480 21330 10532
rect 23308 10520 23336 10628
rect 24486 10616 24492 10668
rect 24544 10616 24550 10668
rect 25317 10659 25375 10665
rect 25317 10625 25329 10659
rect 25363 10656 25375 10659
rect 25593 10659 25651 10665
rect 25593 10656 25605 10659
rect 25363 10628 25605 10656
rect 25363 10625 25375 10628
rect 25317 10619 25375 10625
rect 25593 10625 25605 10628
rect 25639 10625 25651 10659
rect 25593 10619 25651 10625
rect 25835 10659 25893 10665
rect 25835 10625 25847 10659
rect 25881 10656 25893 10659
rect 26050 10656 26056 10668
rect 25881 10628 26056 10656
rect 25881 10625 25893 10628
rect 25835 10619 25893 10625
rect 26050 10616 26056 10628
rect 26108 10616 26114 10668
rect 26252 10665 26280 10696
rect 26329 10693 26341 10696
rect 26375 10724 26387 10727
rect 26418 10724 26424 10736
rect 26375 10696 26424 10724
rect 26375 10693 26387 10696
rect 26329 10687 26387 10693
rect 26418 10684 26424 10696
rect 26476 10724 26482 10736
rect 26970 10724 26976 10736
rect 26476 10696 26832 10724
rect 26931 10696 26976 10724
rect 26476 10684 26482 10696
rect 26237 10659 26295 10665
rect 26237 10625 26249 10659
rect 26283 10625 26295 10659
rect 26237 10619 26295 10625
rect 26513 10659 26571 10665
rect 26513 10625 26525 10659
rect 26559 10625 26571 10659
rect 26694 10656 26700 10668
rect 26655 10628 26700 10656
rect 26513 10619 26571 10625
rect 23382 10548 23388 10600
rect 23440 10588 23446 10600
rect 24857 10591 24915 10597
rect 24857 10588 24869 10591
rect 23440 10560 24869 10588
rect 23440 10548 23446 10560
rect 24857 10557 24869 10560
rect 24903 10557 24915 10591
rect 24857 10551 24915 10557
rect 26145 10591 26203 10597
rect 26145 10557 26157 10591
rect 26191 10588 26203 10591
rect 26326 10588 26332 10600
rect 26191 10560 26332 10588
rect 26191 10557 26203 10560
rect 26145 10551 26203 10557
rect 26326 10548 26332 10560
rect 26384 10548 26390 10600
rect 26528 10588 26556 10619
rect 26694 10616 26700 10628
rect 26752 10616 26758 10668
rect 26804 10656 26832 10696
rect 26970 10684 26976 10696
rect 27028 10684 27034 10736
rect 28350 10724 28356 10736
rect 27540 10696 28356 10724
rect 27540 10665 27568 10696
rect 28350 10684 28356 10696
rect 28408 10684 28414 10736
rect 27158 10659 27216 10665
rect 27158 10656 27170 10659
rect 26804 10628 27170 10656
rect 27158 10625 27170 10628
rect 27204 10625 27216 10659
rect 27158 10619 27216 10625
rect 27525 10659 27583 10665
rect 27525 10625 27537 10659
rect 27571 10625 27583 10659
rect 27890 10656 27896 10668
rect 27851 10628 27896 10656
rect 27525 10619 27583 10625
rect 27540 10588 27568 10619
rect 27890 10616 27896 10628
rect 27948 10616 27954 10668
rect 26528 10560 27568 10588
rect 27617 10591 27675 10597
rect 26712 10532 26740 10560
rect 27617 10557 27629 10591
rect 27663 10557 27675 10591
rect 27617 10551 27675 10557
rect 25498 10520 25504 10532
rect 23308 10492 25504 10520
rect 25498 10480 25504 10492
rect 25556 10480 25562 10532
rect 26694 10480 26700 10532
rect 26752 10480 26758 10532
rect 26786 10480 26792 10532
rect 26844 10520 26850 10532
rect 27632 10520 27660 10551
rect 26844 10492 27660 10520
rect 26844 10480 26850 10492
rect 15841 10455 15899 10461
rect 15841 10452 15853 10455
rect 15804 10424 15853 10452
rect 15804 10412 15810 10424
rect 15841 10421 15853 10424
rect 15887 10421 15899 10455
rect 15841 10415 15899 10421
rect 18417 10455 18475 10461
rect 18417 10421 18429 10455
rect 18463 10421 18475 10455
rect 21542 10452 21548 10464
rect 21503 10424 21548 10452
rect 18417 10415 18475 10421
rect 21542 10412 21548 10424
rect 21600 10412 21606 10464
rect 21634 10412 21640 10464
rect 21692 10452 21698 10464
rect 27522 10452 27528 10464
rect 21692 10424 27528 10452
rect 21692 10412 21698 10424
rect 27522 10412 27528 10424
rect 27580 10412 27586 10464
rect 1104 10362 29532 10384
rect 1104 10310 5688 10362
rect 5740 10310 5752 10362
rect 5804 10310 5816 10362
rect 5868 10310 5880 10362
rect 5932 10310 5944 10362
rect 5996 10310 15163 10362
rect 15215 10310 15227 10362
rect 15279 10310 15291 10362
rect 15343 10310 15355 10362
rect 15407 10310 15419 10362
rect 15471 10310 24639 10362
rect 24691 10310 24703 10362
rect 24755 10310 24767 10362
rect 24819 10310 24831 10362
rect 24883 10310 24895 10362
rect 24947 10310 29532 10362
rect 1104 10288 29532 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 3605 10251 3663 10257
rect 3605 10217 3617 10251
rect 3651 10248 3663 10251
rect 4522 10248 4528 10260
rect 3651 10220 4528 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 4522 10208 4528 10220
rect 4580 10248 4586 10260
rect 4617 10251 4675 10257
rect 4617 10248 4629 10251
rect 4580 10220 4629 10248
rect 4580 10208 4586 10220
rect 4617 10217 4629 10220
rect 4663 10217 4675 10251
rect 4617 10211 4675 10217
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7800 10220 7849 10248
rect 7800 10208 7806 10220
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 10318 10248 10324 10260
rect 10279 10220 10324 10248
rect 7837 10211 7895 10217
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 14185 10251 14243 10257
rect 14185 10217 14197 10251
rect 14231 10248 14243 10251
rect 14826 10248 14832 10260
rect 14231 10220 14832 10248
rect 14231 10217 14243 10220
rect 14185 10211 14243 10217
rect 14826 10208 14832 10220
rect 14884 10208 14890 10260
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 16853 10251 16911 10257
rect 16853 10248 16865 10251
rect 16632 10220 16865 10248
rect 16632 10208 16638 10220
rect 16853 10217 16865 10220
rect 16899 10248 16911 10251
rect 17678 10248 17684 10260
rect 16899 10220 17684 10248
rect 16899 10217 16911 10220
rect 16853 10211 16911 10217
rect 17678 10208 17684 10220
rect 17736 10248 17742 10260
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 17736 10220 18245 10248
rect 17736 10208 17742 10220
rect 18233 10217 18245 10220
rect 18279 10217 18291 10251
rect 18233 10211 18291 10217
rect 24026 10208 24032 10260
rect 24084 10248 24090 10260
rect 24489 10251 24547 10257
rect 24489 10248 24501 10251
rect 24084 10220 24501 10248
rect 24084 10208 24090 10220
rect 24489 10217 24501 10220
rect 24535 10217 24547 10251
rect 24489 10211 24547 10217
rect 26326 10208 26332 10260
rect 26384 10248 26390 10260
rect 26697 10251 26755 10257
rect 26697 10248 26709 10251
rect 26384 10220 26709 10248
rect 26384 10208 26390 10220
rect 26697 10217 26709 10220
rect 26743 10217 26755 10251
rect 26697 10211 26755 10217
rect 3789 10183 3847 10189
rect 3789 10149 3801 10183
rect 3835 10149 3847 10183
rect 3789 10143 3847 10149
rect 1946 10072 1952 10124
rect 2004 10112 2010 10124
rect 2317 10115 2375 10121
rect 2317 10112 2329 10115
rect 2004 10084 2329 10112
rect 2004 10072 2010 10084
rect 2317 10081 2329 10084
rect 2363 10081 2375 10115
rect 2317 10075 2375 10081
rect 2130 10004 2136 10056
rect 2188 10044 2194 10056
rect 2225 10047 2283 10053
rect 2225 10044 2237 10047
rect 2188 10016 2237 10044
rect 2188 10004 2194 10016
rect 2225 10013 2237 10016
rect 2271 10013 2283 10047
rect 2332 10044 2360 10075
rect 2406 10072 2412 10124
rect 2464 10112 2470 10124
rect 3804 10112 3832 10143
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 4028 10152 6132 10180
rect 4028 10140 4034 10152
rect 4430 10112 4436 10124
rect 2464 10084 2509 10112
rect 3344 10084 3832 10112
rect 4391 10084 4436 10112
rect 2464 10072 2470 10084
rect 3344 10053 3372 10084
rect 4430 10072 4436 10084
rect 4488 10112 4494 10124
rect 5169 10115 5227 10121
rect 5169 10112 5181 10115
rect 4488 10084 5181 10112
rect 4488 10072 4494 10084
rect 5169 10081 5181 10084
rect 5215 10081 5227 10115
rect 5994 10112 6000 10124
rect 5955 10084 6000 10112
rect 5169 10075 5227 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 6104 10112 6132 10152
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 10689 10183 10747 10189
rect 10689 10180 10701 10183
rect 10100 10152 10701 10180
rect 10100 10140 10106 10152
rect 10689 10149 10701 10152
rect 10735 10149 10747 10183
rect 12710 10180 12716 10192
rect 12671 10152 12716 10180
rect 10689 10143 10747 10149
rect 12710 10140 12716 10152
rect 12768 10140 12774 10192
rect 21634 10180 21640 10192
rect 16408 10152 21640 10180
rect 8846 10112 8852 10124
rect 6104 10084 6592 10112
rect 3329 10047 3387 10053
rect 3329 10044 3341 10047
rect 2332 10016 3341 10044
rect 2225 10007 2283 10013
rect 3329 10013 3341 10016
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 3467 10016 4108 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 3602 9976 3608 9988
rect 3563 9948 3608 9976
rect 3602 9936 3608 9948
rect 3660 9936 3666 9988
rect 4080 9976 4108 10016
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 5077 10047 5135 10053
rect 5077 10044 5089 10047
rect 4212 10016 5089 10044
rect 4212 10004 4218 10016
rect 5077 10013 5089 10016
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 6086 10044 6092 10056
rect 5859 10016 6092 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 6362 10004 6368 10056
rect 6420 10044 6426 10056
rect 6457 10047 6515 10053
rect 6457 10044 6469 10047
rect 6420 10016 6469 10044
rect 6420 10004 6426 10016
rect 6457 10013 6469 10016
rect 6503 10013 6515 10047
rect 6564 10044 6592 10084
rect 8220 10084 8852 10112
rect 8220 10053 8248 10084
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 10870 10112 10876 10124
rect 10468 10084 10732 10112
rect 10831 10084 10876 10112
rect 10468 10072 10474 10084
rect 8205 10047 8263 10053
rect 6564 10016 8156 10044
rect 6457 10007 6515 10013
rect 4338 9976 4344 9988
rect 4080 9948 4344 9976
rect 4338 9936 4344 9948
rect 4396 9936 4402 9988
rect 4614 9936 4620 9988
rect 4672 9976 4678 9988
rect 5258 9976 5264 9988
rect 4672 9948 5264 9976
rect 4672 9936 4678 9948
rect 5258 9936 5264 9948
rect 5316 9976 5322 9988
rect 5905 9979 5963 9985
rect 5905 9976 5917 9979
rect 5316 9948 5917 9976
rect 5316 9936 5322 9948
rect 5905 9945 5917 9948
rect 5951 9945 5963 9979
rect 5905 9939 5963 9945
rect 6724 9979 6782 9985
rect 6724 9945 6736 9979
rect 6770 9976 6782 9979
rect 8021 9979 8079 9985
rect 8021 9976 8033 9979
rect 6770 9948 8033 9976
rect 6770 9945 6782 9948
rect 6724 9939 6782 9945
rect 8021 9945 8033 9948
rect 8067 9945 8079 9979
rect 8128 9976 8156 10016
rect 8205 10013 8217 10047
rect 8251 10013 8263 10047
rect 8205 10007 8263 10013
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 8478 10044 8484 10056
rect 8435 10016 8484 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8938 10044 8944 10056
rect 8899 10016 8944 10044
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9214 10053 9220 10056
rect 9208 10044 9220 10053
rect 9175 10016 9220 10044
rect 9208 10007 9220 10016
rect 9214 10004 9220 10007
rect 9272 10004 9278 10056
rect 10704 10053 10732 10084
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 10962 10072 10968 10124
rect 11020 10072 11026 10124
rect 16408 10112 16436 10152
rect 21634 10140 21640 10152
rect 21692 10140 21698 10192
rect 11164 10084 14596 10112
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10013 10747 10047
rect 10980 10044 11008 10072
rect 11057 10047 11115 10053
rect 11057 10044 11069 10047
rect 10980 10016 11069 10044
rect 10689 10007 10747 10013
rect 11057 10013 11069 10016
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 10962 9976 10968 9988
rect 8128 9948 10968 9976
rect 8021 9939 8079 9945
rect 10962 9936 10968 9948
rect 11020 9936 11026 9988
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4157 9911 4215 9917
rect 4157 9908 4169 9911
rect 4120 9880 4169 9908
rect 4120 9868 4126 9880
rect 4157 9877 4169 9880
rect 4203 9877 4215 9911
rect 4157 9871 4215 9877
rect 4246 9868 4252 9920
rect 4304 9908 4310 9920
rect 4982 9908 4988 9920
rect 4304 9880 4349 9908
rect 4943 9880 4988 9908
rect 4304 9868 4310 9880
rect 4982 9868 4988 9880
rect 5040 9868 5046 9920
rect 5442 9908 5448 9920
rect 5403 9880 5448 9908
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 7098 9868 7104 9920
rect 7156 9908 7162 9920
rect 11164 9908 11192 10084
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 12713 10047 12771 10053
rect 11296 10016 12434 10044
rect 11296 10004 11302 10016
rect 12406 9976 12434 10016
rect 12713 10013 12725 10047
rect 12759 10013 12771 10047
rect 12894 10044 12900 10056
rect 12855 10016 12900 10044
rect 12713 10007 12771 10013
rect 12728 9976 12756 10007
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10044 13139 10047
rect 13814 10044 13820 10056
rect 13127 10016 13820 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 14568 10044 14596 10084
rect 15488 10084 16436 10112
rect 16577 10115 16635 10121
rect 15488 10044 15516 10084
rect 16577 10081 16589 10115
rect 16623 10112 16635 10115
rect 17310 10112 17316 10124
rect 16623 10084 17316 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 18322 10112 18328 10124
rect 18283 10084 18328 10112
rect 18322 10072 18328 10084
rect 18380 10072 18386 10124
rect 19702 10072 19708 10124
rect 19760 10112 19766 10124
rect 20073 10115 20131 10121
rect 20073 10112 20085 10115
rect 19760 10084 20085 10112
rect 19760 10072 19766 10084
rect 20073 10081 20085 10084
rect 20119 10112 20131 10115
rect 20119 10084 21496 10112
rect 20119 10081 20131 10084
rect 20073 10075 20131 10081
rect 14568 10016 15516 10044
rect 15565 10047 15623 10053
rect 15565 10013 15577 10047
rect 15611 10044 15623 10047
rect 16666 10044 16672 10056
rect 15611 10016 16672 10044
rect 15611 10013 15623 10016
rect 15565 10007 15623 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 12406 9948 12756 9976
rect 15320 9979 15378 9985
rect 15320 9945 15332 9979
rect 15366 9976 15378 9979
rect 15366 9948 15976 9976
rect 15366 9945 15378 9948
rect 15320 9939 15378 9945
rect 7156 9880 11192 9908
rect 7156 9868 7162 9880
rect 11238 9868 11244 9920
rect 11296 9908 11302 9920
rect 11333 9911 11391 9917
rect 11333 9908 11345 9911
rect 11296 9880 11345 9908
rect 11296 9868 11302 9880
rect 11333 9877 11345 9880
rect 11379 9908 11391 9911
rect 11790 9908 11796 9920
rect 11379 9880 11796 9908
rect 11379 9877 11391 9880
rect 11333 9871 11391 9877
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 15948 9917 15976 9948
rect 16022 9936 16028 9988
rect 16080 9976 16086 9988
rect 16776 9976 16804 10007
rect 18138 10004 18144 10056
rect 18196 10044 18202 10056
rect 18233 10047 18291 10053
rect 18233 10044 18245 10047
rect 18196 10016 18245 10044
rect 18196 10004 18202 10016
rect 18233 10013 18245 10016
rect 18279 10013 18291 10047
rect 18877 10047 18935 10053
rect 18877 10044 18889 10047
rect 18233 10007 18291 10013
rect 18616 10016 18889 10044
rect 16080 9948 16804 9976
rect 16080 9936 16086 9948
rect 15933 9911 15991 9917
rect 15933 9877 15945 9911
rect 15979 9877 15991 9911
rect 16298 9908 16304 9920
rect 16259 9880 16304 9908
rect 15933 9871 15991 9877
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 16393 9911 16451 9917
rect 16393 9877 16405 9911
rect 16439 9908 16451 9911
rect 16574 9908 16580 9920
rect 16439 9880 16580 9908
rect 16439 9877 16451 9880
rect 16393 9871 16451 9877
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 18616 9917 18644 10016
rect 18877 10013 18889 10016
rect 18923 10044 18935 10047
rect 19337 10047 19395 10053
rect 19337 10044 19349 10047
rect 18923 10016 19349 10044
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 19337 10013 19349 10016
rect 19383 10013 19395 10047
rect 19794 10044 19800 10056
rect 19755 10016 19800 10044
rect 19337 10007 19395 10013
rect 19794 10004 19800 10016
rect 19852 10004 19858 10056
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 20438 10044 20444 10056
rect 20027 10016 20444 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 19429 9979 19487 9985
rect 19429 9945 19441 9979
rect 19475 9976 19487 9979
rect 19996 9976 20024 10007
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 21358 10044 21364 10056
rect 21319 10016 21364 10044
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 21468 10044 21496 10084
rect 21542 10072 21548 10124
rect 21600 10112 21606 10124
rect 22370 10112 22376 10124
rect 21600 10084 22140 10112
rect 22331 10084 22376 10112
rect 21600 10072 21606 10084
rect 22005 10047 22063 10053
rect 22005 10044 22017 10047
rect 21468 10016 22017 10044
rect 22005 10013 22017 10016
rect 22051 10013 22063 10047
rect 22112 10044 22140 10084
rect 22370 10072 22376 10084
rect 22428 10072 22434 10124
rect 23014 10112 23020 10124
rect 22572 10084 23020 10112
rect 22572 10053 22600 10084
rect 23014 10072 23020 10084
rect 23072 10072 23078 10124
rect 26510 10072 26516 10124
rect 26568 10112 26574 10124
rect 26789 10115 26847 10121
rect 26789 10112 26801 10115
rect 26568 10084 26801 10112
rect 26568 10072 26574 10084
rect 26789 10081 26801 10084
rect 26835 10081 26847 10115
rect 26789 10075 26847 10081
rect 27709 10115 27767 10121
rect 27709 10081 27721 10115
rect 27755 10112 27767 10115
rect 27982 10112 27988 10124
rect 27755 10084 27988 10112
rect 27755 10081 27767 10084
rect 27709 10075 27767 10081
rect 27982 10072 27988 10084
rect 28040 10072 28046 10124
rect 22281 10047 22339 10053
rect 22281 10044 22293 10047
rect 22112 10016 22293 10044
rect 22005 10007 22063 10013
rect 22281 10013 22293 10016
rect 22327 10013 22339 10047
rect 22281 10007 22339 10013
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10013 22615 10047
rect 22738 10044 22744 10056
rect 22699 10016 22744 10044
rect 22557 10007 22615 10013
rect 22738 10004 22744 10016
rect 22796 10004 22802 10056
rect 24486 10004 24492 10056
rect 24544 10044 24550 10056
rect 24673 10047 24731 10053
rect 24673 10044 24685 10047
rect 24544 10016 24685 10044
rect 24544 10004 24550 10016
rect 24673 10013 24685 10016
rect 24719 10013 24731 10047
rect 24854 10044 24860 10056
rect 24815 10016 24860 10044
rect 24673 10007 24731 10013
rect 24854 10004 24860 10016
rect 24912 10004 24918 10056
rect 26694 10044 26700 10056
rect 26655 10016 26700 10044
rect 26694 10004 26700 10016
rect 26752 10004 26758 10056
rect 27893 10047 27951 10053
rect 27893 10013 27905 10047
rect 27939 10013 27951 10047
rect 27893 10007 27951 10013
rect 28077 10047 28135 10053
rect 28077 10013 28089 10047
rect 28123 10044 28135 10047
rect 28261 10047 28319 10053
rect 28261 10044 28273 10047
rect 28123 10016 28273 10044
rect 28123 10013 28135 10016
rect 28077 10007 28135 10013
rect 28261 10013 28273 10016
rect 28307 10013 28319 10047
rect 28261 10007 28319 10013
rect 19475 9948 20024 9976
rect 20165 9979 20223 9985
rect 19475 9945 19487 9948
rect 19429 9939 19487 9945
rect 20165 9945 20177 9979
rect 20211 9945 20223 9979
rect 26970 9976 26976 9988
rect 26931 9948 26976 9976
rect 20165 9939 20223 9945
rect 18601 9911 18659 9917
rect 18601 9877 18613 9911
rect 18647 9877 18659 9911
rect 19058 9908 19064 9920
rect 19019 9880 19064 9908
rect 18601 9871 18659 9877
rect 19058 9868 19064 9880
rect 19116 9868 19122 9920
rect 19610 9868 19616 9920
rect 19668 9908 19674 9920
rect 20180 9908 20208 9939
rect 26970 9936 26976 9948
rect 27028 9936 27034 9988
rect 27614 9936 27620 9988
rect 27672 9976 27678 9988
rect 27908 9976 27936 10007
rect 27672 9948 27936 9976
rect 27672 9936 27678 9948
rect 19668 9880 20208 9908
rect 21545 9911 21603 9917
rect 19668 9868 19674 9880
rect 21545 9877 21557 9911
rect 21591 9908 21603 9911
rect 22278 9908 22284 9920
rect 21591 9880 22284 9908
rect 21591 9877 21603 9880
rect 21545 9871 21603 9877
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 26513 9911 26571 9917
rect 26513 9877 26525 9911
rect 26559 9908 26571 9911
rect 26786 9908 26792 9920
rect 26559 9880 26792 9908
rect 26559 9877 26571 9880
rect 26513 9871 26571 9877
rect 26786 9868 26792 9880
rect 26844 9868 26850 9920
rect 28350 9868 28356 9920
rect 28408 9908 28414 9920
rect 28445 9911 28503 9917
rect 28445 9908 28457 9911
rect 28408 9880 28457 9908
rect 28408 9868 28414 9880
rect 28445 9877 28457 9880
rect 28491 9877 28503 9911
rect 28445 9871 28503 9877
rect 1104 9818 29532 9840
rect 1104 9766 10425 9818
rect 10477 9766 10489 9818
rect 10541 9766 10553 9818
rect 10605 9766 10617 9818
rect 10669 9766 10681 9818
rect 10733 9766 19901 9818
rect 19953 9766 19965 9818
rect 20017 9766 20029 9818
rect 20081 9766 20093 9818
rect 20145 9766 20157 9818
rect 20209 9766 29532 9818
rect 1104 9744 29532 9766
rect 2406 9664 2412 9716
rect 2464 9704 2470 9716
rect 4798 9704 4804 9716
rect 2464 9676 4804 9704
rect 2464 9664 2470 9676
rect 4798 9664 4804 9676
rect 4856 9704 4862 9716
rect 5994 9704 6000 9716
rect 4856 9676 6000 9704
rect 4856 9664 4862 9676
rect 5994 9664 6000 9676
rect 6052 9664 6058 9716
rect 10318 9664 10324 9716
rect 10376 9704 10382 9716
rect 10505 9707 10563 9713
rect 10505 9704 10517 9707
rect 10376 9676 10517 9704
rect 10376 9664 10382 9676
rect 10505 9673 10517 9676
rect 10551 9673 10563 9707
rect 10505 9667 10563 9673
rect 14921 9707 14979 9713
rect 14921 9673 14933 9707
rect 14967 9673 14979 9707
rect 14921 9667 14979 9673
rect 19996 9676 20760 9704
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 6362 9636 6368 9648
rect 1728 9608 6368 9636
rect 1728 9596 1734 9608
rect 2222 9568 2228 9580
rect 2183 9540 2228 9568
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 4724 9577 4752 9608
rect 6362 9596 6368 9608
rect 6420 9596 6426 9648
rect 6733 9639 6791 9645
rect 6733 9605 6745 9639
rect 6779 9636 6791 9639
rect 7926 9636 7932 9648
rect 6779 9608 7932 9636
rect 6779 9605 6791 9608
rect 6733 9599 6791 9605
rect 7926 9596 7932 9608
rect 7984 9596 7990 9648
rect 8938 9596 8944 9648
rect 8996 9636 9002 9648
rect 9582 9636 9588 9648
rect 8996 9608 9588 9636
rect 8996 9596 9002 9608
rect 9582 9596 9588 9608
rect 9640 9636 9646 9648
rect 10689 9639 10747 9645
rect 10689 9636 10701 9639
rect 9640 9608 10701 9636
rect 9640 9596 9646 9608
rect 10689 9605 10701 9608
rect 10735 9605 10747 9639
rect 10689 9599 10747 9605
rect 3697 9571 3755 9577
rect 3697 9568 3709 9571
rect 3476 9540 3709 9568
rect 3476 9528 3482 9540
rect 3697 9537 3709 9540
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 4976 9571 5034 9577
rect 4976 9537 4988 9571
rect 5022 9568 5034 9571
rect 5442 9568 5448 9580
rect 5022 9540 5448 9568
rect 5022 9537 5034 9540
rect 4976 9531 5034 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9568 7251 9571
rect 8110 9568 8116 9580
rect 7239 9540 8116 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 8110 9528 8116 9540
rect 8168 9568 8174 9580
rect 8205 9571 8263 9577
rect 8205 9568 8217 9571
rect 8168 9540 8217 9568
rect 8168 9528 8174 9540
rect 8205 9537 8217 9540
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9537 10379 9571
rect 10704 9568 10732 9599
rect 10778 9596 10784 9648
rect 10836 9636 10842 9648
rect 10873 9639 10931 9645
rect 10873 9636 10885 9639
rect 10836 9608 10885 9636
rect 10836 9596 10842 9608
rect 10873 9605 10885 9608
rect 10919 9605 10931 9639
rect 12621 9639 12679 9645
rect 12621 9636 12633 9639
rect 10873 9599 10931 9605
rect 11992 9608 12633 9636
rect 11992 9580 12020 9608
rect 12621 9605 12633 9608
rect 12667 9605 12679 9639
rect 13906 9636 13912 9648
rect 13867 9608 13912 9636
rect 12621 9599 12679 9605
rect 13906 9596 13912 9608
rect 13964 9636 13970 9648
rect 14461 9639 14519 9645
rect 14461 9636 14473 9639
rect 13964 9608 14473 9636
rect 13964 9596 13970 9608
rect 14461 9605 14473 9608
rect 14507 9605 14519 9639
rect 14461 9599 14519 9605
rect 14550 9596 14556 9648
rect 14608 9636 14614 9648
rect 14645 9639 14703 9645
rect 14645 9636 14657 9639
rect 14608 9608 14657 9636
rect 14608 9596 14614 9608
rect 14645 9605 14657 9608
rect 14691 9636 14703 9639
rect 14936 9636 14964 9667
rect 19996 9648 20024 9676
rect 20732 9648 20760 9676
rect 24854 9664 24860 9716
rect 24912 9704 24918 9716
rect 24912 9676 26372 9704
rect 24912 9664 24918 9676
rect 14691 9608 14964 9636
rect 14691 9605 14703 9608
rect 14645 9599 14703 9605
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 17218 9636 17224 9648
rect 15712 9608 15976 9636
rect 17179 9608 17224 9636
rect 15712 9596 15718 9608
rect 11054 9568 11060 9580
rect 10704 9540 11060 9568
rect 10321 9531 10379 9537
rect 10336 9500 10364 9531
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11195 9540 11713 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 11701 9537 11713 9540
rect 11747 9568 11759 9571
rect 11974 9568 11980 9580
rect 11747 9540 11980 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12066 9528 12072 9580
rect 12124 9568 12130 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 12124 9540 12173 9568
rect 12124 9528 12130 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9537 12495 9571
rect 12710 9568 12716 9580
rect 12671 9540 12716 9568
rect 12437 9531 12495 9537
rect 11517 9503 11575 9509
rect 10336 9472 11376 9500
rect 11348 9444 11376 9472
rect 11517 9469 11529 9503
rect 11563 9469 11575 9503
rect 12452 9500 12480 9531
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 14047 9540 14289 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14918 9528 14924 9580
rect 14976 9568 14982 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14976 9540 15025 9568
rect 14976 9528 14982 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15562 9568 15568 9580
rect 15523 9540 15568 9568
rect 15013 9531 15071 9537
rect 15562 9528 15568 9540
rect 15620 9528 15626 9580
rect 15838 9568 15844 9580
rect 15799 9540 15844 9568
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 13078 9500 13084 9512
rect 12452 9472 13084 9500
rect 11517 9463 11575 9469
rect 1949 9435 2007 9441
rect 1949 9401 1961 9435
rect 1995 9432 2007 9435
rect 2774 9432 2780 9444
rect 1995 9404 2780 9432
rect 1995 9401 2007 9404
rect 1949 9395 2007 9401
rect 2774 9392 2780 9404
rect 2832 9432 2838 9444
rect 3602 9432 3608 9444
rect 2832 9404 3608 9432
rect 2832 9392 2838 9404
rect 3602 9392 3608 9404
rect 3660 9392 3666 9444
rect 6362 9392 6368 9444
rect 6420 9432 6426 9444
rect 6546 9432 6552 9444
rect 6420 9404 6552 9432
rect 6420 9392 6426 9404
rect 6546 9392 6552 9404
rect 6604 9392 6610 9444
rect 7006 9432 7012 9444
rect 6967 9404 7012 9432
rect 7006 9392 7012 9404
rect 7064 9392 7070 9444
rect 11330 9432 11336 9444
rect 11291 9404 11336 9432
rect 11330 9392 11336 9404
rect 11388 9392 11394 9444
rect 1394 9324 1400 9376
rect 1452 9364 1458 9376
rect 1765 9367 1823 9373
rect 1765 9364 1777 9367
rect 1452 9336 1777 9364
rect 1452 9324 1458 9336
rect 1765 9333 1777 9336
rect 1811 9333 1823 9367
rect 3786 9364 3792 9376
rect 3747 9336 3792 9364
rect 1765 9327 1823 9333
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 6086 9364 6092 9376
rect 6047 9336 6092 9364
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 8389 9367 8447 9373
rect 8389 9333 8401 9367
rect 8435 9364 8447 9367
rect 11146 9364 11152 9376
rect 8435 9336 11152 9364
rect 8435 9333 8447 9336
rect 8389 9327 8447 9333
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 11532 9364 11560 9463
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 15470 9500 15476 9512
rect 14200 9472 15476 9500
rect 12161 9435 12219 9441
rect 12161 9401 12173 9435
rect 12207 9432 12219 9435
rect 12250 9432 12256 9444
rect 12207 9404 12256 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 12250 9392 12256 9404
rect 12308 9392 12314 9444
rect 14200 9441 14228 9472
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 15746 9500 15752 9512
rect 15707 9472 15752 9500
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 15948 9509 15976 9608
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 17405 9639 17463 9645
rect 17405 9605 17417 9639
rect 17451 9636 17463 9639
rect 17957 9639 18015 9645
rect 17957 9636 17969 9639
rect 17451 9608 17969 9636
rect 17451 9605 17463 9608
rect 17405 9599 17463 9605
rect 17957 9605 17969 9608
rect 18003 9605 18015 9639
rect 17957 9599 18015 9605
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 16206 9568 16212 9580
rect 16163 9540 16212 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 17126 9568 17132 9580
rect 16540 9540 17132 9568
rect 16540 9528 16546 9540
rect 17126 9528 17132 9540
rect 17184 9568 17190 9580
rect 17420 9568 17448 9599
rect 19150 9596 19156 9648
rect 19208 9636 19214 9648
rect 19245 9639 19303 9645
rect 19245 9636 19257 9639
rect 19208 9608 19257 9636
rect 19208 9596 19214 9608
rect 19245 9605 19257 9608
rect 19291 9605 19303 9639
rect 19794 9636 19800 9648
rect 19755 9608 19800 9636
rect 19245 9599 19303 9605
rect 19794 9596 19800 9608
rect 19852 9596 19858 9648
rect 19978 9596 19984 9648
rect 20036 9596 20042 9648
rect 20254 9596 20260 9648
rect 20312 9636 20318 9648
rect 20312 9608 20668 9636
rect 20312 9596 20318 9608
rect 17184 9540 17448 9568
rect 17681 9571 17739 9577
rect 17184 9528 17190 9540
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 17681 9531 17739 9537
rect 15933 9503 15991 9509
rect 15933 9469 15945 9503
rect 15979 9469 15991 9503
rect 17696 9500 17724 9531
rect 17770 9528 17776 9580
rect 17828 9568 17834 9580
rect 18417 9571 18475 9577
rect 17828 9540 17873 9568
rect 17828 9528 17834 9540
rect 18417 9537 18429 9571
rect 18463 9537 18475 9571
rect 18417 9531 18475 9537
rect 18432 9500 18460 9531
rect 18506 9528 18512 9580
rect 18564 9568 18570 9580
rect 18877 9571 18935 9577
rect 18877 9568 18889 9571
rect 18564 9540 18889 9568
rect 18564 9528 18570 9540
rect 18877 9537 18889 9540
rect 18923 9537 18935 9571
rect 19058 9568 19064 9580
rect 19019 9540 19064 9568
rect 18877 9531 18935 9537
rect 19058 9528 19064 9540
rect 19116 9528 19122 9580
rect 19518 9568 19524 9580
rect 19479 9540 19524 9568
rect 19518 9528 19524 9540
rect 19576 9528 19582 9580
rect 19613 9571 19671 9577
rect 19613 9537 19625 9571
rect 19659 9568 19671 9571
rect 19889 9571 19947 9577
rect 19889 9568 19901 9571
rect 19659 9540 19901 9568
rect 19659 9537 19671 9540
rect 19613 9531 19671 9537
rect 19889 9537 19901 9540
rect 19935 9537 19947 9571
rect 19889 9531 19947 9537
rect 20165 9571 20223 9577
rect 20165 9537 20177 9571
rect 20211 9568 20223 9571
rect 20530 9568 20536 9580
rect 20211 9540 20536 9568
rect 20211 9537 20223 9540
rect 20165 9531 20223 9537
rect 17696 9472 18460 9500
rect 15933 9463 15991 9469
rect 14185 9435 14243 9441
rect 14185 9401 14197 9435
rect 14231 9401 14243 9435
rect 14185 9395 14243 9401
rect 15381 9435 15439 9441
rect 15381 9401 15393 9435
rect 15427 9432 15439 9435
rect 15427 9404 15700 9432
rect 15427 9401 15439 9404
rect 15381 9395 15439 9401
rect 15672 9376 15700 9404
rect 15838 9392 15844 9444
rect 15896 9432 15902 9444
rect 15948 9432 15976 9463
rect 15896 9404 15976 9432
rect 15896 9392 15902 9404
rect 17310 9392 17316 9444
rect 17368 9432 17374 9444
rect 17586 9432 17592 9444
rect 17368 9404 17592 9432
rect 17368 9392 17374 9404
rect 17586 9392 17592 9404
rect 17644 9432 17650 9444
rect 18141 9435 18199 9441
rect 17644 9404 17908 9432
rect 17644 9392 17650 9404
rect 11296 9336 11560 9364
rect 11296 9324 11302 9336
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 11885 9367 11943 9373
rect 11885 9364 11897 9367
rect 11756 9336 11897 9364
rect 11756 9324 11762 9336
rect 11885 9333 11897 9336
rect 11931 9333 11943 9367
rect 11885 9327 11943 9333
rect 14918 9324 14924 9376
rect 14976 9364 14982 9376
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 14976 9336 15577 9364
rect 14976 9324 14982 9336
rect 15565 9333 15577 9336
rect 15611 9333 15623 9367
rect 15565 9327 15623 9333
rect 15654 9324 15660 9376
rect 15712 9324 15718 9376
rect 16114 9324 16120 9376
rect 16172 9364 16178 9376
rect 16301 9367 16359 9373
rect 16301 9364 16313 9367
rect 16172 9336 16313 9364
rect 16172 9324 16178 9336
rect 16301 9333 16313 9336
rect 16347 9333 16359 9367
rect 17402 9364 17408 9376
rect 17363 9336 17408 9364
rect 16301 9327 16359 9333
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 17880 9364 17908 9404
rect 18141 9401 18153 9435
rect 18187 9432 18199 9435
rect 19628 9432 19656 9531
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 20640 9577 20668 9608
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 22278 9636 22284 9648
rect 20772 9608 21128 9636
rect 22239 9608 22284 9636
rect 20772 9596 20778 9608
rect 20625 9571 20683 9577
rect 20625 9537 20637 9571
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 20806 9528 20812 9580
rect 20864 9568 20870 9580
rect 20993 9571 21051 9577
rect 20993 9568 21005 9571
rect 20864 9540 21005 9568
rect 20864 9528 20870 9540
rect 20993 9537 21005 9540
rect 21039 9537 21051 9571
rect 20993 9531 21051 9537
rect 20714 9500 20720 9512
rect 20675 9472 20720 9500
rect 20714 9460 20720 9472
rect 20772 9460 20778 9512
rect 20257 9435 20315 9441
rect 20257 9432 20269 9435
rect 18187 9404 19656 9432
rect 19720 9404 20269 9432
rect 18187 9401 18199 9404
rect 18141 9395 18199 9401
rect 18233 9367 18291 9373
rect 18233 9364 18245 9367
rect 17880 9336 18245 9364
rect 18233 9333 18245 9336
rect 18279 9333 18291 9367
rect 18233 9327 18291 9333
rect 18414 9324 18420 9376
rect 18472 9364 18478 9376
rect 19720 9364 19748 9404
rect 20257 9401 20269 9404
rect 20303 9401 20315 9435
rect 20257 9395 20315 9401
rect 18472 9336 19748 9364
rect 20073 9367 20131 9373
rect 18472 9324 18478 9336
rect 20073 9333 20085 9367
rect 20119 9364 20131 9367
rect 20162 9364 20168 9376
rect 20119 9336 20168 9364
rect 20119 9333 20131 9336
rect 20073 9327 20131 9333
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 21100 9364 21128 9608
rect 22278 9596 22284 9608
rect 22336 9596 22342 9648
rect 26344 9636 26372 9676
rect 27890 9636 27896 9648
rect 25792 9608 26234 9636
rect 26344 9608 27896 9636
rect 21177 9571 21235 9577
rect 21177 9537 21189 9571
rect 21223 9568 21235 9571
rect 22186 9568 22192 9580
rect 21223 9540 21864 9568
rect 22147 9540 22192 9568
rect 21223 9537 21235 9540
rect 21177 9531 21235 9537
rect 21836 9441 21864 9540
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 22554 9528 22560 9580
rect 22612 9568 22618 9580
rect 22741 9571 22799 9577
rect 22741 9568 22753 9571
rect 22612 9540 22753 9568
rect 22612 9528 22618 9540
rect 22741 9537 22753 9540
rect 22787 9537 22799 9571
rect 22741 9531 22799 9537
rect 23106 9528 23112 9580
rect 23164 9568 23170 9580
rect 25792 9577 25820 9608
rect 26206 9580 26234 9608
rect 27890 9596 27896 9608
rect 27948 9596 27954 9648
rect 23477 9571 23535 9577
rect 23477 9568 23489 9571
rect 23164 9540 23489 9568
rect 23164 9528 23170 9540
rect 23477 9537 23489 9540
rect 23523 9537 23535 9571
rect 23477 9531 23535 9537
rect 25777 9571 25835 9577
rect 25777 9537 25789 9571
rect 25823 9537 25835 9571
rect 25958 9568 25964 9580
rect 25919 9540 25964 9568
rect 25777 9531 25835 9537
rect 25958 9528 25964 9540
rect 26016 9528 26022 9580
rect 26206 9540 26240 9580
rect 26234 9528 26240 9540
rect 26292 9568 26298 9580
rect 26510 9568 26516 9580
rect 26292 9540 26337 9568
rect 26471 9540 26516 9568
rect 26292 9528 26298 9540
rect 26510 9528 26516 9540
rect 26568 9528 26574 9580
rect 26605 9571 26663 9577
rect 26605 9537 26617 9571
rect 26651 9537 26663 9571
rect 26605 9531 26663 9537
rect 22002 9460 22008 9512
rect 22060 9500 22066 9512
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 22060 9472 22385 9500
rect 22060 9460 22066 9472
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 25976 9500 26004 9528
rect 22373 9463 22431 9469
rect 22480 9472 26004 9500
rect 21821 9435 21879 9441
rect 21821 9401 21833 9435
rect 21867 9401 21879 9435
rect 21821 9395 21879 9401
rect 21910 9392 21916 9444
rect 21968 9432 21974 9444
rect 22480 9432 22508 9472
rect 26050 9460 26056 9512
rect 26108 9500 26114 9512
rect 26620 9500 26648 9531
rect 26970 9528 26976 9580
rect 27028 9568 27034 9580
rect 27982 9577 27988 9580
rect 27433 9571 27491 9577
rect 27433 9568 27445 9571
rect 27028 9540 27445 9568
rect 27028 9528 27034 9540
rect 27433 9537 27445 9540
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 27976 9531 27988 9577
rect 28040 9568 28046 9580
rect 28040 9540 28076 9568
rect 26108 9472 26648 9500
rect 26108 9460 26114 9472
rect 21968 9404 22508 9432
rect 22925 9435 22983 9441
rect 21968 9392 21974 9404
rect 22925 9401 22937 9435
rect 22971 9432 22983 9435
rect 24854 9432 24860 9444
rect 22971 9404 24860 9432
rect 22971 9401 22983 9404
rect 22925 9395 22983 9401
rect 24854 9392 24860 9404
rect 24912 9392 24918 9444
rect 25685 9435 25743 9441
rect 25685 9401 25697 9435
rect 25731 9432 25743 9435
rect 25774 9432 25780 9444
rect 25731 9404 25780 9432
rect 25731 9401 25743 9404
rect 25685 9395 25743 9401
rect 25774 9392 25780 9404
rect 25832 9392 25838 9444
rect 26697 9435 26755 9441
rect 26697 9401 26709 9435
rect 26743 9432 26755 9435
rect 26970 9432 26976 9444
rect 26743 9404 26976 9432
rect 26743 9401 26755 9404
rect 26697 9395 26755 9401
rect 26970 9392 26976 9404
rect 27028 9392 27034 9444
rect 22738 9364 22744 9376
rect 21100 9336 22744 9364
rect 22738 9324 22744 9336
rect 22796 9364 22802 9376
rect 23017 9367 23075 9373
rect 23017 9364 23029 9367
rect 22796 9336 23029 9364
rect 22796 9324 22802 9336
rect 23017 9333 23029 9336
rect 23063 9333 23075 9367
rect 23017 9327 23075 9333
rect 23661 9367 23719 9373
rect 23661 9333 23673 9367
rect 23707 9364 23719 9367
rect 23750 9364 23756 9376
rect 23707 9336 23756 9364
rect 23707 9333 23719 9336
rect 23661 9327 23719 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 26142 9364 26148 9376
rect 26103 9336 26148 9364
rect 26142 9324 26148 9336
rect 26200 9324 26206 9376
rect 27154 9324 27160 9376
rect 27212 9364 27218 9376
rect 27341 9367 27399 9373
rect 27341 9364 27353 9367
rect 27212 9336 27353 9364
rect 27212 9324 27218 9336
rect 27341 9333 27353 9336
rect 27387 9333 27399 9367
rect 27448 9364 27476 9531
rect 27982 9528 27988 9531
rect 28040 9528 28046 9540
rect 27706 9500 27712 9512
rect 27667 9472 27712 9500
rect 27706 9460 27712 9472
rect 27764 9460 27770 9512
rect 29089 9367 29147 9373
rect 29089 9364 29101 9367
rect 27448 9336 29101 9364
rect 27341 9327 27399 9333
rect 29089 9333 29101 9336
rect 29135 9333 29147 9367
rect 29089 9327 29147 9333
rect 1104 9274 29532 9296
rect 1104 9222 5688 9274
rect 5740 9222 5752 9274
rect 5804 9222 5816 9274
rect 5868 9222 5880 9274
rect 5932 9222 5944 9274
rect 5996 9222 15163 9274
rect 15215 9222 15227 9274
rect 15279 9222 15291 9274
rect 15343 9222 15355 9274
rect 15407 9222 15419 9274
rect 15471 9222 24639 9274
rect 24691 9222 24703 9274
rect 24755 9222 24767 9274
rect 24819 9222 24831 9274
rect 24883 9222 24895 9274
rect 24947 9222 29532 9274
rect 1104 9200 29532 9222
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 3881 9163 3939 9169
rect 3881 9160 3893 9163
rect 3660 9132 3893 9160
rect 3660 9120 3666 9132
rect 3881 9129 3893 9132
rect 3927 9129 3939 9163
rect 3881 9123 3939 9129
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 7616 9132 7757 9160
rect 7616 9120 7622 9132
rect 7745 9129 7757 9132
rect 7791 9129 7803 9163
rect 7745 9123 7803 9129
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 12952 9132 13369 9160
rect 12952 9120 12958 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9160 14243 9163
rect 14918 9160 14924 9172
rect 14231 9132 14924 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 15562 9120 15568 9172
rect 15620 9160 15626 9172
rect 16390 9160 16396 9172
rect 15620 9132 16396 9160
rect 15620 9120 15626 9132
rect 16390 9120 16396 9132
rect 16448 9160 16454 9172
rect 16853 9163 16911 9169
rect 16448 9132 16804 9160
rect 16448 9120 16454 9132
rect 3053 9095 3111 9101
rect 3053 9061 3065 9095
rect 3099 9092 3111 9095
rect 3418 9092 3424 9104
rect 3099 9064 3424 9092
rect 3099 9061 3111 9064
rect 3053 9055 3111 9061
rect 3418 9052 3424 9064
rect 3476 9052 3482 9104
rect 3694 9052 3700 9104
rect 3752 9092 3758 9104
rect 7834 9092 7840 9104
rect 3752 9064 7840 9092
rect 3752 9052 3758 9064
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 16298 9092 16304 9104
rect 16259 9064 16304 9092
rect 16298 9052 16304 9064
rect 16356 9052 16362 9104
rect 1670 9024 1676 9036
rect 1631 8996 1676 9024
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 3786 8984 3792 9036
rect 3844 9024 3850 9036
rect 4019 9027 4077 9033
rect 4019 9024 4031 9027
rect 3844 8996 4031 9024
rect 3844 8984 3850 8996
rect 4019 8993 4031 8996
rect 4065 9024 4077 9027
rect 4525 9027 4583 9033
rect 4525 9024 4537 9027
rect 4065 8996 4537 9024
rect 4065 8993 4077 8996
rect 4019 8987 4077 8993
rect 4525 8993 4537 8996
rect 4571 8993 4583 9027
rect 4525 8987 4583 8993
rect 10318 8984 10324 9036
rect 10376 9024 10382 9036
rect 10781 9027 10839 9033
rect 10781 9024 10793 9027
rect 10376 8996 10793 9024
rect 10376 8984 10382 8996
rect 10781 8993 10793 8996
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 11054 8984 11060 9036
rect 11112 9024 11118 9036
rect 11514 9024 11520 9036
rect 11112 8996 11520 9024
rect 11112 8984 11118 8996
rect 11514 8984 11520 8996
rect 11572 9024 11578 9036
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11572 8996 11989 9024
rect 11572 8984 11578 8996
rect 11977 8993 11989 8996
rect 12023 8993 12035 9027
rect 15565 9027 15623 9033
rect 15565 9024 15577 9027
rect 11977 8987 12035 8993
rect 15488 8996 15577 9024
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 3234 8956 3240 8968
rect 3195 8928 3240 8956
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3418 8956 3424 8968
rect 3379 8928 3424 8956
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8956 7251 8959
rect 7466 8956 7472 8968
rect 7239 8928 7472 8956
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 1946 8897 1952 8900
rect 1940 8851 1952 8897
rect 2004 8888 2010 8900
rect 3602 8888 3608 8900
rect 2004 8860 2040 8888
rect 3563 8860 3608 8888
rect 1946 8848 1952 8851
rect 2004 8848 2010 8860
rect 3602 8848 3608 8860
rect 3660 8848 3666 8900
rect 4172 8888 4200 8919
rect 7466 8916 7472 8928
rect 7524 8956 7530 8968
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7524 8928 7573 8956
rect 7524 8916 7530 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 10597 8959 10655 8965
rect 10597 8925 10609 8959
rect 10643 8956 10655 8959
rect 10870 8956 10876 8968
rect 10643 8928 10876 8956
rect 10643 8925 10655 8928
rect 10597 8919 10655 8925
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 11330 8956 11336 8968
rect 11291 8928 11336 8956
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11606 8956 11612 8968
rect 11567 8928 11612 8956
rect 11425 8919 11483 8925
rect 4430 8888 4436 8900
rect 4172 8860 4436 8888
rect 4430 8848 4436 8860
rect 4488 8888 4494 8900
rect 5074 8888 5080 8900
rect 4488 8860 5080 8888
rect 4488 8848 4494 8860
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 7009 8891 7067 8897
rect 7009 8857 7021 8891
rect 7055 8888 7067 8891
rect 7098 8888 7104 8900
rect 7055 8860 7104 8888
rect 7055 8857 7067 8860
rect 7009 8851 7067 8857
rect 7098 8848 7104 8860
rect 7156 8848 7162 8900
rect 7377 8891 7435 8897
rect 7377 8857 7389 8891
rect 7423 8888 7435 8891
rect 8018 8888 8024 8900
rect 7423 8860 8024 8888
rect 7423 8857 7435 8860
rect 7377 8851 7435 8857
rect 8018 8848 8024 8860
rect 8076 8848 8082 8900
rect 10689 8891 10747 8897
rect 10689 8857 10701 8891
rect 10735 8888 10747 8891
rect 11440 8888 11468 8919
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 12250 8965 12256 8968
rect 12244 8956 12256 8965
rect 11756 8928 11801 8956
rect 12211 8928 12256 8956
rect 11756 8916 11762 8928
rect 12244 8919 12256 8928
rect 12250 8916 12256 8919
rect 12308 8916 12314 8968
rect 15010 8916 15016 8968
rect 15068 8956 15074 8968
rect 15488 8956 15516 8996
rect 15565 8993 15577 8996
rect 15611 9024 15623 9027
rect 16666 9024 16672 9036
rect 15611 8996 16672 9024
rect 15611 8993 15623 8996
rect 15565 8987 15623 8993
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 15654 8956 15660 8968
rect 15068 8928 15516 8956
rect 15615 8928 15660 8956
rect 15068 8916 15074 8928
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 15930 8956 15936 8968
rect 15891 8928 15936 8956
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 16114 8956 16120 8968
rect 16075 8928 16120 8956
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16482 8956 16488 8968
rect 16443 8928 16488 8956
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 16776 8965 16804 9132
rect 16853 9129 16865 9163
rect 16899 9160 16911 9163
rect 17218 9160 17224 9172
rect 16899 9132 17224 9160
rect 16899 9129 16911 9132
rect 16853 9123 16911 9129
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 17862 9160 17868 9172
rect 17368 9132 17868 9160
rect 17368 9120 17374 9132
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 19334 9160 19340 9172
rect 18248 9132 19340 9160
rect 18138 9092 18144 9104
rect 17503 9064 18144 9092
rect 17503 9024 17531 9064
rect 18138 9052 18144 9064
rect 18196 9052 18202 9104
rect 17144 8996 17531 9024
rect 16761 8959 16819 8965
rect 16632 8928 16677 8956
rect 16632 8916 16638 8928
rect 16761 8925 16773 8959
rect 16807 8956 16819 8959
rect 17144 8956 17172 8996
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 17644 8996 17689 9024
rect 17644 8984 17650 8996
rect 18138 8956 18144 8968
rect 16807 8928 17172 8956
rect 18099 8928 18144 8956
rect 16807 8925 16819 8928
rect 16761 8919 16819 8925
rect 18138 8916 18144 8928
rect 18196 8916 18202 8968
rect 18248 8965 18276 9132
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 20073 9163 20131 9169
rect 20073 9160 20085 9163
rect 19576 9132 20085 9160
rect 19576 9120 19582 9132
rect 20073 9129 20085 9132
rect 20119 9129 20131 9163
rect 20714 9160 20720 9172
rect 20675 9132 20720 9160
rect 20073 9123 20131 9129
rect 18325 9095 18383 9101
rect 18325 9061 18337 9095
rect 18371 9061 18383 9095
rect 19245 9095 19303 9101
rect 19245 9092 19257 9095
rect 18325 9055 18383 9061
rect 18892 9064 19257 9092
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 12158 8888 12164 8900
rect 10735 8860 12164 8888
rect 10735 8857 10747 8860
rect 10689 8851 10747 8857
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 15320 8891 15378 8897
rect 15320 8857 15332 8891
rect 15366 8888 15378 8891
rect 17405 8891 17463 8897
rect 15366 8860 17080 8888
rect 15366 8857 15378 8860
rect 15320 8851 15378 8857
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 2222 8820 2228 8832
rect 1627 8792 2228 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 2222 8780 2228 8792
rect 2280 8780 2286 8832
rect 10042 8780 10048 8832
rect 10100 8820 10106 8832
rect 10229 8823 10287 8829
rect 10229 8820 10241 8823
rect 10100 8792 10241 8820
rect 10100 8780 10106 8792
rect 10229 8789 10241 8792
rect 10275 8789 10287 8823
rect 10229 8783 10287 8789
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 17052 8829 17080 8860
rect 17405 8857 17417 8891
rect 17451 8888 17463 8891
rect 18340 8888 18368 9055
rect 18892 9033 18920 9064
rect 19245 9061 19257 9064
rect 19291 9061 19303 9095
rect 20088 9092 20116 9123
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 23106 9160 23112 9172
rect 23067 9132 23112 9160
rect 23106 9120 23112 9132
rect 23164 9120 23170 9172
rect 27614 9160 27620 9172
rect 27575 9132 27620 9160
rect 27614 9120 27620 9132
rect 27672 9120 27678 9172
rect 27893 9163 27951 9169
rect 27893 9129 27905 9163
rect 27939 9160 27951 9163
rect 27982 9160 27988 9172
rect 27939 9132 27988 9160
rect 27939 9129 27951 9132
rect 27893 9123 27951 9129
rect 27982 9120 27988 9132
rect 28040 9120 28046 9172
rect 20625 9095 20683 9101
rect 20625 9092 20637 9095
rect 20088 9064 20637 9092
rect 19245 9055 19303 9061
rect 20625 9061 20637 9064
rect 20671 9061 20683 9095
rect 21542 9092 21548 9104
rect 21503 9064 21548 9092
rect 20625 9055 20683 9061
rect 21542 9052 21548 9064
rect 21600 9052 21606 9104
rect 23382 9092 23388 9104
rect 23124 9064 23388 9092
rect 23124 9036 23152 9064
rect 23382 9052 23388 9064
rect 23440 9092 23446 9104
rect 23440 9064 23888 9092
rect 23440 9052 23446 9064
rect 18877 9027 18935 9033
rect 18877 8993 18889 9027
rect 18923 8993 18935 9027
rect 18877 8987 18935 8993
rect 19610 8984 19616 9036
rect 19668 9024 19674 9036
rect 19889 9027 19947 9033
rect 19889 9024 19901 9027
rect 19668 8996 19901 9024
rect 19668 8984 19674 8996
rect 19889 8993 19901 8996
rect 19935 9024 19947 9027
rect 21361 9027 21419 9033
rect 21361 9024 21373 9027
rect 19935 8996 21373 9024
rect 19935 8993 19947 8996
rect 19889 8987 19947 8993
rect 21361 8993 21373 8996
rect 21407 9024 21419 9027
rect 21910 9024 21916 9036
rect 21407 8996 21916 9024
rect 21407 8993 21419 8996
rect 21361 8987 21419 8993
rect 21910 8984 21916 8996
rect 21968 9024 21974 9036
rect 22097 9027 22155 9033
rect 22097 9024 22109 9027
rect 21968 8996 22109 9024
rect 21968 8984 21974 8996
rect 22097 8993 22109 8996
rect 22143 8993 22155 9027
rect 22738 9024 22744 9036
rect 22699 8996 22744 9024
rect 22097 8987 22155 8993
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 23106 8984 23112 9036
rect 23164 8984 23170 9036
rect 23750 9024 23756 9036
rect 23711 8996 23756 9024
rect 23750 8984 23756 8996
rect 23808 8984 23814 9036
rect 23860 9033 23888 9064
rect 26234 9052 26240 9104
rect 26292 9092 26298 9104
rect 26881 9095 26939 9101
rect 26881 9092 26893 9095
rect 26292 9064 26893 9092
rect 26292 9052 26298 9064
rect 26881 9061 26893 9064
rect 26927 9061 26939 9095
rect 26881 9055 26939 9061
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 8993 23903 9027
rect 27706 9024 27712 9036
rect 23845 8987 23903 8993
rect 25884 8996 27712 9024
rect 18598 8956 18604 8968
rect 18559 8928 18604 8956
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 19058 8956 19064 8968
rect 18971 8928 19064 8956
rect 19058 8916 19064 8928
rect 19116 8916 19122 8968
rect 20625 8959 20683 8965
rect 20625 8925 20637 8959
rect 20671 8956 20683 8959
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 20671 8928 22017 8956
rect 20671 8925 20683 8928
rect 20625 8919 20683 8925
rect 22005 8925 22017 8928
rect 22051 8956 22063 8959
rect 22370 8956 22376 8968
rect 22051 8928 22376 8956
rect 22051 8925 22063 8928
rect 22005 8919 22063 8925
rect 22370 8916 22376 8928
rect 22428 8916 22434 8968
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8956 22983 8959
rect 22971 8928 23704 8956
rect 22971 8925 22983 8928
rect 22925 8919 22983 8925
rect 17451 8860 18368 8888
rect 19076 8888 19104 8916
rect 20714 8888 20720 8900
rect 19076 8860 20720 8888
rect 17451 8857 17463 8860
rect 17405 8851 17463 8857
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 21177 8891 21235 8897
rect 21177 8888 21189 8891
rect 20824 8860 21189 8888
rect 11149 8823 11207 8829
rect 11149 8820 11161 8823
rect 10928 8792 11161 8820
rect 10928 8780 10934 8792
rect 11149 8789 11161 8792
rect 11195 8789 11207 8823
rect 11149 8783 11207 8789
rect 17037 8823 17095 8829
rect 17037 8789 17049 8823
rect 17083 8789 17095 8823
rect 17037 8783 17095 8789
rect 17218 8780 17224 8832
rect 17276 8820 17282 8832
rect 17494 8820 17500 8832
rect 17276 8792 17500 8820
rect 17276 8780 17282 8792
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 19242 8780 19248 8832
rect 19300 8820 19306 8832
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 19300 8792 19625 8820
rect 19300 8780 19306 8792
rect 19613 8789 19625 8792
rect 19659 8789 19671 8823
rect 19613 8783 19671 8789
rect 19702 8780 19708 8832
rect 19760 8820 19766 8832
rect 20824 8820 20852 8860
rect 21177 8857 21189 8860
rect 21223 8888 21235 8891
rect 21818 8888 21824 8900
rect 21223 8860 21824 8888
rect 21223 8857 21235 8860
rect 21177 8851 21235 8857
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 22186 8888 22192 8900
rect 22066 8860 22192 8888
rect 21082 8820 21088 8832
rect 19760 8792 20852 8820
rect 21043 8792 21088 8820
rect 19760 8780 19766 8792
rect 21082 8780 21088 8792
rect 21140 8820 21146 8832
rect 21913 8823 21971 8829
rect 21913 8820 21925 8823
rect 21140 8792 21925 8820
rect 21140 8780 21146 8792
rect 21913 8789 21925 8792
rect 21959 8820 21971 8823
rect 22066 8820 22094 8860
rect 22186 8848 22192 8860
rect 22244 8848 22250 8900
rect 23676 8832 23704 8928
rect 22554 8820 22560 8832
rect 21959 8792 22094 8820
rect 22515 8792 22560 8820
rect 21959 8789 21971 8792
rect 21913 8783 21971 8789
rect 22554 8780 22560 8792
rect 22612 8780 22618 8832
rect 23293 8823 23351 8829
rect 23293 8789 23305 8823
rect 23339 8820 23351 8823
rect 23382 8820 23388 8832
rect 23339 8792 23388 8820
rect 23339 8789 23351 8792
rect 23293 8783 23351 8789
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 23658 8820 23664 8832
rect 23619 8792 23664 8820
rect 23658 8780 23664 8792
rect 23716 8780 23722 8832
rect 23860 8820 23888 8987
rect 24857 8959 24915 8965
rect 24857 8925 24869 8959
rect 24903 8956 24915 8959
rect 24946 8956 24952 8968
rect 24903 8928 24952 8956
rect 24903 8925 24915 8928
rect 24857 8919 24915 8925
rect 24946 8916 24952 8928
rect 25004 8956 25010 8968
rect 25884 8956 25912 8996
rect 27706 8984 27712 8996
rect 27764 8984 27770 9036
rect 28350 9024 28356 9036
rect 28311 8996 28356 9024
rect 28350 8984 28356 8996
rect 28408 8984 28414 9036
rect 28442 8984 28448 9036
rect 28500 9024 28506 9036
rect 28500 8996 28545 9024
rect 28500 8984 28506 8996
rect 25004 8928 25912 8956
rect 25004 8916 25010 8928
rect 26050 8916 26056 8968
rect 26108 8956 26114 8968
rect 26421 8959 26479 8965
rect 26421 8956 26433 8959
rect 26108 8928 26433 8956
rect 26108 8916 26114 8928
rect 26421 8925 26433 8928
rect 26467 8925 26479 8959
rect 26421 8919 26479 8925
rect 26510 8916 26516 8968
rect 26568 8956 26574 8968
rect 26605 8959 26663 8965
rect 26605 8956 26617 8959
rect 26568 8928 26617 8956
rect 26568 8916 26574 8928
rect 26605 8925 26617 8928
rect 26651 8925 26663 8959
rect 26970 8956 26976 8968
rect 26931 8928 26976 8956
rect 26605 8919 26663 8925
rect 26970 8916 26976 8928
rect 27028 8916 27034 8968
rect 27154 8956 27160 8968
rect 27115 8928 27160 8956
rect 27154 8916 27160 8928
rect 27212 8916 27218 8968
rect 27341 8959 27399 8965
rect 27341 8925 27353 8959
rect 27387 8925 27399 8959
rect 27341 8919 27399 8925
rect 25124 8891 25182 8897
rect 25124 8857 25136 8891
rect 25170 8888 25182 8891
rect 25314 8888 25320 8900
rect 25170 8860 25320 8888
rect 25170 8857 25182 8860
rect 25124 8851 25182 8857
rect 25314 8848 25320 8860
rect 25372 8848 25378 8900
rect 25866 8820 25872 8832
rect 23860 8792 25872 8820
rect 25866 8780 25872 8792
rect 25924 8780 25930 8832
rect 26237 8823 26295 8829
rect 26237 8789 26249 8823
rect 26283 8820 26295 8823
rect 26528 8820 26556 8916
rect 26988 8888 27016 8916
rect 27356 8888 27384 8919
rect 27614 8916 27620 8968
rect 27672 8956 27678 8968
rect 28261 8959 28319 8965
rect 28261 8956 28273 8959
rect 27672 8928 28273 8956
rect 27672 8916 27678 8928
rect 28261 8925 28273 8928
rect 28307 8925 28319 8959
rect 28261 8919 28319 8925
rect 26988 8860 27384 8888
rect 27709 8891 27767 8897
rect 27709 8857 27721 8891
rect 27755 8857 27767 8891
rect 27709 8851 27767 8857
rect 26283 8792 26556 8820
rect 26283 8789 26295 8792
rect 26237 8783 26295 8789
rect 27614 8780 27620 8832
rect 27672 8820 27678 8832
rect 27724 8820 27752 8851
rect 27672 8792 27752 8820
rect 27672 8780 27678 8792
rect 1104 8730 29532 8752
rect 1104 8678 10425 8730
rect 10477 8678 10489 8730
rect 10541 8678 10553 8730
rect 10605 8678 10617 8730
rect 10669 8678 10681 8730
rect 10733 8678 19901 8730
rect 19953 8678 19965 8730
rect 20017 8678 20029 8730
rect 20081 8678 20093 8730
rect 20145 8678 20157 8730
rect 20209 8678 29532 8730
rect 1104 8656 29532 8678
rect 1857 8619 1915 8625
rect 1857 8585 1869 8619
rect 1903 8616 1915 8619
rect 1946 8616 1952 8628
rect 1903 8588 1952 8616
rect 1903 8585 1915 8588
rect 1857 8579 1915 8585
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 2222 8616 2228 8628
rect 2183 8588 2228 8616
rect 2222 8576 2228 8588
rect 2280 8576 2286 8628
rect 2317 8619 2375 8625
rect 2317 8585 2329 8619
rect 2363 8616 2375 8619
rect 2774 8616 2780 8628
rect 2363 8588 2780 8616
rect 2363 8585 2375 8588
rect 2317 8579 2375 8585
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 5316 8588 6224 8616
rect 5316 8576 5322 8588
rect 3418 8508 3424 8560
rect 3476 8548 3482 8560
rect 4065 8551 4123 8557
rect 3476 8520 3556 8548
rect 3476 8508 3482 8520
rect 3528 8489 3556 8520
rect 4065 8517 4077 8551
rect 4111 8548 4123 8551
rect 4246 8548 4252 8560
rect 4111 8520 4252 8548
rect 4111 8517 4123 8520
rect 4065 8511 4123 8517
rect 4246 8508 4252 8520
rect 4304 8508 4310 8560
rect 5353 8551 5411 8557
rect 5353 8517 5365 8551
rect 5399 8548 5411 8551
rect 5534 8548 5540 8560
rect 5399 8520 5540 8548
rect 5399 8517 5411 8520
rect 5353 8511 5411 8517
rect 5534 8508 5540 8520
rect 5592 8548 5598 8560
rect 5997 8551 6055 8557
rect 5997 8548 6009 8551
rect 5592 8520 6009 8548
rect 5592 8508 5598 8520
rect 5997 8517 6009 8520
rect 6043 8548 6055 8551
rect 6086 8548 6092 8560
rect 6043 8520 6092 8548
rect 6043 8517 6055 8520
rect 5997 8511 6055 8517
rect 6086 8508 6092 8520
rect 6144 8508 6150 8560
rect 6196 8557 6224 8588
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 9640 8588 9812 8616
rect 9640 8576 9646 8588
rect 6181 8551 6239 8557
rect 6181 8517 6193 8551
rect 6227 8517 6239 8551
rect 6546 8548 6552 8560
rect 6181 8511 6239 8517
rect 6380 8520 6552 8548
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 3823 8483 3881 8489
rect 3823 8480 3835 8483
rect 3660 8452 3835 8480
rect 3660 8440 3666 8452
rect 3823 8449 3835 8452
rect 3869 8480 3881 8483
rect 4154 8480 4160 8492
rect 3869 8452 4016 8480
rect 4115 8452 4160 8480
rect 3869 8449 3881 8452
rect 3823 8443 3881 8449
rect 2406 8412 2412 8424
rect 2367 8384 2412 8412
rect 2406 8372 2412 8384
rect 2464 8372 2470 8424
rect 3234 8372 3240 8424
rect 3292 8412 3298 8424
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 3292 8384 3433 8412
rect 3292 8372 3298 8384
rect 3421 8381 3433 8384
rect 3467 8381 3479 8415
rect 3988 8412 4016 8452
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 4430 8489 4436 8492
rect 4399 8483 4436 8489
rect 4399 8449 4411 8483
rect 4399 8443 4436 8449
rect 4430 8440 4436 8443
rect 4488 8440 4494 8492
rect 6380 8489 6408 8520
rect 6546 8508 6552 8520
rect 6604 8548 6610 8560
rect 8294 8548 8300 8560
rect 6604 8520 8300 8548
rect 6604 8508 6610 8520
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 9340 8551 9398 8557
rect 9340 8517 9352 8551
rect 9386 8548 9398 8551
rect 9677 8551 9735 8557
rect 9677 8548 9689 8551
rect 9386 8520 9689 8548
rect 9386 8517 9398 8520
rect 9340 8511 9398 8517
rect 9677 8517 9689 8520
rect 9723 8517 9735 8551
rect 9677 8511 9735 8517
rect 6638 8489 6644 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 4632 8452 5825 8480
rect 4632 8412 4660 8452
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6632 8443 6644 8489
rect 6696 8480 6702 8492
rect 9596 8483 9654 8489
rect 6696 8452 6732 8480
rect 8220 8452 9536 8480
rect 3988 8384 4660 8412
rect 4689 8415 4747 8421
rect 3421 8375 3479 8381
rect 4689 8381 4701 8415
rect 4735 8412 4747 8415
rect 4801 8415 4859 8421
rect 4735 8381 4752 8412
rect 4689 8375 4752 8381
rect 4801 8381 4813 8415
rect 4847 8412 4859 8415
rect 5258 8412 5264 8424
rect 4847 8384 5264 8412
rect 4847 8381 4859 8384
rect 4801 8375 4859 8381
rect 4724 8344 4752 8375
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 5442 8412 5448 8424
rect 5403 8384 5448 8412
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8381 5687 8415
rect 5828 8412 5856 8443
rect 6638 8440 6644 8443
rect 6696 8440 6702 8452
rect 6086 8412 6092 8424
rect 5828 8384 6092 8412
rect 5629 8375 5687 8381
rect 4890 8344 4896 8356
rect 4724 8316 4896 8344
rect 4890 8304 4896 8316
rect 4948 8304 4954 8356
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 4985 8279 5043 8285
rect 4985 8276 4997 8279
rect 4672 8248 4997 8276
rect 4672 8236 4678 8248
rect 4985 8245 4997 8248
rect 5031 8245 5043 8279
rect 4985 8239 5043 8245
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5644 8276 5672 8375
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 7834 8304 7840 8356
rect 7892 8344 7898 8356
rect 8220 8353 8248 8452
rect 9508 8412 9536 8452
rect 9596 8449 9608 8483
rect 9642 8480 9654 8483
rect 9784 8480 9812 8588
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11112 8588 11805 8616
rect 11112 8576 11118 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 12066 8616 12072 8628
rect 12027 8588 12072 8616
rect 11793 8579 11851 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 15841 8619 15899 8625
rect 15841 8616 15853 8619
rect 15804 8588 15853 8616
rect 15804 8576 15810 8588
rect 15841 8585 15853 8588
rect 15887 8585 15899 8619
rect 16206 8616 16212 8628
rect 16167 8588 16212 8616
rect 15841 8579 15899 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 17770 8616 17776 8628
rect 16868 8588 17776 8616
rect 10042 8508 10048 8560
rect 10100 8548 10106 8560
rect 11609 8551 11667 8557
rect 11609 8548 11621 8551
rect 10100 8520 10640 8548
rect 10100 8508 10106 8520
rect 9642 8452 9812 8480
rect 9861 8483 9919 8489
rect 9642 8449 9654 8452
rect 9596 8443 9654 8449
rect 9861 8449 9873 8483
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 9876 8412 9904 8443
rect 9950 8440 9956 8492
rect 10008 8480 10014 8492
rect 10230 8483 10288 8489
rect 10230 8480 10242 8483
rect 10008 8452 10242 8480
rect 10008 8440 10014 8452
rect 10230 8449 10242 8452
rect 10276 8449 10288 8483
rect 10230 8443 10288 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 10505 8483 10563 8489
rect 10505 8480 10517 8483
rect 10459 8452 10517 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 10505 8449 10517 8452
rect 10551 8449 10563 8483
rect 10612 8480 10640 8520
rect 10796 8520 11621 8548
rect 10796 8489 10824 8520
rect 11609 8517 11621 8520
rect 11655 8517 11667 8551
rect 11609 8511 11667 8517
rect 11698 8508 11704 8560
rect 11756 8548 11762 8560
rect 11756 8520 12388 8548
rect 11756 8508 11762 8520
rect 10670 8483 10728 8489
rect 10670 8480 10682 8483
rect 10612 8452 10682 8480
rect 10505 8443 10563 8449
rect 10670 8449 10682 8452
rect 10716 8449 10728 8483
rect 10670 8443 10728 8449
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10042 8412 10048 8424
rect 9508 8384 9904 8412
rect 10003 8384 10048 8412
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10137 8415 10195 8421
rect 10137 8381 10149 8415
rect 10183 8412 10195 8415
rect 10318 8412 10324 8424
rect 10183 8384 10324 8412
rect 10183 8381 10195 8384
rect 10137 8375 10195 8381
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 8205 8347 8263 8353
rect 8205 8344 8217 8347
rect 7892 8316 8217 8344
rect 7892 8304 7898 8316
rect 8205 8313 8217 8316
rect 8251 8313 8263 8347
rect 8205 8307 8263 8313
rect 9766 8304 9772 8356
rect 9824 8344 9830 8356
rect 10428 8344 10456 8443
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 10928 8452 10973 8480
rect 10928 8440 10934 8452
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11517 8483 11575 8489
rect 11112 8452 11157 8480
rect 11112 8440 11118 8452
rect 11517 8449 11529 8483
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 10888 8412 10916 8440
rect 11532 8412 11560 8443
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 12360 8489 12388 8520
rect 15930 8508 15936 8560
rect 15988 8548 15994 8560
rect 16868 8548 16896 8588
rect 17494 8548 17500 8560
rect 15988 8520 16896 8548
rect 17455 8520 17500 8548
rect 15988 8508 15994 8520
rect 12253 8483 12311 8489
rect 12253 8480 12265 8483
rect 12216 8452 12265 8480
rect 12216 8440 12222 8452
rect 12253 8449 12265 8452
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8449 12403 8483
rect 12710 8480 12716 8492
rect 12345 8443 12403 8449
rect 12544 8452 12716 8480
rect 10888 8384 11560 8412
rect 9824 8316 10456 8344
rect 11241 8347 11299 8353
rect 9824 8304 9830 8316
rect 11241 8313 11253 8347
rect 11287 8344 11299 8347
rect 11330 8344 11336 8356
rect 11287 8316 11336 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 12268 8344 12296 8443
rect 12544 8421 12572 8452
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12894 8480 12900 8492
rect 12855 8452 12900 8480
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 17126 8466 17132 8518
rect 17184 8506 17190 8518
rect 17494 8508 17500 8520
rect 17552 8508 17558 8560
rect 17696 8557 17724 8588
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 19061 8619 19119 8625
rect 19061 8616 19073 8619
rect 18196 8588 19073 8616
rect 18196 8576 18202 8588
rect 19061 8585 19073 8588
rect 19107 8585 19119 8619
rect 19061 8579 19119 8585
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 20346 8616 20352 8628
rect 19392 8588 20352 8616
rect 19392 8576 19398 8588
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 20530 8616 20536 8628
rect 20491 8588 20536 8616
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 22370 8616 22376 8628
rect 20640 8588 22376 8616
rect 17681 8551 17739 8557
rect 17681 8517 17693 8551
rect 17727 8517 17739 8551
rect 17681 8511 17739 8517
rect 19521 8551 19579 8557
rect 19521 8517 19533 8551
rect 19567 8548 19579 8551
rect 19981 8551 20039 8557
rect 19981 8548 19993 8551
rect 19567 8520 19993 8548
rect 19567 8517 19579 8520
rect 19521 8511 19579 8517
rect 19981 8517 19993 8520
rect 20027 8548 20039 8551
rect 20640 8548 20668 8588
rect 22370 8576 22376 8588
rect 22428 8616 22434 8628
rect 23017 8619 23075 8625
rect 23017 8616 23029 8619
rect 22428 8588 23029 8616
rect 22428 8576 22434 8588
rect 23017 8585 23029 8588
rect 23063 8616 23075 8619
rect 23201 8619 23259 8625
rect 23201 8616 23213 8619
rect 23063 8588 23213 8616
rect 23063 8585 23075 8588
rect 23017 8579 23075 8585
rect 23201 8585 23213 8588
rect 23247 8616 23259 8619
rect 25314 8616 25320 8628
rect 23247 8588 25084 8616
rect 25275 8588 25320 8616
rect 23247 8585 23259 8588
rect 23201 8579 23259 8585
rect 24946 8548 24952 8560
rect 20027 8520 20668 8548
rect 20732 8520 21680 8548
rect 20027 8517 20039 8520
rect 19981 8511 20039 8517
rect 17184 8489 17264 8506
rect 17184 8483 17279 8489
rect 17184 8478 17233 8483
rect 17184 8466 17190 8478
rect 17221 8449 17233 8478
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 12529 8415 12587 8421
rect 12529 8381 12541 8415
rect 12575 8381 12587 8415
rect 12529 8375 12587 8381
rect 12621 8415 12679 8421
rect 12621 8381 12633 8415
rect 12667 8412 12679 8415
rect 12912 8412 12940 8440
rect 12667 8384 12940 8412
rect 15657 8415 15715 8421
rect 12667 8381 12679 8384
rect 12621 8375 12679 8381
rect 15657 8381 15669 8415
rect 15703 8381 15715 8415
rect 15657 8375 15715 8381
rect 12805 8347 12863 8353
rect 12805 8344 12817 8347
rect 12268 8316 12817 8344
rect 12805 8313 12817 8316
rect 12851 8313 12863 8347
rect 15672 8344 15700 8375
rect 15746 8372 15752 8424
rect 15804 8412 15810 8424
rect 15804 8384 15849 8412
rect 15804 8372 15810 8384
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 17129 8415 17187 8421
rect 16448 8384 16988 8412
rect 16448 8372 16454 8384
rect 16022 8344 16028 8356
rect 15672 8316 16028 8344
rect 12805 8307 12863 8313
rect 16022 8304 16028 8316
rect 16080 8344 16086 8356
rect 16080 8316 16436 8344
rect 16080 8304 16086 8316
rect 6730 8276 6736 8288
rect 5132 8248 6736 8276
rect 5132 8236 5138 8248
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 7742 8276 7748 8288
rect 7703 8248 7748 8276
rect 7742 8236 7748 8248
rect 7800 8236 7806 8288
rect 16408 8276 16436 8316
rect 16482 8304 16488 8356
rect 16540 8344 16546 8356
rect 16960 8344 16988 8384
rect 17129 8381 17141 8415
rect 17175 8381 17187 8415
rect 17129 8375 17187 8381
rect 17144 8344 17172 8375
rect 16540 8316 16896 8344
rect 16960 8316 17172 8344
rect 16540 8304 16546 8316
rect 16758 8276 16764 8288
rect 16408 8248 16764 8276
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 16868 8285 16896 8316
rect 16853 8279 16911 8285
rect 16853 8245 16865 8279
rect 16899 8276 16911 8279
rect 17126 8276 17132 8288
rect 16899 8248 17132 8276
rect 16899 8245 16911 8248
rect 16853 8239 16911 8245
rect 17126 8236 17132 8248
rect 17184 8236 17190 8288
rect 17221 8279 17279 8285
rect 17221 8245 17233 8279
rect 17267 8276 17279 8279
rect 17328 8276 17356 8443
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 19242 8480 19248 8492
rect 18288 8452 19248 8480
rect 18288 8440 18294 8452
rect 19242 8440 19248 8452
rect 19300 8480 19306 8492
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 19300 8452 19441 8480
rect 19300 8440 19306 8452
rect 19429 8449 19441 8452
rect 19475 8449 19487 8483
rect 19702 8480 19708 8492
rect 19429 8443 19487 8449
rect 19536 8452 19708 8480
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 19536 8412 19564 8452
rect 19702 8440 19708 8452
rect 19760 8440 19766 8492
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8480 20223 8483
rect 20254 8480 20260 8492
rect 20211 8452 20260 8480
rect 20211 8449 20223 8452
rect 20165 8443 20223 8449
rect 20254 8440 20260 8452
rect 20312 8440 20318 8492
rect 20732 8489 20760 8520
rect 20717 8483 20775 8489
rect 20717 8449 20729 8483
rect 20763 8449 20775 8483
rect 20717 8443 20775 8449
rect 20806 8440 20812 8492
rect 20864 8480 20870 8492
rect 21085 8483 21143 8489
rect 20864 8452 20909 8480
rect 20864 8440 20870 8452
rect 21085 8449 21097 8483
rect 21131 8480 21143 8483
rect 21542 8480 21548 8492
rect 21131 8452 21548 8480
rect 21131 8449 21143 8452
rect 21085 8443 21143 8449
rect 21542 8440 21548 8452
rect 21600 8440 21606 8492
rect 21652 8489 21680 8520
rect 23308 8520 24952 8548
rect 21637 8483 21695 8489
rect 21637 8449 21649 8483
rect 21683 8480 21695 8483
rect 22373 8483 22431 8489
rect 22373 8480 22385 8483
rect 21683 8452 22385 8480
rect 21683 8449 21695 8452
rect 21637 8443 21695 8449
rect 22373 8449 22385 8452
rect 22419 8480 22431 8483
rect 22554 8480 22560 8492
rect 22419 8452 22560 8480
rect 22419 8449 22431 8452
rect 22373 8443 22431 8449
rect 22554 8440 22560 8452
rect 22612 8440 22618 8492
rect 22649 8483 22707 8489
rect 22649 8449 22661 8483
rect 22695 8449 22707 8483
rect 22649 8443 22707 8449
rect 17828 8384 19564 8412
rect 17828 8372 17834 8384
rect 19610 8372 19616 8424
rect 19668 8412 19674 8424
rect 20824 8412 20852 8440
rect 22664 8412 22692 8443
rect 22922 8440 22928 8492
rect 22980 8480 22986 8492
rect 23308 8489 23336 8520
rect 24946 8508 24952 8520
rect 25004 8508 25010 8560
rect 25056 8548 25084 8588
rect 25314 8576 25320 8588
rect 25372 8576 25378 8628
rect 25685 8619 25743 8625
rect 25685 8585 25697 8619
rect 25731 8616 25743 8619
rect 26142 8616 26148 8628
rect 25731 8588 26148 8616
rect 25731 8585 25743 8588
rect 25685 8579 25743 8585
rect 26142 8576 26148 8588
rect 26200 8576 26206 8628
rect 25774 8548 25780 8560
rect 25056 8520 25360 8548
rect 25735 8520 25780 8548
rect 23293 8483 23351 8489
rect 23293 8480 23305 8483
rect 22980 8452 23305 8480
rect 22980 8440 22986 8452
rect 23293 8449 23305 8452
rect 23339 8449 23351 8483
rect 23293 8443 23351 8449
rect 23382 8440 23388 8492
rect 23440 8480 23446 8492
rect 23549 8483 23607 8489
rect 23549 8480 23561 8483
rect 23440 8452 23561 8480
rect 23440 8440 23446 8452
rect 23549 8449 23561 8452
rect 23595 8449 23607 8483
rect 23549 8443 23607 8449
rect 19668 8384 19713 8412
rect 20824 8384 22692 8412
rect 19668 8372 19674 8384
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 20993 8347 21051 8353
rect 20993 8344 21005 8347
rect 18656 8316 21005 8344
rect 18656 8304 18662 8316
rect 20993 8313 21005 8316
rect 21039 8313 21051 8347
rect 20993 8307 21051 8313
rect 22741 8347 22799 8353
rect 22741 8313 22753 8347
rect 22787 8344 22799 8347
rect 23106 8344 23112 8356
rect 22787 8316 23112 8344
rect 22787 8313 22799 8316
rect 22741 8307 22799 8313
rect 23106 8304 23112 8316
rect 23164 8304 23170 8356
rect 24673 8347 24731 8353
rect 24673 8313 24685 8347
rect 24719 8344 24731 8347
rect 25222 8344 25228 8356
rect 24719 8316 25228 8344
rect 24719 8313 24731 8316
rect 24673 8307 24731 8313
rect 25222 8304 25228 8316
rect 25280 8304 25286 8356
rect 25332 8344 25360 8520
rect 25774 8508 25780 8520
rect 25832 8508 25838 8560
rect 27890 8480 27896 8492
rect 27851 8452 27896 8480
rect 27890 8440 27896 8452
rect 27948 8440 27954 8492
rect 28074 8480 28080 8492
rect 28035 8452 28080 8480
rect 28074 8440 28080 8452
rect 28132 8440 28138 8492
rect 28261 8483 28319 8489
rect 28261 8449 28273 8483
rect 28307 8480 28319 8483
rect 28629 8483 28687 8489
rect 28629 8480 28641 8483
rect 28307 8452 28641 8480
rect 28307 8449 28319 8452
rect 28261 8443 28319 8449
rect 28629 8449 28641 8452
rect 28675 8449 28687 8483
rect 28629 8443 28687 8449
rect 25866 8412 25872 8424
rect 25827 8384 25872 8412
rect 25866 8372 25872 8384
rect 25924 8412 25930 8424
rect 28534 8412 28540 8424
rect 25924 8384 28540 8412
rect 25924 8372 25930 8384
rect 28534 8372 28540 8384
rect 28592 8372 28598 8424
rect 28997 8415 29055 8421
rect 28997 8381 29009 8415
rect 29043 8381 29055 8415
rect 28997 8375 29055 8381
rect 26510 8344 26516 8356
rect 25332 8316 26516 8344
rect 26510 8304 26516 8316
rect 26568 8304 26574 8356
rect 18046 8276 18052 8288
rect 17267 8248 18052 8276
rect 17267 8245 17279 8248
rect 17221 8239 17279 8245
rect 18046 8236 18052 8248
rect 18104 8276 18110 8288
rect 21082 8276 21088 8288
rect 18104 8248 21088 8276
rect 18104 8236 18110 8248
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 21266 8236 21272 8288
rect 21324 8276 21330 8288
rect 21545 8279 21603 8285
rect 21545 8276 21557 8279
rect 21324 8248 21557 8276
rect 21324 8236 21330 8248
rect 21545 8245 21557 8248
rect 21591 8245 21603 8279
rect 21545 8239 21603 8245
rect 22557 8279 22615 8285
rect 22557 8245 22569 8279
rect 22603 8276 22615 8279
rect 22830 8276 22836 8288
rect 22603 8248 22836 8276
rect 22603 8245 22615 8248
rect 22557 8239 22615 8245
rect 22830 8236 22836 8248
rect 22888 8236 22894 8288
rect 28442 8276 28448 8288
rect 28403 8248 28448 8276
rect 28442 8236 28448 8248
rect 28500 8236 28506 8288
rect 29012 8276 29040 8375
rect 29086 8276 29092 8288
rect 29012 8248 29092 8276
rect 29086 8236 29092 8248
rect 29144 8236 29150 8288
rect 1104 8186 29532 8208
rect 1104 8134 5688 8186
rect 5740 8134 5752 8186
rect 5804 8134 5816 8186
rect 5868 8134 5880 8186
rect 5932 8134 5944 8186
rect 5996 8134 15163 8186
rect 15215 8134 15227 8186
rect 15279 8134 15291 8186
rect 15343 8134 15355 8186
rect 15407 8134 15419 8186
rect 15471 8134 24639 8186
rect 24691 8134 24703 8186
rect 24755 8134 24767 8186
rect 24819 8134 24831 8186
rect 24883 8134 24895 8186
rect 24947 8134 29532 8186
rect 1104 8112 29532 8134
rect 2774 8072 2780 8084
rect 2608 8044 2780 8072
rect 2608 8013 2636 8044
rect 2774 8032 2780 8044
rect 2832 8072 2838 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 2832 8044 3801 8072
rect 2832 8032 2838 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 4157 8075 4215 8081
rect 4157 8041 4169 8075
rect 4203 8072 4215 8075
rect 4338 8072 4344 8084
rect 4203 8044 4344 8072
rect 4203 8041 4215 8044
rect 4157 8035 4215 8041
rect 4338 8032 4344 8044
rect 4396 8032 4402 8084
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 5442 8072 5448 8084
rect 5123 8044 5448 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 6638 8032 6644 8084
rect 6696 8072 6702 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6696 8044 6745 8072
rect 6696 8032 6702 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 6733 8035 6791 8041
rect 9401 8075 9459 8081
rect 9401 8041 9413 8075
rect 9447 8072 9459 8075
rect 9950 8072 9956 8084
rect 9447 8044 9956 8072
rect 9447 8041 9459 8044
rect 9401 8035 9459 8041
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 17586 8072 17592 8084
rect 17547 8044 17592 8072
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 21818 8072 21824 8084
rect 21779 8044 21824 8072
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 22830 8032 22836 8084
rect 22888 8072 22894 8084
rect 22925 8075 22983 8081
rect 22925 8072 22937 8075
rect 22888 8044 22937 8072
rect 22888 8032 22894 8044
rect 22925 8041 22937 8044
rect 22971 8041 22983 8075
rect 22925 8035 22983 8041
rect 23658 8032 23664 8084
rect 23716 8072 23722 8084
rect 23937 8075 23995 8081
rect 23937 8072 23949 8075
rect 23716 8044 23949 8072
rect 23716 8032 23722 8044
rect 23937 8041 23949 8044
rect 23983 8041 23995 8075
rect 23937 8035 23995 8041
rect 2593 8007 2651 8013
rect 2593 7973 2605 8007
rect 2639 7973 2651 8007
rect 2593 7967 2651 7973
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 8570 8004 8576 8016
rect 4120 7976 8576 8004
rect 4120 7964 4126 7976
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 26053 8007 26111 8013
rect 26053 8004 26065 8007
rect 24964 7976 26065 8004
rect 2130 7896 2136 7948
rect 2188 7936 2194 7948
rect 2225 7939 2283 7945
rect 2225 7936 2237 7939
rect 2188 7908 2237 7936
rect 2188 7896 2194 7908
rect 2225 7905 2237 7908
rect 2271 7905 2283 7939
rect 5534 7936 5540 7948
rect 5495 7908 5540 7936
rect 2225 7899 2283 7905
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 6086 7936 6092 7948
rect 5675 7908 6092 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 7190 7896 7196 7948
rect 7248 7936 7254 7948
rect 7285 7939 7343 7945
rect 7285 7936 7297 7939
rect 7248 7908 7297 7936
rect 7248 7896 7254 7908
rect 7285 7905 7297 7908
rect 7331 7936 7343 7939
rect 7650 7936 7656 7948
rect 7331 7908 7656 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 7650 7896 7656 7908
rect 7708 7896 7714 7948
rect 17402 7896 17408 7948
rect 17460 7936 17466 7948
rect 17681 7939 17739 7945
rect 17681 7936 17693 7939
rect 17460 7908 17693 7936
rect 17460 7896 17466 7908
rect 17681 7905 17693 7908
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 21266 7896 21272 7948
rect 21324 7936 21330 7948
rect 21324 7908 21680 7936
rect 21324 7896 21330 7908
rect 3786 7868 3792 7880
rect 3747 7840 3792 7868
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4614 7868 4620 7880
rect 4019 7840 4620 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 5258 7877 5264 7880
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7868 4767 7871
rect 5227 7871 5264 7877
rect 5227 7868 5239 7871
rect 4755 7840 5239 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 5227 7837 5239 7840
rect 5227 7831 5264 7837
rect 5258 7828 5264 7831
rect 5316 7828 5322 7880
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 6972 7840 7757 7868
rect 6972 7828 6978 7840
rect 7745 7837 7757 7840
rect 7791 7837 7803 7871
rect 8018 7868 8024 7880
rect 7979 7840 8024 7868
rect 7745 7831 7803 7837
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7868 9551 7871
rect 10042 7868 10048 7880
rect 9539 7840 10048 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 11330 7828 11336 7880
rect 11388 7877 11394 7880
rect 11388 7868 11400 7877
rect 11388 7840 11433 7868
rect 11388 7831 11400 7840
rect 11388 7828 11394 7831
rect 11514 7828 11520 7880
rect 11572 7868 11578 7880
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11572 7840 11621 7868
rect 11572 7828 11578 7840
rect 11609 7837 11621 7840
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 17494 7828 17500 7880
rect 17552 7868 17558 7880
rect 17589 7871 17647 7877
rect 17589 7868 17601 7871
rect 17552 7840 17601 7868
rect 17552 7828 17558 7840
rect 17589 7837 17601 7840
rect 17635 7837 17647 7871
rect 19058 7868 19064 7880
rect 19019 7840 19064 7868
rect 17589 7831 17647 7837
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7868 20959 7871
rect 21358 7868 21364 7880
rect 20947 7840 21364 7868
rect 20947 7837 20959 7840
rect 20901 7831 20959 7837
rect 21358 7828 21364 7840
rect 21416 7828 21422 7880
rect 21652 7877 21680 7908
rect 21637 7871 21695 7877
rect 21637 7837 21649 7871
rect 21683 7837 21695 7871
rect 21637 7831 21695 7837
rect 22738 7828 22744 7880
rect 22796 7868 22802 7880
rect 23109 7871 23167 7877
rect 23109 7868 23121 7871
rect 22796 7840 23121 7868
rect 22796 7828 22802 7840
rect 23109 7837 23121 7840
rect 23155 7837 23167 7871
rect 23842 7868 23848 7880
rect 23803 7840 23848 7868
rect 23109 7831 23167 7837
rect 23842 7828 23848 7840
rect 23900 7828 23906 7880
rect 24121 7871 24179 7877
rect 24121 7837 24133 7871
rect 24167 7868 24179 7871
rect 24489 7871 24547 7877
rect 24489 7868 24501 7871
rect 24167 7840 24501 7868
rect 24167 7837 24179 7840
rect 24121 7831 24179 7837
rect 24489 7837 24501 7840
rect 24535 7837 24547 7871
rect 24489 7831 24547 7837
rect 24731 7871 24789 7877
rect 24731 7837 24743 7871
rect 24777 7868 24789 7871
rect 24964 7868 24992 7976
rect 26053 7973 26065 7976
rect 26099 8004 26111 8007
rect 26878 8004 26884 8016
rect 26099 7976 26884 8004
rect 26099 7973 26111 7976
rect 26053 7967 26111 7973
rect 26878 7964 26884 7976
rect 26936 7964 26942 8016
rect 28813 8007 28871 8013
rect 28813 7973 28825 8007
rect 28859 7973 28871 8007
rect 28813 7967 28871 7973
rect 25041 7939 25099 7945
rect 25041 7905 25053 7939
rect 25087 7936 25099 7939
rect 25222 7936 25228 7948
rect 25087 7908 25228 7936
rect 25087 7905 25099 7908
rect 25041 7899 25099 7905
rect 25222 7896 25228 7908
rect 25280 7896 25286 7948
rect 26694 7896 26700 7948
rect 26752 7936 26758 7948
rect 27341 7939 27399 7945
rect 27341 7936 27353 7939
rect 26752 7908 27353 7936
rect 26752 7896 26758 7908
rect 27341 7905 27353 7908
rect 27387 7936 27399 7939
rect 27430 7936 27436 7948
rect 27387 7908 27436 7936
rect 27387 7905 27399 7908
rect 27341 7899 27399 7905
rect 27430 7896 27436 7908
rect 27488 7896 27494 7948
rect 28442 7936 28448 7948
rect 28403 7908 28448 7936
rect 28442 7896 28448 7908
rect 28500 7896 28506 7948
rect 28534 7896 28540 7948
rect 28592 7936 28598 7948
rect 28592 7908 28637 7936
rect 28592 7896 28598 7908
rect 24777 7840 24992 7868
rect 24777 7837 24789 7840
rect 24731 7831 24789 7837
rect 25130 7828 25136 7880
rect 25188 7868 25194 7880
rect 25188 7840 25233 7868
rect 25188 7828 25194 7840
rect 26234 7828 26240 7880
rect 26292 7868 26298 7880
rect 26786 7868 26792 7880
rect 26292 7840 26337 7868
rect 26747 7840 26792 7868
rect 26292 7828 26298 7840
rect 26786 7828 26792 7840
rect 26844 7828 26850 7880
rect 26878 7828 26884 7880
rect 26936 7868 26942 7880
rect 26973 7871 27031 7877
rect 26973 7868 26985 7871
rect 26936 7840 26985 7868
rect 26936 7828 26942 7840
rect 26973 7837 26985 7840
rect 27019 7837 27031 7871
rect 26973 7831 27031 7837
rect 27157 7871 27215 7877
rect 27157 7837 27169 7871
rect 27203 7868 27215 7871
rect 27614 7868 27620 7880
rect 27203 7840 27620 7868
rect 27203 7837 27215 7840
rect 27157 7831 27215 7837
rect 27614 7828 27620 7840
rect 27672 7868 27678 7880
rect 27709 7871 27767 7877
rect 27709 7868 27721 7871
rect 27672 7840 27721 7868
rect 27672 7828 27678 7840
rect 27709 7837 27721 7840
rect 27755 7868 27767 7871
rect 27890 7868 27896 7880
rect 27755 7840 27896 7868
rect 27755 7837 27767 7840
rect 27709 7831 27767 7837
rect 27890 7828 27896 7840
rect 27948 7828 27954 7880
rect 28074 7828 28080 7880
rect 28132 7868 28138 7880
rect 28353 7871 28411 7877
rect 28353 7868 28365 7871
rect 28132 7840 28365 7868
rect 28132 7828 28138 7840
rect 28353 7837 28365 7840
rect 28399 7868 28411 7871
rect 28828 7868 28856 7967
rect 28994 7868 29000 7880
rect 28399 7840 28856 7868
rect 28955 7840 29000 7868
rect 28399 7837 28411 7840
rect 28353 7831 28411 7837
rect 28994 7828 29000 7840
rect 29052 7828 29058 7880
rect 4338 7800 4344 7812
rect 4299 7772 4344 7800
rect 4338 7760 4344 7772
rect 4396 7760 4402 7812
rect 4525 7803 4583 7809
rect 4525 7769 4537 7803
rect 4571 7800 4583 7803
rect 4890 7800 4896 7812
rect 4571 7772 4896 7800
rect 4571 7769 4583 7772
rect 4525 7763 4583 7769
rect 4890 7760 4896 7772
rect 4948 7760 4954 7812
rect 7098 7800 7104 7812
rect 7059 7772 7104 7800
rect 7098 7760 7104 7772
rect 7156 7760 7162 7812
rect 7193 7803 7251 7809
rect 7193 7769 7205 7803
rect 7239 7800 7251 7803
rect 21085 7803 21143 7809
rect 7239 7772 7880 7800
rect 7239 7769 7251 7772
rect 7193 7763 7251 7769
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7732 2743 7735
rect 3326 7732 3332 7744
rect 2731 7704 3332 7732
rect 2731 7701 2743 7704
rect 2685 7695 2743 7701
rect 3326 7692 3332 7704
rect 3384 7692 3390 7744
rect 7116 7732 7144 7760
rect 7852 7741 7880 7772
rect 21085 7769 21097 7803
rect 21131 7800 21143 7803
rect 21174 7800 21180 7812
rect 21131 7772 21180 7800
rect 21131 7769 21143 7772
rect 21085 7763 21143 7769
rect 21174 7760 21180 7772
rect 21232 7760 21238 7812
rect 21269 7803 21327 7809
rect 21269 7769 21281 7803
rect 21315 7769 21327 7803
rect 27522 7800 27528 7812
rect 27483 7772 27528 7800
rect 21269 7763 21327 7769
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7116 7704 7573 7732
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 7837 7735 7895 7741
rect 7837 7701 7849 7735
rect 7883 7701 7895 7735
rect 7837 7695 7895 7701
rect 9766 7692 9772 7744
rect 9824 7732 9830 7744
rect 10229 7735 10287 7741
rect 10229 7732 10241 7735
rect 9824 7704 10241 7732
rect 9824 7692 9830 7704
rect 10229 7701 10241 7704
rect 10275 7732 10287 7735
rect 11054 7732 11060 7744
rect 10275 7704 11060 7732
rect 10275 7701 10287 7704
rect 10229 7695 10287 7701
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 17957 7735 18015 7741
rect 17957 7701 17969 7735
rect 18003 7732 18015 7735
rect 18230 7732 18236 7744
rect 18003 7704 18236 7732
rect 18003 7701 18015 7704
rect 17957 7695 18015 7701
rect 18230 7692 18236 7704
rect 18288 7692 18294 7744
rect 18322 7692 18328 7744
rect 18380 7732 18386 7744
rect 18877 7735 18935 7741
rect 18877 7732 18889 7735
rect 18380 7704 18889 7732
rect 18380 7692 18386 7704
rect 18877 7701 18889 7704
rect 18923 7701 18935 7735
rect 18877 7695 18935 7701
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 21284 7732 21312 7763
rect 27522 7760 27528 7772
rect 27580 7760 27586 7812
rect 23290 7732 23296 7744
rect 20864 7704 21312 7732
rect 23251 7704 23296 7732
rect 20864 7692 20870 7704
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 23382 7692 23388 7744
rect 23440 7732 23446 7744
rect 23661 7735 23719 7741
rect 23661 7732 23673 7735
rect 23440 7704 23673 7732
rect 23440 7692 23446 7704
rect 23661 7701 23673 7704
rect 23707 7701 23719 7735
rect 27982 7732 27988 7744
rect 27943 7704 27988 7732
rect 23661 7695 23719 7701
rect 27982 7692 27988 7704
rect 28040 7692 28046 7744
rect 1104 7642 29532 7664
rect 1104 7590 10425 7642
rect 10477 7590 10489 7642
rect 10541 7590 10553 7642
rect 10605 7590 10617 7642
rect 10669 7590 10681 7642
rect 10733 7590 19901 7642
rect 19953 7590 19965 7642
rect 20017 7590 20029 7642
rect 20081 7590 20093 7642
rect 20145 7590 20157 7642
rect 20209 7590 29532 7642
rect 1104 7568 29532 7590
rect 2685 7531 2743 7537
rect 2685 7497 2697 7531
rect 2731 7528 2743 7531
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 2731 7500 3157 7528
rect 2731 7497 2743 7500
rect 2685 7491 2743 7497
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 15838 7528 15844 7540
rect 3145 7491 3203 7497
rect 14844 7500 15844 7528
rect 1581 7463 1639 7469
rect 1581 7429 1593 7463
rect 1627 7460 1639 7463
rect 2130 7460 2136 7472
rect 1627 7432 2136 7460
rect 1627 7429 1639 7432
rect 1581 7423 1639 7429
rect 2130 7420 2136 7432
rect 2188 7420 2194 7472
rect 2774 7420 2780 7472
rect 2832 7460 2838 7472
rect 6914 7460 6920 7472
rect 2832 7432 2877 7460
rect 6875 7432 6920 7460
rect 2832 7420 2838 7432
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 3326 7392 3332 7404
rect 2746 7364 2912 7392
rect 3287 7364 3332 7392
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 2746 7324 2774 7364
rect 2884 7333 2912 7364
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 6546 7392 6552 7404
rect 6507 7364 6552 7392
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 6730 7392 6736 7404
rect 6691 7364 6736 7392
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 7190 7392 7196 7404
rect 7103 7364 7196 7392
rect 7190 7352 7196 7364
rect 7248 7392 7254 7404
rect 7742 7392 7748 7404
rect 7248 7364 7748 7392
rect 7248 7352 7254 7364
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7392 8263 7395
rect 8294 7392 8300 7404
rect 8251 7364 8300 7392
rect 8251 7361 8263 7364
rect 8205 7355 8263 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 8472 7395 8530 7401
rect 8472 7361 8484 7395
rect 8518 7392 8530 7395
rect 8754 7392 8760 7404
rect 8518 7364 8760 7392
rect 8518 7361 8530 7364
rect 8472 7355 8530 7361
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 14844 7401 14872 7500
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 17313 7531 17371 7537
rect 17313 7497 17325 7531
rect 17359 7528 17371 7531
rect 17494 7528 17500 7540
rect 17359 7500 17500 7528
rect 17359 7497 17371 7500
rect 17313 7491 17371 7497
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 18322 7528 18328 7540
rect 18283 7500 18328 7528
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 19518 7488 19524 7540
rect 19576 7528 19582 7540
rect 20254 7528 20260 7540
rect 19576 7500 20260 7528
rect 19576 7488 19582 7500
rect 20254 7488 20260 7500
rect 20312 7528 20318 7540
rect 22738 7528 22744 7540
rect 20312 7500 21036 7528
rect 22699 7500 22744 7528
rect 20312 7488 20318 7500
rect 15930 7460 15936 7472
rect 15396 7432 15936 7460
rect 15396 7401 15424 7432
rect 15930 7420 15936 7432
rect 15988 7420 15994 7472
rect 18230 7420 18236 7472
rect 18288 7460 18294 7472
rect 20806 7460 20812 7472
rect 18288 7432 20812 7460
rect 18288 7420 18294 7432
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7361 15623 7395
rect 15565 7355 15623 7361
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7361 15899 7395
rect 16022 7392 16028 7404
rect 15983 7364 16028 7392
rect 15841 7355 15899 7361
rect 2464 7296 2774 7324
rect 2869 7327 2927 7333
rect 2464 7284 2470 7296
rect 2869 7293 2881 7327
rect 2915 7293 2927 7327
rect 2869 7287 2927 7293
rect 1949 7259 2007 7265
rect 1949 7225 1961 7259
rect 1995 7256 2007 7259
rect 2130 7256 2136 7268
rect 1995 7228 2136 7256
rect 1995 7225 2007 7228
rect 1949 7219 2007 7225
rect 2130 7216 2136 7228
rect 2188 7216 2194 7268
rect 14936 7256 14964 7355
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7324 15163 7327
rect 15580 7324 15608 7355
rect 15151 7296 15608 7324
rect 15151 7293 15163 7296
rect 15105 7287 15163 7293
rect 15654 7284 15660 7336
rect 15712 7324 15718 7336
rect 15856 7324 15884 7355
rect 16022 7352 16028 7364
rect 16080 7352 16086 7404
rect 16393 7395 16451 7401
rect 16393 7361 16405 7395
rect 16439 7392 16451 7395
rect 16666 7392 16672 7404
rect 16439 7364 16672 7392
rect 16439 7361 16451 7364
rect 16393 7355 16451 7361
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 16761 7395 16819 7401
rect 16761 7361 16773 7395
rect 16807 7361 16819 7395
rect 16761 7355 16819 7361
rect 17405 7395 17463 7401
rect 17405 7361 17417 7395
rect 17451 7392 17463 7395
rect 17494 7392 17500 7404
rect 17451 7364 17500 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 15930 7324 15936 7336
rect 15712 7296 15757 7324
rect 15856 7296 15936 7324
rect 15712 7284 15718 7296
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 15746 7256 15752 7268
rect 14936 7228 15752 7256
rect 15746 7216 15752 7228
rect 15804 7216 15810 7268
rect 16574 7216 16580 7268
rect 16632 7256 16638 7268
rect 16776 7256 16804 7355
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 18782 7392 18788 7404
rect 18743 7364 18788 7392
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 19245 7395 19303 7401
rect 19245 7361 19257 7395
rect 19291 7392 19303 7395
rect 19518 7392 19524 7404
rect 19291 7364 19524 7392
rect 19291 7361 19303 7364
rect 19245 7355 19303 7361
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 19628 7401 19656 7432
rect 20806 7420 20812 7432
rect 20864 7420 20870 7472
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7361 19671 7395
rect 19794 7392 19800 7404
rect 19755 7364 19800 7392
rect 19613 7355 19671 7361
rect 19794 7352 19800 7364
rect 19852 7352 19858 7404
rect 20073 7395 20131 7401
rect 20073 7361 20085 7395
rect 20119 7361 20131 7395
rect 20438 7392 20444 7404
rect 20399 7364 20444 7392
rect 20073 7355 20131 7361
rect 17221 7327 17279 7333
rect 17221 7293 17233 7327
rect 17267 7324 17279 7327
rect 17310 7324 17316 7336
rect 17267 7296 17316 7324
rect 17267 7293 17279 7296
rect 17221 7287 17279 7293
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 18064 7256 18092 7287
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18233 7327 18291 7333
rect 18233 7324 18245 7327
rect 18196 7296 18245 7324
rect 18196 7284 18202 7296
rect 18233 7293 18245 7296
rect 18279 7293 18291 7327
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 18233 7287 18291 7293
rect 18708 7296 18981 7324
rect 18322 7256 18328 7268
rect 16632 7228 18328 7256
rect 16632 7216 16638 7228
rect 18322 7216 18328 7228
rect 18380 7216 18386 7268
rect 18708 7265 18736 7296
rect 18969 7293 18981 7296
rect 19015 7293 19027 7327
rect 18969 7287 19027 7293
rect 19702 7284 19708 7336
rect 19760 7324 19766 7336
rect 20088 7324 20116 7355
rect 20438 7352 20444 7364
rect 20496 7352 20502 7404
rect 21008 7401 21036 7500
rect 22738 7488 22744 7500
rect 22796 7488 22802 7540
rect 23842 7488 23848 7540
rect 23900 7528 23906 7540
rect 24581 7531 24639 7537
rect 24581 7528 24593 7531
rect 23900 7500 24593 7528
rect 23900 7488 23906 7500
rect 24581 7497 24593 7500
rect 24627 7497 24639 7531
rect 24581 7491 24639 7497
rect 25222 7488 25228 7540
rect 25280 7528 25286 7540
rect 27246 7528 27252 7540
rect 25280 7500 25912 7528
rect 27207 7500 27252 7528
rect 25280 7488 25286 7500
rect 23382 7460 23388 7472
rect 22572 7432 23388 7460
rect 20533 7395 20591 7401
rect 20533 7361 20545 7395
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 20993 7395 21051 7401
rect 20993 7361 21005 7395
rect 21039 7361 21051 7395
rect 21358 7392 21364 7404
rect 21319 7364 21364 7392
rect 20993 7355 21051 7361
rect 19760 7296 20116 7324
rect 20257 7327 20315 7333
rect 19760 7284 19766 7296
rect 20257 7293 20269 7327
rect 20303 7293 20315 7327
rect 20257 7287 20315 7293
rect 20349 7327 20407 7333
rect 20349 7293 20361 7327
rect 20395 7324 20407 7327
rect 20548 7324 20576 7355
rect 21358 7352 21364 7364
rect 21416 7352 21422 7404
rect 21542 7392 21548 7404
rect 21503 7364 21548 7392
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 22572 7401 22600 7432
rect 23382 7420 23388 7432
rect 23440 7420 23446 7472
rect 25130 7460 25136 7472
rect 25043 7432 25136 7460
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7361 22615 7395
rect 22922 7392 22928 7404
rect 22883 7364 22928 7392
rect 22557 7355 22615 7361
rect 22922 7352 22928 7364
rect 22980 7352 22986 7404
rect 23014 7352 23020 7404
rect 23072 7392 23078 7404
rect 23181 7395 23239 7401
rect 23181 7392 23193 7395
rect 23072 7364 23193 7392
rect 23072 7352 23078 7364
rect 23181 7361 23193 7364
rect 23227 7361 23239 7395
rect 23181 7355 23239 7361
rect 24731 7395 24789 7401
rect 24731 7361 24743 7395
rect 24777 7392 24789 7395
rect 25056 7392 25084 7432
rect 25130 7420 25136 7432
rect 25188 7460 25194 7472
rect 25884 7469 25912 7500
rect 27246 7488 27252 7500
rect 27304 7488 27310 7540
rect 28445 7531 28503 7537
rect 28445 7497 28457 7531
rect 28491 7528 28503 7531
rect 28994 7528 29000 7540
rect 28491 7500 29000 7528
rect 28491 7497 28503 7500
rect 28445 7491 28503 7497
rect 28994 7488 29000 7500
rect 29052 7488 29058 7540
rect 25593 7463 25651 7469
rect 25593 7460 25605 7463
rect 25188 7432 25605 7460
rect 25188 7420 25194 7432
rect 25593 7429 25605 7432
rect 25639 7460 25651 7463
rect 25685 7463 25743 7469
rect 25685 7460 25697 7463
rect 25639 7432 25697 7460
rect 25639 7429 25651 7432
rect 25593 7423 25651 7429
rect 25685 7429 25697 7432
rect 25731 7429 25743 7463
rect 25685 7423 25743 7429
rect 25869 7463 25927 7469
rect 25869 7429 25881 7463
rect 25915 7429 25927 7463
rect 25869 7423 25927 7429
rect 26786 7420 26792 7472
rect 26844 7460 26850 7472
rect 26844 7432 27292 7460
rect 26844 7420 26850 7432
rect 24777 7364 25084 7392
rect 25225 7395 25283 7401
rect 24777 7361 24789 7364
rect 24731 7355 24789 7361
rect 25225 7361 25237 7395
rect 25271 7361 25283 7395
rect 25225 7355 25283 7361
rect 25409 7395 25467 7401
rect 25409 7361 25421 7395
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 26053 7395 26111 7401
rect 26053 7361 26065 7395
rect 26099 7392 26111 7395
rect 26234 7392 26240 7404
rect 26099 7364 26240 7392
rect 26099 7361 26111 7364
rect 26053 7355 26111 7361
rect 21082 7324 21088 7336
rect 20395 7296 20576 7324
rect 21043 7296 21088 7324
rect 20395 7293 20407 7296
rect 20349 7287 20407 7293
rect 18693 7259 18751 7265
rect 18693 7225 18705 7259
rect 18739 7225 18751 7259
rect 19426 7256 19432 7268
rect 19387 7228 19432 7256
rect 18693 7219 18751 7225
rect 19426 7216 19432 7228
rect 19484 7216 19490 7268
rect 20272 7256 20300 7287
rect 21082 7284 21088 7296
rect 21140 7284 21146 7336
rect 22373 7327 22431 7333
rect 22373 7293 22385 7327
rect 22419 7324 22431 7327
rect 22830 7324 22836 7336
rect 22419 7296 22836 7324
rect 22419 7293 22431 7296
rect 22373 7287 22431 7293
rect 22830 7284 22836 7296
rect 22888 7284 22894 7336
rect 25041 7327 25099 7333
rect 25041 7293 25053 7327
rect 25087 7293 25099 7327
rect 25041 7287 25099 7293
rect 21174 7256 21180 7268
rect 20272 7228 20392 7256
rect 21135 7228 21180 7256
rect 2038 7188 2044 7200
rect 1999 7160 2044 7188
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 2222 7148 2228 7200
rect 2280 7188 2286 7200
rect 2317 7191 2375 7197
rect 2317 7188 2329 7191
rect 2280 7160 2329 7188
rect 2280 7148 2286 7160
rect 2317 7157 2329 7160
rect 2363 7157 2375 7191
rect 7098 7188 7104 7200
rect 7059 7160 7104 7188
rect 2317 7151 2375 7157
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 9582 7188 9588 7200
rect 9543 7160 9588 7188
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 16206 7188 16212 7200
rect 16167 7160 16212 7188
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 16853 7191 16911 7197
rect 16853 7188 16865 7191
rect 16816 7160 16865 7188
rect 16816 7148 16822 7160
rect 16853 7157 16865 7160
rect 16899 7188 16911 7191
rect 17402 7188 17408 7200
rect 16899 7160 17408 7188
rect 16899 7157 16911 7160
rect 16853 7151 16911 7157
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 17678 7148 17684 7200
rect 17736 7188 17742 7200
rect 17773 7191 17831 7197
rect 17773 7188 17785 7191
rect 17736 7160 17785 7188
rect 17736 7148 17742 7160
rect 17773 7157 17785 7160
rect 17819 7157 17831 7191
rect 20364 7188 20392 7228
rect 21174 7216 21180 7228
rect 21232 7216 21238 7268
rect 24305 7259 24363 7265
rect 24305 7225 24317 7259
rect 24351 7256 24363 7259
rect 25056 7256 25084 7287
rect 25130 7284 25136 7336
rect 25188 7324 25194 7336
rect 25240 7324 25268 7355
rect 25188 7296 25268 7324
rect 25188 7284 25194 7296
rect 25222 7256 25228 7268
rect 24351 7228 25228 7256
rect 24351 7225 24363 7228
rect 24305 7219 24363 7225
rect 25222 7216 25228 7228
rect 25280 7256 25286 7268
rect 25424 7256 25452 7355
rect 26234 7352 26240 7364
rect 26292 7392 26298 7404
rect 27264 7401 27292 7432
rect 27430 7420 27436 7472
rect 27488 7460 27494 7472
rect 27488 7432 27844 7460
rect 27488 7420 27494 7432
rect 27065 7395 27123 7401
rect 27065 7392 27077 7395
rect 26292 7364 27077 7392
rect 26292 7352 26298 7364
rect 27065 7361 27077 7364
rect 27111 7361 27123 7395
rect 27065 7355 27123 7361
rect 27249 7395 27307 7401
rect 27249 7361 27261 7395
rect 27295 7361 27307 7395
rect 27249 7355 27307 7361
rect 27338 7352 27344 7404
rect 27396 7392 27402 7404
rect 27525 7395 27583 7401
rect 27525 7392 27537 7395
rect 27396 7364 27537 7392
rect 27396 7352 27402 7364
rect 27525 7361 27537 7364
rect 27571 7361 27583 7395
rect 27525 7355 27583 7361
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27816 7392 27844 7432
rect 28295 7395 28353 7401
rect 28295 7392 28307 7395
rect 27816 7364 28307 7392
rect 27709 7355 27767 7361
rect 28295 7361 28307 7364
rect 28341 7361 28353 7395
rect 28295 7355 28353 7361
rect 27154 7284 27160 7336
rect 27212 7324 27218 7336
rect 27430 7324 27436 7336
rect 27212 7296 27436 7324
rect 27212 7284 27218 7296
rect 27430 7284 27436 7296
rect 27488 7284 27494 7336
rect 25280 7228 25452 7256
rect 25280 7216 25286 7228
rect 26326 7216 26332 7268
rect 26384 7256 26390 7268
rect 27522 7256 27528 7268
rect 26384 7228 27528 7256
rect 26384 7216 26390 7228
rect 27522 7216 27528 7228
rect 27580 7256 27586 7268
rect 27724 7256 27752 7355
rect 27890 7324 27896 7336
rect 27851 7296 27896 7324
rect 27890 7284 27896 7296
rect 27948 7284 27954 7336
rect 27985 7327 28043 7333
rect 27985 7293 27997 7327
rect 28031 7293 28043 7327
rect 27985 7287 28043 7293
rect 28000 7256 28028 7287
rect 27580 7228 28028 7256
rect 27580 7216 27586 7228
rect 21910 7188 21916 7200
rect 20364 7160 21916 7188
rect 17773 7151 17831 7157
rect 21910 7148 21916 7160
rect 21968 7148 21974 7200
rect 27614 7148 27620 7200
rect 27672 7188 27678 7200
rect 28534 7188 28540 7200
rect 27672 7160 28540 7188
rect 27672 7148 27678 7160
rect 28534 7148 28540 7160
rect 28592 7148 28598 7200
rect 1104 7098 29532 7120
rect 1104 7046 5688 7098
rect 5740 7046 5752 7098
rect 5804 7046 5816 7098
rect 5868 7046 5880 7098
rect 5932 7046 5944 7098
rect 5996 7046 15163 7098
rect 15215 7046 15227 7098
rect 15279 7046 15291 7098
rect 15343 7046 15355 7098
rect 15407 7046 15419 7098
rect 15471 7046 24639 7098
rect 24691 7046 24703 7098
rect 24755 7046 24767 7098
rect 24819 7046 24831 7098
rect 24883 7046 24895 7098
rect 24947 7046 29532 7098
rect 1104 7024 29532 7046
rect 2130 6944 2136 6996
rect 2188 6984 2194 6996
rect 3786 6984 3792 6996
rect 2188 6956 3792 6984
rect 2188 6944 2194 6956
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 6457 6987 6515 6993
rect 6457 6953 6469 6987
rect 6503 6984 6515 6987
rect 6546 6984 6552 6996
rect 6503 6956 6552 6984
rect 6503 6953 6515 6956
rect 6457 6947 6515 6953
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 6914 6984 6920 6996
rect 6827 6956 6920 6984
rect 6914 6944 6920 6956
rect 6972 6984 6978 6996
rect 7190 6984 7196 6996
rect 6972 6956 7196 6984
rect 6972 6944 6978 6956
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 8754 6984 8760 6996
rect 8715 6956 8760 6984
rect 8754 6944 8760 6956
rect 8812 6944 8818 6996
rect 15746 6984 15752 6996
rect 15707 6956 15752 6984
rect 15746 6944 15752 6956
rect 15804 6944 15810 6996
rect 17494 6944 17500 6996
rect 17552 6984 17558 6996
rect 18141 6987 18199 6993
rect 18141 6984 18153 6987
rect 17552 6956 18153 6984
rect 17552 6944 17558 6956
rect 18141 6953 18153 6956
rect 18187 6953 18199 6987
rect 18141 6947 18199 6953
rect 18509 6987 18567 6993
rect 18509 6953 18521 6987
rect 18555 6984 18567 6987
rect 18782 6984 18788 6996
rect 18555 6956 18788 6984
rect 18555 6953 18567 6956
rect 18509 6947 18567 6953
rect 18782 6944 18788 6956
rect 18840 6944 18846 6996
rect 19702 6984 19708 6996
rect 18892 6956 19708 6984
rect 6730 6916 6736 6928
rect 4356 6888 6736 6916
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2130 6848 2136 6860
rect 2087 6820 2136 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6848 2283 6851
rect 2406 6848 2412 6860
rect 2271 6820 2412 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 2406 6808 2412 6820
rect 2464 6808 2470 6860
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 4356 6857 4384 6888
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 9677 6919 9735 6925
rect 9677 6885 9689 6919
rect 9723 6916 9735 6919
rect 10226 6916 10232 6928
rect 9723 6888 10232 6916
rect 9723 6885 9735 6888
rect 9677 6879 9735 6885
rect 10226 6876 10232 6888
rect 10284 6876 10290 6928
rect 17402 6876 17408 6928
rect 17460 6916 17466 6928
rect 18892 6916 18920 6956
rect 19702 6944 19708 6956
rect 19760 6944 19766 6996
rect 19794 6944 19800 6996
rect 19852 6984 19858 6996
rect 19889 6987 19947 6993
rect 19889 6984 19901 6987
rect 19852 6956 19901 6984
rect 19852 6944 19858 6956
rect 19889 6953 19901 6956
rect 19935 6953 19947 6987
rect 19889 6947 19947 6953
rect 21082 6944 21088 6996
rect 21140 6984 21146 6996
rect 21361 6987 21419 6993
rect 21361 6984 21373 6987
rect 21140 6956 21373 6984
rect 21140 6944 21146 6956
rect 21361 6953 21373 6956
rect 21407 6953 21419 6987
rect 21361 6947 21419 6953
rect 22925 6987 22983 6993
rect 22925 6953 22937 6987
rect 22971 6984 22983 6987
rect 23014 6984 23020 6996
rect 22971 6956 23020 6984
rect 22971 6953 22983 6956
rect 22925 6947 22983 6953
rect 23014 6944 23020 6956
rect 23072 6944 23078 6996
rect 25041 6987 25099 6993
rect 25041 6953 25053 6987
rect 25087 6984 25099 6987
rect 25314 6984 25320 6996
rect 25087 6956 25320 6984
rect 25087 6953 25099 6956
rect 25041 6947 25099 6953
rect 25314 6944 25320 6956
rect 25372 6944 25378 6996
rect 26605 6987 26663 6993
rect 26605 6953 26617 6987
rect 26651 6984 26663 6987
rect 26651 6956 26924 6984
rect 26651 6953 26663 6956
rect 26605 6947 26663 6953
rect 19058 6916 19064 6928
rect 17460 6888 18920 6916
rect 19019 6888 19064 6916
rect 17460 6876 17466 6888
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 26786 6916 26792 6928
rect 26528 6888 26792 6916
rect 4341 6851 4399 6857
rect 4341 6848 4353 6851
rect 4212 6820 4353 6848
rect 4212 6808 4218 6820
rect 4341 6817 4353 6820
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6848 7067 6851
rect 7190 6848 7196 6860
rect 7055 6820 7196 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 7190 6808 7196 6820
rect 7248 6808 7254 6860
rect 7650 6808 7656 6860
rect 7708 6848 7714 6860
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 7708 6820 8217 6848
rect 7708 6808 7714 6820
rect 8205 6817 8217 6820
rect 8251 6817 8263 6851
rect 8205 6811 8263 6817
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 9769 6851 9827 6857
rect 9769 6848 9781 6851
rect 9640 6820 9781 6848
rect 9640 6808 9646 6820
rect 9769 6817 9781 6820
rect 9815 6817 9827 6851
rect 9769 6811 9827 6817
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 16393 6851 16451 6857
rect 9916 6820 16344 6848
rect 9916 6808 9922 6820
rect 1854 6740 1860 6792
rect 1912 6780 1918 6792
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 1912 6752 2605 6780
rect 1912 6740 1918 6752
rect 2593 6749 2605 6752
rect 2639 6749 2651 6783
rect 5902 6780 5908 6792
rect 5863 6752 5908 6780
rect 2593 6743 2651 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6178 6780 6184 6792
rect 6135 6752 6184 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6749 6791 6783
rect 7282 6780 7288 6792
rect 7243 6752 7288 6780
rect 6733 6743 6791 6749
rect 1949 6715 2007 6721
rect 1949 6681 1961 6715
rect 1995 6712 2007 6715
rect 1995 6684 2452 6712
rect 1995 6681 2007 6684
rect 1949 6675 2007 6681
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 1670 6644 1676 6656
rect 1627 6616 1676 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1670 6604 1676 6616
rect 1728 6604 1734 6656
rect 2424 6653 2452 6684
rect 2958 6672 2964 6724
rect 3016 6712 3022 6724
rect 4249 6715 4307 6721
rect 4249 6712 4261 6715
rect 3016 6684 4261 6712
rect 3016 6672 3022 6684
rect 4249 6681 4261 6684
rect 4295 6681 4307 6715
rect 5920 6712 5948 6740
rect 6656 6712 6684 6743
rect 5920 6684 6684 6712
rect 6748 6712 6776 6743
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 8478 6780 8484 6792
rect 7975 6752 8484 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 7098 6712 7104 6724
rect 6748 6684 7104 6712
rect 4249 6675 4307 6681
rect 7098 6672 7104 6684
rect 7156 6672 7162 6724
rect 7576 6712 7604 6743
rect 8478 6740 8484 6752
rect 8536 6780 8542 6792
rect 9307 6783 9365 6789
rect 8536 6752 9168 6780
rect 8536 6740 8542 6752
rect 7837 6715 7895 6721
rect 7837 6712 7849 6715
rect 7576 6684 7849 6712
rect 7837 6681 7849 6684
rect 7883 6712 7895 6715
rect 8389 6715 8447 6721
rect 8389 6712 8401 6715
rect 7883 6684 8401 6712
rect 7883 6681 7895 6684
rect 7837 6675 7895 6681
rect 8389 6681 8401 6684
rect 8435 6681 8447 6715
rect 8389 6675 8447 6681
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6613 2467 6647
rect 2409 6607 2467 6613
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 4157 6647 4215 6653
rect 4157 6644 4169 6647
rect 3384 6616 4169 6644
rect 3384 6604 3390 6616
rect 4157 6613 4169 6616
rect 4203 6613 4215 6647
rect 4157 6607 4215 6613
rect 5997 6647 6055 6653
rect 5997 6613 6009 6647
rect 6043 6644 6055 6647
rect 6086 6644 6092 6656
rect 6043 6616 6092 6644
rect 6043 6613 6055 6616
rect 5997 6607 6055 6613
rect 6086 6604 6092 6616
rect 6144 6604 6150 6656
rect 6730 6604 6736 6656
rect 6788 6644 6794 6656
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 6788 6616 7297 6644
rect 6788 6604 6794 6616
rect 7285 6613 7297 6616
rect 7331 6613 7343 6647
rect 8294 6644 8300 6656
rect 8255 6616 8300 6644
rect 7285 6607 7343 6613
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 9140 6653 9168 6752
rect 9307 6749 9319 6783
rect 9353 6780 9365 6783
rect 9600 6780 9628 6808
rect 9353 6752 9628 6780
rect 10689 6783 10747 6789
rect 9353 6749 9365 6752
rect 9307 6743 9365 6749
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 11422 6780 11428 6792
rect 10735 6752 11428 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6780 16175 6783
rect 16206 6780 16212 6792
rect 16163 6752 16212 6780
rect 16163 6749 16175 6752
rect 16117 6743 16175 6749
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 16316 6780 16344 6820
rect 16393 6817 16405 6851
rect 16439 6848 16451 6851
rect 16574 6848 16580 6860
rect 16439 6820 16580 6848
rect 16439 6817 16451 6820
rect 16393 6811 16451 6817
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 16945 6851 17003 6857
rect 16945 6848 16957 6851
rect 16724 6820 16957 6848
rect 16724 6808 16730 6820
rect 16945 6817 16957 6820
rect 16991 6817 17003 6851
rect 16945 6811 17003 6817
rect 17310 6808 17316 6860
rect 17368 6848 17374 6860
rect 18233 6851 18291 6857
rect 18233 6848 18245 6851
rect 17368 6820 18245 6848
rect 17368 6808 17374 6820
rect 18233 6817 18245 6820
rect 18279 6817 18291 6851
rect 21358 6848 21364 6860
rect 18233 6811 18291 6817
rect 20824 6820 21364 6848
rect 17218 6780 17224 6792
rect 16316 6752 17224 6780
rect 17218 6740 17224 6752
rect 17276 6740 17282 6792
rect 18138 6780 18144 6792
rect 18051 6752 18144 6780
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 20824 6789 20852 6820
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 21818 6808 21824 6860
rect 21876 6848 21882 6860
rect 21913 6851 21971 6857
rect 21913 6848 21925 6851
rect 21876 6820 21925 6848
rect 21876 6808 21882 6820
rect 21913 6817 21925 6820
rect 21959 6817 21971 6851
rect 21913 6811 21971 6817
rect 23106 6808 23112 6860
rect 23164 6848 23170 6860
rect 23477 6851 23535 6857
rect 23477 6848 23489 6851
rect 23164 6820 23489 6848
rect 23164 6808 23170 6820
rect 23477 6817 23489 6820
rect 23523 6817 23535 6851
rect 23477 6811 23535 6817
rect 24486 6808 24492 6860
rect 24544 6848 24550 6860
rect 26528 6857 26556 6888
rect 26786 6876 26792 6888
rect 26844 6876 26850 6928
rect 24857 6851 24915 6857
rect 24857 6848 24869 6851
rect 24544 6820 24869 6848
rect 24544 6808 24550 6820
rect 24857 6817 24869 6820
rect 24903 6817 24915 6851
rect 24857 6811 24915 6817
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 26694 6848 26700 6860
rect 26559 6820 26593 6848
rect 26655 6820 26700 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 26694 6808 26700 6820
rect 26752 6808 26758 6860
rect 26896 6792 26924 6956
rect 27522 6944 27528 6996
rect 27580 6984 27586 6996
rect 29089 6987 29147 6993
rect 29089 6984 29101 6987
rect 27580 6956 29101 6984
rect 27580 6944 27586 6956
rect 29089 6953 29101 6956
rect 29135 6953 29147 6987
rect 29089 6947 29147 6953
rect 27246 6848 27252 6860
rect 27207 6820 27252 6848
rect 27246 6808 27252 6820
rect 27304 6808 27310 6860
rect 27706 6848 27712 6860
rect 27667 6820 27712 6848
rect 27706 6808 27712 6820
rect 27764 6808 27770 6860
rect 20809 6783 20867 6789
rect 20809 6749 20821 6783
rect 20855 6749 20867 6783
rect 20809 6743 20867 6749
rect 20898 6740 20904 6792
rect 20956 6780 20962 6792
rect 21266 6780 21272 6792
rect 20956 6752 21001 6780
rect 21227 6752 21272 6780
rect 20956 6740 20962 6752
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 21542 6740 21548 6792
rect 21600 6780 21606 6792
rect 21729 6783 21787 6789
rect 21729 6780 21741 6783
rect 21600 6752 21741 6780
rect 21600 6740 21606 6752
rect 21729 6749 21741 6752
rect 21775 6749 21787 6783
rect 21729 6743 21787 6749
rect 22094 6740 22100 6792
rect 22152 6780 22158 6792
rect 22281 6783 22339 6789
rect 22281 6780 22293 6783
rect 22152 6752 22293 6780
rect 22152 6740 22158 6752
rect 22281 6749 22293 6752
rect 22327 6749 22339 6783
rect 22462 6780 22468 6792
rect 22423 6752 22468 6780
rect 22281 6743 22339 6749
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 23293 6783 23351 6789
rect 23293 6749 23305 6783
rect 23339 6780 23351 6783
rect 23382 6780 23388 6792
rect 23339 6752 23388 6780
rect 23339 6749 23351 6752
rect 23293 6743 23351 6749
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 25041 6783 25099 6789
rect 25041 6749 25053 6783
rect 25087 6780 25099 6783
rect 25222 6780 25228 6792
rect 25087 6752 25228 6780
rect 25087 6749 25099 6752
rect 25041 6743 25099 6749
rect 25222 6740 25228 6752
rect 25280 6740 25286 6792
rect 26326 6780 26332 6792
rect 26287 6752 26332 6780
rect 26326 6740 26332 6752
rect 26384 6740 26390 6792
rect 26878 6780 26884 6792
rect 26839 6752 26884 6780
rect 26878 6740 26884 6752
rect 26936 6780 26942 6792
rect 27338 6780 27344 6792
rect 26936 6752 27344 6780
rect 26936 6740 26942 6752
rect 27338 6740 27344 6752
rect 27396 6740 27402 6792
rect 27982 6789 27988 6792
rect 27976 6743 27988 6789
rect 28040 6780 28046 6792
rect 28040 6752 28076 6780
rect 27982 6740 27988 6743
rect 28040 6740 28046 6752
rect 16022 6672 16028 6724
rect 16080 6712 16086 6724
rect 16390 6712 16396 6724
rect 16080 6684 16396 6712
rect 16080 6672 16086 6684
rect 9125 6647 9183 6653
rect 9125 6613 9137 6647
rect 9171 6613 9183 6647
rect 9125 6607 9183 6613
rect 9309 6647 9367 6653
rect 9309 6613 9321 6647
rect 9355 6644 9367 6647
rect 10226 6644 10232 6656
rect 9355 6616 10232 6644
rect 9355 6613 9367 6616
rect 9309 6607 9367 6613
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 10318 6604 10324 6656
rect 10376 6644 10382 6656
rect 16224 6653 16252 6684
rect 16390 6672 16396 6684
rect 16448 6712 16454 6724
rect 16577 6715 16635 6721
rect 16577 6712 16589 6715
rect 16448 6684 16589 6712
rect 16448 6672 16454 6684
rect 16577 6681 16589 6684
rect 16623 6681 16635 6715
rect 16577 6675 16635 6681
rect 16758 6672 16764 6724
rect 16816 6712 16822 6724
rect 18156 6712 18184 6740
rect 18690 6712 18696 6724
rect 16816 6684 17816 6712
rect 18156 6684 18696 6712
rect 16816 6672 16822 6684
rect 17788 6656 17816 6684
rect 18690 6672 18696 6684
rect 18748 6672 18754 6724
rect 18877 6715 18935 6721
rect 18877 6681 18889 6715
rect 18923 6712 18935 6715
rect 21821 6715 21879 6721
rect 18923 6684 21128 6712
rect 18923 6681 18935 6684
rect 18877 6675 18935 6681
rect 10505 6647 10563 6653
rect 10505 6644 10517 6647
rect 10376 6616 10517 6644
rect 10376 6604 10382 6616
rect 10505 6613 10517 6616
rect 10551 6613 10563 6647
rect 10505 6607 10563 6613
rect 16209 6647 16267 6653
rect 16209 6613 16221 6647
rect 16255 6613 16267 6647
rect 16209 6607 16267 6613
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 18892 6644 18920 6675
rect 20622 6644 20628 6656
rect 17828 6616 18920 6644
rect 20583 6616 20628 6644
rect 17828 6604 17834 6616
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 21100 6653 21128 6684
rect 21821 6681 21833 6715
rect 21867 6712 21879 6715
rect 22189 6715 22247 6721
rect 22189 6712 22201 6715
rect 21867 6684 22201 6712
rect 21867 6681 21879 6684
rect 21821 6675 21879 6681
rect 22189 6681 22201 6684
rect 22235 6681 22247 6715
rect 22189 6675 22247 6681
rect 24394 6672 24400 6724
rect 24452 6712 24458 6724
rect 24765 6715 24823 6721
rect 24765 6712 24777 6715
rect 24452 6684 24777 6712
rect 24452 6672 24458 6684
rect 24765 6681 24777 6684
rect 24811 6681 24823 6715
rect 26605 6715 26663 6721
rect 26605 6712 26617 6715
rect 24765 6675 24823 6681
rect 25240 6684 26617 6712
rect 21085 6647 21143 6653
rect 21085 6613 21097 6647
rect 21131 6613 21143 6647
rect 21085 6607 21143 6613
rect 23290 6604 23296 6656
rect 23348 6644 23354 6656
rect 25240 6653 25268 6684
rect 26605 6681 26617 6684
rect 26651 6681 26663 6715
rect 26605 6675 26663 6681
rect 23385 6647 23443 6653
rect 23385 6644 23397 6647
rect 23348 6616 23397 6644
rect 23348 6604 23354 6616
rect 23385 6613 23397 6616
rect 23431 6613 23443 6647
rect 23385 6607 23443 6613
rect 25225 6647 25283 6653
rect 25225 6613 25237 6647
rect 25271 6613 25283 6647
rect 26142 6644 26148 6656
rect 26103 6616 26148 6644
rect 25225 6607 25283 6613
rect 26142 6604 26148 6616
rect 26200 6604 26206 6656
rect 27154 6644 27160 6656
rect 27115 6616 27160 6644
rect 27154 6604 27160 6616
rect 27212 6604 27218 6656
rect 1104 6554 29532 6576
rect 1104 6502 10425 6554
rect 10477 6502 10489 6554
rect 10541 6502 10553 6554
rect 10605 6502 10617 6554
rect 10669 6502 10681 6554
rect 10733 6502 19901 6554
rect 19953 6502 19965 6554
rect 20017 6502 20029 6554
rect 20081 6502 20093 6554
rect 20145 6502 20157 6554
rect 20209 6502 29532 6554
rect 1104 6480 29532 6502
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3513 6443 3571 6449
rect 3513 6440 3525 6443
rect 2832 6412 3525 6440
rect 2832 6400 2838 6412
rect 3513 6409 3525 6412
rect 3559 6409 3571 6443
rect 4338 6440 4344 6452
rect 3513 6403 3571 6409
rect 3712 6412 4344 6440
rect 2958 6372 2964 6384
rect 2919 6344 2964 6372
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6273 3203 6307
rect 3326 6304 3332 6316
rect 3287 6276 3332 6304
rect 3145 6267 3203 6273
rect 3160 6236 3188 6267
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3712 6304 3740 6412
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6089 6443 6147 6449
rect 6089 6440 6101 6443
rect 5960 6412 6101 6440
rect 5960 6400 5966 6412
rect 6089 6409 6101 6412
rect 6135 6440 6147 6443
rect 7009 6443 7067 6449
rect 6135 6412 6592 6440
rect 6135 6409 6147 6412
rect 6089 6403 6147 6409
rect 6564 6384 6592 6412
rect 7009 6409 7021 6443
rect 7055 6440 7067 6443
rect 7282 6440 7288 6452
rect 7055 6412 7288 6440
rect 7055 6409 7067 6412
rect 7009 6403 7067 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 8294 6440 8300 6452
rect 8255 6412 8300 6440
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 18690 6400 18696 6452
rect 18748 6440 18754 6452
rect 19153 6443 19211 6449
rect 19153 6440 19165 6443
rect 18748 6412 19165 6440
rect 18748 6400 18754 6412
rect 19153 6409 19165 6412
rect 19199 6409 19211 6443
rect 19153 6403 19211 6409
rect 21726 6400 21732 6452
rect 21784 6440 21790 6452
rect 25406 6440 25412 6452
rect 21784 6412 25412 6440
rect 21784 6400 21790 6412
rect 25406 6400 25412 6412
rect 25464 6400 25470 6452
rect 26697 6443 26755 6449
rect 26697 6409 26709 6443
rect 26743 6440 26755 6443
rect 26878 6440 26884 6452
rect 26743 6412 26884 6440
rect 26743 6409 26755 6412
rect 26697 6403 26755 6409
rect 26878 6400 26884 6412
rect 26936 6400 26942 6452
rect 6546 6372 6552 6384
rect 6459 6344 6552 6372
rect 6546 6332 6552 6344
rect 6604 6332 6610 6384
rect 6733 6375 6791 6381
rect 6733 6341 6745 6375
rect 6779 6372 6791 6375
rect 6914 6372 6920 6384
rect 6779 6344 6920 6372
rect 6779 6341 6791 6344
rect 6733 6335 6791 6341
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 7024 6344 7604 6372
rect 3878 6304 3884 6316
rect 3467 6276 3740 6304
rect 3839 6276 3884 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3878 6264 3884 6276
rect 3936 6264 3942 6316
rect 4522 6304 4528 6316
rect 4483 6276 4528 6304
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 4976 6307 5034 6313
rect 4976 6273 4988 6307
rect 5022 6304 5034 6307
rect 5350 6304 5356 6316
rect 5022 6276 5356 6304
rect 5022 6273 5034 6276
rect 4976 6267 5034 6273
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 7024 6304 7052 6344
rect 7576 6316 7604 6344
rect 17494 6332 17500 6384
rect 17552 6372 17558 6384
rect 17589 6375 17647 6381
rect 17589 6372 17601 6375
rect 17552 6344 17601 6372
rect 17552 6332 17558 6344
rect 17589 6341 17601 6344
rect 17635 6372 17647 6375
rect 18782 6372 18788 6384
rect 17635 6344 18788 6372
rect 17635 6341 17647 6344
rect 17589 6335 17647 6341
rect 18782 6332 18788 6344
rect 18840 6332 18846 6384
rect 24673 6375 24731 6381
rect 24673 6372 24685 6375
rect 23584 6344 24685 6372
rect 23584 6316 23612 6344
rect 24673 6341 24685 6344
rect 24719 6341 24731 6375
rect 24673 6335 24731 6341
rect 24857 6375 24915 6381
rect 24857 6341 24869 6375
rect 24903 6372 24915 6375
rect 25130 6372 25136 6384
rect 24903 6344 25136 6372
rect 24903 6341 24915 6344
rect 24857 6335 24915 6341
rect 25130 6332 25136 6344
rect 25188 6332 25194 6384
rect 25866 6372 25872 6384
rect 25240 6344 25872 6372
rect 7190 6304 7196 6316
rect 6236 6276 7052 6304
rect 7151 6276 7196 6304
rect 6236 6264 6242 6276
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 7616 6276 8033 6304
rect 7616 6264 7622 6276
rect 8021 6273 8033 6276
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6304 8355 6307
rect 8478 6304 8484 6316
rect 8343 6276 8484 6304
rect 8343 6273 8355 6276
rect 8297 6267 8355 6273
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 11054 6304 11060 6316
rect 11112 6313 11118 6316
rect 11024 6276 11060 6304
rect 11054 6264 11060 6276
rect 11112 6267 11124 6313
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6304 11391 6307
rect 11514 6304 11520 6316
rect 11379 6276 11520 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11112 6264 11118 6267
rect 11514 6264 11520 6276
rect 11572 6304 11578 6316
rect 12894 6304 12900 6316
rect 11572 6276 12900 6304
rect 11572 6264 11578 6276
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16390 6304 16396 6316
rect 15979 6276 16396 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 17770 6304 17776 6316
rect 17731 6276 17776 6304
rect 17770 6264 17776 6276
rect 17828 6264 17834 6316
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6304 18015 6307
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 18003 6276 18061 6304
rect 18003 6273 18015 6276
rect 17957 6267 18015 6273
rect 18049 6273 18061 6276
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 19245 6307 19303 6313
rect 19245 6273 19257 6307
rect 19291 6304 19303 6307
rect 19518 6304 19524 6316
rect 19291 6276 19524 6304
rect 19291 6273 19303 6276
rect 19245 6267 19303 6273
rect 19518 6264 19524 6276
rect 19576 6264 19582 6316
rect 21266 6264 21272 6316
rect 21324 6304 21330 6316
rect 21821 6307 21879 6313
rect 21821 6304 21833 6307
rect 21324 6276 21833 6304
rect 21324 6264 21330 6276
rect 21821 6273 21833 6276
rect 21867 6273 21879 6307
rect 23566 6304 23572 6316
rect 23527 6276 23572 6304
rect 21821 6267 21879 6273
rect 23566 6264 23572 6276
rect 23624 6264 23630 6316
rect 23753 6307 23811 6313
rect 23753 6273 23765 6307
rect 23799 6273 23811 6307
rect 23753 6267 23811 6273
rect 3970 6236 3976 6248
rect 3160 6208 3832 6236
rect 3931 6208 3976 6236
rect 3804 6112 3832 6208
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 4154 6236 4160 6248
rect 4111 6208 4160 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 7282 6236 7288 6248
rect 7243 6208 7288 6236
rect 4709 6199 4767 6205
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 4433 6103 4491 6109
rect 4433 6100 4445 6103
rect 3844 6072 4445 6100
rect 3844 6060 3850 6072
rect 4433 6069 4445 6072
rect 4479 6069 4491 6103
rect 4724 6100 4752 6199
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 23768 6236 23796 6267
rect 24394 6264 24400 6316
rect 24452 6304 24458 6316
rect 24489 6307 24547 6313
rect 24489 6304 24501 6307
rect 24452 6276 24501 6304
rect 24452 6264 24458 6276
rect 24489 6273 24501 6276
rect 24535 6273 24547 6307
rect 25240 6304 25268 6344
rect 25866 6332 25872 6344
rect 25924 6372 25930 6384
rect 25924 6344 26234 6372
rect 25924 6332 25930 6344
rect 24489 6267 24547 6273
rect 24964 6276 25268 6304
rect 25584 6307 25642 6313
rect 24964 6236 24992 6276
rect 25584 6273 25596 6307
rect 25630 6304 25642 6307
rect 25958 6304 25964 6316
rect 25630 6276 25964 6304
rect 25630 6273 25642 6276
rect 25584 6267 25642 6273
rect 25958 6264 25964 6276
rect 26016 6264 26022 6316
rect 26206 6304 26234 6344
rect 26973 6307 27031 6313
rect 26973 6304 26985 6307
rect 26206 6276 26985 6304
rect 26973 6273 26985 6276
rect 27019 6273 27031 6307
rect 27154 6304 27160 6316
rect 27115 6276 27160 6304
rect 26973 6267 27031 6273
rect 27154 6264 27160 6276
rect 27212 6264 27218 6316
rect 23768 6208 24992 6236
rect 25038 6196 25044 6248
rect 25096 6236 25102 6248
rect 25314 6236 25320 6248
rect 25096 6208 25320 6236
rect 25096 6196 25102 6208
rect 25314 6196 25320 6208
rect 25372 6196 25378 6248
rect 6362 6168 6368 6180
rect 6323 6140 6368 6168
rect 6362 6128 6368 6140
rect 6420 6128 6426 6180
rect 8386 6168 8392 6180
rect 6472 6140 8392 6168
rect 6472 6100 6500 6140
rect 8386 6128 8392 6140
rect 8444 6128 8450 6180
rect 23474 6168 23480 6180
rect 23435 6140 23480 6168
rect 23474 6128 23480 6140
rect 23532 6128 23538 6180
rect 26418 6128 26424 6180
rect 26476 6168 26482 6180
rect 27249 6171 27307 6177
rect 27249 6168 27261 6171
rect 26476 6140 27261 6168
rect 26476 6128 26482 6140
rect 27249 6137 27261 6140
rect 27295 6137 27307 6171
rect 27249 6131 27307 6137
rect 4724 6072 6500 6100
rect 4433 6063 4491 6069
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7193 6103 7251 6109
rect 7193 6100 7205 6103
rect 6972 6072 7205 6100
rect 6972 6060 6978 6072
rect 7193 6069 7205 6072
rect 7239 6069 7251 6103
rect 9950 6100 9956 6112
rect 9911 6072 9956 6100
rect 7193 6063 7251 6069
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 15838 6100 15844 6112
rect 15799 6072 15844 6100
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 18233 6103 18291 6109
rect 18233 6069 18245 6103
rect 18279 6100 18291 6103
rect 18690 6100 18696 6112
rect 18279 6072 18696 6100
rect 18279 6069 18291 6072
rect 18233 6063 18291 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 22002 6100 22008 6112
rect 21915 6072 22008 6100
rect 22002 6060 22008 6072
rect 22060 6100 22066 6112
rect 22462 6100 22468 6112
rect 22060 6072 22468 6100
rect 22060 6060 22066 6072
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 1104 6010 29532 6032
rect 1104 5958 5688 6010
rect 5740 5958 5752 6010
rect 5804 5958 5816 6010
rect 5868 5958 5880 6010
rect 5932 5958 5944 6010
rect 5996 5958 15163 6010
rect 15215 5958 15227 6010
rect 15279 5958 15291 6010
rect 15343 5958 15355 6010
rect 15407 5958 15419 6010
rect 15471 5958 24639 6010
rect 24691 5958 24703 6010
rect 24755 5958 24767 6010
rect 24819 5958 24831 6010
rect 24883 5958 24895 6010
rect 24947 5958 29532 6010
rect 1104 5936 29532 5958
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 3326 5896 3332 5908
rect 2823 5868 3332 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4341 5899 4399 5905
rect 4341 5896 4353 5899
rect 4028 5868 4353 5896
rect 4028 5856 4034 5868
rect 4341 5865 4353 5868
rect 4387 5865 4399 5899
rect 5350 5896 5356 5908
rect 5311 5868 5356 5896
rect 4341 5859 4399 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 9858 5896 9864 5908
rect 5460 5868 9864 5896
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 5460 5828 5488 5868
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10318 5856 10324 5908
rect 10376 5856 10382 5908
rect 10965 5899 11023 5905
rect 10965 5865 10977 5899
rect 11011 5896 11023 5899
rect 11054 5896 11060 5908
rect 11011 5868 11060 5896
rect 11011 5865 11023 5868
rect 10965 5859 11023 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11422 5896 11428 5908
rect 11383 5868 11428 5896
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 15838 5856 15844 5908
rect 15896 5896 15902 5908
rect 19245 5899 19303 5905
rect 19245 5896 19257 5899
rect 15896 5868 19257 5896
rect 15896 5856 15902 5868
rect 19245 5865 19257 5868
rect 19291 5865 19303 5899
rect 20622 5896 20628 5908
rect 19245 5859 19303 5865
rect 19628 5868 20628 5896
rect 6086 5828 6092 5840
rect 4120 5800 5488 5828
rect 5828 5800 6092 5828
rect 4120 5788 4126 5800
rect 3878 5760 3884 5772
rect 3436 5732 3884 5760
rect 3436 5704 3464 5732
rect 3878 5720 3884 5732
rect 3936 5760 3942 5772
rect 3936 5732 4108 5760
rect 3936 5720 3942 5732
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 1670 5701 1676 5704
rect 1664 5655 1676 5701
rect 1728 5692 1734 5704
rect 3418 5692 3424 5704
rect 1728 5664 1764 5692
rect 3379 5664 3424 5692
rect 1670 5652 1676 5655
rect 1728 5652 1734 5664
rect 3418 5652 3424 5664
rect 3476 5652 3482 5704
rect 3786 5692 3792 5704
rect 3747 5664 3792 5692
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4080 5701 4108 5732
rect 4522 5720 4528 5772
rect 4580 5720 4586 5772
rect 5828 5769 5856 5800
rect 6086 5788 6092 5800
rect 6144 5788 6150 5840
rect 10336 5828 10364 5856
rect 15856 5828 15884 5856
rect 19628 5828 19656 5868
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 23106 5856 23112 5908
rect 23164 5896 23170 5908
rect 23382 5896 23388 5908
rect 23164 5868 23388 5896
rect 23164 5856 23170 5868
rect 23382 5856 23388 5868
rect 23440 5856 23446 5908
rect 23566 5856 23572 5908
rect 23624 5896 23630 5908
rect 23845 5899 23903 5905
rect 23845 5896 23857 5899
rect 23624 5868 23857 5896
rect 23624 5856 23630 5868
rect 23845 5865 23857 5868
rect 23891 5865 23903 5899
rect 23845 5859 23903 5865
rect 8956 5800 10160 5828
rect 10336 5800 10548 5828
rect 8956 5772 8984 5800
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5729 5871 5763
rect 5813 5723 5871 5729
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5760 6055 5763
rect 7650 5760 7656 5772
rect 6043 5732 7656 5760
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 7650 5720 7656 5732
rect 7708 5760 7714 5772
rect 8938 5760 8944 5772
rect 7708 5732 8944 5760
rect 7708 5720 7714 5732
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 9723 5732 10057 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 10132 5760 10160 5800
rect 10318 5760 10324 5772
rect 10132 5732 10324 5760
rect 10045 5723 10103 5729
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 10520 5769 10548 5800
rect 15396 5800 15884 5828
rect 16224 5800 19656 5828
rect 15396 5769 15424 5800
rect 10505 5763 10563 5769
rect 10505 5729 10517 5763
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 15381 5763 15439 5769
rect 15381 5729 15393 5763
rect 15427 5729 15439 5763
rect 15562 5760 15568 5772
rect 15523 5732 15568 5760
rect 15381 5723 15439 5729
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 16114 5760 16120 5772
rect 16075 5732 16120 5760
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4209 5695 4267 5701
rect 4209 5661 4221 5695
rect 4255 5692 4267 5695
rect 4540 5692 4568 5720
rect 4893 5695 4951 5701
rect 4893 5692 4905 5695
rect 4255 5664 4905 5692
rect 4255 5661 4267 5664
rect 4209 5655 4267 5661
rect 4893 5661 4905 5664
rect 4939 5661 4951 5695
rect 6546 5692 6552 5704
rect 6507 5664 6552 5692
rect 4893 5655 4951 5661
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 7558 5652 7564 5704
rect 7616 5692 7622 5704
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 7616 5664 7849 5692
rect 7616 5652 7622 5664
rect 7837 5661 7849 5664
rect 7883 5661 7895 5695
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 7837 5655 7895 5661
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 9490 5692 9496 5704
rect 9451 5664 9496 5692
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 9950 5692 9956 5704
rect 9911 5664 9956 5692
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 11146 5692 11152 5704
rect 10928 5664 11152 5692
rect 10928 5652 10934 5664
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5692 15347 5695
rect 15654 5692 15660 5704
rect 15335 5664 15660 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 3513 5627 3571 5633
rect 3513 5593 3525 5627
rect 3559 5624 3571 5627
rect 3973 5627 4031 5633
rect 3973 5624 3985 5627
rect 3559 5596 3985 5624
rect 3559 5593 3571 5596
rect 3513 5587 3571 5593
rect 3973 5593 3985 5596
rect 4019 5593 4031 5627
rect 3973 5587 4031 5593
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 4525 5627 4583 5633
rect 4525 5624 4537 5627
rect 4396 5596 4537 5624
rect 4396 5584 4402 5596
rect 4525 5593 4537 5596
rect 4571 5593 4583 5627
rect 4525 5587 4583 5593
rect 4709 5627 4767 5633
rect 4709 5593 4721 5627
rect 4755 5593 4767 5627
rect 4709 5587 4767 5593
rect 5721 5627 5779 5633
rect 5721 5593 5733 5627
rect 5767 5624 5779 5627
rect 6457 5627 6515 5633
rect 6457 5624 6469 5627
rect 5767 5596 6469 5624
rect 5767 5593 5779 5596
rect 5721 5587 5779 5593
rect 6457 5593 6469 5596
rect 6503 5624 6515 5627
rect 7190 5624 7196 5636
rect 6503 5596 7196 5624
rect 6503 5593 6515 5596
rect 6457 5587 6515 5593
rect 3329 5559 3387 5565
rect 3329 5525 3341 5559
rect 3375 5556 3387 5559
rect 4724 5556 4752 5587
rect 7190 5584 7196 5596
rect 7248 5584 7254 5636
rect 8205 5627 8263 5633
rect 8205 5593 8217 5627
rect 8251 5624 8263 5627
rect 8846 5624 8852 5636
rect 8251 5596 8852 5624
rect 8251 5593 8263 5596
rect 8205 5587 8263 5593
rect 8846 5584 8852 5596
rect 8904 5584 8910 5636
rect 9769 5627 9827 5633
rect 9769 5593 9781 5627
rect 9815 5593 9827 5627
rect 9769 5587 9827 5593
rect 9861 5627 9919 5633
rect 9861 5593 9873 5627
rect 9907 5624 9919 5627
rect 10226 5624 10232 5636
rect 9907 5596 10232 5624
rect 9907 5593 9919 5596
rect 9861 5587 9919 5593
rect 3375 5528 4752 5556
rect 9784 5556 9812 5587
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 11256 5624 11284 5655
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 10612 5596 11284 5624
rect 15856 5624 15884 5655
rect 15930 5652 15936 5704
rect 15988 5692 15994 5704
rect 16025 5695 16083 5701
rect 16025 5692 16037 5695
rect 15988 5664 16037 5692
rect 15988 5652 15994 5664
rect 16025 5661 16037 5664
rect 16071 5692 16083 5695
rect 16224 5692 16252 5800
rect 16758 5720 16764 5772
rect 16816 5720 16822 5772
rect 16071 5664 16252 5692
rect 16301 5695 16359 5701
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 16301 5661 16313 5695
rect 16347 5661 16359 5695
rect 16301 5655 16359 5661
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5692 16543 5695
rect 16574 5692 16580 5704
rect 16531 5664 16580 5692
rect 16531 5661 16543 5664
rect 16485 5655 16543 5661
rect 16206 5624 16212 5636
rect 15856 5596 16212 5624
rect 10612 5565 10640 5596
rect 16206 5584 16212 5596
rect 16264 5584 16270 5636
rect 10597 5559 10655 5565
rect 10597 5556 10609 5559
rect 9784 5528 10609 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 10597 5525 10609 5528
rect 10643 5525 10655 5559
rect 14918 5556 14924 5568
rect 14879 5528 14924 5556
rect 10597 5519 10655 5525
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 16316 5556 16344 5655
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 16776 5692 16804 5720
rect 16853 5695 16911 5701
rect 16853 5692 16865 5695
rect 16776 5664 16865 5692
rect 16853 5661 16865 5664
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 17037 5695 17095 5701
rect 17037 5661 17049 5695
rect 17083 5692 17095 5695
rect 17313 5695 17371 5701
rect 17313 5692 17325 5695
rect 17083 5664 17325 5692
rect 17083 5661 17095 5664
rect 17037 5655 17095 5661
rect 17313 5661 17325 5664
rect 17359 5661 17371 5695
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17313 5655 17371 5661
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 17604 5692 17632 5800
rect 19702 5788 19708 5840
rect 19760 5828 19766 5840
rect 19760 5800 19805 5828
rect 19760 5788 19766 5800
rect 19886 5788 19892 5840
rect 19944 5828 19950 5840
rect 20346 5828 20352 5840
rect 19944 5800 20352 5828
rect 19944 5788 19950 5800
rect 20346 5788 20352 5800
rect 20404 5828 20410 5840
rect 20404 5800 20668 5828
rect 20404 5788 20410 5800
rect 17770 5760 17776 5772
rect 17731 5732 17776 5760
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 18969 5763 19027 5769
rect 18969 5760 18981 5763
rect 18380 5732 18981 5760
rect 18380 5720 18386 5732
rect 18969 5729 18981 5732
rect 19015 5729 19027 5763
rect 19334 5760 19340 5772
rect 19295 5732 19340 5760
rect 18969 5723 19027 5729
rect 17681 5695 17739 5701
rect 17681 5692 17693 5695
rect 17604 5664 17693 5692
rect 17681 5661 17693 5664
rect 17727 5661 17739 5695
rect 17681 5655 17739 5661
rect 17957 5695 18015 5701
rect 17957 5661 17969 5695
rect 18003 5661 18015 5695
rect 18141 5695 18199 5701
rect 18141 5688 18153 5695
rect 17957 5655 18015 5661
rect 18044 5661 18153 5688
rect 18187 5661 18199 5695
rect 18044 5660 18199 5661
rect 16669 5627 16727 5633
rect 16669 5593 16681 5627
rect 16715 5624 16727 5627
rect 16758 5624 16764 5636
rect 16715 5596 16764 5624
rect 16715 5593 16727 5596
rect 16669 5587 16727 5593
rect 16758 5584 16764 5596
rect 16816 5584 16822 5636
rect 17972 5624 18000 5655
rect 16960 5596 18000 5624
rect 18044 5624 18072 5660
rect 18141 5655 18199 5660
rect 18230 5652 18236 5704
rect 18288 5692 18294 5704
rect 18690 5692 18696 5704
rect 18288 5664 18552 5692
rect 18651 5664 18696 5692
rect 18288 5652 18294 5664
rect 18524 5624 18552 5664
rect 18690 5652 18696 5664
rect 18748 5652 18754 5704
rect 18984 5692 19012 5723
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 20530 5760 20536 5772
rect 19444 5732 19840 5760
rect 20491 5732 20536 5760
rect 19444 5692 19472 5732
rect 18984 5664 19472 5692
rect 19521 5695 19579 5701
rect 19521 5661 19533 5695
rect 19567 5692 19579 5695
rect 19610 5692 19616 5704
rect 19567 5664 19616 5692
rect 19567 5661 19579 5664
rect 19521 5655 19579 5661
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 19245 5627 19303 5633
rect 18044 5596 18368 5624
rect 18524 5596 18920 5624
rect 16960 5556 16988 5596
rect 17126 5556 17132 5568
rect 16316 5528 16988 5556
rect 17087 5528 17132 5556
rect 17126 5516 17132 5528
rect 17184 5516 17190 5568
rect 17972 5556 18000 5596
rect 18230 5556 18236 5568
rect 17972 5528 18236 5556
rect 18230 5516 18236 5528
rect 18288 5516 18294 5568
rect 18340 5565 18368 5596
rect 18325 5559 18383 5565
rect 18325 5525 18337 5559
rect 18371 5525 18383 5559
rect 18782 5556 18788 5568
rect 18743 5528 18788 5556
rect 18325 5519 18383 5525
rect 18782 5516 18788 5528
rect 18840 5516 18846 5568
rect 18892 5556 18920 5596
rect 19245 5593 19257 5627
rect 19291 5624 19303 5627
rect 19702 5624 19708 5636
rect 19291 5596 19708 5624
rect 19291 5593 19303 5596
rect 19245 5587 19303 5593
rect 19702 5584 19708 5596
rect 19760 5584 19766 5636
rect 19812 5624 19840 5732
rect 20530 5720 20536 5732
rect 20588 5720 20594 5772
rect 20640 5760 20668 5800
rect 21637 5763 21695 5769
rect 21637 5760 21649 5763
rect 20640 5732 20760 5760
rect 19978 5652 19984 5704
rect 20036 5692 20042 5704
rect 20073 5695 20131 5701
rect 20073 5692 20085 5695
rect 20036 5664 20085 5692
rect 20036 5652 20042 5664
rect 20073 5661 20085 5664
rect 20119 5661 20131 5695
rect 20073 5655 20131 5661
rect 20165 5695 20223 5701
rect 20165 5661 20177 5695
rect 20211 5692 20223 5695
rect 20441 5695 20499 5701
rect 20211 5664 20392 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 20364 5624 20392 5664
rect 20441 5661 20453 5695
rect 20487 5692 20499 5695
rect 20622 5692 20628 5704
rect 20487 5664 20628 5692
rect 20487 5661 20499 5664
rect 20441 5655 20499 5661
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 20732 5701 20760 5732
rect 21008 5732 21649 5760
rect 20717 5695 20775 5701
rect 20717 5661 20729 5695
rect 20763 5661 20775 5695
rect 20898 5692 20904 5704
rect 20859 5664 20904 5692
rect 20717 5655 20775 5661
rect 20898 5652 20904 5664
rect 20956 5652 20962 5704
rect 20806 5624 20812 5636
rect 19812 5596 19932 5624
rect 20364 5596 20812 5624
rect 19794 5556 19800 5568
rect 18892 5528 19800 5556
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 19904 5565 19932 5596
rect 20806 5584 20812 5596
rect 20864 5584 20870 5636
rect 21008 5624 21036 5732
rect 21637 5729 21649 5732
rect 21683 5729 21695 5763
rect 21637 5723 21695 5729
rect 21174 5652 21180 5704
rect 21232 5692 21238 5704
rect 21453 5695 21511 5701
rect 21453 5692 21465 5695
rect 21232 5664 21465 5692
rect 21232 5652 21238 5664
rect 21453 5661 21465 5664
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 21542 5652 21548 5704
rect 21600 5692 21606 5704
rect 21913 5695 21971 5701
rect 21913 5692 21925 5695
rect 21600 5664 21925 5692
rect 21600 5652 21606 5664
rect 21913 5661 21925 5664
rect 21959 5661 21971 5695
rect 21913 5655 21971 5661
rect 22094 5652 22100 5704
rect 22152 5692 22158 5704
rect 22189 5695 22247 5701
rect 22189 5692 22201 5695
rect 22152 5664 22201 5692
rect 22152 5652 22158 5664
rect 22189 5661 22201 5664
rect 22235 5661 22247 5695
rect 22189 5655 22247 5661
rect 22465 5695 22523 5701
rect 22465 5661 22477 5695
rect 22511 5692 22523 5695
rect 23198 5692 23204 5704
rect 22511 5664 23204 5692
rect 22511 5661 22523 5664
rect 22465 5655 22523 5661
rect 22940 5636 22968 5664
rect 23198 5652 23204 5664
rect 23256 5652 23262 5704
rect 23860 5692 23888 5859
rect 24394 5856 24400 5908
rect 24452 5896 24458 5908
rect 24949 5899 25007 5905
rect 24949 5896 24961 5899
rect 24452 5868 24961 5896
rect 24452 5856 24458 5868
rect 24949 5865 24961 5868
rect 24995 5896 25007 5899
rect 25958 5896 25964 5908
rect 24995 5868 25452 5896
rect 25919 5868 25964 5896
rect 24995 5865 25007 5868
rect 24949 5859 25007 5865
rect 24688 5800 25176 5828
rect 24688 5701 24716 5800
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 23860 5664 24685 5692
rect 24673 5661 24685 5664
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 24765 5695 24823 5701
rect 24765 5661 24777 5695
rect 24811 5661 24823 5695
rect 24765 5655 24823 5661
rect 20916 5596 21036 5624
rect 22732 5627 22790 5633
rect 19889 5559 19947 5565
rect 19889 5525 19901 5559
rect 19935 5525 19947 5559
rect 19889 5519 19947 5525
rect 20438 5516 20444 5568
rect 20496 5556 20502 5568
rect 20916 5556 20944 5596
rect 22732 5593 22744 5627
rect 22778 5624 22790 5627
rect 22830 5624 22836 5636
rect 22778 5596 22836 5624
rect 22778 5593 22790 5596
rect 22732 5587 22790 5593
rect 22830 5584 22836 5596
rect 22888 5584 22894 5636
rect 22922 5584 22928 5636
rect 22980 5584 22986 5636
rect 24780 5624 24808 5655
rect 24854 5652 24860 5704
rect 24912 5692 24918 5704
rect 25148 5701 25176 5800
rect 25424 5701 25452 5868
rect 25958 5856 25964 5868
rect 26016 5856 26022 5908
rect 26418 5760 26424 5772
rect 26379 5732 26424 5760
rect 26418 5720 26424 5732
rect 26476 5720 26482 5772
rect 26605 5763 26663 5769
rect 26605 5729 26617 5763
rect 26651 5760 26663 5763
rect 27522 5760 27528 5772
rect 26651 5732 27528 5760
rect 26651 5729 26663 5732
rect 26605 5723 26663 5729
rect 27522 5720 27528 5732
rect 27580 5720 27586 5772
rect 25041 5695 25099 5701
rect 25041 5692 25053 5695
rect 24912 5664 25053 5692
rect 24912 5652 24918 5664
rect 25041 5661 25053 5664
rect 25087 5661 25099 5695
rect 25041 5655 25099 5661
rect 25133 5695 25191 5701
rect 25133 5661 25145 5695
rect 25179 5661 25191 5695
rect 25133 5655 25191 5661
rect 25409 5695 25467 5701
rect 25409 5661 25421 5695
rect 25455 5661 25467 5695
rect 25409 5655 25467 5661
rect 26973 5695 27031 5701
rect 26973 5661 26985 5695
rect 27019 5692 27031 5695
rect 27154 5692 27160 5704
rect 27019 5664 27160 5692
rect 27019 5661 27031 5664
rect 26973 5655 27031 5661
rect 27154 5652 27160 5664
rect 27212 5652 27218 5704
rect 25501 5627 25559 5633
rect 25501 5624 25513 5627
rect 24780 5596 25513 5624
rect 25501 5593 25513 5596
rect 25547 5593 25559 5627
rect 25501 5587 25559 5593
rect 26329 5627 26387 5633
rect 26329 5593 26341 5627
rect 26375 5624 26387 5627
rect 26881 5627 26939 5633
rect 26881 5624 26893 5627
rect 26375 5596 26893 5624
rect 26375 5593 26387 5596
rect 26329 5587 26387 5593
rect 26881 5593 26893 5596
rect 26927 5593 26939 5627
rect 26881 5587 26939 5593
rect 21082 5556 21088 5568
rect 20496 5528 20944 5556
rect 21043 5528 21088 5556
rect 20496 5516 20502 5528
rect 21082 5516 21088 5528
rect 21140 5516 21146 5568
rect 21358 5516 21364 5568
rect 21416 5556 21422 5568
rect 21545 5559 21603 5565
rect 21545 5556 21557 5559
rect 21416 5528 21557 5556
rect 21416 5516 21422 5528
rect 21545 5525 21557 5528
rect 21591 5556 21603 5559
rect 21910 5556 21916 5568
rect 21591 5528 21916 5556
rect 21591 5525 21603 5528
rect 21545 5519 21603 5525
rect 21910 5516 21916 5528
rect 21968 5556 21974 5568
rect 22005 5559 22063 5565
rect 22005 5556 22017 5559
rect 21968 5528 22017 5556
rect 21968 5516 21974 5528
rect 22005 5525 22017 5528
rect 22051 5525 22063 5559
rect 22370 5556 22376 5568
rect 22331 5528 22376 5556
rect 22005 5519 22063 5525
rect 22370 5516 22376 5528
rect 22428 5516 22434 5568
rect 24486 5556 24492 5568
rect 24447 5528 24492 5556
rect 24486 5516 24492 5528
rect 24544 5516 24550 5568
rect 24762 5516 24768 5568
rect 24820 5556 24826 5568
rect 25225 5559 25283 5565
rect 25225 5556 25237 5559
rect 24820 5528 25237 5556
rect 24820 5516 24826 5528
rect 25225 5525 25237 5528
rect 25271 5525 25283 5559
rect 25225 5519 25283 5525
rect 1104 5466 29532 5488
rect 1104 5414 10425 5466
rect 10477 5414 10489 5466
rect 10541 5414 10553 5466
rect 10605 5414 10617 5466
rect 10669 5414 10681 5466
rect 10733 5414 19901 5466
rect 19953 5414 19965 5466
rect 20017 5414 20029 5466
rect 20081 5414 20093 5466
rect 20145 5414 20157 5466
rect 20209 5414 29532 5466
rect 1104 5392 29532 5414
rect 3329 5355 3387 5361
rect 3329 5321 3341 5355
rect 3375 5352 3387 5355
rect 3418 5352 3424 5364
rect 3375 5324 3424 5352
rect 3375 5321 3387 5324
rect 3329 5315 3387 5321
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 8389 5355 8447 5361
rect 8389 5352 8401 5355
rect 8220 5324 8401 5352
rect 2222 5293 2228 5296
rect 2216 5284 2228 5293
rect 2183 5256 2228 5284
rect 2216 5247 2228 5256
rect 2222 5244 2228 5247
rect 2280 5244 2286 5296
rect 6362 5284 6368 5296
rect 6323 5256 6368 5284
rect 6362 5244 6368 5256
rect 6420 5244 6426 5296
rect 8052 5287 8110 5293
rect 8052 5253 8064 5287
rect 8098 5284 8110 5287
rect 8220 5284 8248 5324
rect 8389 5321 8401 5324
rect 8435 5321 8447 5355
rect 8846 5352 8852 5364
rect 8807 5324 8852 5352
rect 8389 5315 8447 5321
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 9214 5312 9220 5364
rect 9272 5352 9278 5364
rect 10226 5352 10232 5364
rect 9272 5324 9812 5352
rect 10187 5324 10232 5352
rect 9272 5312 9278 5324
rect 8098 5256 8248 5284
rect 8098 5253 8110 5256
rect 8052 5247 8110 5253
rect 1394 5176 1400 5228
rect 1452 5216 1458 5228
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1452 5188 1961 5216
rect 1452 5176 1458 5188
rect 1949 5185 1961 5188
rect 1995 5216 2007 5219
rect 4062 5216 4068 5228
rect 1995 5188 4068 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4430 5216 4436 5228
rect 4387 5188 4436 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4430 5176 4436 5188
rect 4488 5216 4494 5228
rect 4982 5216 4988 5228
rect 4488 5188 4844 5216
rect 4943 5188 4988 5216
rect 4488 5176 4494 5188
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5117 4583 5151
rect 4525 5111 4583 5117
rect 3786 4972 3792 5024
rect 3844 5012 3850 5024
rect 4157 5015 4215 5021
rect 4157 5012 4169 5015
rect 3844 4984 4169 5012
rect 3844 4972 3850 4984
rect 4157 4981 4169 4984
rect 4203 4981 4215 5015
rect 4540 5012 4568 5111
rect 4816 5089 4844 5188
rect 4982 5176 4988 5188
rect 5040 5176 5046 5228
rect 6546 5216 6552 5228
rect 6507 5188 6552 5216
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8260 5188 8769 5216
rect 8260 5176 8266 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 9217 5219 9275 5225
rect 9217 5185 9229 5219
rect 9263 5216 9275 5219
rect 9490 5216 9496 5228
rect 9263 5188 9496 5216
rect 9263 5185 9275 5188
rect 9217 5179 9275 5185
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 9784 5225 9812 5324
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 11977 5355 12035 5361
rect 11977 5321 11989 5355
rect 12023 5352 12035 5355
rect 12345 5355 12403 5361
rect 12345 5352 12357 5355
rect 12023 5324 12357 5352
rect 12023 5321 12035 5324
rect 11977 5315 12035 5321
rect 12345 5321 12357 5324
rect 12391 5321 12403 5355
rect 12345 5315 12403 5321
rect 15749 5355 15807 5361
rect 15749 5321 15761 5355
rect 15795 5352 15807 5355
rect 16114 5352 16120 5364
rect 15795 5324 16120 5352
rect 15795 5321 15807 5324
rect 15749 5315 15807 5321
rect 16114 5312 16120 5324
rect 16172 5312 16178 5364
rect 16574 5312 16580 5364
rect 16632 5352 16638 5364
rect 16669 5355 16727 5361
rect 16669 5352 16681 5355
rect 16632 5324 16681 5352
rect 16632 5312 16638 5324
rect 16669 5321 16681 5324
rect 16715 5321 16727 5355
rect 17126 5352 17132 5364
rect 17087 5324 17132 5352
rect 16669 5315 16727 5321
rect 17126 5312 17132 5324
rect 17184 5312 17190 5364
rect 17770 5312 17776 5364
rect 17828 5352 17834 5364
rect 17957 5355 18015 5361
rect 17957 5352 17969 5355
rect 17828 5324 17969 5352
rect 17828 5312 17834 5324
rect 17957 5321 17969 5324
rect 18003 5321 18015 5355
rect 17957 5315 18015 5321
rect 18785 5355 18843 5361
rect 18785 5321 18797 5355
rect 18831 5352 18843 5355
rect 19242 5352 19248 5364
rect 18831 5324 19248 5352
rect 18831 5321 18843 5324
rect 18785 5315 18843 5321
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 20165 5355 20223 5361
rect 20165 5321 20177 5355
rect 20211 5352 20223 5355
rect 20530 5352 20536 5364
rect 20211 5324 20536 5352
rect 20211 5321 20223 5324
rect 20165 5315 20223 5321
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 20898 5312 20904 5364
rect 20956 5352 20962 5364
rect 21821 5355 21879 5361
rect 21821 5352 21833 5355
rect 20956 5324 21833 5352
rect 20956 5312 20962 5324
rect 21821 5321 21833 5324
rect 21867 5321 21879 5355
rect 21821 5315 21879 5321
rect 22281 5355 22339 5361
rect 22281 5321 22293 5355
rect 22327 5352 22339 5355
rect 22370 5352 22376 5364
rect 22327 5324 22376 5352
rect 22327 5321 22339 5324
rect 22281 5315 22339 5321
rect 22370 5312 22376 5324
rect 22428 5312 22434 5364
rect 22830 5312 22836 5364
rect 22888 5352 22894 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22888 5324 23029 5352
rect 22888 5312 22894 5324
rect 23017 5321 23029 5324
rect 23063 5321 23075 5355
rect 23474 5352 23480 5364
rect 23435 5324 23480 5352
rect 23017 5315 23075 5321
rect 23474 5312 23480 5324
rect 23532 5312 23538 5364
rect 11241 5287 11299 5293
rect 11241 5253 11253 5287
rect 11287 5284 11299 5287
rect 15841 5287 15899 5293
rect 11287 5256 12434 5284
rect 11287 5253 11299 5256
rect 11241 5247 11299 5253
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5216 9827 5219
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9815 5188 9873 5216
rect 9815 5185 9827 5188
rect 9769 5179 9827 5185
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 8297 5151 8355 5157
rect 8297 5117 8309 5151
rect 8343 5148 8355 5151
rect 8386 5148 8392 5160
rect 8343 5120 8392 5148
rect 8343 5117 8355 5120
rect 8297 5111 8355 5117
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 8938 5148 8944 5160
rect 8720 5120 8944 5148
rect 8720 5108 8726 5120
rect 8938 5108 8944 5120
rect 8996 5108 9002 5160
rect 9600 5148 9628 5179
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10870 5216 10876 5228
rect 10192 5188 10876 5216
rect 10192 5176 10198 5188
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11054 5216 11060 5228
rect 10967 5188 11060 5216
rect 11054 5176 11060 5188
rect 11112 5216 11118 5228
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11112 5188 11897 5216
rect 11112 5176 11118 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 12406 5216 12434 5256
rect 15841 5253 15853 5287
rect 15887 5284 15899 5287
rect 16301 5287 16359 5293
rect 16301 5284 16313 5287
rect 15887 5256 16313 5284
rect 15887 5253 15899 5256
rect 15841 5247 15899 5253
rect 16301 5253 16313 5256
rect 16347 5284 16359 5287
rect 19337 5287 19395 5293
rect 16347 5256 18460 5284
rect 16347 5253 16359 5256
rect 16301 5247 16359 5253
rect 12529 5219 12587 5225
rect 12529 5216 12541 5219
rect 12406 5188 12541 5216
rect 11885 5179 11943 5185
rect 12529 5185 12541 5188
rect 12575 5185 12587 5219
rect 16206 5216 16212 5228
rect 16119 5188 16212 5216
rect 12529 5179 12587 5185
rect 16206 5176 16212 5188
rect 16264 5216 16270 5228
rect 16758 5216 16764 5228
rect 16264 5188 16764 5216
rect 16264 5176 16270 5188
rect 16758 5176 16764 5188
rect 16816 5216 16822 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16816 5188 17049 5216
rect 16816 5176 16822 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 17678 5216 17684 5228
rect 17037 5179 17095 5185
rect 17236 5188 17684 5216
rect 9950 5148 9956 5160
rect 9600 5120 9956 5148
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 10318 5108 10324 5160
rect 10376 5148 10382 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 10376 5120 12081 5148
rect 10376 5108 10382 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 15562 5108 15568 5160
rect 15620 5148 15626 5160
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15620 5120 16037 5148
rect 15620 5108 15626 5120
rect 16025 5117 16037 5120
rect 16071 5148 16083 5151
rect 17236 5148 17264 5188
rect 17678 5176 17684 5188
rect 17736 5216 17742 5228
rect 18432 5225 18460 5256
rect 19337 5253 19349 5287
rect 19383 5284 19395 5287
rect 19426 5284 19432 5296
rect 19383 5256 19432 5284
rect 19383 5253 19395 5256
rect 19337 5247 19395 5253
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 19702 5244 19708 5296
rect 19760 5284 19766 5296
rect 20257 5287 20315 5293
rect 20257 5284 20269 5287
rect 19760 5256 20269 5284
rect 19760 5244 19766 5256
rect 20257 5253 20269 5256
rect 20303 5284 20315 5287
rect 20717 5287 20775 5293
rect 20717 5284 20729 5287
rect 20303 5256 20729 5284
rect 20303 5253 20315 5256
rect 20257 5247 20315 5253
rect 20717 5253 20729 5256
rect 20763 5253 20775 5287
rect 21637 5287 21695 5293
rect 20717 5247 20775 5253
rect 21284 5256 21588 5284
rect 18417 5219 18475 5225
rect 17736 5188 18276 5216
rect 17736 5176 17742 5188
rect 16071 5120 17264 5148
rect 17313 5151 17371 5157
rect 16071 5117 16083 5120
rect 16025 5111 16083 5117
rect 17313 5117 17325 5151
rect 17359 5148 17371 5151
rect 17402 5148 17408 5160
rect 17359 5120 17408 5148
rect 17359 5117 17371 5120
rect 17313 5111 17371 5117
rect 17402 5108 17408 5120
rect 17460 5108 17466 5160
rect 18248 5157 18276 5188
rect 18417 5185 18429 5219
rect 18463 5185 18475 5219
rect 18417 5179 18475 5185
rect 18601 5219 18659 5225
rect 18601 5185 18613 5219
rect 18647 5216 18659 5219
rect 20806 5216 20812 5228
rect 18647 5188 20668 5216
rect 20767 5188 20812 5216
rect 18647 5185 18659 5188
rect 18601 5179 18659 5185
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 18233 5151 18291 5157
rect 18233 5117 18245 5151
rect 18279 5117 18291 5151
rect 19426 5148 19432 5160
rect 19387 5120 19432 5148
rect 18233 5111 18291 5117
rect 4801 5083 4859 5089
rect 4801 5049 4813 5083
rect 4847 5049 4859 5083
rect 7006 5080 7012 5092
rect 4801 5043 4859 5049
rect 4908 5052 7012 5080
rect 4908 5024 4936 5052
rect 7006 5040 7012 5052
rect 7064 5040 7070 5092
rect 9309 5083 9367 5089
rect 9309 5049 9321 5083
rect 9355 5049 9367 5083
rect 9309 5043 9367 5049
rect 4890 5012 4896 5024
rect 4540 4984 4896 5012
rect 4157 4975 4215 4981
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 6641 5015 6699 5021
rect 6641 5012 6653 5015
rect 6144 4984 6653 5012
rect 6144 4972 6150 4984
rect 6641 4981 6653 4984
rect 6687 4981 6699 5015
rect 6914 5012 6920 5024
rect 6875 4984 6920 5012
rect 6641 4975 6699 4981
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 8110 4972 8116 5024
rect 8168 5012 8174 5024
rect 9324 5012 9352 5043
rect 9398 5040 9404 5092
rect 9456 5080 9462 5092
rect 17034 5080 17040 5092
rect 9456 5052 17040 5080
rect 9456 5040 9462 5052
rect 17034 5040 17040 5052
rect 17092 5040 17098 5092
rect 18064 5024 18092 5111
rect 18248 5080 18276 5111
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 19613 5151 19671 5157
rect 19613 5117 19625 5151
rect 19659 5148 19671 5151
rect 20438 5148 20444 5160
rect 19659 5120 20444 5148
rect 19659 5117 19671 5120
rect 19613 5111 19671 5117
rect 18248 5052 19196 5080
rect 9858 5012 9864 5024
rect 8168 4984 9352 5012
rect 9819 4984 9864 5012
rect 8168 4972 8174 4984
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 11514 5012 11520 5024
rect 11475 4984 11520 5012
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 15381 5015 15439 5021
rect 15381 4981 15393 5015
rect 15427 5012 15439 5015
rect 15562 5012 15568 5024
rect 15427 4984 15568 5012
rect 15427 4981 15439 4984
rect 15381 4975 15439 4981
rect 15562 4972 15568 4984
rect 15620 4972 15626 5024
rect 17494 4972 17500 5024
rect 17552 5012 17558 5024
rect 17589 5015 17647 5021
rect 17589 5012 17601 5015
rect 17552 4984 17601 5012
rect 17552 4972 17558 4984
rect 17589 4981 17601 4984
rect 17635 4981 17647 5015
rect 18046 5012 18052 5024
rect 17959 4984 18052 5012
rect 17589 4975 17647 4981
rect 18046 4972 18052 4984
rect 18104 5012 18110 5024
rect 18417 5015 18475 5021
rect 18417 5012 18429 5015
rect 18104 4984 18429 5012
rect 18104 4972 18110 4984
rect 18417 4981 18429 4984
rect 18463 4981 18475 5015
rect 18417 4975 18475 4981
rect 18969 5015 19027 5021
rect 18969 4981 18981 5015
rect 19015 5012 19027 5015
rect 19058 5012 19064 5024
rect 19015 4984 19064 5012
rect 19015 4981 19027 4984
rect 18969 4975 19027 4981
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 19168 5012 19196 5052
rect 19628 5012 19656 5111
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 20640 5148 20668 5188
rect 20806 5176 20812 5188
rect 20864 5216 20870 5228
rect 21174 5216 21180 5228
rect 20864 5188 21180 5216
rect 20864 5176 20870 5188
rect 21174 5176 21180 5188
rect 21232 5216 21238 5228
rect 21284 5225 21312 5256
rect 21269 5219 21327 5225
rect 21269 5216 21281 5219
rect 21232 5188 21281 5216
rect 21232 5176 21238 5188
rect 21269 5185 21281 5188
rect 21315 5185 21327 5219
rect 21269 5179 21327 5185
rect 21453 5219 21511 5225
rect 21453 5185 21465 5219
rect 21499 5185 21511 5219
rect 21560 5216 21588 5256
rect 21637 5253 21649 5287
rect 21683 5284 21695 5287
rect 22094 5284 22100 5296
rect 21683 5256 22100 5284
rect 21683 5253 21695 5256
rect 21637 5247 21695 5253
rect 22094 5244 22100 5256
rect 22152 5244 22158 5296
rect 23385 5287 23443 5293
rect 23385 5253 23397 5287
rect 23431 5284 23443 5287
rect 24762 5284 24768 5296
rect 23431 5256 24768 5284
rect 23431 5253 23443 5256
rect 23385 5247 23443 5253
rect 24762 5244 24768 5256
rect 24820 5244 24826 5296
rect 22189 5219 22247 5225
rect 22189 5216 22201 5219
rect 21560 5188 22201 5216
rect 21453 5179 21511 5185
rect 22189 5185 22201 5188
rect 22235 5185 22247 5219
rect 22189 5179 22247 5185
rect 21358 5148 21364 5160
rect 20640 5120 21364 5148
rect 21358 5108 21364 5120
rect 21416 5108 21422 5160
rect 21468 5080 21496 5179
rect 23934 5176 23940 5228
rect 23992 5216 23998 5228
rect 25409 5219 25467 5225
rect 25409 5216 25421 5219
rect 23992 5188 25421 5216
rect 23992 5176 23998 5188
rect 25409 5185 25421 5188
rect 25455 5185 25467 5219
rect 25409 5179 25467 5185
rect 25685 5219 25743 5225
rect 25685 5185 25697 5219
rect 25731 5216 25743 5219
rect 26053 5219 26111 5225
rect 26053 5216 26065 5219
rect 25731 5188 26065 5216
rect 25731 5185 25743 5188
rect 25685 5179 25743 5185
rect 26053 5185 26065 5188
rect 26099 5216 26111 5219
rect 28166 5216 28172 5228
rect 26099 5188 28172 5216
rect 26099 5185 26111 5188
rect 26053 5179 26111 5185
rect 28166 5176 28172 5188
rect 28224 5176 28230 5228
rect 21818 5108 21824 5160
rect 21876 5148 21882 5160
rect 22373 5151 22431 5157
rect 22373 5148 22385 5151
rect 21876 5120 22385 5148
rect 21876 5108 21882 5120
rect 22373 5117 22385 5120
rect 22419 5117 22431 5151
rect 22373 5111 22431 5117
rect 23382 5108 23388 5160
rect 23440 5148 23446 5160
rect 23569 5151 23627 5157
rect 23569 5148 23581 5151
rect 23440 5120 23581 5148
rect 23440 5108 23446 5120
rect 23569 5117 23581 5120
rect 23615 5117 23627 5151
rect 23569 5111 23627 5117
rect 22002 5080 22008 5092
rect 21468 5052 22008 5080
rect 22002 5040 22008 5052
rect 22060 5080 22066 5092
rect 23934 5080 23940 5092
rect 22060 5052 23940 5080
rect 22060 5040 22066 5052
rect 23934 5040 23940 5052
rect 23992 5040 23998 5092
rect 25406 5040 25412 5092
rect 25464 5080 25470 5092
rect 25685 5083 25743 5089
rect 25685 5080 25697 5083
rect 25464 5052 25697 5080
rect 25464 5040 25470 5052
rect 25685 5049 25697 5052
rect 25731 5049 25743 5083
rect 25685 5043 25743 5049
rect 19794 5012 19800 5024
rect 19168 4984 19656 5012
rect 19755 4984 19800 5012
rect 19794 4972 19800 4984
rect 19852 4972 19858 5024
rect 25498 4972 25504 5024
rect 25556 5012 25562 5024
rect 25961 5015 26019 5021
rect 25961 5012 25973 5015
rect 25556 4984 25973 5012
rect 25556 4972 25562 4984
rect 25961 4981 25973 4984
rect 26007 4981 26019 5015
rect 25961 4975 26019 4981
rect 1104 4922 29532 4944
rect 1104 4870 5688 4922
rect 5740 4870 5752 4922
rect 5804 4870 5816 4922
rect 5868 4870 5880 4922
rect 5932 4870 5944 4922
rect 5996 4870 15163 4922
rect 15215 4870 15227 4922
rect 15279 4870 15291 4922
rect 15343 4870 15355 4922
rect 15407 4870 15419 4922
rect 15471 4870 24639 4922
rect 24691 4870 24703 4922
rect 24755 4870 24767 4922
rect 24819 4870 24831 4922
rect 24883 4870 24895 4922
rect 24947 4870 29532 4922
rect 1104 4848 29532 4870
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5721 4811 5779 4817
rect 5721 4808 5733 4811
rect 5040 4780 5733 4808
rect 5040 4768 5046 4780
rect 5721 4777 5733 4780
rect 5767 4777 5779 4811
rect 5721 4771 5779 4777
rect 6733 4811 6791 4817
rect 6733 4777 6745 4811
rect 6779 4777 6791 4811
rect 6733 4771 6791 4777
rect 6917 4811 6975 4817
rect 6917 4777 6929 4811
rect 6963 4808 6975 4811
rect 7282 4808 7288 4820
rect 6963 4780 7288 4808
rect 6963 4777 6975 4780
rect 6917 4771 6975 4777
rect 5445 4743 5503 4749
rect 5445 4709 5457 4743
rect 5491 4740 5503 4743
rect 6748 4740 6776 4771
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 8202 4808 8208 4820
rect 8163 4780 8208 4808
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 9858 4808 9864 4820
rect 8864 4780 9864 4808
rect 8864 4740 8892 4780
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10597 4811 10655 4817
rect 10597 4777 10609 4811
rect 10643 4777 10655 4811
rect 11054 4808 11060 4820
rect 11015 4780 11060 4808
rect 10597 4771 10655 4777
rect 9950 4740 9956 4752
rect 5491 4712 6224 4740
rect 6748 4712 8892 4740
rect 8956 4712 9956 4740
rect 5491 4709 5503 4712
rect 5445 4703 5503 4709
rect 3786 4604 3792 4616
rect 3747 4576 3792 4604
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 4062 4604 4068 4616
rect 4023 4576 4068 4604
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 5871 4607 5929 4613
rect 4264 4576 4660 4604
rect 3878 4496 3884 4548
rect 3936 4536 3942 4548
rect 4264 4536 4292 4576
rect 4338 4545 4344 4548
rect 3936 4508 4292 4536
rect 3936 4496 3942 4508
rect 4332 4499 4344 4545
rect 4396 4536 4402 4548
rect 4396 4508 4432 4536
rect 4338 4496 4344 4499
rect 4396 4496 4402 4508
rect 3973 4471 4031 4477
rect 3973 4437 3985 4471
rect 4019 4468 4031 4471
rect 4522 4468 4528 4480
rect 4019 4440 4528 4468
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 4632 4468 4660 4576
rect 5871 4573 5883 4607
rect 5917 4604 5929 4607
rect 6086 4604 6092 4616
rect 5917 4576 6092 4604
rect 5917 4573 5929 4576
rect 5871 4567 5929 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 6196 4613 6224 4712
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 6362 4672 6368 4684
rect 6319 4644 6368 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 6546 4672 6552 4684
rect 6507 4644 6552 4672
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 8956 4672 8984 4712
rect 9950 4700 9956 4712
rect 10008 4700 10014 4752
rect 10612 4740 10640 4771
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 18046 4808 18052 4820
rect 18007 4780 18052 4808
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 21174 4808 21180 4820
rect 21135 4780 21180 4808
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 21542 4768 21548 4820
rect 21600 4808 21606 4820
rect 21821 4811 21879 4817
rect 21821 4808 21833 4811
rect 21600 4780 21833 4808
rect 21600 4768 21606 4780
rect 21821 4777 21833 4780
rect 21867 4777 21879 4811
rect 27522 4808 27528 4820
rect 21821 4771 21879 4777
rect 22066 4780 27528 4808
rect 10962 4740 10968 4752
rect 10612 4712 10968 4740
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 20346 4700 20352 4752
rect 20404 4740 20410 4752
rect 22066 4740 22094 4780
rect 27522 4768 27528 4780
rect 27580 4768 27586 4820
rect 28166 4808 28172 4820
rect 28127 4780 28172 4808
rect 28166 4768 28172 4780
rect 28224 4768 28230 4820
rect 20404 4712 22094 4740
rect 20404 4700 20410 4712
rect 6932 4644 8984 4672
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4604 6239 4607
rect 6564 4604 6592 4632
rect 6932 4616 6960 4644
rect 6227 4576 6592 4604
rect 6733 4607 6791 4613
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 6733 4573 6745 4607
rect 6779 4604 6791 4607
rect 6914 4604 6920 4616
rect 6779 4576 6920 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 6914 4564 6920 4576
rect 6972 4564 6978 4616
rect 8110 4604 8116 4616
rect 8071 4576 8116 4604
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8956 4613 8984 4644
rect 9309 4675 9367 4681
rect 9309 4641 9321 4675
rect 9355 4672 9367 4675
rect 9490 4672 9496 4684
rect 9355 4644 9496 4672
rect 9355 4641 9367 4644
rect 9309 4635 9367 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 12894 4672 12900 4684
rect 12855 4644 12900 4672
rect 12894 4632 12900 4644
rect 12952 4632 12958 4684
rect 22370 4672 22376 4684
rect 22331 4644 22376 4672
rect 22370 4632 22376 4644
rect 22428 4632 22434 4684
rect 23382 4632 23388 4684
rect 23440 4672 23446 4684
rect 25225 4675 25283 4681
rect 25225 4672 25237 4675
rect 23440 4644 25237 4672
rect 23440 4632 23446 4644
rect 25225 4641 25237 4644
rect 25271 4641 25283 4675
rect 25225 4635 25283 4641
rect 25314 4632 25320 4684
rect 25372 4672 25378 4684
rect 25961 4675 26019 4681
rect 25961 4672 25973 4675
rect 25372 4644 25973 4672
rect 25372 4632 25378 4644
rect 25961 4641 25973 4644
rect 26007 4641 26019 4675
rect 25961 4635 26019 4641
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4573 8999 4607
rect 9214 4604 9220 4616
rect 9175 4576 9220 4604
rect 8941 4567 8999 4573
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 10042 4564 10048 4616
rect 10100 4604 10106 4616
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 10100 4576 10425 4604
rect 10100 4564 10106 4576
rect 10413 4573 10425 4576
rect 10459 4573 10471 4607
rect 10413 4567 10471 4573
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10870 4604 10876 4616
rect 10831 4576 10876 4604
rect 10597 4567 10655 4573
rect 6454 4536 6460 4548
rect 6415 4508 6460 4536
rect 6454 4496 6460 4508
rect 6512 4496 6518 4548
rect 10612 4536 10640 4567
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 11514 4564 11520 4616
rect 11572 4604 11578 4616
rect 12630 4607 12688 4613
rect 12630 4604 12642 4607
rect 11572 4576 12642 4604
rect 11572 4564 11578 4576
rect 12630 4573 12642 4576
rect 12676 4573 12688 4607
rect 15930 4604 15936 4616
rect 15891 4576 15936 4604
rect 12630 4567 12688 4573
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 18138 4604 18144 4616
rect 18099 4576 18144 4604
rect 18138 4564 18144 4576
rect 18196 4564 18202 4616
rect 21358 4604 21364 4616
rect 21319 4576 21364 4604
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 23934 4604 23940 4616
rect 23895 4576 23940 4604
rect 23934 4564 23940 4576
rect 23992 4564 23998 4616
rect 24397 4607 24455 4613
rect 24397 4573 24409 4607
rect 24443 4604 24455 4607
rect 24486 4604 24492 4616
rect 24443 4576 24492 4604
rect 24443 4573 24455 4576
rect 24397 4567 24455 4573
rect 24486 4564 24492 4576
rect 24544 4564 24550 4616
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4604 24823 4607
rect 25041 4607 25099 4613
rect 25041 4604 25053 4607
rect 24811 4576 25053 4604
rect 24811 4573 24823 4576
rect 24765 4567 24823 4573
rect 25041 4573 25053 4576
rect 25087 4573 25099 4607
rect 25406 4604 25412 4616
rect 25367 4576 25412 4604
rect 25041 4567 25099 4573
rect 25406 4564 25412 4576
rect 25464 4564 25470 4616
rect 25498 4564 25504 4616
rect 25556 4604 25562 4616
rect 25556 4576 25601 4604
rect 25556 4564 25562 4576
rect 27246 4564 27252 4616
rect 27304 4604 27310 4616
rect 27617 4607 27675 4613
rect 27617 4604 27629 4607
rect 27304 4576 27629 4604
rect 27304 4564 27310 4576
rect 27617 4573 27629 4576
rect 27663 4604 27675 4607
rect 27893 4607 27951 4613
rect 27893 4604 27905 4607
rect 27663 4576 27905 4604
rect 27663 4573 27675 4576
rect 27617 4567 27675 4573
rect 27893 4573 27905 4576
rect 27939 4573 27951 4607
rect 28005 4607 28063 4613
rect 28005 4604 28017 4607
rect 27893 4567 27951 4573
rect 28000 4573 28017 4604
rect 28051 4573 28063 4607
rect 28000 4567 28063 4573
rect 10778 4536 10784 4548
rect 10612 4508 10784 4536
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 22189 4539 22247 4545
rect 22189 4505 22201 4539
rect 22235 4536 22247 4539
rect 22646 4536 22652 4548
rect 22235 4508 22652 4536
rect 22235 4505 22247 4508
rect 22189 4499 22247 4505
rect 22646 4496 22652 4508
rect 22704 4496 22710 4548
rect 23750 4536 23756 4548
rect 23711 4508 23756 4536
rect 23750 4496 23756 4508
rect 23808 4496 23814 4548
rect 24121 4539 24179 4545
rect 24121 4505 24133 4539
rect 24167 4505 24179 4539
rect 24578 4536 24584 4548
rect 24539 4508 24584 4536
rect 24121 4499 24179 4505
rect 9398 4468 9404 4480
rect 4632 4440 9404 4468
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 10226 4468 10232 4480
rect 10187 4440 10232 4468
rect 10226 4428 10232 4440
rect 10284 4428 10290 4480
rect 10962 4428 10968 4480
rect 11020 4468 11026 4480
rect 11517 4471 11575 4477
rect 11517 4468 11529 4471
rect 11020 4440 11529 4468
rect 11020 4428 11026 4440
rect 11517 4437 11529 4440
rect 11563 4437 11575 4471
rect 16022 4468 16028 4480
rect 15983 4440 16028 4468
rect 11517 4431 11575 4437
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 22278 4428 22284 4480
rect 22336 4468 22342 4480
rect 22336 4440 22381 4468
rect 22336 4428 22342 4440
rect 23842 4428 23848 4480
rect 23900 4468 23906 4480
rect 24136 4468 24164 4499
rect 24578 4496 24584 4508
rect 24636 4496 24642 4548
rect 26206 4539 26264 4545
rect 26206 4505 26218 4539
rect 26252 4505 26264 4539
rect 26206 4499 26264 4505
rect 27525 4539 27583 4545
rect 27525 4505 27537 4539
rect 27571 4536 27583 4539
rect 28000 4536 28028 4567
rect 27571 4508 28028 4536
rect 27571 4505 27583 4508
rect 27525 4499 27583 4505
rect 24857 4471 24915 4477
rect 24857 4468 24869 4471
rect 23900 4440 24869 4468
rect 23900 4428 23906 4440
rect 24857 4437 24869 4440
rect 24903 4437 24915 4471
rect 24857 4431 24915 4437
rect 25869 4471 25927 4477
rect 25869 4437 25881 4471
rect 25915 4468 25927 4471
rect 26206 4468 26234 4499
rect 25915 4440 26234 4468
rect 27341 4471 27399 4477
rect 25915 4437 25927 4440
rect 25869 4431 25927 4437
rect 27341 4437 27353 4471
rect 27387 4468 27399 4471
rect 27540 4468 27568 4499
rect 27387 4440 27568 4468
rect 27387 4437 27399 4440
rect 27341 4431 27399 4437
rect 1104 4378 29532 4400
rect 1104 4326 10425 4378
rect 10477 4326 10489 4378
rect 10541 4326 10553 4378
rect 10605 4326 10617 4378
rect 10669 4326 10681 4378
rect 10733 4326 19901 4378
rect 19953 4326 19965 4378
rect 20017 4326 20029 4378
rect 20081 4326 20093 4378
rect 20145 4326 20157 4378
rect 20209 4326 29532 4378
rect 1104 4304 29532 4326
rect 4430 4264 4436 4276
rect 4391 4236 4436 4264
rect 4430 4224 4436 4236
rect 4488 4224 4494 4276
rect 10505 4267 10563 4273
rect 10505 4233 10517 4267
rect 10551 4264 10563 4267
rect 10870 4264 10876 4276
rect 10551 4236 10876 4264
rect 10551 4233 10563 4236
rect 10505 4227 10563 4233
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 15657 4267 15715 4273
rect 15657 4233 15669 4267
rect 15703 4264 15715 4267
rect 15930 4264 15936 4276
rect 15703 4236 15936 4264
rect 15703 4233 15715 4236
rect 15657 4227 15715 4233
rect 15930 4224 15936 4236
rect 15988 4264 15994 4276
rect 16758 4264 16764 4276
rect 15988 4236 16252 4264
rect 16719 4236 16764 4264
rect 15988 4224 15994 4236
rect 8110 4156 8116 4208
rect 8168 4196 8174 4208
rect 8389 4199 8447 4205
rect 8389 4196 8401 4199
rect 8168 4168 8401 4196
rect 8168 4156 8174 4168
rect 8389 4165 8401 4168
rect 8435 4165 8447 4199
rect 8389 4159 8447 4165
rect 1854 4128 1860 4140
rect 1815 4100 1860 4128
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 4522 4088 4528 4140
rect 4580 4128 4586 4140
rect 6362 4128 6368 4140
rect 4580 4100 4625 4128
rect 6323 4100 6368 4128
rect 4580 4088 4586 4100
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 6546 4128 6552 4140
rect 6507 4100 6552 4128
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 7524 4100 8217 4128
rect 7524 4088 7530 4100
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4128 8631 4131
rect 9214 4128 9220 4140
rect 8619 4100 9220 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 4706 4060 4712 4072
rect 4667 4032 4712 4060
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 8220 4060 8248 4091
rect 9214 4088 9220 4100
rect 9272 4128 9278 4140
rect 9402 4131 9460 4137
rect 9402 4128 9414 4131
rect 9272 4100 9414 4128
rect 9272 4088 9278 4100
rect 9402 4097 9414 4100
rect 9448 4097 9460 4131
rect 9402 4091 9460 4097
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4128 9919 4131
rect 10226 4128 10232 4140
rect 9907 4100 10232 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 10226 4088 10232 4100
rect 10284 4128 10290 4140
rect 10598 4131 10656 4137
rect 10598 4128 10610 4131
rect 10284 4100 10610 4128
rect 10284 4088 10290 4100
rect 10598 4097 10610 4100
rect 10644 4097 10656 4131
rect 10962 4128 10968 4140
rect 10923 4100 10968 4128
rect 10598 4091 10656 4097
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 12894 4088 12900 4140
rect 12952 4128 12958 4140
rect 14277 4131 14335 4137
rect 14277 4128 14289 4131
rect 12952 4100 14289 4128
rect 12952 4088 12958 4100
rect 14277 4097 14289 4100
rect 14323 4097 14335 4131
rect 14277 4091 14335 4097
rect 14544 4131 14602 4137
rect 14544 4097 14556 4131
rect 14590 4128 14602 4131
rect 14918 4128 14924 4140
rect 14590 4100 14924 4128
rect 14590 4097 14602 4100
rect 14544 4091 14602 4097
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 16224 4137 16252 4236
rect 16758 4224 16764 4236
rect 16816 4224 16822 4276
rect 18138 4224 18144 4276
rect 18196 4264 18202 4276
rect 18601 4267 18659 4273
rect 18601 4264 18613 4267
rect 18196 4236 18613 4264
rect 18196 4224 18202 4236
rect 18601 4233 18613 4236
rect 18647 4264 18659 4267
rect 18782 4264 18788 4276
rect 18647 4236 18788 4264
rect 18647 4233 18659 4236
rect 18601 4227 18659 4233
rect 18782 4224 18788 4236
rect 18840 4224 18846 4276
rect 21358 4224 21364 4276
rect 21416 4264 21422 4276
rect 21913 4267 21971 4273
rect 21913 4264 21925 4267
rect 21416 4236 21925 4264
rect 21416 4224 21422 4236
rect 21913 4233 21925 4236
rect 21959 4233 21971 4267
rect 24578 4264 24584 4276
rect 21913 4227 21971 4233
rect 22572 4236 24584 4264
rect 16393 4199 16451 4205
rect 16393 4165 16405 4199
rect 16439 4196 16451 4199
rect 16666 4196 16672 4208
rect 16439 4168 16672 4196
rect 16439 4165 16451 4168
rect 16393 4159 16451 4165
rect 16666 4156 16672 4168
rect 16724 4156 16730 4208
rect 17129 4199 17187 4205
rect 17129 4165 17141 4199
rect 17175 4196 17187 4199
rect 18046 4196 18052 4208
rect 17175 4168 18052 4196
rect 17175 4165 17187 4168
rect 17129 4159 17187 4165
rect 18046 4156 18052 4168
rect 18104 4156 18110 4208
rect 18233 4199 18291 4205
rect 18233 4165 18245 4199
rect 18279 4196 18291 4199
rect 18506 4196 18512 4208
rect 18279 4168 18512 4196
rect 18279 4165 18291 4168
rect 18233 4159 18291 4165
rect 18506 4156 18512 4168
rect 18564 4156 18570 4208
rect 19696 4199 19754 4205
rect 19696 4165 19708 4199
rect 19742 4196 19754 4199
rect 19794 4196 19800 4208
rect 19742 4168 19800 4196
rect 19742 4165 19754 4168
rect 19696 4159 19754 4165
rect 19794 4156 19800 4168
rect 19852 4156 19858 4208
rect 22094 4156 22100 4208
rect 22152 4196 22158 4208
rect 22370 4196 22376 4208
rect 22152 4168 22376 4196
rect 22152 4156 22158 4168
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4128 16267 4131
rect 16298 4128 16304 4140
rect 16255 4100 16304 4128
rect 16255 4097 16267 4100
rect 16209 4091 16267 4097
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 22204 4137 22232 4168
rect 22370 4156 22376 4168
rect 22428 4196 22434 4208
rect 22465 4199 22523 4205
rect 22465 4196 22477 4199
rect 22428 4168 22477 4196
rect 22428 4156 22434 4168
rect 22465 4165 22477 4168
rect 22511 4196 22523 4199
rect 22572 4196 22600 4236
rect 24578 4224 24584 4236
rect 24636 4264 24642 4276
rect 25869 4267 25927 4273
rect 25869 4264 25881 4267
rect 24636 4236 25881 4264
rect 24636 4224 24642 4236
rect 25869 4233 25881 4236
rect 25915 4233 25927 4267
rect 25869 4227 25927 4233
rect 23750 4196 23756 4208
rect 22511 4168 22600 4196
rect 23032 4168 23756 4196
rect 22511 4165 22523 4168
rect 22465 4159 22523 4165
rect 22189 4131 22247 4137
rect 22189 4128 22201 4131
rect 18380 4100 22201 4128
rect 18380 4088 18386 4100
rect 22189 4097 22201 4100
rect 22235 4097 22247 4131
rect 22557 4131 22615 4137
rect 22557 4128 22569 4131
rect 22189 4091 22247 4097
rect 22296 4100 22569 4128
rect 9582 4060 9588 4072
rect 8220 4032 9588 4060
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 9769 4063 9827 4069
rect 9769 4029 9781 4063
rect 9815 4060 9827 4063
rect 9950 4060 9956 4072
rect 9815 4032 9956 4060
rect 9815 4029 9827 4032
rect 9769 4023 9827 4029
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 11054 4060 11060 4072
rect 11015 4032 11060 4060
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 16942 4060 16948 4072
rect 15304 4032 16948 4060
rect 4065 3995 4123 4001
rect 4065 3961 4077 3995
rect 4111 3992 4123 3995
rect 4338 3992 4344 4004
rect 4111 3964 4344 3992
rect 4111 3961 4123 3964
rect 4065 3955 4123 3961
rect 4338 3952 4344 3964
rect 4396 3952 4402 4004
rect 11238 3992 11244 4004
rect 6196 3964 11244 3992
rect 842 3884 848 3936
rect 900 3924 906 3936
rect 6196 3924 6224 3964
rect 11238 3952 11244 3964
rect 11296 3952 11302 4004
rect 6362 3924 6368 3936
rect 900 3896 6224 3924
rect 6323 3896 6368 3924
rect 900 3884 906 3896
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 6914 3924 6920 3936
rect 6779 3896 6920 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 6914 3884 6920 3896
rect 6972 3924 6978 3936
rect 8110 3924 8116 3936
rect 6972 3896 8116 3924
rect 6972 3884 6978 3896
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 9309 3927 9367 3933
rect 9309 3893 9321 3927
rect 9355 3924 9367 3927
rect 9674 3924 9680 3936
rect 9355 3896 9680 3924
rect 9355 3893 9367 3896
rect 9309 3887 9367 3893
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 15304 3924 15332 4032
rect 16942 4020 16948 4032
rect 17000 4020 17006 4072
rect 17218 4060 17224 4072
rect 17179 4032 17224 4060
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4060 17371 4063
rect 17770 4060 17776 4072
rect 17359 4032 17776 4060
rect 17359 4029 17371 4032
rect 17313 4023 17371 4029
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 17328 3992 17356 4023
rect 17770 4020 17776 4032
rect 17828 4060 17834 4072
rect 17957 4063 18015 4069
rect 17957 4060 17969 4063
rect 17828 4032 17969 4060
rect 17828 4020 17834 4032
rect 17957 4029 17969 4032
rect 18003 4029 18015 4063
rect 17957 4023 18015 4029
rect 18138 4020 18144 4072
rect 18196 4060 18202 4072
rect 19429 4063 19487 4069
rect 18196 4032 18241 4060
rect 18196 4020 18202 4032
rect 19429 4029 19441 4063
rect 19475 4029 19487 4063
rect 22077 4063 22135 4069
rect 22077 4060 22089 4063
rect 19429 4023 19487 4029
rect 20824 4032 22089 4060
rect 15988 3964 17356 3992
rect 15988 3952 15994 3964
rect 17862 3952 17868 4004
rect 17920 3992 17926 4004
rect 19444 3992 19472 4023
rect 20824 4004 20852 4032
rect 22077 4029 22089 4032
rect 22123 4060 22135 4063
rect 22296 4060 22324 4100
rect 22557 4097 22569 4100
rect 22603 4097 22615 4131
rect 22557 4091 22615 4097
rect 22925 4131 22983 4137
rect 22925 4097 22937 4131
rect 22971 4128 22983 4131
rect 23032 4128 23060 4168
rect 23750 4156 23756 4168
rect 23808 4156 23814 4208
rect 23198 4128 23204 4140
rect 22971 4100 23060 4128
rect 23159 4100 23204 4128
rect 22971 4097 22983 4100
rect 22925 4091 22983 4097
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 23474 4137 23480 4140
rect 23468 4091 23480 4137
rect 23532 4128 23538 4140
rect 23532 4100 23568 4128
rect 23474 4088 23480 4091
rect 23532 4088 23538 4100
rect 25498 4088 25504 4140
rect 25556 4128 25562 4140
rect 25777 4131 25835 4137
rect 25777 4128 25789 4131
rect 25556 4100 25789 4128
rect 25556 4088 25562 4100
rect 25777 4097 25789 4100
rect 25823 4097 25835 4131
rect 25777 4091 25835 4097
rect 26053 4131 26111 4137
rect 26053 4097 26065 4131
rect 26099 4128 26111 4131
rect 26142 4128 26148 4140
rect 26099 4100 26148 4128
rect 26099 4097 26111 4100
rect 26053 4091 26111 4097
rect 26142 4088 26148 4100
rect 26200 4088 26206 4140
rect 22123 4032 22324 4060
rect 22123 4029 22135 4032
rect 22077 4023 22135 4029
rect 20806 3992 20812 4004
rect 17920 3964 19472 3992
rect 20719 3964 20812 3992
rect 17920 3952 17926 3964
rect 14700 3896 15332 3924
rect 16117 3927 16175 3933
rect 14700 3884 14706 3896
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 16666 3924 16672 3936
rect 16163 3896 16672 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 17770 3884 17776 3936
rect 17828 3924 17834 3936
rect 18138 3924 18144 3936
rect 17828 3896 18144 3924
rect 17828 3884 17834 3896
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 19444 3924 19472 3964
rect 20806 3952 20812 3964
rect 20864 3952 20870 4004
rect 24394 3952 24400 4004
rect 24452 3992 24458 4004
rect 24581 3995 24639 4001
rect 24581 3992 24593 3995
rect 24452 3964 24593 3992
rect 24452 3952 24458 3964
rect 24581 3961 24593 3964
rect 24627 3961 24639 3995
rect 24581 3955 24639 3961
rect 20530 3924 20536 3936
rect 19444 3896 20536 3924
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 23109 3927 23167 3933
rect 23109 3893 23121 3927
rect 23155 3924 23167 3927
rect 23934 3924 23940 3936
rect 23155 3896 23940 3924
rect 23155 3893 23167 3896
rect 23109 3887 23167 3893
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 1104 3834 29532 3856
rect 1104 3782 5688 3834
rect 5740 3782 5752 3834
rect 5804 3782 5816 3834
rect 5868 3782 5880 3834
rect 5932 3782 5944 3834
rect 5996 3782 15163 3834
rect 15215 3782 15227 3834
rect 15279 3782 15291 3834
rect 15343 3782 15355 3834
rect 15407 3782 15419 3834
rect 15471 3782 24639 3834
rect 24691 3782 24703 3834
rect 24755 3782 24767 3834
rect 24819 3782 24831 3834
rect 24883 3782 24895 3834
rect 24947 3782 29532 3834
rect 1104 3760 29532 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 2556 3692 2774 3720
rect 2556 3680 2562 3692
rect 2746 3448 2774 3692
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 7834 3720 7840 3732
rect 4304 3692 7840 3720
rect 4304 3680 4310 3692
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 9861 3723 9919 3729
rect 9861 3720 9873 3723
rect 9640 3692 9873 3720
rect 9640 3680 9646 3692
rect 9861 3689 9873 3692
rect 9907 3689 9919 3723
rect 9861 3683 9919 3689
rect 10321 3723 10379 3729
rect 10321 3689 10333 3723
rect 10367 3720 10379 3723
rect 10962 3720 10968 3732
rect 10367 3692 10968 3720
rect 10367 3689 10379 3692
rect 10321 3683 10379 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 14642 3720 14648 3732
rect 11204 3692 14648 3720
rect 11204 3680 11210 3692
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 17770 3720 17776 3732
rect 17731 3692 17776 3720
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 18874 3720 18880 3732
rect 18156 3692 18552 3720
rect 18835 3692 18880 3720
rect 6914 3652 6920 3664
rect 5736 3624 6920 3652
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3584 4859 3587
rect 4890 3584 4896 3596
rect 4847 3556 4896 3584
rect 4847 3553 4859 3556
rect 4801 3547 4859 3553
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 4614 3516 4620 3528
rect 4575 3488 4620 3516
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 5736 3525 5764 3624
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 8573 3655 8631 3661
rect 8573 3652 8585 3655
rect 7944 3624 8585 3652
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 5687 3519 5764 3525
rect 5687 3485 5699 3519
rect 5733 3488 5764 3519
rect 5733 3485 5745 3488
rect 5687 3479 5745 3485
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5868 3488 6009 3516
rect 5868 3476 5874 3488
rect 5997 3485 6009 3488
rect 6043 3516 6055 3519
rect 6362 3516 6368 3528
rect 6043 3488 6368 3516
rect 6043 3485 6055 3488
rect 5997 3479 6055 3485
rect 6362 3476 6368 3488
rect 6420 3476 6426 3528
rect 6730 3516 6736 3528
rect 6691 3488 6736 3516
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 6917 3519 6975 3525
rect 6917 3485 6929 3519
rect 6963 3516 6975 3519
rect 7006 3516 7012 3528
rect 6963 3488 7012 3516
rect 6963 3485 6975 3488
rect 6917 3479 6975 3485
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3516 7251 3519
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 7239 3488 7481 3516
rect 7239 3485 7251 3488
rect 7193 3479 7251 3485
rect 7469 3485 7481 3488
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 7711 3519 7769 3525
rect 7711 3485 7723 3519
rect 7757 3516 7769 3519
rect 7944 3516 7972 3624
rect 8573 3621 8585 3624
rect 8619 3652 8631 3655
rect 10778 3652 10784 3664
rect 8619 3624 10784 3652
rect 8619 3621 8631 3624
rect 8573 3615 8631 3621
rect 10778 3612 10784 3624
rect 10836 3652 10842 3664
rect 11238 3652 11244 3664
rect 10836 3624 11244 3652
rect 10836 3612 10842 3624
rect 11238 3612 11244 3624
rect 11296 3612 11302 3664
rect 11422 3612 11428 3664
rect 11480 3652 11486 3664
rect 12710 3652 12716 3664
rect 11480 3624 12716 3652
rect 11480 3612 11486 3624
rect 12710 3612 12716 3624
rect 12768 3612 12774 3664
rect 16666 3612 16672 3664
rect 16724 3652 16730 3664
rect 16724 3624 16988 3652
rect 16724 3612 16730 3624
rect 8110 3584 8116 3596
rect 8071 3556 8116 3584
rect 8110 3544 8116 3556
rect 8168 3584 8174 3596
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 8168 3556 8248 3584
rect 8168 3544 8174 3556
rect 7757 3488 7972 3516
rect 7757 3485 7769 3488
rect 7711 3479 7769 3485
rect 8018 3476 8024 3528
rect 8076 3518 8082 3528
rect 8220 3525 8248 3556
rect 8404 3556 10149 3584
rect 8404 3525 8432 3556
rect 10137 3553 10149 3556
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 11054 3544 11060 3596
rect 11112 3584 11118 3596
rect 11793 3587 11851 3593
rect 11793 3584 11805 3587
rect 11112 3556 11805 3584
rect 11112 3544 11118 3556
rect 8205 3519 8263 3525
rect 8076 3516 8095 3518
rect 8076 3488 8169 3516
rect 8076 3476 8082 3488
rect 8128 3448 8156 3488
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 9214 3516 9220 3528
rect 9175 3488 9220 3516
rect 8389 3479 8447 3485
rect 8404 3448 8432 3479
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3485 9459 3519
rect 9674 3516 9680 3528
rect 9635 3488 9680 3516
rect 9401 3479 9459 3485
rect 2746 3420 7880 3448
rect 8128 3420 8432 3448
rect 9416 3448 9444 3479
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 10042 3516 10048 3528
rect 10003 3488 10048 3516
rect 10042 3476 10048 3488
rect 10100 3516 10106 3528
rect 10931 3519 10989 3525
rect 10100 3488 10824 3516
rect 10100 3476 10106 3488
rect 9416 3420 9628 3448
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 4433 3383 4491 3389
rect 4433 3380 4445 3383
rect 3936 3352 4445 3380
rect 3936 3340 3942 3352
rect 4433 3349 4445 3352
rect 4479 3349 4491 3383
rect 4433 3343 4491 3349
rect 5537 3383 5595 3389
rect 5537 3349 5549 3383
rect 5583 3380 5595 3383
rect 5902 3380 5908 3392
rect 5583 3352 5908 3380
rect 5583 3349 5595 3352
rect 5537 3343 5595 3349
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 5994 3340 6000 3392
rect 6052 3380 6058 3392
rect 6549 3383 6607 3389
rect 6549 3380 6561 3383
rect 6052 3352 6561 3380
rect 6052 3340 6058 3352
rect 6549 3349 6561 3352
rect 6595 3349 6607 3383
rect 6549 3343 6607 3349
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6788 3352 7021 3380
rect 6788 3340 6794 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 7852 3380 7880 3420
rect 8202 3380 8208 3392
rect 7852 3352 8208 3380
rect 7009 3343 7067 3349
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 9033 3383 9091 3389
rect 9033 3380 9045 3383
rect 8352 3352 9045 3380
rect 8352 3340 8358 3352
rect 9033 3349 9045 3352
rect 9079 3349 9091 3383
rect 9033 3343 9091 3349
rect 9214 3340 9220 3392
rect 9272 3380 9278 3392
rect 9493 3383 9551 3389
rect 9493 3380 9505 3383
rect 9272 3352 9505 3380
rect 9272 3340 9278 3352
rect 9493 3349 9505 3352
rect 9539 3349 9551 3383
rect 9600 3380 9628 3420
rect 9950 3408 9956 3460
rect 10008 3448 10014 3460
rect 10321 3451 10379 3457
rect 10321 3448 10333 3451
rect 10008 3420 10333 3448
rect 10008 3408 10014 3420
rect 10321 3417 10333 3420
rect 10367 3417 10379 3451
rect 10796 3448 10824 3488
rect 10931 3485 10943 3519
rect 10977 3516 10989 3519
rect 11164 3516 11192 3556
rect 11793 3553 11805 3556
rect 11839 3553 11851 3587
rect 15930 3584 15936 3596
rect 15891 3556 15936 3584
rect 11793 3547 11851 3553
rect 15930 3544 15936 3556
rect 15988 3544 15994 3596
rect 16298 3544 16304 3596
rect 16356 3584 16362 3596
rect 16356 3556 16896 3584
rect 16356 3544 16362 3556
rect 10977 3488 11192 3516
rect 11241 3519 11299 3525
rect 10977 3485 10989 3488
rect 10931 3479 10989 3485
rect 11241 3485 11253 3519
rect 11287 3485 11299 3519
rect 11241 3479 11299 3485
rect 11256 3448 11284 3479
rect 11330 3476 11336 3528
rect 11388 3516 11394 3528
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 11388 3488 11437 3516
rect 11388 3476 11394 3488
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 11882 3516 11888 3528
rect 11843 3488 11888 3516
rect 11425 3479 11483 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16209 3519 16267 3525
rect 16209 3516 16221 3519
rect 16080 3488 16221 3516
rect 16080 3476 16086 3488
rect 16209 3485 16221 3488
rect 16255 3485 16267 3519
rect 16209 3479 16267 3485
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3516 16727 3519
rect 16758 3516 16764 3528
rect 16715 3488 16764 3516
rect 16715 3485 16727 3488
rect 16669 3479 16727 3485
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 16868 3525 16896 3556
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3485 16911 3519
rect 16960 3516 16988 3624
rect 17221 3587 17279 3593
rect 17221 3553 17233 3587
rect 17267 3584 17279 3587
rect 17405 3587 17463 3593
rect 17405 3584 17417 3587
rect 17267 3556 17417 3584
rect 17267 3553 17279 3556
rect 17221 3547 17279 3553
rect 17405 3553 17417 3556
rect 17451 3584 17463 3587
rect 18156 3584 18184 3692
rect 18524 3661 18552 3692
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 19613 3723 19671 3729
rect 19613 3720 19625 3723
rect 19484 3692 19625 3720
rect 19484 3680 19490 3692
rect 19613 3689 19625 3692
rect 19659 3689 19671 3723
rect 22094 3720 22100 3732
rect 19613 3683 19671 3689
rect 20364 3692 22100 3720
rect 18509 3655 18567 3661
rect 18509 3621 18521 3655
rect 18555 3621 18567 3655
rect 18509 3615 18567 3621
rect 18966 3612 18972 3664
rect 19024 3652 19030 3664
rect 19024 3624 19380 3652
rect 19024 3612 19030 3624
rect 18233 3587 18291 3593
rect 18233 3584 18245 3587
rect 17451 3556 18245 3584
rect 17451 3553 17463 3556
rect 17405 3547 17463 3553
rect 18233 3553 18245 3556
rect 18279 3553 18291 3587
rect 18233 3547 18291 3553
rect 18325 3587 18383 3593
rect 18325 3553 18337 3587
rect 18371 3584 18383 3587
rect 18782 3584 18788 3596
rect 18371 3556 18788 3584
rect 18371 3553 18383 3556
rect 18325 3547 18383 3553
rect 18782 3544 18788 3556
rect 18840 3584 18846 3596
rect 18840 3556 19288 3584
rect 18840 3544 18846 3556
rect 17313 3519 17371 3525
rect 17313 3516 17325 3519
rect 16960 3488 17325 3516
rect 16853 3479 16911 3485
rect 17313 3485 17325 3488
rect 17359 3485 17371 3519
rect 17313 3479 17371 3485
rect 18029 3519 18087 3525
rect 18029 3485 18041 3519
rect 18075 3516 18087 3519
rect 18416 3519 18474 3525
rect 18075 3488 18368 3516
rect 18075 3485 18087 3488
rect 18029 3479 18087 3485
rect 11609 3451 11667 3457
rect 11609 3448 11621 3451
rect 10796 3420 11621 3448
rect 10321 3411 10379 3417
rect 10980 3392 11008 3420
rect 11609 3417 11621 3420
rect 11655 3417 11667 3451
rect 11609 3411 11667 3417
rect 16117 3451 16175 3457
rect 16117 3417 16129 3451
rect 16163 3448 16175 3451
rect 16163 3420 16896 3448
rect 16163 3417 16175 3420
rect 16117 3411 16175 3417
rect 10134 3380 10140 3392
rect 9600 3352 10140 3380
rect 9493 3343 9551 3349
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 10778 3380 10784 3392
rect 10739 3352 10784 3380
rect 10778 3340 10784 3352
rect 10836 3340 10842 3392
rect 10962 3340 10968 3392
rect 11020 3340 11026 3392
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 12069 3383 12127 3389
rect 12069 3380 12081 3383
rect 12032 3352 12081 3380
rect 12032 3340 12038 3352
rect 12069 3349 12081 3352
rect 12115 3349 12127 3383
rect 12069 3343 12127 3349
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 16868 3389 16896 3420
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 17773 3451 17831 3457
rect 17773 3448 17785 3451
rect 17092 3420 17785 3448
rect 17092 3408 17098 3420
rect 17773 3417 17785 3420
rect 17819 3448 17831 3451
rect 18340 3448 18368 3488
rect 18416 3485 18428 3519
rect 18462 3518 18474 3519
rect 18598 3518 18604 3528
rect 18462 3490 18604 3518
rect 18462 3485 18474 3490
rect 18416 3479 18474 3485
rect 18598 3476 18604 3490
rect 18656 3476 18662 3528
rect 18690 3476 18696 3528
rect 18748 3516 18754 3528
rect 19260 3525 19288 3556
rect 19245 3519 19303 3525
rect 18748 3488 18793 3516
rect 18748 3476 18754 3488
rect 19245 3485 19257 3519
rect 19291 3485 19303 3519
rect 19352 3516 19380 3624
rect 20257 3587 20315 3593
rect 20257 3553 20269 3587
rect 20303 3584 20315 3587
rect 20364 3584 20392 3692
rect 22094 3680 22100 3692
rect 22152 3680 22158 3732
rect 22189 3723 22247 3729
rect 22189 3689 22201 3723
rect 22235 3720 22247 3723
rect 22278 3720 22284 3732
rect 22235 3692 22284 3720
rect 22235 3689 22247 3692
rect 22189 3683 22247 3689
rect 22278 3680 22284 3692
rect 22336 3680 22342 3732
rect 23474 3720 23480 3732
rect 23435 3692 23480 3720
rect 23474 3680 23480 3692
rect 23532 3680 23538 3732
rect 23382 3612 23388 3664
rect 23440 3652 23446 3664
rect 23440 3624 24072 3652
rect 23440 3612 23446 3624
rect 20530 3584 20536 3596
rect 20303 3556 20392 3584
rect 20491 3556 20536 3584
rect 20303 3553 20315 3556
rect 20257 3547 20315 3553
rect 20530 3544 20536 3556
rect 20588 3544 20594 3596
rect 22557 3587 22615 3593
rect 22557 3584 22569 3587
rect 21560 3556 22569 3584
rect 20800 3519 20858 3525
rect 19352 3488 20576 3516
rect 19245 3479 19303 3485
rect 18506 3448 18512 3460
rect 17819 3420 18276 3448
rect 18340 3420 18512 3448
rect 17819 3417 17831 3420
rect 17773 3411 17831 3417
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 16448 3352 16589 3380
rect 16448 3340 16454 3352
rect 16577 3349 16589 3352
rect 16623 3349 16635 3383
rect 16577 3343 16635 3349
rect 16853 3383 16911 3389
rect 16853 3349 16865 3383
rect 16899 3349 16911 3383
rect 16853 3343 16911 3349
rect 18046 3340 18052 3392
rect 18104 3380 18110 3392
rect 18141 3383 18199 3389
rect 18141 3380 18153 3383
rect 18104 3352 18153 3380
rect 18104 3340 18110 3352
rect 18141 3349 18153 3352
rect 18187 3349 18199 3383
rect 18248 3380 18276 3420
rect 18506 3408 18512 3420
rect 18564 3448 18570 3460
rect 19337 3451 19395 3457
rect 19337 3448 19349 3451
rect 18564 3420 19349 3448
rect 18564 3408 18570 3420
rect 19337 3417 19349 3420
rect 19383 3417 19395 3451
rect 19337 3411 19395 3417
rect 19981 3451 20039 3457
rect 19981 3417 19993 3451
rect 20027 3448 20039 3451
rect 20254 3448 20260 3460
rect 20027 3420 20260 3448
rect 20027 3417 20039 3420
rect 19981 3411 20039 3417
rect 20254 3408 20260 3420
rect 20312 3408 20318 3460
rect 18690 3380 18696 3392
rect 18248 3352 18696 3380
rect 18141 3343 18199 3349
rect 18690 3340 18696 3352
rect 18748 3340 18754 3392
rect 20073 3383 20131 3389
rect 20073 3349 20085 3383
rect 20119 3380 20131 3383
rect 20438 3380 20444 3392
rect 20119 3352 20444 3380
rect 20119 3349 20131 3352
rect 20073 3343 20131 3349
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 20548 3380 20576 3488
rect 20800 3485 20812 3519
rect 20846 3516 20858 3519
rect 21082 3516 21088 3528
rect 20846 3488 21088 3516
rect 20846 3485 20858 3488
rect 20800 3479 20858 3485
rect 21082 3476 21088 3488
rect 21140 3476 21146 3528
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 21560 3448 21588 3556
rect 22557 3553 22569 3556
rect 22603 3584 22615 3587
rect 22833 3587 22891 3593
rect 22833 3584 22845 3587
rect 22603 3556 22845 3584
rect 22603 3553 22615 3556
rect 22557 3547 22615 3553
rect 22833 3553 22845 3556
rect 22879 3553 22891 3587
rect 23934 3584 23940 3596
rect 23895 3556 23940 3584
rect 22833 3547 22891 3553
rect 23934 3544 23940 3556
rect 23992 3544 23998 3596
rect 24044 3593 24072 3624
rect 24029 3587 24087 3593
rect 24029 3553 24041 3587
rect 24075 3553 24087 3587
rect 24029 3547 24087 3553
rect 22370 3516 22376 3528
rect 22331 3488 22376 3516
rect 22370 3476 22376 3488
rect 22428 3476 22434 3528
rect 22646 3516 22652 3528
rect 22607 3488 22652 3516
rect 22646 3476 22652 3488
rect 22704 3476 22710 3528
rect 22741 3519 22799 3525
rect 22741 3485 22753 3519
rect 22787 3485 22799 3519
rect 23842 3516 23848 3528
rect 23803 3488 23848 3516
rect 22741 3479 22799 3485
rect 20680 3420 21588 3448
rect 21652 3420 22140 3448
rect 20680 3408 20686 3420
rect 21652 3380 21680 3420
rect 20548 3352 21680 3380
rect 21913 3383 21971 3389
rect 21913 3349 21925 3383
rect 21959 3380 21971 3383
rect 22002 3380 22008 3392
rect 21959 3352 22008 3380
rect 21959 3349 21971 3352
rect 21913 3343 21971 3349
rect 22002 3340 22008 3352
rect 22060 3340 22066 3392
rect 22112 3380 22140 3420
rect 22186 3408 22192 3460
rect 22244 3448 22250 3460
rect 22756 3448 22784 3479
rect 23842 3476 23848 3488
rect 23900 3476 23906 3528
rect 29641 3519 29699 3525
rect 29641 3485 29653 3519
rect 29687 3516 29699 3519
rect 29822 3516 29828 3528
rect 29687 3488 29828 3516
rect 29687 3485 29699 3488
rect 29641 3479 29699 3485
rect 29822 3476 29828 3488
rect 29880 3476 29886 3528
rect 22244 3420 22784 3448
rect 22244 3408 22250 3420
rect 22738 3380 22744 3392
rect 22112 3352 22744 3380
rect 22738 3340 22744 3352
rect 22796 3340 22802 3392
rect 1104 3290 29532 3312
rect 1104 3238 10425 3290
rect 10477 3238 10489 3290
rect 10541 3238 10553 3290
rect 10605 3238 10617 3290
rect 10669 3238 10681 3290
rect 10733 3238 19901 3290
rect 19953 3238 19965 3290
rect 20017 3238 20029 3290
rect 20081 3238 20093 3290
rect 20145 3238 20157 3290
rect 20209 3238 29532 3290
rect 1104 3216 29532 3238
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 4672 3148 5733 3176
rect 4672 3136 4678 3148
rect 5721 3145 5733 3148
rect 5767 3145 5779 3179
rect 5721 3139 5779 3145
rect 7745 3179 7803 3185
rect 7745 3145 7757 3179
rect 7791 3176 7803 3179
rect 8018 3176 8024 3188
rect 7791 3148 8024 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 8202 3136 8208 3188
rect 8260 3176 8266 3188
rect 9766 3176 9772 3188
rect 8260 3148 9772 3176
rect 8260 3136 8266 3148
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 9950 3176 9956 3188
rect 9911 3148 9956 3176
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 11241 3179 11299 3185
rect 11241 3145 11253 3179
rect 11287 3176 11299 3179
rect 11882 3176 11888 3188
rect 11287 3148 11888 3176
rect 11287 3145 11299 3148
rect 11241 3139 11299 3145
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 16206 3136 16212 3188
rect 16264 3176 16270 3188
rect 18230 3176 18236 3188
rect 16264 3148 18236 3176
rect 16264 3136 16270 3148
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 18601 3179 18659 3185
rect 18601 3145 18613 3179
rect 18647 3176 18659 3179
rect 18782 3176 18788 3188
rect 18647 3148 18788 3176
rect 18647 3145 18659 3148
rect 18601 3139 18659 3145
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 18874 3136 18880 3188
rect 18932 3176 18938 3188
rect 19794 3176 19800 3188
rect 18932 3148 19800 3176
rect 18932 3136 18938 3148
rect 19794 3136 19800 3148
rect 19852 3136 19858 3188
rect 20165 3179 20223 3185
rect 20165 3145 20177 3179
rect 20211 3176 20223 3179
rect 20254 3176 20260 3188
rect 20211 3148 20260 3176
rect 20211 3145 20223 3148
rect 20165 3139 20223 3145
rect 20254 3136 20260 3148
rect 20312 3176 20318 3188
rect 22373 3179 22431 3185
rect 20312 3148 20944 3176
rect 20312 3136 20318 3148
rect 8386 3108 8392 3120
rect 4356 3080 8392 3108
rect 3878 3040 3884 3052
rect 3839 3012 3884 3040
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 4356 3040 4384 3080
rect 4430 3049 4436 3052
rect 4264 3012 4384 3040
rect 4062 2932 4068 2984
rect 4120 2972 4126 2984
rect 4157 2975 4215 2981
rect 4157 2972 4169 2975
rect 4120 2944 4169 2972
rect 4120 2932 4126 2944
rect 4157 2941 4169 2944
rect 4203 2972 4215 2975
rect 4264 2972 4292 3012
rect 4424 3003 4436 3049
rect 4488 3040 4494 3052
rect 5902 3040 5908 3052
rect 4488 3012 4524 3040
rect 5863 3012 5908 3040
rect 4430 3000 4436 3003
rect 4488 3000 4494 3012
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 5994 3000 6000 3052
rect 6052 3040 6058 3052
rect 6380 3049 6408 3080
rect 8386 3068 8392 3080
rect 8444 3108 8450 3120
rect 14458 3108 14464 3120
rect 8444 3080 8616 3108
rect 8444 3068 8450 3080
rect 6365 3043 6423 3049
rect 6052 3012 6097 3040
rect 6052 3000 6058 3012
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6621 3043 6679 3049
rect 6621 3040 6633 3043
rect 6512 3012 6633 3040
rect 6512 3000 6518 3012
rect 6621 3009 6633 3012
rect 6667 3009 6679 3043
rect 8294 3040 8300 3052
rect 8255 3012 8300 3040
rect 6621 3003 6679 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8588 3049 8616 3080
rect 8680 3080 14464 3108
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 4203 2944 4292 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 7650 2932 7656 2984
rect 7708 2972 7714 2984
rect 8680 2972 8708 3080
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 17862 3108 17868 3120
rect 15028 3080 17868 3108
rect 15028 3052 15056 3080
rect 8846 3049 8852 3052
rect 8840 3003 8852 3049
rect 8904 3040 8910 3052
rect 10597 3043 10655 3049
rect 8904 3012 8940 3040
rect 8846 3000 8852 3003
rect 8904 3000 8910 3012
rect 10597 3009 10609 3043
rect 10643 3040 10655 3043
rect 10778 3040 10784 3052
rect 10643 3012 10784 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11057 3043 11115 3049
rect 11057 3009 11069 3043
rect 11103 3009 11115 3043
rect 11057 3003 11115 3009
rect 7708 2944 8708 2972
rect 7708 2932 7714 2944
rect 10134 2932 10140 2984
rect 10192 2972 10198 2984
rect 10873 2975 10931 2981
rect 10873 2972 10885 2975
rect 10192 2944 10885 2972
rect 10192 2932 10198 2944
rect 10873 2941 10885 2944
rect 10919 2941 10931 2975
rect 10873 2935 10931 2941
rect 11072 2916 11100 3003
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12722 3043 12780 3049
rect 12722 3040 12734 3043
rect 12492 3012 12734 3040
rect 12492 3000 12498 3012
rect 12722 3009 12734 3012
rect 12768 3009 12780 3043
rect 12722 3003 12780 3009
rect 12894 3000 12900 3052
rect 12952 3040 12958 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12952 3012 13001 3040
rect 12952 3000 12958 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 15010 3040 15016 3052
rect 14971 3012 15016 3040
rect 12989 3003 13047 3009
rect 15010 3000 15016 3012
rect 15068 3000 15074 3052
rect 15280 3043 15338 3049
rect 15280 3009 15292 3043
rect 15326 3040 15338 3043
rect 15562 3040 15568 3052
rect 15326 3012 15568 3040
rect 15326 3009 15338 3012
rect 15280 3003 15338 3009
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 17034 3040 17040 3052
rect 16995 3012 17040 3040
rect 16853 3003 16911 3009
rect 16868 2972 16896 3003
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 17236 3049 17264 3080
rect 17862 3068 17868 3080
rect 17920 3108 17926 3120
rect 19702 3108 19708 3120
rect 17920 3080 18828 3108
rect 17920 3068 17926 3080
rect 17494 3049 17500 3052
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3009 17279 3043
rect 17488 3040 17500 3049
rect 17455 3012 17500 3040
rect 17221 3003 17279 3009
rect 17488 3003 17500 3012
rect 17494 3000 17500 3003
rect 17552 3000 17558 3052
rect 18800 3049 18828 3080
rect 18892 3080 19708 3108
rect 18785 3043 18843 3049
rect 18785 3009 18797 3043
rect 18831 3009 18843 3043
rect 18785 3003 18843 3009
rect 16942 2972 16948 2984
rect 16408 2944 16948 2972
rect 5537 2907 5595 2913
rect 5537 2873 5549 2907
rect 5583 2904 5595 2907
rect 5810 2904 5816 2916
rect 5583 2876 5816 2904
rect 5583 2873 5595 2876
rect 5537 2867 5595 2873
rect 5810 2864 5816 2876
rect 5868 2864 5874 2916
rect 7374 2864 7380 2916
rect 7432 2904 7438 2916
rect 10781 2907 10839 2913
rect 7432 2876 8616 2904
rect 7432 2864 7438 2876
rect 4065 2839 4123 2845
rect 4065 2805 4077 2839
rect 4111 2836 4123 2839
rect 4798 2836 4804 2848
rect 4111 2808 4804 2836
rect 4111 2805 4123 2808
rect 4065 2799 4123 2805
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 6178 2836 6184 2848
rect 6139 2808 6184 2836
rect 6178 2796 6184 2808
rect 6236 2796 6242 2848
rect 8478 2836 8484 2848
rect 8439 2808 8484 2836
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 8588 2836 8616 2876
rect 10781 2873 10793 2907
rect 10827 2904 10839 2907
rect 11054 2904 11060 2916
rect 10827 2876 11060 2904
rect 10827 2873 10839 2876
rect 10781 2867 10839 2873
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 16408 2913 16436 2944
rect 16942 2932 16948 2944
rect 17000 2932 17006 2984
rect 18230 2932 18236 2984
rect 18288 2972 18294 2984
rect 18892 2972 18920 3080
rect 19702 3068 19708 3080
rect 19760 3068 19766 3120
rect 20438 3108 20444 3120
rect 20399 3080 20444 3108
rect 20438 3068 20444 3080
rect 20496 3068 20502 3120
rect 20806 3108 20812 3120
rect 20767 3080 20812 3108
rect 20806 3068 20812 3080
rect 20864 3068 20870 3120
rect 20916 3117 20944 3148
rect 22373 3145 22385 3179
rect 22419 3176 22431 3179
rect 22646 3176 22652 3188
rect 22419 3148 22652 3176
rect 22419 3145 22431 3148
rect 22373 3139 22431 3145
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 20901 3111 20959 3117
rect 20901 3077 20913 3111
rect 20947 3108 20959 3111
rect 20993 3111 21051 3117
rect 20993 3108 21005 3111
rect 20947 3080 21005 3108
rect 20947 3077 20959 3080
rect 20901 3071 20959 3077
rect 20993 3077 21005 3080
rect 21039 3077 21051 3111
rect 21818 3108 21824 3120
rect 21779 3080 21824 3108
rect 20993 3071 21051 3077
rect 21818 3068 21824 3080
rect 21876 3068 21882 3120
rect 22002 3108 22008 3120
rect 21963 3080 22008 3108
rect 22002 3068 22008 3080
rect 22060 3108 22066 3120
rect 22060 3080 22324 3108
rect 22060 3068 22066 3080
rect 19058 3049 19064 3052
rect 19052 3040 19064 3049
rect 19019 3012 19064 3040
rect 19052 3003 19064 3012
rect 19058 3000 19064 3003
rect 19116 3000 19122 3052
rect 20622 3040 20628 3052
rect 20583 3012 20628 3040
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 20824 3040 20852 3068
rect 21177 3043 21235 3049
rect 21177 3040 21189 3043
rect 20824 3012 21189 3040
rect 21177 3009 21189 3012
rect 21223 3009 21235 3043
rect 21177 3003 21235 3009
rect 21361 3043 21419 3049
rect 21361 3009 21373 3043
rect 21407 3040 21419 3043
rect 22186 3040 22192 3052
rect 21407 3012 22192 3040
rect 21407 3009 21419 3012
rect 21361 3003 21419 3009
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 22296 3049 22324 3080
rect 22281 3043 22339 3049
rect 22281 3009 22293 3043
rect 22327 3009 22339 3043
rect 22281 3003 22339 3009
rect 18288 2944 18920 2972
rect 18288 2932 18294 2944
rect 22002 2932 22008 2984
rect 22060 2972 22066 2984
rect 22370 2972 22376 2984
rect 22060 2944 22376 2972
rect 22060 2932 22066 2944
rect 22370 2932 22376 2944
rect 22428 2932 22434 2984
rect 16393 2907 16451 2913
rect 16393 2873 16405 2907
rect 16439 2873 16451 2907
rect 21726 2904 21732 2916
rect 16393 2867 16451 2873
rect 19720 2876 21732 2904
rect 9306 2836 9312 2848
rect 8588 2808 9312 2836
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 10962 2796 10968 2848
rect 11020 2836 11026 2848
rect 11609 2839 11667 2845
rect 11609 2836 11621 2839
rect 11020 2808 11621 2836
rect 11020 2796 11026 2808
rect 11609 2805 11621 2808
rect 11655 2805 11667 2839
rect 11609 2799 11667 2805
rect 14458 2796 14464 2848
rect 14516 2836 14522 2848
rect 19720 2836 19748 2876
rect 21726 2864 21732 2876
rect 21784 2864 21790 2916
rect 14516 2808 19748 2836
rect 14516 2796 14522 2808
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 21818 2836 21824 2848
rect 19852 2808 21824 2836
rect 19852 2796 19858 2808
rect 21818 2796 21824 2808
rect 21876 2796 21882 2848
rect 1104 2746 29532 2768
rect 1104 2694 5688 2746
rect 5740 2694 5752 2746
rect 5804 2694 5816 2746
rect 5868 2694 5880 2746
rect 5932 2694 5944 2746
rect 5996 2694 15163 2746
rect 15215 2694 15227 2746
rect 15279 2694 15291 2746
rect 15343 2694 15355 2746
rect 15407 2694 15419 2746
rect 15471 2694 24639 2746
rect 24691 2694 24703 2746
rect 24755 2694 24767 2746
rect 24819 2694 24831 2746
rect 24883 2694 24895 2746
rect 24947 2694 29532 2746
rect 1104 2672 29532 2694
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2632 4399 2635
rect 4430 2632 4436 2644
rect 4387 2604 4436 2632
rect 4387 2601 4399 2604
rect 4341 2595 4399 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 6454 2632 6460 2644
rect 6415 2604 6460 2632
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 8846 2592 8852 2644
rect 8904 2632 8910 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8904 2604 8953 2632
rect 8904 2592 8910 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 11517 2635 11575 2641
rect 11517 2601 11529 2635
rect 11563 2632 11575 2635
rect 12434 2632 12440 2644
rect 11563 2604 12440 2632
rect 11563 2601 11575 2604
rect 11517 2595 11575 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 17037 2635 17095 2641
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 18046 2632 18052 2644
rect 17083 2604 18052 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 4706 2524 4712 2576
rect 4764 2564 4770 2576
rect 8662 2564 8668 2576
rect 4764 2536 8668 2564
rect 4764 2524 4770 2536
rect 4798 2496 4804 2508
rect 4759 2468 4804 2496
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 5000 2505 5028 2536
rect 4985 2499 5043 2505
rect 4985 2465 4997 2499
rect 5031 2465 5043 2499
rect 4985 2459 5043 2465
rect 6178 2456 6184 2508
rect 6236 2496 6242 2508
rect 7116 2505 7144 2536
rect 8662 2524 8668 2536
rect 8720 2564 8726 2576
rect 8720 2536 12112 2564
rect 8720 2524 8726 2536
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6236 2468 6929 2496
rect 6236 2456 6242 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 7101 2499 7159 2505
rect 7101 2465 7113 2499
rect 7147 2496 7159 2499
rect 7147 2468 7181 2496
rect 7147 2465 7159 2468
rect 7101 2459 7159 2465
rect 8478 2456 8484 2508
rect 8536 2496 8542 2508
rect 9600 2505 9628 2536
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 8536 2468 9413 2496
rect 8536 2456 8542 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2465 9643 2499
rect 11974 2496 11980 2508
rect 11935 2468 11980 2496
rect 9585 2459 9643 2465
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 12084 2505 12112 2536
rect 12069 2499 12127 2505
rect 12069 2465 12081 2499
rect 12115 2465 12127 2499
rect 12069 2459 12127 2465
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4672 2400 4721 2428
rect 4672 2388 4678 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6788 2400 6837 2428
rect 6788 2388 6794 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9272 2400 9321 2428
rect 9272 2388 9278 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11112 2400 11897 2428
rect 11112 2388 11118 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 16942 2428 16948 2440
rect 16903 2400 16948 2428
rect 11885 2391 11943 2397
rect 16942 2388 16948 2400
rect 17000 2388 17006 2440
rect 3418 2320 3424 2372
rect 3476 2360 3482 2372
rect 9122 2360 9128 2372
rect 3476 2332 9128 2360
rect 3476 2320 3482 2332
rect 9122 2320 9128 2332
rect 9180 2320 9186 2372
rect 1104 2202 29532 2224
rect 1104 2150 10425 2202
rect 10477 2150 10489 2202
rect 10541 2150 10553 2202
rect 10605 2150 10617 2202
rect 10669 2150 10681 2202
rect 10733 2150 19901 2202
rect 19953 2150 19965 2202
rect 20017 2150 20029 2202
rect 20081 2150 20093 2202
rect 20145 2150 20157 2202
rect 20209 2150 29532 2202
rect 1104 2128 29532 2150
rect 3142 1300 3148 1352
rect 3200 1340 3206 1352
rect 9030 1340 9036 1352
rect 3200 1312 9036 1340
rect 3200 1300 3206 1312
rect 9030 1300 9036 1312
rect 9088 1300 9094 1352
rect 16850 1300 16856 1352
rect 16908 1340 16914 1352
rect 27522 1340 27528 1352
rect 16908 1312 27528 1340
rect 16908 1300 16914 1312
rect 27522 1300 27528 1312
rect 27580 1300 27586 1352
<< via1 >>
rect 11152 30676 11204 30728
rect 11612 30676 11664 30728
rect 3884 30608 3936 30660
rect 13912 30608 13964 30660
rect 15292 30608 15344 30660
rect 16028 30608 16080 30660
rect 10784 30540 10836 30592
rect 16488 30540 16540 30592
rect 10425 30438 10477 30490
rect 10489 30438 10541 30490
rect 10553 30438 10605 30490
rect 10617 30438 10669 30490
rect 10681 30438 10733 30490
rect 19901 30438 19953 30490
rect 19965 30438 20017 30490
rect 20029 30438 20081 30490
rect 20093 30438 20145 30490
rect 20157 30438 20209 30490
rect 4068 30336 4120 30388
rect 10784 30268 10836 30320
rect 9036 30200 9088 30252
rect 10140 30243 10192 30252
rect 10140 30209 10149 30243
rect 10149 30209 10183 30243
rect 10183 30209 10192 30243
rect 11704 30243 11756 30252
rect 10140 30200 10192 30209
rect 11704 30209 11713 30243
rect 11713 30209 11747 30243
rect 11747 30209 11756 30243
rect 11704 30200 11756 30209
rect 9680 30132 9732 30184
rect 9864 30175 9916 30184
rect 9864 30141 9873 30175
rect 9873 30141 9907 30175
rect 9907 30141 9916 30175
rect 12532 30200 12584 30252
rect 13268 30200 13320 30252
rect 14464 30243 14516 30252
rect 14464 30209 14473 30243
rect 14473 30209 14507 30243
rect 14507 30209 14516 30243
rect 14464 30200 14516 30209
rect 14740 30243 14792 30252
rect 14740 30209 14749 30243
rect 14749 30209 14783 30243
rect 14783 30209 14792 30243
rect 15016 30243 15068 30252
rect 14740 30200 14792 30209
rect 15016 30209 15025 30243
rect 15025 30209 15059 30243
rect 15059 30209 15068 30243
rect 15016 30200 15068 30209
rect 9864 30132 9916 30141
rect 4068 30064 4120 30116
rect 11980 30175 12032 30184
rect 11980 30141 11989 30175
rect 11989 30141 12023 30175
rect 12023 30141 12032 30175
rect 14832 30175 14884 30184
rect 11980 30132 12032 30141
rect 14832 30141 14841 30175
rect 14841 30141 14875 30175
rect 14875 30141 14884 30175
rect 14832 30132 14884 30141
rect 16948 30243 17000 30252
rect 16948 30209 16957 30243
rect 16957 30209 16991 30243
rect 16991 30209 17000 30243
rect 16948 30200 17000 30209
rect 17592 30200 17644 30252
rect 27528 30200 27580 30252
rect 12900 30064 12952 30116
rect 17132 30064 17184 30116
rect 9496 30039 9548 30048
rect 9496 30005 9505 30039
rect 9505 30005 9539 30039
rect 9539 30005 9548 30039
rect 9496 29996 9548 30005
rect 11612 30039 11664 30048
rect 11612 30005 11621 30039
rect 11621 30005 11655 30039
rect 11655 30005 11664 30039
rect 11612 29996 11664 30005
rect 16120 29996 16172 30048
rect 17040 29996 17092 30048
rect 17684 29996 17736 30048
rect 5688 29894 5740 29946
rect 5752 29894 5804 29946
rect 5816 29894 5868 29946
rect 5880 29894 5932 29946
rect 5944 29894 5996 29946
rect 15163 29894 15215 29946
rect 15227 29894 15279 29946
rect 15291 29894 15343 29946
rect 15355 29894 15407 29946
rect 15419 29894 15471 29946
rect 24639 29894 24691 29946
rect 24703 29894 24755 29946
rect 24767 29894 24819 29946
rect 24831 29894 24883 29946
rect 24895 29894 24947 29946
rect 14832 29792 14884 29844
rect 17040 29792 17092 29844
rect 17592 29767 17644 29776
rect 17592 29733 17601 29767
rect 17601 29733 17635 29767
rect 17635 29733 17644 29767
rect 17592 29724 17644 29733
rect 2964 29699 3016 29708
rect 2964 29665 2973 29699
rect 2973 29665 3007 29699
rect 3007 29665 3016 29699
rect 2964 29656 3016 29665
rect 4252 29699 4304 29708
rect 4252 29665 4261 29699
rect 4261 29665 4295 29699
rect 4295 29665 4304 29699
rect 4252 29656 4304 29665
rect 6644 29699 6696 29708
rect 6644 29665 6653 29699
rect 6653 29665 6687 29699
rect 6687 29665 6696 29699
rect 6644 29656 6696 29665
rect 11980 29656 12032 29708
rect 6368 29588 6420 29640
rect 9588 29588 9640 29640
rect 11520 29588 11572 29640
rect 12900 29631 12952 29640
rect 8024 29520 8076 29572
rect 9496 29520 9548 29572
rect 11612 29520 11664 29572
rect 12900 29597 12909 29631
rect 12909 29597 12943 29631
rect 12943 29597 12952 29631
rect 12900 29588 12952 29597
rect 13268 29631 13320 29640
rect 13268 29597 13277 29631
rect 13277 29597 13311 29631
rect 13311 29597 13320 29631
rect 13268 29588 13320 29597
rect 13636 29520 13688 29572
rect 14280 29520 14332 29572
rect 8300 29452 8352 29504
rect 9036 29495 9088 29504
rect 9036 29461 9045 29495
rect 9045 29461 9079 29495
rect 9079 29461 9088 29495
rect 9036 29452 9088 29461
rect 11704 29452 11756 29504
rect 12164 29452 12216 29504
rect 12624 29495 12676 29504
rect 12624 29461 12633 29495
rect 12633 29461 12667 29495
rect 12667 29461 12676 29495
rect 12624 29452 12676 29461
rect 14372 29452 14424 29504
rect 15660 29452 15712 29504
rect 16488 29520 16540 29572
rect 16764 29520 16816 29572
rect 17684 29520 17736 29572
rect 21456 29452 21508 29504
rect 10425 29350 10477 29402
rect 10489 29350 10541 29402
rect 10553 29350 10605 29402
rect 10617 29350 10669 29402
rect 10681 29350 10733 29402
rect 19901 29350 19953 29402
rect 19965 29350 20017 29402
rect 20029 29350 20081 29402
rect 20093 29350 20145 29402
rect 20157 29350 20209 29402
rect 8024 29291 8076 29300
rect 8024 29257 8033 29291
rect 8033 29257 8067 29291
rect 8067 29257 8076 29291
rect 8024 29248 8076 29257
rect 13636 29291 13688 29300
rect 8300 29180 8352 29232
rect 7564 28976 7616 29028
rect 9864 29180 9916 29232
rect 10232 29180 10284 29232
rect 9772 29112 9824 29164
rect 9956 29155 10008 29164
rect 9956 29121 9990 29155
rect 9990 29121 10008 29155
rect 9956 29112 10008 29121
rect 8760 29044 8812 29096
rect 9588 29044 9640 29096
rect 572 28908 624 28960
rect 1308 28908 1360 28960
rect 6460 28908 6512 28960
rect 9680 28908 9732 28960
rect 10048 28908 10100 28960
rect 11060 28951 11112 28960
rect 11060 28917 11069 28951
rect 11069 28917 11103 28951
rect 11103 28917 11112 28951
rect 11060 28908 11112 28917
rect 13636 29257 13645 29291
rect 13645 29257 13679 29291
rect 13679 29257 13688 29291
rect 13636 29248 13688 29257
rect 13912 29291 13964 29300
rect 13912 29257 13921 29291
rect 13921 29257 13955 29291
rect 13955 29257 13964 29291
rect 13912 29248 13964 29257
rect 14280 29248 14332 29300
rect 16764 29291 16816 29300
rect 16764 29257 16773 29291
rect 16773 29257 16807 29291
rect 16807 29257 16816 29291
rect 16764 29248 16816 29257
rect 12624 29180 12676 29232
rect 14372 29112 14424 29164
rect 14556 29180 14608 29232
rect 16120 29223 16172 29232
rect 16120 29189 16138 29223
rect 16138 29189 16172 29223
rect 16120 29180 16172 29189
rect 17408 29248 17460 29300
rect 11520 29044 11572 29096
rect 14740 29044 14792 29096
rect 14648 28976 14700 29028
rect 14832 28976 14884 29028
rect 15016 29019 15068 29028
rect 15016 28985 15025 29019
rect 15025 28985 15059 29019
rect 15059 28985 15068 29019
rect 15016 28976 15068 28985
rect 15660 29112 15712 29164
rect 17224 29155 17276 29164
rect 17224 29121 17234 29155
rect 17234 29121 17268 29155
rect 17268 29121 17276 29155
rect 17224 29112 17276 29121
rect 16488 29044 16540 29096
rect 17040 29087 17092 29096
rect 17040 29053 17049 29087
rect 17049 29053 17083 29087
rect 17083 29053 17092 29087
rect 17040 29044 17092 29053
rect 17132 29087 17184 29096
rect 17132 29053 17141 29087
rect 17141 29053 17175 29087
rect 17175 29053 17184 29087
rect 17132 29044 17184 29053
rect 14004 28908 14056 28960
rect 16580 28976 16632 29028
rect 17316 28976 17368 29028
rect 28816 28976 28868 29028
rect 30012 28908 30064 28960
rect 5688 28806 5740 28858
rect 5752 28806 5804 28858
rect 5816 28806 5868 28858
rect 5880 28806 5932 28858
rect 5944 28806 5996 28858
rect 15163 28806 15215 28858
rect 15227 28806 15279 28858
rect 15291 28806 15343 28858
rect 15355 28806 15407 28858
rect 15419 28806 15471 28858
rect 24639 28806 24691 28858
rect 24703 28806 24755 28858
rect 24767 28806 24819 28858
rect 24831 28806 24883 28858
rect 24895 28806 24947 28858
rect 9956 28704 10008 28756
rect 10048 28704 10100 28756
rect 12440 28747 12492 28756
rect 12440 28713 12449 28747
rect 12449 28713 12483 28747
rect 12483 28713 12492 28747
rect 12440 28704 12492 28713
rect 12900 28704 12952 28756
rect 14648 28704 14700 28756
rect 14740 28704 14792 28756
rect 7932 28500 7984 28552
rect 9864 28500 9916 28552
rect 11060 28636 11112 28688
rect 10048 28568 10100 28620
rect 17776 28636 17828 28688
rect 10232 28543 10284 28552
rect 10232 28509 10241 28543
rect 10241 28509 10275 28543
rect 10275 28509 10284 28543
rect 10232 28500 10284 28509
rect 12808 28568 12860 28620
rect 16120 28611 16172 28620
rect 10784 28543 10836 28552
rect 9772 28432 9824 28484
rect 10784 28509 10793 28543
rect 10793 28509 10827 28543
rect 10827 28509 10836 28543
rect 10784 28500 10836 28509
rect 12624 28543 12676 28552
rect 10600 28432 10652 28484
rect 12624 28509 12633 28543
rect 12633 28509 12667 28543
rect 12667 28509 12676 28543
rect 14740 28543 14792 28552
rect 12624 28500 12676 28509
rect 14740 28509 14749 28543
rect 14749 28509 14783 28543
rect 14783 28509 14792 28543
rect 14740 28500 14792 28509
rect 16120 28577 16129 28611
rect 16129 28577 16163 28611
rect 16163 28577 16172 28611
rect 16120 28568 16172 28577
rect 9864 28364 9916 28416
rect 10232 28364 10284 28416
rect 11244 28432 11296 28484
rect 17776 28500 17828 28552
rect 12256 28364 12308 28416
rect 14832 28364 14884 28416
rect 15568 28407 15620 28416
rect 15568 28373 15577 28407
rect 15577 28373 15611 28407
rect 15611 28373 15620 28407
rect 15568 28364 15620 28373
rect 15936 28407 15988 28416
rect 15936 28373 15945 28407
rect 15945 28373 15979 28407
rect 15979 28373 15988 28407
rect 15936 28364 15988 28373
rect 17040 28364 17092 28416
rect 17132 28364 17184 28416
rect 26332 28364 26384 28416
rect 10425 28262 10477 28314
rect 10489 28262 10541 28314
rect 10553 28262 10605 28314
rect 10617 28262 10669 28314
rect 10681 28262 10733 28314
rect 19901 28262 19953 28314
rect 19965 28262 20017 28314
rect 20029 28262 20081 28314
rect 20093 28262 20145 28314
rect 20157 28262 20209 28314
rect 4068 28092 4120 28144
rect 5540 28024 5592 28076
rect 5724 28067 5776 28076
rect 5724 28033 5733 28067
rect 5733 28033 5767 28067
rect 5767 28033 5776 28067
rect 5724 28024 5776 28033
rect 5172 27956 5224 28008
rect 7656 28160 7708 28212
rect 9772 28160 9824 28212
rect 6368 28067 6420 28076
rect 6368 28033 6377 28067
rect 6377 28033 6411 28067
rect 6411 28033 6420 28067
rect 6368 28024 6420 28033
rect 8944 28024 8996 28076
rect 9404 28024 9456 28076
rect 12072 28160 12124 28212
rect 14556 28160 14608 28212
rect 11980 28092 12032 28144
rect 12256 28092 12308 28144
rect 14188 28092 14240 28144
rect 5356 27888 5408 27940
rect 5724 27888 5776 27940
rect 6276 27820 6328 27872
rect 9128 27956 9180 28008
rect 13820 28024 13872 28076
rect 16488 28092 16540 28144
rect 14740 28067 14792 28076
rect 14740 28033 14749 28067
rect 14749 28033 14783 28067
rect 14783 28033 14792 28067
rect 14740 28024 14792 28033
rect 15844 28024 15896 28076
rect 16580 28024 16632 28076
rect 16948 28067 17000 28076
rect 16948 28033 16957 28067
rect 16957 28033 16991 28067
rect 16991 28033 17000 28067
rect 16948 28024 17000 28033
rect 17132 28067 17184 28076
rect 17132 28033 17140 28067
rect 17140 28033 17174 28067
rect 17174 28033 17184 28067
rect 17132 28024 17184 28033
rect 17224 28067 17276 28076
rect 17224 28033 17233 28067
rect 17233 28033 17267 28067
rect 17267 28033 17276 28067
rect 17224 28024 17276 28033
rect 20812 28067 20864 28076
rect 20812 28033 20821 28067
rect 20821 28033 20855 28067
rect 20855 28033 20864 28067
rect 20812 28024 20864 28033
rect 8668 27820 8720 27872
rect 9128 27820 9180 27872
rect 10140 27863 10192 27872
rect 10140 27829 10149 27863
rect 10149 27829 10183 27863
rect 10183 27829 10192 27863
rect 10140 27820 10192 27829
rect 10876 27820 10928 27872
rect 11520 27999 11572 28008
rect 11520 27965 11529 27999
rect 11529 27965 11563 27999
rect 11563 27965 11572 27999
rect 16488 27999 16540 28008
rect 11520 27956 11572 27965
rect 16488 27965 16497 27999
rect 16497 27965 16531 27999
rect 16531 27965 16540 27999
rect 16488 27956 16540 27965
rect 16856 27956 16908 28008
rect 12440 27820 12492 27872
rect 12992 27820 13044 27872
rect 13176 27863 13228 27872
rect 13176 27829 13185 27863
rect 13185 27829 13219 27863
rect 13219 27829 13228 27863
rect 13176 27820 13228 27829
rect 14924 27863 14976 27872
rect 14924 27829 14933 27863
rect 14933 27829 14967 27863
rect 14967 27829 14976 27863
rect 14924 27820 14976 27829
rect 15752 27820 15804 27872
rect 18880 27820 18932 27872
rect 22100 27820 22152 27872
rect 5688 27718 5740 27770
rect 5752 27718 5804 27770
rect 5816 27718 5868 27770
rect 5880 27718 5932 27770
rect 5944 27718 5996 27770
rect 15163 27718 15215 27770
rect 15227 27718 15279 27770
rect 15291 27718 15343 27770
rect 15355 27718 15407 27770
rect 15419 27718 15471 27770
rect 24639 27718 24691 27770
rect 24703 27718 24755 27770
rect 24767 27718 24819 27770
rect 24831 27718 24883 27770
rect 24895 27718 24947 27770
rect 5540 27616 5592 27668
rect 6460 27616 6512 27668
rect 9220 27616 9272 27668
rect 9864 27616 9916 27668
rect 10784 27616 10836 27668
rect 10876 27616 10928 27668
rect 14648 27616 14700 27668
rect 14924 27616 14976 27668
rect 8944 27591 8996 27600
rect 8944 27557 8953 27591
rect 8953 27557 8987 27591
rect 8987 27557 8996 27591
rect 8944 27548 8996 27557
rect 7472 27523 7524 27532
rect 7472 27489 7481 27523
rect 7481 27489 7515 27523
rect 7515 27489 7524 27523
rect 7472 27480 7524 27489
rect 7656 27523 7708 27532
rect 7656 27489 7665 27523
rect 7665 27489 7699 27523
rect 7699 27489 7708 27523
rect 7656 27480 7708 27489
rect 9680 27548 9732 27600
rect 9128 27455 9180 27464
rect 9128 27421 9137 27455
rect 9137 27421 9171 27455
rect 9171 27421 9180 27455
rect 9128 27412 9180 27421
rect 9220 27412 9272 27464
rect 10232 27480 10284 27532
rect 11060 27548 11112 27600
rect 11244 27591 11296 27600
rect 11244 27557 11253 27591
rect 11253 27557 11287 27591
rect 11287 27557 11296 27591
rect 11244 27548 11296 27557
rect 11980 27548 12032 27600
rect 9680 27455 9732 27464
rect 9680 27421 9689 27455
rect 9689 27421 9723 27455
rect 9723 27421 9732 27455
rect 9864 27455 9916 27464
rect 9680 27412 9732 27421
rect 9864 27421 9873 27455
rect 9873 27421 9907 27455
rect 9907 27421 9916 27455
rect 9864 27412 9916 27421
rect 10968 27412 11020 27464
rect 12992 27548 13044 27600
rect 13820 27548 13872 27600
rect 13268 27480 13320 27532
rect 14832 27548 14884 27600
rect 15292 27548 15344 27600
rect 14280 27523 14332 27532
rect 12532 27412 12584 27464
rect 12900 27412 12952 27464
rect 13176 27412 13228 27464
rect 13728 27455 13780 27464
rect 13728 27421 13737 27455
rect 13737 27421 13771 27455
rect 13771 27421 13780 27455
rect 13728 27412 13780 27421
rect 14280 27489 14289 27523
rect 14289 27489 14323 27523
rect 14323 27489 14332 27523
rect 14280 27480 14332 27489
rect 14556 27480 14608 27532
rect 15844 27591 15896 27600
rect 15844 27557 15853 27591
rect 15853 27557 15887 27591
rect 15887 27557 15896 27591
rect 15844 27548 15896 27557
rect 15384 27455 15436 27464
rect 15384 27421 15393 27455
rect 15393 27421 15427 27455
rect 15427 27421 15436 27455
rect 15752 27480 15804 27532
rect 16856 27548 16908 27600
rect 15384 27412 15436 27421
rect 16580 27455 16632 27464
rect 16580 27421 16589 27455
rect 16589 27421 16623 27455
rect 16623 27421 16632 27455
rect 16580 27412 16632 27421
rect 16672 27412 16724 27464
rect 7104 27344 7156 27396
rect 4068 27276 4120 27328
rect 6736 27276 6788 27328
rect 7748 27319 7800 27328
rect 7748 27285 7757 27319
rect 7757 27285 7791 27319
rect 7791 27285 7800 27319
rect 7748 27276 7800 27285
rect 8852 27276 8904 27328
rect 9588 27276 9640 27328
rect 12532 27276 12584 27328
rect 12900 27276 12952 27328
rect 13268 27319 13320 27328
rect 13268 27285 13277 27319
rect 13277 27285 13311 27319
rect 13311 27285 13320 27319
rect 13268 27276 13320 27285
rect 13360 27276 13412 27328
rect 14740 27276 14792 27328
rect 16396 27344 16448 27396
rect 17040 27412 17092 27464
rect 22652 27548 22704 27600
rect 20260 27480 20312 27532
rect 20444 27480 20496 27532
rect 18880 27455 18932 27464
rect 18880 27421 18889 27455
rect 18889 27421 18923 27455
rect 18923 27421 18932 27455
rect 18880 27412 18932 27421
rect 21088 27455 21140 27464
rect 21088 27421 21097 27455
rect 21097 27421 21131 27455
rect 21131 27421 21140 27455
rect 21088 27412 21140 27421
rect 17224 27344 17276 27396
rect 18788 27344 18840 27396
rect 19248 27344 19300 27396
rect 20720 27344 20772 27396
rect 21548 27344 21600 27396
rect 22100 27344 22152 27396
rect 27436 27276 27488 27328
rect 10425 27174 10477 27226
rect 10489 27174 10541 27226
rect 10553 27174 10605 27226
rect 10617 27174 10669 27226
rect 10681 27174 10733 27226
rect 19901 27174 19953 27226
rect 19965 27174 20017 27226
rect 20029 27174 20081 27226
rect 20093 27174 20145 27226
rect 20157 27174 20209 27226
rect 6092 27115 6144 27124
rect 6092 27081 6101 27115
rect 6101 27081 6135 27115
rect 6135 27081 6144 27115
rect 6092 27072 6144 27081
rect 7104 27115 7156 27124
rect 7104 27081 7113 27115
rect 7113 27081 7147 27115
rect 7147 27081 7156 27115
rect 7104 27072 7156 27081
rect 8852 27115 8904 27124
rect 8852 27081 8861 27115
rect 8861 27081 8895 27115
rect 8895 27081 8904 27115
rect 8852 27072 8904 27081
rect 12072 27072 12124 27124
rect 14464 27115 14516 27124
rect 14464 27081 14473 27115
rect 14473 27081 14507 27115
rect 14507 27081 14516 27115
rect 15844 27115 15896 27124
rect 14464 27072 14516 27081
rect 15844 27081 15853 27115
rect 15853 27081 15887 27115
rect 15887 27081 15896 27115
rect 15844 27072 15896 27081
rect 16948 27072 17000 27124
rect 4160 27004 4212 27056
rect 4620 26936 4672 26988
rect 6368 27004 6420 27056
rect 5540 26936 5592 26988
rect 7472 27004 7524 27056
rect 9128 27004 9180 27056
rect 6736 26936 6788 26988
rect 9404 26936 9456 26988
rect 10048 26936 10100 26988
rect 10968 26936 11020 26988
rect 12256 26979 12308 26988
rect 12256 26945 12265 26979
rect 12265 26945 12299 26979
rect 12299 26945 12308 26979
rect 12256 26936 12308 26945
rect 12348 26936 12400 26988
rect 15936 27004 15988 27056
rect 4988 26732 5040 26784
rect 8576 26868 8628 26920
rect 9588 26868 9640 26920
rect 12072 26911 12124 26920
rect 12072 26877 12081 26911
rect 12081 26877 12115 26911
rect 12115 26877 12124 26911
rect 12072 26868 12124 26877
rect 12532 26868 12584 26920
rect 16304 26936 16356 26988
rect 20812 27072 20864 27124
rect 20444 27047 20496 27056
rect 20444 27013 20453 27047
rect 20453 27013 20487 27047
rect 20487 27013 20496 27047
rect 20444 27004 20496 27013
rect 20352 26979 20404 26988
rect 20352 26945 20356 26979
rect 20356 26945 20390 26979
rect 20390 26945 20404 26979
rect 20352 26936 20404 26945
rect 20536 26979 20588 26988
rect 20536 26945 20545 26979
rect 20545 26945 20579 26979
rect 20579 26945 20588 26979
rect 20536 26936 20588 26945
rect 20812 26936 20864 26988
rect 14280 26868 14332 26920
rect 14832 26868 14884 26920
rect 16120 26868 16172 26920
rect 16856 26868 16908 26920
rect 27528 27072 27580 27124
rect 22652 27004 22704 27056
rect 20996 26979 21048 26988
rect 20996 26945 21005 26979
rect 21005 26945 21039 26979
rect 21039 26945 21048 26979
rect 21180 26979 21232 26988
rect 20996 26936 21048 26945
rect 21180 26945 21189 26979
rect 21189 26945 21223 26979
rect 21223 26945 21232 26979
rect 21180 26936 21232 26945
rect 21456 26979 21508 26988
rect 21456 26945 21459 26979
rect 21459 26945 21508 26979
rect 21456 26936 21508 26945
rect 11980 26800 12032 26852
rect 18972 26800 19024 26852
rect 20720 26800 20772 26852
rect 21548 26843 21600 26852
rect 21548 26809 21557 26843
rect 21557 26809 21591 26843
rect 21591 26809 21600 26843
rect 21548 26800 21600 26809
rect 9680 26775 9732 26784
rect 9680 26741 9689 26775
rect 9689 26741 9723 26775
rect 9723 26741 9732 26775
rect 9680 26732 9732 26741
rect 9864 26775 9916 26784
rect 9864 26741 9873 26775
rect 9873 26741 9907 26775
rect 9907 26741 9916 26775
rect 9864 26732 9916 26741
rect 10232 26732 10284 26784
rect 12532 26732 12584 26784
rect 13728 26732 13780 26784
rect 14004 26775 14056 26784
rect 14004 26741 14013 26775
rect 14013 26741 14047 26775
rect 14047 26741 14056 26775
rect 14004 26732 14056 26741
rect 15752 26732 15804 26784
rect 16672 26732 16724 26784
rect 17592 26732 17644 26784
rect 20260 26732 20312 26784
rect 20536 26732 20588 26784
rect 5688 26630 5740 26682
rect 5752 26630 5804 26682
rect 5816 26630 5868 26682
rect 5880 26630 5932 26682
rect 5944 26630 5996 26682
rect 15163 26630 15215 26682
rect 15227 26630 15279 26682
rect 15291 26630 15343 26682
rect 15355 26630 15407 26682
rect 15419 26630 15471 26682
rect 24639 26630 24691 26682
rect 24703 26630 24755 26682
rect 24767 26630 24819 26682
rect 24831 26630 24883 26682
rect 24895 26630 24947 26682
rect 4620 26528 4672 26580
rect 5540 26528 5592 26580
rect 7288 26528 7340 26580
rect 7748 26528 7800 26580
rect 10232 26528 10284 26580
rect 16856 26528 16908 26580
rect 17592 26528 17644 26580
rect 23848 26528 23900 26580
rect 5356 26460 5408 26512
rect 6184 26460 6236 26512
rect 6368 26460 6420 26512
rect 4988 26367 5040 26376
rect 4988 26333 4997 26367
rect 4997 26333 5031 26367
rect 5031 26333 5040 26367
rect 4988 26324 5040 26333
rect 5172 26367 5224 26376
rect 5172 26333 5181 26367
rect 5181 26333 5215 26367
rect 5215 26333 5224 26367
rect 5172 26324 5224 26333
rect 6920 26392 6972 26444
rect 12348 26460 12400 26512
rect 9588 26435 9640 26444
rect 9588 26401 9597 26435
rect 9597 26401 9631 26435
rect 9631 26401 9640 26435
rect 9588 26392 9640 26401
rect 12072 26392 12124 26444
rect 13176 26392 13228 26444
rect 14832 26392 14884 26444
rect 15108 26392 15160 26444
rect 15660 26435 15712 26444
rect 15660 26401 15669 26435
rect 15669 26401 15703 26435
rect 15703 26401 15712 26435
rect 15660 26392 15712 26401
rect 5724 26324 5776 26376
rect 6092 26367 6144 26376
rect 6092 26333 6101 26367
rect 6101 26333 6135 26367
rect 6135 26333 6144 26367
rect 6368 26367 6420 26376
rect 6092 26324 6144 26333
rect 6368 26333 6377 26367
rect 6377 26333 6411 26367
rect 6411 26333 6420 26367
rect 6368 26324 6420 26333
rect 6460 26367 6512 26376
rect 6460 26333 6470 26367
rect 6470 26333 6504 26367
rect 6504 26333 6512 26367
rect 6460 26324 6512 26333
rect 6736 26324 6788 26376
rect 9036 26324 9088 26376
rect 9864 26324 9916 26376
rect 19248 26503 19300 26512
rect 16396 26392 16448 26444
rect 16948 26435 17000 26444
rect 16948 26401 16957 26435
rect 16957 26401 16991 26435
rect 16991 26401 17000 26435
rect 19248 26469 19257 26503
rect 19257 26469 19291 26503
rect 19291 26469 19300 26503
rect 19248 26460 19300 26469
rect 20352 26460 20404 26512
rect 21548 26460 21600 26512
rect 16948 26392 17000 26401
rect 16580 26367 16632 26376
rect 16580 26333 16589 26367
rect 16589 26333 16623 26367
rect 16623 26333 16632 26367
rect 16580 26324 16632 26333
rect 16764 26367 16816 26376
rect 16764 26333 16772 26367
rect 16772 26333 16806 26367
rect 16806 26333 16816 26367
rect 16764 26324 16816 26333
rect 18972 26392 19024 26444
rect 22100 26392 22152 26444
rect 23480 26435 23532 26444
rect 23480 26401 23489 26435
rect 23489 26401 23523 26435
rect 23523 26401 23532 26435
rect 23480 26392 23532 26401
rect 18880 26367 18932 26376
rect 7380 26256 7432 26308
rect 7656 26256 7708 26308
rect 12716 26256 12768 26308
rect 13728 26256 13780 26308
rect 16304 26256 16356 26308
rect 16396 26256 16448 26308
rect 18880 26333 18889 26367
rect 18889 26333 18923 26367
rect 18923 26333 18932 26367
rect 18880 26324 18932 26333
rect 5724 26188 5776 26240
rect 6276 26188 6328 26240
rect 9680 26188 9732 26240
rect 9864 26188 9916 26240
rect 16120 26231 16172 26240
rect 16120 26197 16129 26231
rect 16129 26197 16163 26231
rect 16163 26197 16172 26231
rect 16120 26188 16172 26197
rect 17960 26256 18012 26308
rect 19524 26299 19576 26308
rect 19524 26265 19533 26299
rect 19533 26265 19567 26299
rect 19567 26265 19576 26299
rect 19524 26256 19576 26265
rect 21088 26188 21140 26240
rect 24492 26324 24544 26376
rect 21916 26256 21968 26308
rect 23020 26256 23072 26308
rect 23388 26188 23440 26240
rect 24400 26231 24452 26240
rect 24400 26197 24409 26231
rect 24409 26197 24443 26231
rect 24443 26197 24452 26231
rect 24400 26188 24452 26197
rect 10425 26086 10477 26138
rect 10489 26086 10541 26138
rect 10553 26086 10605 26138
rect 10617 26086 10669 26138
rect 10681 26086 10733 26138
rect 19901 26086 19953 26138
rect 19965 26086 20017 26138
rect 20029 26086 20081 26138
rect 20093 26086 20145 26138
rect 20157 26086 20209 26138
rect 5356 25984 5408 26036
rect 5448 25984 5500 26036
rect 6460 25984 6512 26036
rect 7380 26027 7432 26036
rect 7380 25993 7389 26027
rect 7389 25993 7423 26027
rect 7423 25993 7432 26027
rect 7380 25984 7432 25993
rect 8300 25984 8352 26036
rect 4804 25891 4856 25900
rect 4804 25857 4813 25891
rect 4813 25857 4847 25891
rect 4847 25857 4856 25891
rect 4804 25848 4856 25857
rect 4252 25644 4304 25696
rect 7104 25916 7156 25968
rect 12164 25959 12216 25968
rect 5724 25848 5776 25900
rect 6736 25891 6788 25900
rect 6736 25857 6745 25891
rect 6745 25857 6779 25891
rect 6779 25857 6788 25891
rect 6736 25848 6788 25857
rect 7288 25891 7340 25900
rect 7288 25857 7297 25891
rect 7297 25857 7331 25891
rect 7331 25857 7340 25891
rect 7288 25848 7340 25857
rect 7932 25848 7984 25900
rect 6092 25780 6144 25832
rect 6368 25780 6420 25832
rect 8576 25823 8628 25832
rect 5172 25712 5224 25764
rect 6920 25712 6972 25764
rect 8576 25789 8585 25823
rect 8585 25789 8619 25823
rect 8619 25789 8628 25823
rect 8576 25780 8628 25789
rect 9128 25712 9180 25764
rect 10600 25848 10652 25900
rect 9772 25780 9824 25832
rect 12164 25925 12173 25959
rect 12173 25925 12207 25959
rect 12207 25925 12216 25959
rect 12164 25916 12216 25925
rect 15016 26027 15068 26036
rect 15016 25993 15025 26027
rect 15025 25993 15059 26027
rect 15059 25993 15068 26027
rect 15016 25984 15068 25993
rect 19340 26027 19392 26036
rect 19340 25993 19349 26027
rect 19349 25993 19383 26027
rect 19383 25993 19392 26027
rect 19340 25984 19392 25993
rect 22100 25984 22152 26036
rect 20076 25916 20128 25968
rect 27528 25984 27580 26036
rect 24400 25916 24452 25968
rect 12348 25848 12400 25900
rect 16396 25848 16448 25900
rect 21640 25848 21692 25900
rect 22284 25891 22336 25900
rect 12072 25823 12124 25832
rect 12072 25789 12081 25823
rect 12081 25789 12115 25823
rect 12115 25789 12124 25823
rect 12072 25780 12124 25789
rect 12808 25780 12860 25832
rect 14280 25823 14332 25832
rect 14280 25789 14289 25823
rect 14289 25789 14323 25823
rect 14323 25789 14332 25823
rect 15108 25823 15160 25832
rect 14280 25780 14332 25789
rect 15108 25789 15117 25823
rect 15117 25789 15151 25823
rect 15151 25789 15160 25823
rect 15108 25780 15160 25789
rect 20812 25823 20864 25832
rect 20812 25789 20821 25823
rect 20821 25789 20855 25823
rect 20855 25789 20864 25823
rect 20812 25780 20864 25789
rect 21088 25823 21140 25832
rect 21088 25789 21097 25823
rect 21097 25789 21131 25823
rect 21131 25789 21140 25823
rect 21088 25780 21140 25789
rect 4712 25687 4764 25696
rect 4712 25653 4721 25687
rect 4721 25653 4755 25687
rect 4755 25653 4764 25687
rect 4712 25644 4764 25653
rect 6736 25644 6788 25696
rect 8944 25644 8996 25696
rect 11520 25644 11572 25696
rect 19524 25712 19576 25764
rect 21916 25755 21968 25764
rect 21916 25721 21925 25755
rect 21925 25721 21959 25755
rect 21959 25721 21968 25755
rect 21916 25712 21968 25721
rect 22284 25857 22293 25891
rect 22293 25857 22327 25891
rect 22327 25857 22336 25891
rect 22284 25848 22336 25857
rect 22744 25848 22796 25900
rect 23388 25891 23440 25900
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23388 25848 23440 25857
rect 13820 25644 13872 25696
rect 13912 25644 13964 25696
rect 14832 25644 14884 25696
rect 16028 25644 16080 25696
rect 16764 25644 16816 25696
rect 17592 25644 17644 25696
rect 22008 25644 22060 25696
rect 5688 25542 5740 25594
rect 5752 25542 5804 25594
rect 5816 25542 5868 25594
rect 5880 25542 5932 25594
rect 5944 25542 5996 25594
rect 15163 25542 15215 25594
rect 15227 25542 15279 25594
rect 15291 25542 15343 25594
rect 15355 25542 15407 25594
rect 15419 25542 15471 25594
rect 24639 25542 24691 25594
rect 24703 25542 24755 25594
rect 24767 25542 24819 25594
rect 24831 25542 24883 25594
rect 24895 25542 24947 25594
rect 4068 25440 4120 25492
rect 7564 25440 7616 25492
rect 7932 25483 7984 25492
rect 7932 25449 7941 25483
rect 7941 25449 7975 25483
rect 7975 25449 7984 25483
rect 7932 25440 7984 25449
rect 10600 25483 10652 25492
rect 10600 25449 10609 25483
rect 10609 25449 10643 25483
rect 10643 25449 10652 25483
rect 10600 25440 10652 25449
rect 12256 25440 12308 25492
rect 5172 25372 5224 25424
rect 9680 25372 9732 25424
rect 4160 25347 4212 25356
rect 4160 25313 4169 25347
rect 4169 25313 4203 25347
rect 4203 25313 4212 25347
rect 4160 25304 4212 25313
rect 7472 25304 7524 25356
rect 4712 25236 4764 25288
rect 9864 25236 9916 25288
rect 14648 25440 14700 25492
rect 20076 25440 20128 25492
rect 20812 25440 20864 25492
rect 23020 25483 23072 25492
rect 23020 25449 23029 25483
rect 23029 25449 23063 25483
rect 23063 25449 23072 25483
rect 23020 25440 23072 25449
rect 23480 25440 23532 25492
rect 24492 25440 24544 25492
rect 14832 25372 14884 25424
rect 19524 25372 19576 25424
rect 11336 25347 11388 25356
rect 11336 25313 11345 25347
rect 11345 25313 11379 25347
rect 11379 25313 11388 25347
rect 11336 25304 11388 25313
rect 11520 25347 11572 25356
rect 11520 25313 11529 25347
rect 11529 25313 11563 25347
rect 11563 25313 11572 25347
rect 11520 25304 11572 25313
rect 12808 25347 12860 25356
rect 12808 25313 12817 25347
rect 12817 25313 12851 25347
rect 12851 25313 12860 25347
rect 12808 25304 12860 25313
rect 13636 25304 13688 25356
rect 14372 25347 14424 25356
rect 4804 25168 4856 25220
rect 8668 25168 8720 25220
rect 9588 25168 9640 25220
rect 10324 25279 10376 25288
rect 10324 25245 10333 25279
rect 10333 25245 10367 25279
rect 10367 25245 10376 25279
rect 10324 25236 10376 25245
rect 14372 25313 14381 25347
rect 14381 25313 14415 25347
rect 14415 25313 14424 25347
rect 14372 25304 14424 25313
rect 16488 25304 16540 25356
rect 17960 25304 18012 25356
rect 19340 25304 19392 25356
rect 14280 25236 14332 25288
rect 16580 25236 16632 25288
rect 19616 25279 19668 25288
rect 19616 25245 19625 25279
rect 19625 25245 19659 25279
rect 19659 25245 19668 25279
rect 19616 25236 19668 25245
rect 6828 25100 6880 25152
rect 7748 25100 7800 25152
rect 9312 25100 9364 25152
rect 9864 25143 9916 25152
rect 9864 25109 9873 25143
rect 9873 25109 9907 25143
rect 9907 25109 9916 25143
rect 9864 25100 9916 25109
rect 9956 25100 10008 25152
rect 10232 25100 10284 25152
rect 13084 25143 13136 25152
rect 13084 25109 13093 25143
rect 13093 25109 13127 25143
rect 13127 25109 13136 25143
rect 15476 25211 15528 25220
rect 15476 25177 15485 25211
rect 15485 25177 15519 25211
rect 15519 25177 15528 25211
rect 15476 25168 15528 25177
rect 17408 25211 17460 25220
rect 17408 25177 17417 25211
rect 17417 25177 17451 25211
rect 17451 25177 17460 25211
rect 17408 25168 17460 25177
rect 19800 25168 19852 25220
rect 13084 25100 13136 25109
rect 14832 25143 14884 25152
rect 14832 25109 14841 25143
rect 14841 25109 14875 25143
rect 14875 25109 14884 25143
rect 14832 25100 14884 25109
rect 18052 25100 18104 25152
rect 21640 25304 21692 25356
rect 21916 25236 21968 25288
rect 22560 25279 22612 25288
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 22560 25236 22612 25245
rect 22100 25100 22152 25152
rect 22560 25100 22612 25152
rect 24400 25279 24452 25288
rect 24400 25245 24409 25279
rect 24409 25245 24443 25279
rect 24443 25245 24452 25279
rect 24400 25236 24452 25245
rect 10425 24998 10477 25050
rect 10489 24998 10541 25050
rect 10553 24998 10605 25050
rect 10617 24998 10669 25050
rect 10681 24998 10733 25050
rect 19901 24998 19953 25050
rect 19965 24998 20017 25050
rect 20029 24998 20081 25050
rect 20093 24998 20145 25050
rect 20157 24998 20209 25050
rect 9864 24896 9916 24948
rect 10324 24896 10376 24948
rect 13084 24896 13136 24948
rect 16580 24896 16632 24948
rect 19800 24896 19852 24948
rect 2688 24828 2740 24880
rect 4160 24828 4212 24880
rect 4620 24828 4672 24880
rect 1400 24692 1452 24744
rect 3700 24735 3752 24744
rect 3700 24701 3709 24735
rect 3709 24701 3743 24735
rect 3743 24701 3752 24735
rect 3700 24692 3752 24701
rect 3976 24692 4028 24744
rect 3700 24556 3752 24608
rect 5540 24760 5592 24812
rect 6644 24803 6696 24812
rect 6644 24769 6678 24803
rect 6678 24769 6696 24803
rect 6644 24760 6696 24769
rect 6920 24760 6972 24812
rect 9496 24760 9548 24812
rect 12256 24828 12308 24880
rect 13452 24828 13504 24880
rect 14556 24871 14608 24880
rect 14556 24837 14565 24871
rect 14565 24837 14599 24871
rect 14599 24837 14608 24871
rect 14556 24828 14608 24837
rect 14648 24871 14700 24880
rect 14648 24837 14657 24871
rect 14657 24837 14691 24871
rect 14691 24837 14700 24871
rect 14648 24828 14700 24837
rect 14924 24828 14976 24880
rect 10324 24803 10376 24812
rect 8668 24735 8720 24744
rect 8668 24701 8677 24735
rect 8677 24701 8711 24735
rect 8711 24701 8720 24735
rect 8668 24692 8720 24701
rect 10324 24769 10333 24803
rect 10333 24769 10367 24803
rect 10367 24769 10376 24803
rect 10324 24760 10376 24769
rect 11336 24692 11388 24744
rect 12072 24735 12124 24744
rect 12072 24701 12081 24735
rect 12081 24701 12115 24735
rect 12115 24701 12124 24735
rect 12072 24692 12124 24701
rect 7748 24599 7800 24608
rect 7748 24565 7757 24599
rect 7757 24565 7791 24599
rect 7791 24565 7800 24599
rect 7748 24556 7800 24565
rect 9680 24624 9732 24676
rect 10232 24624 10284 24676
rect 10600 24624 10652 24676
rect 11428 24624 11480 24676
rect 14372 24624 14424 24676
rect 8852 24556 8904 24608
rect 15108 24803 15160 24812
rect 15108 24769 15117 24803
rect 15117 24769 15151 24803
rect 15151 24769 15160 24803
rect 15108 24760 15160 24769
rect 15660 24760 15712 24812
rect 22560 24828 22612 24880
rect 16212 24760 16264 24812
rect 16672 24760 16724 24812
rect 18052 24760 18104 24812
rect 18236 24803 18288 24812
rect 18236 24769 18270 24803
rect 18270 24769 18288 24803
rect 18236 24760 18288 24769
rect 19708 24760 19760 24812
rect 17960 24735 18012 24744
rect 17960 24701 17969 24735
rect 17969 24701 18003 24735
rect 18003 24701 18012 24735
rect 17960 24692 18012 24701
rect 15476 24624 15528 24676
rect 17408 24624 17460 24676
rect 19432 24624 19484 24676
rect 21272 24692 21324 24744
rect 21456 24803 21508 24812
rect 21456 24769 21465 24803
rect 21465 24769 21499 24803
rect 21499 24769 21508 24803
rect 21456 24760 21508 24769
rect 22192 24760 22244 24812
rect 21640 24667 21692 24676
rect 21640 24633 21649 24667
rect 21649 24633 21683 24667
rect 21683 24633 21692 24667
rect 21640 24624 21692 24633
rect 21732 24624 21784 24676
rect 22008 24667 22060 24676
rect 22008 24633 22017 24667
rect 22017 24633 22051 24667
rect 22051 24633 22060 24667
rect 22008 24624 22060 24633
rect 24400 24760 24452 24812
rect 24492 24692 24544 24744
rect 15016 24556 15068 24608
rect 17684 24556 17736 24608
rect 19248 24556 19300 24608
rect 20260 24556 20312 24608
rect 20904 24556 20956 24608
rect 21916 24556 21968 24608
rect 23756 24556 23808 24608
rect 25320 24599 25372 24608
rect 25320 24565 25329 24599
rect 25329 24565 25363 24599
rect 25363 24565 25372 24599
rect 25320 24556 25372 24565
rect 25872 24599 25924 24608
rect 25872 24565 25881 24599
rect 25881 24565 25915 24599
rect 25915 24565 25924 24599
rect 25872 24556 25924 24565
rect 5688 24454 5740 24506
rect 5752 24454 5804 24506
rect 5816 24454 5868 24506
rect 5880 24454 5932 24506
rect 5944 24454 5996 24506
rect 15163 24454 15215 24506
rect 15227 24454 15279 24506
rect 15291 24454 15343 24506
rect 15355 24454 15407 24506
rect 15419 24454 15471 24506
rect 24639 24454 24691 24506
rect 24703 24454 24755 24506
rect 24767 24454 24819 24506
rect 24831 24454 24883 24506
rect 24895 24454 24947 24506
rect 2688 24395 2740 24404
rect 2688 24361 2697 24395
rect 2697 24361 2731 24395
rect 2731 24361 2740 24395
rect 2688 24352 2740 24361
rect 6092 24352 6144 24404
rect 6368 24395 6420 24404
rect 6368 24361 6377 24395
rect 6377 24361 6411 24395
rect 6411 24361 6420 24395
rect 6368 24352 6420 24361
rect 6644 24352 6696 24404
rect 8300 24352 8352 24404
rect 9496 24352 9548 24404
rect 9772 24327 9824 24336
rect 2320 24148 2372 24200
rect 7748 24216 7800 24268
rect 6828 24191 6880 24200
rect 6828 24157 6837 24191
rect 6837 24157 6871 24191
rect 6871 24157 6880 24191
rect 6828 24148 6880 24157
rect 6368 24080 6420 24132
rect 6736 24080 6788 24132
rect 9772 24293 9781 24327
rect 9781 24293 9815 24327
rect 9815 24293 9824 24327
rect 9772 24284 9824 24293
rect 9220 24259 9272 24268
rect 9220 24225 9229 24259
rect 9229 24225 9263 24259
rect 9263 24225 9272 24259
rect 9220 24216 9272 24225
rect 9312 24259 9364 24268
rect 9312 24225 9321 24259
rect 9321 24225 9355 24259
rect 9355 24225 9364 24259
rect 9312 24216 9364 24225
rect 9588 24216 9640 24268
rect 8944 24183 8996 24200
rect 8944 24149 8950 24183
rect 8950 24149 8984 24183
rect 8984 24149 8996 24183
rect 8944 24148 8996 24149
rect 9036 24145 9088 24197
rect 9680 24148 9732 24200
rect 10048 24352 10100 24404
rect 10784 24352 10836 24404
rect 11428 24395 11480 24404
rect 11428 24361 11437 24395
rect 11437 24361 11471 24395
rect 11471 24361 11480 24395
rect 11428 24352 11480 24361
rect 14372 24352 14424 24404
rect 16672 24395 16724 24404
rect 14464 24284 14516 24336
rect 16672 24361 16681 24395
rect 16681 24361 16715 24395
rect 16715 24361 16724 24395
rect 16672 24352 16724 24361
rect 18236 24352 18288 24404
rect 21916 24352 21968 24404
rect 26148 24352 26200 24404
rect 26884 24352 26936 24404
rect 27436 24352 27488 24404
rect 10600 24148 10652 24200
rect 10784 24080 10836 24132
rect 4068 24012 4120 24064
rect 6920 24012 6972 24064
rect 7380 24055 7432 24064
rect 7380 24021 7389 24055
rect 7389 24021 7423 24055
rect 7423 24021 7432 24055
rect 7380 24012 7432 24021
rect 8484 24012 8536 24064
rect 8852 24012 8904 24064
rect 13452 24191 13504 24200
rect 12164 24080 12216 24132
rect 12256 24012 12308 24064
rect 13452 24157 13461 24191
rect 13461 24157 13495 24191
rect 13495 24157 13504 24191
rect 13452 24148 13504 24157
rect 13912 24148 13964 24200
rect 14096 24191 14148 24200
rect 14096 24157 14105 24191
rect 14105 24157 14139 24191
rect 14139 24157 14148 24191
rect 14096 24148 14148 24157
rect 14924 24216 14976 24268
rect 18236 24216 18288 24268
rect 14832 24191 14884 24200
rect 13544 24123 13596 24132
rect 13544 24089 13553 24123
rect 13553 24089 13587 24123
rect 13587 24089 13596 24123
rect 14832 24157 14841 24191
rect 14841 24157 14875 24191
rect 14875 24157 14884 24191
rect 14832 24148 14884 24157
rect 16672 24148 16724 24200
rect 17408 24148 17460 24200
rect 17868 24148 17920 24200
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 19432 24191 19484 24200
rect 19432 24157 19441 24191
rect 19441 24157 19475 24191
rect 19475 24157 19484 24191
rect 19432 24148 19484 24157
rect 21364 24148 21416 24200
rect 21732 24148 21784 24200
rect 13544 24080 13596 24089
rect 17684 24080 17736 24132
rect 14096 24012 14148 24064
rect 14556 24012 14608 24064
rect 18144 24012 18196 24064
rect 19800 24080 19852 24132
rect 21824 24123 21876 24132
rect 21824 24089 21833 24123
rect 21833 24089 21867 24123
rect 21867 24089 21876 24123
rect 21824 24080 21876 24089
rect 22008 24284 22060 24336
rect 23664 24216 23716 24268
rect 25228 24216 25280 24268
rect 19524 24055 19576 24064
rect 19524 24021 19533 24055
rect 19533 24021 19567 24055
rect 19567 24021 19576 24055
rect 19524 24012 19576 24021
rect 19708 24012 19760 24064
rect 20628 24012 20680 24064
rect 21272 24055 21324 24064
rect 21272 24021 21281 24055
rect 21281 24021 21315 24055
rect 21315 24021 21324 24055
rect 21272 24012 21324 24021
rect 21548 24012 21600 24064
rect 21640 24012 21692 24064
rect 23756 24148 23808 24200
rect 26056 24148 26108 24200
rect 26700 24191 26752 24200
rect 26700 24157 26709 24191
rect 26709 24157 26743 24191
rect 26743 24157 26752 24191
rect 26700 24148 26752 24157
rect 27344 24191 27396 24200
rect 24032 24080 24084 24132
rect 25320 24080 25372 24132
rect 26792 24123 26844 24132
rect 25596 24012 25648 24064
rect 26148 24055 26200 24064
rect 26148 24021 26157 24055
rect 26157 24021 26191 24055
rect 26191 24021 26200 24055
rect 26148 24012 26200 24021
rect 26792 24089 26801 24123
rect 26801 24089 26835 24123
rect 26835 24089 26844 24123
rect 26792 24080 26844 24089
rect 27344 24157 27353 24191
rect 27353 24157 27387 24191
rect 27387 24157 27396 24191
rect 27344 24148 27396 24157
rect 27620 24123 27672 24132
rect 27620 24089 27629 24123
rect 27629 24089 27663 24123
rect 27663 24089 27672 24123
rect 27620 24080 27672 24089
rect 28632 24080 28684 24132
rect 27068 24055 27120 24064
rect 27068 24021 27077 24055
rect 27077 24021 27111 24055
rect 27111 24021 27120 24055
rect 27068 24012 27120 24021
rect 10425 23910 10477 23962
rect 10489 23910 10541 23962
rect 10553 23910 10605 23962
rect 10617 23910 10669 23962
rect 10681 23910 10733 23962
rect 19901 23910 19953 23962
rect 19965 23910 20017 23962
rect 20029 23910 20081 23962
rect 20093 23910 20145 23962
rect 20157 23910 20209 23962
rect 1400 23808 1452 23860
rect 4620 23808 4672 23860
rect 6092 23808 6144 23860
rect 7656 23851 7708 23860
rect 7656 23817 7665 23851
rect 7665 23817 7699 23851
rect 7699 23817 7708 23851
rect 7656 23808 7708 23817
rect 8484 23808 8536 23860
rect 9036 23808 9088 23860
rect 9220 23808 9272 23860
rect 11796 23808 11848 23860
rect 12164 23851 12216 23860
rect 12164 23817 12173 23851
rect 12173 23817 12207 23851
rect 12207 23817 12216 23851
rect 12164 23808 12216 23817
rect 14188 23808 14240 23860
rect 15844 23808 15896 23860
rect 2872 23740 2924 23792
rect 3424 23672 3476 23724
rect 4620 23715 4672 23724
rect 1400 23604 1452 23656
rect 4620 23681 4629 23715
rect 4629 23681 4663 23715
rect 4663 23681 4672 23715
rect 4620 23672 4672 23681
rect 4896 23715 4948 23724
rect 4896 23681 4930 23715
rect 4930 23681 4948 23715
rect 7288 23715 7340 23724
rect 4896 23672 4948 23681
rect 7288 23681 7297 23715
rect 7297 23681 7331 23715
rect 7331 23681 7340 23715
rect 7288 23672 7340 23681
rect 9404 23672 9456 23724
rect 9772 23672 9824 23724
rect 10048 23715 10100 23724
rect 10048 23681 10057 23715
rect 10057 23681 10091 23715
rect 10091 23681 10100 23715
rect 10048 23672 10100 23681
rect 3976 23604 4028 23656
rect 7472 23604 7524 23656
rect 9956 23604 10008 23656
rect 11428 23672 11480 23724
rect 11704 23715 11756 23724
rect 9588 23536 9640 23588
rect 9772 23579 9824 23588
rect 9772 23545 9781 23579
rect 9781 23545 9815 23579
rect 9815 23545 9824 23579
rect 9772 23536 9824 23545
rect 9864 23536 9916 23588
rect 10232 23536 10284 23588
rect 10692 23536 10744 23588
rect 11244 23604 11296 23656
rect 11704 23681 11712 23715
rect 11712 23681 11746 23715
rect 11746 23681 11756 23715
rect 11704 23672 11756 23681
rect 11888 23715 11940 23724
rect 11888 23681 11897 23715
rect 11897 23681 11931 23715
rect 11931 23681 11940 23715
rect 11888 23672 11940 23681
rect 12256 23672 12308 23724
rect 11796 23647 11848 23656
rect 11796 23613 11805 23647
rect 11805 23613 11839 23647
rect 11839 23613 11848 23647
rect 11796 23604 11848 23613
rect 3424 23468 3476 23520
rect 8024 23468 8076 23520
rect 10600 23468 10652 23520
rect 10968 23511 11020 23520
rect 10968 23477 10977 23511
rect 10977 23477 11011 23511
rect 11011 23477 11020 23511
rect 10968 23468 11020 23477
rect 11704 23468 11756 23520
rect 12440 23511 12492 23520
rect 12440 23477 12449 23511
rect 12449 23477 12483 23511
rect 12483 23477 12492 23511
rect 12440 23468 12492 23477
rect 13636 23672 13688 23724
rect 14004 23715 14056 23724
rect 14004 23681 14013 23715
rect 14013 23681 14047 23715
rect 14047 23681 14056 23715
rect 14004 23672 14056 23681
rect 14924 23536 14976 23588
rect 14096 23468 14148 23520
rect 16488 23715 16540 23724
rect 16488 23681 16497 23715
rect 16497 23681 16531 23715
rect 16531 23681 16540 23715
rect 16488 23672 16540 23681
rect 16672 23715 16724 23724
rect 16672 23681 16681 23715
rect 16681 23681 16715 23715
rect 16715 23681 16724 23715
rect 19432 23783 19484 23792
rect 19432 23749 19441 23783
rect 19441 23749 19475 23783
rect 19475 23749 19484 23783
rect 19432 23740 19484 23749
rect 16672 23672 16724 23681
rect 17868 23715 17920 23724
rect 17868 23681 17872 23715
rect 17872 23681 17906 23715
rect 17906 23681 17920 23715
rect 17868 23672 17920 23681
rect 16212 23647 16264 23656
rect 16212 23613 16221 23647
rect 16221 23613 16255 23647
rect 16255 23613 16264 23647
rect 16212 23604 16264 23613
rect 17500 23604 17552 23656
rect 18144 23672 18196 23724
rect 18236 23715 18288 23724
rect 18236 23681 18245 23715
rect 18245 23681 18279 23715
rect 18279 23681 18288 23715
rect 18512 23715 18564 23724
rect 18236 23672 18288 23681
rect 18512 23681 18521 23715
rect 18521 23681 18555 23715
rect 18555 23681 18564 23715
rect 18512 23672 18564 23681
rect 19340 23672 19392 23724
rect 19800 23851 19852 23860
rect 19800 23817 19817 23851
rect 19817 23817 19851 23851
rect 19851 23817 19852 23851
rect 19800 23808 19852 23817
rect 21088 23808 21140 23860
rect 22008 23808 22060 23860
rect 23664 23808 23716 23860
rect 24492 23808 24544 23860
rect 20260 23740 20312 23792
rect 24860 23740 24912 23792
rect 20168 23715 20220 23724
rect 20168 23681 20177 23715
rect 20177 23681 20211 23715
rect 20211 23681 20220 23715
rect 20168 23672 20220 23681
rect 20628 23672 20680 23724
rect 17684 23511 17736 23520
rect 17684 23477 17693 23511
rect 17693 23477 17727 23511
rect 17727 23477 17736 23511
rect 17684 23468 17736 23477
rect 19248 23468 19300 23520
rect 22836 23604 22888 23656
rect 23020 23672 23072 23724
rect 24124 23672 24176 23724
rect 23480 23604 23532 23656
rect 23664 23604 23716 23656
rect 27344 23808 27396 23860
rect 27436 23808 27488 23860
rect 28632 23808 28684 23860
rect 25228 23783 25280 23792
rect 25228 23749 25237 23783
rect 25237 23749 25271 23783
rect 25271 23749 25280 23783
rect 25228 23740 25280 23749
rect 25872 23740 25924 23792
rect 26976 23740 27028 23792
rect 26608 23672 26660 23724
rect 26700 23647 26752 23656
rect 19984 23579 20036 23588
rect 19984 23545 19993 23579
rect 19993 23545 20027 23579
rect 20027 23545 20036 23579
rect 19984 23536 20036 23545
rect 21180 23536 21232 23588
rect 22192 23579 22244 23588
rect 19432 23468 19484 23520
rect 20444 23511 20496 23520
rect 20444 23477 20453 23511
rect 20453 23477 20487 23511
rect 20487 23477 20496 23511
rect 20444 23468 20496 23477
rect 22192 23545 22201 23579
rect 22201 23545 22235 23579
rect 22235 23545 22244 23579
rect 22192 23536 22244 23545
rect 26700 23613 26709 23647
rect 26709 23613 26743 23647
rect 26743 23613 26752 23647
rect 26700 23604 26752 23613
rect 27160 23604 27212 23656
rect 28172 23672 28224 23724
rect 27620 23579 27672 23588
rect 26792 23468 26844 23520
rect 27252 23468 27304 23520
rect 27620 23545 27629 23579
rect 27629 23545 27663 23579
rect 27663 23545 27672 23579
rect 27620 23536 27672 23545
rect 28172 23468 28224 23520
rect 5688 23366 5740 23418
rect 5752 23366 5804 23418
rect 5816 23366 5868 23418
rect 5880 23366 5932 23418
rect 5944 23366 5996 23418
rect 15163 23366 15215 23418
rect 15227 23366 15279 23418
rect 15291 23366 15343 23418
rect 15355 23366 15407 23418
rect 15419 23366 15471 23418
rect 24639 23366 24691 23418
rect 24703 23366 24755 23418
rect 24767 23366 24819 23418
rect 24831 23366 24883 23418
rect 24895 23366 24947 23418
rect 2872 23264 2924 23316
rect 3976 23264 4028 23316
rect 4896 23307 4948 23316
rect 4896 23273 4905 23307
rect 4905 23273 4939 23307
rect 4939 23273 4948 23307
rect 4896 23264 4948 23273
rect 2228 23103 2280 23112
rect 2228 23069 2237 23103
rect 2237 23069 2271 23103
rect 2271 23069 2280 23103
rect 2228 23060 2280 23069
rect 2320 23060 2372 23112
rect 3608 23060 3660 23112
rect 6092 23264 6144 23316
rect 9680 23264 9732 23316
rect 10048 23264 10100 23316
rect 12716 23264 12768 23316
rect 16212 23264 16264 23316
rect 5540 23196 5592 23248
rect 5172 23171 5224 23180
rect 5172 23137 5181 23171
rect 5181 23137 5215 23171
rect 5215 23137 5224 23171
rect 5172 23128 5224 23137
rect 5632 23128 5684 23180
rect 9312 23196 9364 23248
rect 8300 23171 8352 23180
rect 8300 23137 8309 23171
rect 8309 23137 8343 23171
rect 8343 23137 8352 23171
rect 8300 23128 8352 23137
rect 5356 23103 5408 23112
rect 5356 23069 5366 23103
rect 5366 23069 5400 23103
rect 5400 23069 5408 23103
rect 5356 23060 5408 23069
rect 8024 23103 8076 23112
rect 8024 23069 8033 23103
rect 8033 23069 8067 23103
rect 8067 23069 8076 23103
rect 8024 23060 8076 23069
rect 9588 23128 9640 23180
rect 9956 23128 10008 23180
rect 10968 23196 11020 23248
rect 18512 23264 18564 23316
rect 19524 23264 19576 23316
rect 27436 23264 27488 23316
rect 22100 23196 22152 23248
rect 24308 23196 24360 23248
rect 25688 23196 25740 23248
rect 26976 23196 27028 23248
rect 11888 23128 11940 23180
rect 12072 23128 12124 23180
rect 9312 23060 9364 23112
rect 10600 23060 10652 23112
rect 11244 23103 11296 23112
rect 11244 23069 11253 23103
rect 11253 23069 11287 23103
rect 11287 23069 11296 23103
rect 11244 23060 11296 23069
rect 11428 23103 11480 23112
rect 11428 23069 11436 23103
rect 11436 23069 11470 23103
rect 11470 23069 11480 23103
rect 11428 23060 11480 23069
rect 11704 23060 11756 23112
rect 12440 23060 12492 23112
rect 14096 23103 14148 23112
rect 14096 23069 14105 23103
rect 14105 23069 14139 23103
rect 14139 23069 14148 23103
rect 14096 23060 14148 23069
rect 17316 23128 17368 23180
rect 19248 23128 19300 23180
rect 14740 23103 14792 23112
rect 5724 22992 5776 23044
rect 6460 23035 6512 23044
rect 6460 23001 6494 23035
rect 6494 23001 6512 23035
rect 6460 22992 6512 23001
rect 10048 22992 10100 23044
rect 13636 22992 13688 23044
rect 14740 23069 14749 23103
rect 14749 23069 14783 23103
rect 14783 23069 14792 23103
rect 14740 23060 14792 23069
rect 15016 23103 15068 23112
rect 15016 23069 15025 23103
rect 15025 23069 15059 23103
rect 15059 23069 15068 23103
rect 15016 23060 15068 23069
rect 15476 23103 15528 23112
rect 15476 23069 15479 23103
rect 15479 23069 15528 23103
rect 15476 23060 15528 23069
rect 15660 23060 15712 23112
rect 15844 23060 15896 23112
rect 18144 23060 18196 23112
rect 14924 22992 14976 23044
rect 17684 22992 17736 23044
rect 19708 23128 19760 23180
rect 27344 23171 27396 23180
rect 20168 23103 20220 23112
rect 20168 23069 20177 23103
rect 20177 23069 20211 23103
rect 20211 23069 20220 23103
rect 20168 23060 20220 23069
rect 2412 22967 2464 22976
rect 2412 22933 2421 22967
rect 2421 22933 2455 22967
rect 2455 22933 2464 22967
rect 2412 22924 2464 22933
rect 6644 22924 6696 22976
rect 7288 22924 7340 22976
rect 7840 22967 7892 22976
rect 7840 22933 7849 22967
rect 7849 22933 7883 22967
rect 7883 22933 7892 22967
rect 7840 22924 7892 22933
rect 8208 22924 8260 22976
rect 9588 22924 9640 22976
rect 11888 22967 11940 22976
rect 11888 22933 11897 22967
rect 11897 22933 11931 22967
rect 11931 22933 11940 22967
rect 11888 22924 11940 22933
rect 15844 22967 15896 22976
rect 15844 22933 15853 22967
rect 15853 22933 15887 22967
rect 15887 22933 15896 22967
rect 15844 22924 15896 22933
rect 17224 22924 17276 22976
rect 19340 22924 19392 22976
rect 21088 23060 21140 23112
rect 20812 22992 20864 23044
rect 20628 22924 20680 22976
rect 21640 22924 21692 22976
rect 24492 23060 24544 23112
rect 25044 22992 25096 23044
rect 25688 22992 25740 23044
rect 27344 23137 27353 23171
rect 27353 23137 27387 23171
rect 27387 23137 27396 23171
rect 27344 23128 27396 23137
rect 26608 23103 26660 23112
rect 26608 23069 26617 23103
rect 26617 23069 26651 23103
rect 26651 23069 26660 23103
rect 26608 23060 26660 23069
rect 27160 23060 27212 23112
rect 26792 23035 26844 23044
rect 26792 23001 26801 23035
rect 26801 23001 26835 23035
rect 26835 23001 26844 23035
rect 26792 22992 26844 23001
rect 22376 22967 22428 22976
rect 22376 22933 22385 22967
rect 22385 22933 22419 22967
rect 22419 22933 22428 22967
rect 22376 22924 22428 22933
rect 24676 22924 24728 22976
rect 25504 22967 25556 22976
rect 25504 22933 25513 22967
rect 25513 22933 25547 22967
rect 25547 22933 25556 22967
rect 25504 22924 25556 22933
rect 28632 22992 28684 23044
rect 10425 22822 10477 22874
rect 10489 22822 10541 22874
rect 10553 22822 10605 22874
rect 10617 22822 10669 22874
rect 10681 22822 10733 22874
rect 19901 22822 19953 22874
rect 19965 22822 20017 22874
rect 20029 22822 20081 22874
rect 20093 22822 20145 22874
rect 20157 22822 20209 22874
rect 6460 22763 6512 22772
rect 2412 22652 2464 22704
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 6460 22729 6469 22763
rect 6469 22729 6503 22763
rect 6503 22729 6512 22763
rect 6460 22720 6512 22729
rect 6828 22720 6880 22772
rect 9312 22763 9364 22772
rect 9312 22729 9321 22763
rect 9321 22729 9355 22763
rect 9355 22729 9364 22763
rect 9312 22720 9364 22729
rect 9496 22720 9548 22772
rect 9956 22720 10008 22772
rect 12164 22720 12216 22772
rect 13636 22720 13688 22772
rect 14096 22720 14148 22772
rect 1676 22559 1728 22568
rect 1676 22525 1685 22559
rect 1685 22525 1719 22559
rect 1719 22525 1728 22559
rect 1676 22516 1728 22525
rect 2320 22516 2372 22568
rect 5080 22516 5132 22568
rect 6644 22584 6696 22636
rect 6828 22627 6880 22636
rect 6828 22593 6837 22627
rect 6837 22593 6871 22627
rect 6871 22593 6880 22627
rect 6828 22584 6880 22593
rect 8208 22627 8260 22636
rect 8208 22593 8242 22627
rect 8242 22593 8260 22627
rect 6276 22448 6328 22500
rect 3056 22380 3108 22432
rect 5172 22423 5224 22432
rect 5172 22389 5181 22423
rect 5181 22389 5215 22423
rect 5215 22389 5224 22423
rect 5172 22380 5224 22389
rect 8208 22584 8260 22593
rect 9588 22584 9640 22636
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 10048 22627 10100 22636
rect 9772 22584 9824 22593
rect 10048 22593 10057 22627
rect 10057 22593 10091 22627
rect 10091 22593 10100 22627
rect 10048 22584 10100 22593
rect 11888 22652 11940 22704
rect 15844 22652 15896 22704
rect 13544 22627 13596 22636
rect 13544 22593 13553 22627
rect 13553 22593 13587 22627
rect 13587 22593 13596 22627
rect 13544 22584 13596 22593
rect 14004 22627 14056 22636
rect 14004 22593 14013 22627
rect 14013 22593 14047 22627
rect 14047 22593 14056 22627
rect 14004 22584 14056 22593
rect 15016 22627 15068 22636
rect 15016 22593 15025 22627
rect 15025 22593 15059 22627
rect 15059 22593 15068 22627
rect 15016 22584 15068 22593
rect 15476 22627 15528 22636
rect 15476 22593 15479 22627
rect 15479 22593 15528 22627
rect 10232 22516 10284 22568
rect 14832 22516 14884 22568
rect 15476 22584 15528 22593
rect 15660 22584 15712 22636
rect 16488 22652 16540 22704
rect 16120 22627 16172 22636
rect 16120 22593 16134 22627
rect 16134 22593 16168 22627
rect 16168 22593 16172 22627
rect 16672 22627 16724 22636
rect 16120 22584 16172 22593
rect 16672 22593 16681 22627
rect 16681 22593 16715 22627
rect 16715 22593 16724 22627
rect 16672 22584 16724 22593
rect 20260 22720 20312 22772
rect 17316 22652 17368 22704
rect 17408 22627 17460 22636
rect 17408 22593 17417 22627
rect 17417 22593 17451 22627
rect 17451 22593 17460 22627
rect 17408 22584 17460 22593
rect 17868 22627 17920 22636
rect 17868 22593 17871 22627
rect 17871 22593 17920 22627
rect 17500 22516 17552 22568
rect 9312 22448 9364 22500
rect 9588 22448 9640 22500
rect 9680 22448 9732 22500
rect 14924 22448 14976 22500
rect 17868 22584 17920 22593
rect 18144 22627 18196 22636
rect 18144 22593 18153 22627
rect 18153 22593 18187 22627
rect 18187 22593 18196 22627
rect 18144 22584 18196 22593
rect 19248 22652 19300 22704
rect 19708 22627 19760 22636
rect 19708 22593 19717 22627
rect 19717 22593 19751 22627
rect 19751 22593 19760 22627
rect 19708 22584 19760 22593
rect 22284 22720 22336 22772
rect 22560 22720 22612 22772
rect 22100 22627 22152 22636
rect 9036 22380 9088 22432
rect 10140 22423 10192 22432
rect 10140 22389 10149 22423
rect 10149 22389 10183 22423
rect 10183 22389 10192 22423
rect 10140 22380 10192 22389
rect 12440 22380 12492 22432
rect 16028 22380 16080 22432
rect 16304 22423 16356 22432
rect 16304 22389 16313 22423
rect 16313 22389 16347 22423
rect 16347 22389 16356 22423
rect 16304 22380 16356 22389
rect 17040 22380 17092 22432
rect 19984 22423 20036 22432
rect 19984 22389 19993 22423
rect 19993 22389 20027 22423
rect 20027 22389 20036 22423
rect 19984 22380 20036 22389
rect 20168 22448 20220 22500
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 22376 22652 22428 22704
rect 26148 22720 26200 22772
rect 28632 22763 28684 22772
rect 28632 22729 28641 22763
rect 28641 22729 28675 22763
rect 28675 22729 28684 22763
rect 28632 22720 28684 22729
rect 24676 22652 24728 22704
rect 25504 22652 25556 22704
rect 23296 22627 23348 22636
rect 23296 22593 23310 22627
rect 23310 22593 23344 22627
rect 23344 22593 23348 22627
rect 23664 22627 23716 22636
rect 23296 22584 23348 22593
rect 23664 22593 23673 22627
rect 23673 22593 23707 22627
rect 23707 22593 23716 22627
rect 23664 22584 23716 22593
rect 25596 22627 25648 22636
rect 25596 22593 25605 22627
rect 25605 22593 25639 22627
rect 25639 22593 25648 22627
rect 25596 22584 25648 22593
rect 25688 22584 25740 22636
rect 26056 22627 26108 22636
rect 26056 22593 26059 22627
rect 26059 22593 26108 22627
rect 26056 22584 26108 22593
rect 26516 22627 26568 22636
rect 26516 22593 26525 22627
rect 26525 22593 26559 22627
rect 26559 22593 26568 22627
rect 26516 22584 26568 22593
rect 28172 22584 28224 22636
rect 23204 22516 23256 22568
rect 23940 22559 23992 22568
rect 23940 22525 23949 22559
rect 23949 22525 23983 22559
rect 23983 22525 23992 22559
rect 23940 22516 23992 22525
rect 25412 22559 25464 22568
rect 25412 22525 25421 22559
rect 25421 22525 25455 22559
rect 25455 22525 25464 22559
rect 25412 22516 25464 22525
rect 20352 22423 20404 22432
rect 20352 22389 20361 22423
rect 20361 22389 20395 22423
rect 20395 22389 20404 22423
rect 20352 22380 20404 22389
rect 20536 22380 20588 22432
rect 20720 22380 20772 22432
rect 21916 22423 21968 22432
rect 21916 22389 21925 22423
rect 21925 22389 21959 22423
rect 21959 22389 21968 22423
rect 21916 22380 21968 22389
rect 24032 22380 24084 22432
rect 26148 22423 26200 22432
rect 26148 22389 26157 22423
rect 26157 22389 26191 22423
rect 26191 22389 26200 22423
rect 26148 22380 26200 22389
rect 26332 22423 26384 22432
rect 26332 22389 26341 22423
rect 26341 22389 26375 22423
rect 26375 22389 26384 22423
rect 26332 22380 26384 22389
rect 5688 22278 5740 22330
rect 5752 22278 5804 22330
rect 5816 22278 5868 22330
rect 5880 22278 5932 22330
rect 5944 22278 5996 22330
rect 15163 22278 15215 22330
rect 15227 22278 15279 22330
rect 15291 22278 15343 22330
rect 15355 22278 15407 22330
rect 15419 22278 15471 22330
rect 24639 22278 24691 22330
rect 24703 22278 24755 22330
rect 24767 22278 24819 22330
rect 24831 22278 24883 22330
rect 24895 22278 24947 22330
rect 1676 22176 1728 22228
rect 2228 22176 2280 22228
rect 3976 22176 4028 22228
rect 1400 22040 1452 22092
rect 2320 22015 2372 22024
rect 2320 21981 2329 22015
rect 2329 21981 2363 22015
rect 2363 21981 2372 22015
rect 2320 21972 2372 21981
rect 3608 21904 3660 21956
rect 3056 21836 3108 21888
rect 4160 21947 4212 21956
rect 4160 21913 4169 21947
rect 4169 21913 4203 21947
rect 4203 21913 4212 21947
rect 4160 21904 4212 21913
rect 5172 21904 5224 21956
rect 8208 22108 8260 22160
rect 12164 22108 12216 22160
rect 6552 22083 6604 22092
rect 6552 22049 6561 22083
rect 6561 22049 6595 22083
rect 6595 22049 6604 22083
rect 6552 22040 6604 22049
rect 14832 22108 14884 22160
rect 17224 22151 17276 22160
rect 17224 22117 17233 22151
rect 17233 22117 17267 22151
rect 17267 22117 17276 22151
rect 17224 22108 17276 22117
rect 17684 22108 17736 22160
rect 20076 22176 20128 22228
rect 20536 22176 20588 22228
rect 20812 22176 20864 22228
rect 22100 22176 22152 22228
rect 23940 22219 23992 22228
rect 23940 22185 23949 22219
rect 23949 22185 23983 22219
rect 23983 22185 23992 22219
rect 23940 22176 23992 22185
rect 24492 22176 24544 22228
rect 26148 22176 26200 22228
rect 6644 22015 6696 22024
rect 6644 21981 6653 22015
rect 6653 21981 6687 22015
rect 6687 21981 6696 22015
rect 6644 21972 6696 21981
rect 9220 21904 9272 21956
rect 9588 21972 9640 22024
rect 10140 21947 10192 21956
rect 5632 21879 5684 21888
rect 5632 21845 5641 21879
rect 5641 21845 5675 21879
rect 5675 21845 5684 21879
rect 5632 21836 5684 21845
rect 6184 21836 6236 21888
rect 8668 21836 8720 21888
rect 9772 21836 9824 21888
rect 10140 21913 10158 21947
rect 10158 21913 10192 21947
rect 10140 21904 10192 21913
rect 14004 22040 14056 22092
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 13544 22015 13596 22024
rect 10784 21947 10836 21956
rect 10784 21913 10818 21947
rect 10818 21913 10836 21947
rect 10784 21904 10836 21913
rect 13544 21981 13553 22015
rect 13553 21981 13587 22015
rect 13587 21981 13596 22015
rect 13544 21972 13596 21981
rect 13820 22015 13872 22024
rect 13820 21981 13829 22015
rect 13829 21981 13863 22015
rect 13863 21981 13872 22015
rect 13820 21972 13872 21981
rect 14464 22015 14516 22024
rect 14464 21981 14473 22015
rect 14473 21981 14507 22015
rect 14507 21981 14516 22015
rect 14464 21972 14516 21981
rect 15292 22015 15344 22024
rect 15292 21981 15301 22015
rect 15301 21981 15335 22015
rect 15335 21981 15344 22015
rect 15292 21972 15344 21981
rect 17408 22040 17460 22092
rect 18236 22040 18288 22092
rect 18880 22040 18932 22092
rect 19800 22040 19852 22092
rect 20076 22040 20128 22092
rect 11888 21879 11940 21888
rect 11888 21845 11897 21879
rect 11897 21845 11931 21879
rect 11931 21845 11940 21879
rect 11888 21836 11940 21845
rect 12348 21836 12400 21888
rect 12440 21879 12492 21888
rect 12440 21845 12449 21879
rect 12449 21845 12483 21879
rect 12483 21845 12492 21879
rect 12440 21836 12492 21845
rect 14004 21836 14056 21888
rect 14648 21836 14700 21888
rect 19708 21972 19760 22024
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 20352 22015 20404 22024
rect 16028 21904 16080 21956
rect 17040 21904 17092 21956
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 20536 22015 20588 22024
rect 20536 21981 20550 22015
rect 20550 21981 20584 22015
rect 20584 21981 20588 22015
rect 21088 22040 21140 22092
rect 25504 22108 25556 22160
rect 23296 22040 23348 22092
rect 22836 22015 22888 22024
rect 20536 21972 20588 21981
rect 22836 21981 22845 22015
rect 22845 21981 22879 22015
rect 22879 21981 22888 22015
rect 22836 21972 22888 21981
rect 23204 21972 23256 22024
rect 24492 21972 24544 22024
rect 27160 22015 27212 22024
rect 27160 21981 27169 22015
rect 27169 21981 27203 22015
rect 27203 21981 27212 22015
rect 27160 21972 27212 21981
rect 20260 21904 20312 21956
rect 20996 21904 21048 21956
rect 21916 21904 21968 21956
rect 23020 21947 23072 21956
rect 15844 21836 15896 21888
rect 17960 21836 18012 21888
rect 19616 21836 19668 21888
rect 22652 21836 22704 21888
rect 23020 21913 23029 21947
rect 23029 21913 23063 21947
rect 23063 21913 23072 21947
rect 23020 21904 23072 21913
rect 25412 21904 25464 21956
rect 26332 21904 26384 21956
rect 24032 21836 24084 21888
rect 24308 21836 24360 21888
rect 25964 21836 26016 21888
rect 26516 21836 26568 21888
rect 10425 21734 10477 21786
rect 10489 21734 10541 21786
rect 10553 21734 10605 21786
rect 10617 21734 10669 21786
rect 10681 21734 10733 21786
rect 19901 21734 19953 21786
rect 19965 21734 20017 21786
rect 20029 21734 20081 21786
rect 20093 21734 20145 21786
rect 20157 21734 20209 21786
rect 3424 21675 3476 21684
rect 3424 21641 3433 21675
rect 3433 21641 3467 21675
rect 3467 21641 3476 21675
rect 3424 21632 3476 21641
rect 4160 21632 4212 21684
rect 5080 21632 5132 21684
rect 4528 21564 4580 21616
rect 5632 21564 5684 21616
rect 7564 21564 7616 21616
rect 8392 21564 8444 21616
rect 7012 21496 7064 21548
rect 10324 21564 10376 21616
rect 10784 21632 10836 21684
rect 15292 21632 15344 21684
rect 16212 21632 16264 21684
rect 16672 21632 16724 21684
rect 14004 21564 14056 21616
rect 15384 21607 15436 21616
rect 15384 21573 15393 21607
rect 15393 21573 15427 21607
rect 15427 21573 15436 21607
rect 15384 21564 15436 21573
rect 17868 21632 17920 21684
rect 19708 21632 19760 21684
rect 22100 21632 22152 21684
rect 22652 21632 22704 21684
rect 9128 21496 9180 21548
rect 9404 21539 9456 21548
rect 9404 21505 9413 21539
rect 9413 21505 9447 21539
rect 9447 21505 9456 21539
rect 9404 21496 9456 21505
rect 9864 21539 9916 21548
rect 9864 21505 9873 21539
rect 9873 21505 9907 21539
rect 9907 21505 9916 21539
rect 9864 21496 9916 21505
rect 3148 21471 3200 21480
rect 3148 21437 3157 21471
rect 3157 21437 3191 21471
rect 3191 21437 3200 21471
rect 3148 21428 3200 21437
rect 3240 21428 3292 21480
rect 3608 21428 3660 21480
rect 6184 21428 6236 21480
rect 8300 21471 8352 21480
rect 8300 21437 8309 21471
rect 8309 21437 8343 21471
rect 8343 21437 8352 21471
rect 8300 21428 8352 21437
rect 8576 21471 8628 21480
rect 8576 21437 8585 21471
rect 8585 21437 8619 21471
rect 8619 21437 8628 21471
rect 8576 21428 8628 21437
rect 8944 21428 8996 21480
rect 10232 21539 10284 21548
rect 10232 21505 10241 21539
rect 10241 21505 10275 21539
rect 10275 21505 10284 21539
rect 10232 21496 10284 21505
rect 11888 21496 11940 21548
rect 12532 21496 12584 21548
rect 12624 21496 12676 21548
rect 13084 21496 13136 21548
rect 13544 21496 13596 21548
rect 14096 21539 14148 21548
rect 14096 21505 14105 21539
rect 14105 21505 14139 21539
rect 14139 21505 14148 21539
rect 14096 21496 14148 21505
rect 14464 21496 14516 21548
rect 14740 21496 14792 21548
rect 10140 21471 10192 21480
rect 10140 21437 10149 21471
rect 10149 21437 10183 21471
rect 10183 21437 10192 21471
rect 10140 21428 10192 21437
rect 10508 21428 10560 21480
rect 15936 21496 15988 21548
rect 17132 21539 17184 21548
rect 17132 21505 17141 21539
rect 17141 21505 17175 21539
rect 17175 21505 17184 21539
rect 17132 21496 17184 21505
rect 18144 21564 18196 21616
rect 19800 21564 19852 21616
rect 23020 21564 23072 21616
rect 25596 21564 25648 21616
rect 1492 21360 1544 21412
rect 3516 21292 3568 21344
rect 6736 21292 6788 21344
rect 12348 21360 12400 21412
rect 12624 21403 12676 21412
rect 12624 21369 12633 21403
rect 12633 21369 12667 21403
rect 12667 21369 12676 21403
rect 12624 21360 12676 21369
rect 8668 21335 8720 21344
rect 8668 21301 8677 21335
rect 8677 21301 8711 21335
rect 8711 21301 8720 21335
rect 8668 21292 8720 21301
rect 9036 21335 9088 21344
rect 9036 21301 9045 21335
rect 9045 21301 9079 21335
rect 9079 21301 9088 21335
rect 9036 21292 9088 21301
rect 9220 21292 9272 21344
rect 16120 21428 16172 21480
rect 18144 21428 18196 21480
rect 19800 21360 19852 21412
rect 12900 21335 12952 21344
rect 12900 21301 12909 21335
rect 12909 21301 12943 21335
rect 12943 21301 12952 21335
rect 12900 21292 12952 21301
rect 13268 21292 13320 21344
rect 14924 21292 14976 21344
rect 15660 21292 15712 21344
rect 16856 21292 16908 21344
rect 18972 21292 19024 21344
rect 20260 21496 20312 21548
rect 20720 21539 20772 21548
rect 20720 21505 20729 21539
rect 20729 21505 20763 21539
rect 20763 21505 20772 21539
rect 20720 21496 20772 21505
rect 22836 21539 22888 21548
rect 20352 21428 20404 21480
rect 20536 21428 20588 21480
rect 22836 21505 22845 21539
rect 22845 21505 22879 21539
rect 22879 21505 22888 21539
rect 22836 21496 22888 21505
rect 24216 21496 24268 21548
rect 24492 21496 24544 21548
rect 26240 21564 26292 21616
rect 27344 21632 27396 21684
rect 28816 21675 28868 21684
rect 28816 21641 28825 21675
rect 28825 21641 28859 21675
rect 28859 21641 28868 21675
rect 28816 21632 28868 21641
rect 27988 21564 28040 21616
rect 20996 21403 21048 21412
rect 20996 21369 21005 21403
rect 21005 21369 21039 21403
rect 21039 21369 21048 21403
rect 20996 21360 21048 21369
rect 24308 21360 24360 21412
rect 21088 21292 21140 21344
rect 22652 21335 22704 21344
rect 22652 21301 22661 21335
rect 22661 21301 22695 21335
rect 22695 21301 22704 21335
rect 22652 21292 22704 21301
rect 24492 21335 24544 21344
rect 24492 21301 24501 21335
rect 24501 21301 24535 21335
rect 24535 21301 24544 21335
rect 24492 21292 24544 21301
rect 25044 21292 25096 21344
rect 25964 21428 26016 21480
rect 26240 21428 26292 21480
rect 27068 21471 27120 21480
rect 27068 21437 27077 21471
rect 27077 21437 27111 21471
rect 27111 21437 27120 21471
rect 27068 21428 27120 21437
rect 26332 21292 26384 21344
rect 5688 21190 5740 21242
rect 5752 21190 5804 21242
rect 5816 21190 5868 21242
rect 5880 21190 5932 21242
rect 5944 21190 5996 21242
rect 15163 21190 15215 21242
rect 15227 21190 15279 21242
rect 15291 21190 15343 21242
rect 15355 21190 15407 21242
rect 15419 21190 15471 21242
rect 24639 21190 24691 21242
rect 24703 21190 24755 21242
rect 24767 21190 24819 21242
rect 24831 21190 24883 21242
rect 24895 21190 24947 21242
rect 4068 21088 4120 21140
rect 3240 21020 3292 21072
rect 8300 21020 8352 21072
rect 8576 21088 8628 21140
rect 9588 21088 9640 21140
rect 12440 21088 12492 21140
rect 8944 21020 8996 21072
rect 9128 21063 9180 21072
rect 9128 21029 9137 21063
rect 9137 21029 9171 21063
rect 9171 21029 9180 21063
rect 9128 21020 9180 21029
rect 10784 21020 10836 21072
rect 3424 20952 3476 21004
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 3240 20927 3292 20936
rect 3240 20893 3249 20927
rect 3249 20893 3283 20927
rect 3283 20893 3292 20927
rect 3240 20884 3292 20893
rect 3332 20927 3384 20936
rect 3332 20893 3341 20927
rect 3341 20893 3375 20927
rect 3375 20893 3384 20927
rect 3608 20927 3660 20936
rect 3332 20884 3384 20893
rect 3608 20893 3617 20927
rect 3617 20893 3651 20927
rect 3651 20893 3660 20927
rect 3608 20884 3660 20893
rect 4620 20884 4672 20936
rect 4068 20859 4120 20868
rect 4068 20825 4102 20859
rect 4102 20825 4120 20859
rect 4068 20816 4120 20825
rect 3884 20748 3936 20800
rect 6736 20995 6788 21004
rect 6736 20961 6745 20995
rect 6745 20961 6779 20995
rect 6779 20961 6788 20995
rect 6736 20952 6788 20961
rect 6644 20927 6696 20936
rect 6644 20893 6653 20927
rect 6653 20893 6687 20927
rect 6687 20893 6696 20927
rect 6644 20884 6696 20893
rect 9128 20884 9180 20936
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 9404 20816 9456 20868
rect 10324 20884 10376 20936
rect 10508 20884 10560 20936
rect 11336 20952 11388 21004
rect 13268 20952 13320 21004
rect 14832 20952 14884 21004
rect 16488 21088 16540 21140
rect 19800 21088 19852 21140
rect 22192 21088 22244 21140
rect 23296 21088 23348 21140
rect 24124 21131 24176 21140
rect 24124 21097 24133 21131
rect 24133 21097 24167 21131
rect 24167 21097 24176 21131
rect 24124 21088 24176 21097
rect 24400 21088 24452 21140
rect 15660 21063 15712 21072
rect 15660 21029 15669 21063
rect 15669 21029 15703 21063
rect 15703 21029 15712 21063
rect 15660 21020 15712 21029
rect 17960 21020 18012 21072
rect 18328 21020 18380 21072
rect 19248 21020 19300 21072
rect 20536 21063 20588 21072
rect 15844 20995 15896 21004
rect 10968 20927 11020 20936
rect 10968 20893 10977 20927
rect 10977 20893 11011 20927
rect 11011 20893 11020 20927
rect 10968 20884 11020 20893
rect 11060 20884 11112 20936
rect 12440 20927 12492 20936
rect 12440 20893 12449 20927
rect 12449 20893 12483 20927
rect 12483 20893 12492 20927
rect 12440 20884 12492 20893
rect 14924 20884 14976 20936
rect 15108 20927 15160 20936
rect 15108 20893 15117 20927
rect 15117 20893 15151 20927
rect 15151 20893 15160 20927
rect 15108 20884 15160 20893
rect 15844 20961 15853 20995
rect 15853 20961 15887 20995
rect 15887 20961 15896 20995
rect 15844 20952 15896 20961
rect 16488 20952 16540 21004
rect 17316 20952 17368 21004
rect 17684 20952 17736 21004
rect 20536 21029 20545 21063
rect 20545 21029 20579 21063
rect 20579 21029 20588 21063
rect 20536 21020 20588 21029
rect 24216 21063 24268 21072
rect 22008 20952 22060 21004
rect 24216 21029 24225 21063
rect 24225 21029 24259 21063
rect 24259 21029 24268 21063
rect 24216 21020 24268 21029
rect 24308 20952 24360 21004
rect 26240 20995 26292 21004
rect 26240 20961 26249 20995
rect 26249 20961 26283 20995
rect 26283 20961 26292 20995
rect 26240 20952 26292 20961
rect 15752 20884 15804 20936
rect 18144 20884 18196 20936
rect 18696 20884 18748 20936
rect 18972 20927 19024 20936
rect 18972 20893 18981 20927
rect 18981 20893 19015 20927
rect 19015 20893 19024 20927
rect 18972 20884 19024 20893
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 19800 20927 19852 20936
rect 19800 20893 19809 20927
rect 19809 20893 19843 20927
rect 19843 20893 19852 20927
rect 19800 20884 19852 20893
rect 20076 20884 20128 20936
rect 20168 20927 20220 20936
rect 20168 20893 20177 20927
rect 20177 20893 20211 20927
rect 20211 20893 20220 20927
rect 20168 20884 20220 20893
rect 20352 20927 20404 20936
rect 20352 20893 20366 20927
rect 20366 20893 20400 20927
rect 20400 20893 20404 20927
rect 20352 20884 20404 20893
rect 21088 20884 21140 20936
rect 23664 20927 23716 20936
rect 23664 20893 23673 20927
rect 23673 20893 23707 20927
rect 23707 20893 23716 20927
rect 23664 20884 23716 20893
rect 26608 21088 26660 21140
rect 27988 21131 28040 21140
rect 27988 21097 27997 21131
rect 27997 21097 28031 21131
rect 28031 21097 28040 21131
rect 27988 21088 28040 21097
rect 26424 20952 26476 21004
rect 26516 20927 26568 20936
rect 26516 20893 26525 20927
rect 26525 20893 26559 20927
rect 26559 20893 26568 20927
rect 26516 20884 26568 20893
rect 12072 20816 12124 20868
rect 12900 20816 12952 20868
rect 13820 20816 13872 20868
rect 14372 20816 14424 20868
rect 15844 20816 15896 20868
rect 5172 20791 5224 20800
rect 5172 20757 5181 20791
rect 5181 20757 5215 20791
rect 5215 20757 5224 20791
rect 5172 20748 5224 20757
rect 5632 20748 5684 20800
rect 9496 20748 9548 20800
rect 9864 20791 9916 20800
rect 9864 20757 9873 20791
rect 9873 20757 9907 20791
rect 9907 20757 9916 20791
rect 9864 20748 9916 20757
rect 10232 20748 10284 20800
rect 12348 20748 12400 20800
rect 15752 20748 15804 20800
rect 16856 20816 16908 20868
rect 17500 20748 17552 20800
rect 17868 20791 17920 20800
rect 17868 20757 17877 20791
rect 17877 20757 17911 20791
rect 17911 20757 17920 20791
rect 17868 20748 17920 20757
rect 18696 20748 18748 20800
rect 18880 20748 18932 20800
rect 19524 20748 19576 20800
rect 21180 20816 21232 20868
rect 22652 20816 22704 20868
rect 23388 20816 23440 20868
rect 24400 20816 24452 20868
rect 24952 20816 25004 20868
rect 20352 20748 20404 20800
rect 22376 20748 22428 20800
rect 23848 20748 23900 20800
rect 24584 20748 24636 20800
rect 26424 20791 26476 20800
rect 26424 20757 26433 20791
rect 26433 20757 26467 20791
rect 26467 20757 26476 20791
rect 26424 20748 26476 20757
rect 10425 20646 10477 20698
rect 10489 20646 10541 20698
rect 10553 20646 10605 20698
rect 10617 20646 10669 20698
rect 10681 20646 10733 20698
rect 19901 20646 19953 20698
rect 19965 20646 20017 20698
rect 20029 20646 20081 20698
rect 20093 20646 20145 20698
rect 20157 20646 20209 20698
rect 3056 20587 3108 20596
rect 3056 20553 3065 20587
rect 3065 20553 3099 20587
rect 3099 20553 3108 20587
rect 3056 20544 3108 20553
rect 3608 20544 3660 20596
rect 4068 20587 4120 20596
rect 4068 20553 4077 20587
rect 4077 20553 4111 20587
rect 4111 20553 4120 20587
rect 4068 20544 4120 20553
rect 3332 20476 3384 20528
rect 3516 20451 3568 20460
rect 3516 20417 3525 20451
rect 3525 20417 3559 20451
rect 3559 20417 3568 20451
rect 3516 20408 3568 20417
rect 5264 20476 5316 20528
rect 5540 20476 5592 20528
rect 9404 20544 9456 20596
rect 10140 20544 10192 20596
rect 11060 20544 11112 20596
rect 12440 20544 12492 20596
rect 15016 20544 15068 20596
rect 17132 20544 17184 20596
rect 17776 20544 17828 20596
rect 19800 20587 19852 20596
rect 10784 20476 10836 20528
rect 13544 20476 13596 20528
rect 17500 20476 17552 20528
rect 18696 20476 18748 20528
rect 19248 20476 19300 20528
rect 19800 20553 19809 20587
rect 19809 20553 19843 20587
rect 19843 20553 19852 20587
rect 19800 20544 19852 20553
rect 20260 20544 20312 20596
rect 22008 20587 22060 20596
rect 22008 20553 22017 20587
rect 22017 20553 22051 20587
rect 22051 20553 22060 20587
rect 22008 20544 22060 20553
rect 22836 20544 22888 20596
rect 5172 20408 5224 20460
rect 7288 20451 7340 20460
rect 7288 20417 7297 20451
rect 7297 20417 7331 20451
rect 7331 20417 7340 20451
rect 7288 20408 7340 20417
rect 7748 20451 7800 20460
rect 7748 20417 7757 20451
rect 7757 20417 7791 20451
rect 7791 20417 7800 20451
rect 7748 20408 7800 20417
rect 9128 20408 9180 20460
rect 2964 20383 3016 20392
rect 2964 20349 2973 20383
rect 2973 20349 3007 20383
rect 3007 20349 3016 20383
rect 2964 20340 3016 20349
rect 3148 20272 3200 20324
rect 3884 20272 3936 20324
rect 4620 20272 4672 20324
rect 8760 20272 8812 20324
rect 9772 20340 9824 20392
rect 11060 20383 11112 20392
rect 11060 20349 11069 20383
rect 11069 20349 11103 20383
rect 11103 20349 11112 20383
rect 11060 20340 11112 20349
rect 11336 20383 11388 20392
rect 11336 20349 11345 20383
rect 11345 20349 11379 20383
rect 11379 20349 11388 20383
rect 11336 20340 11388 20349
rect 3516 20204 3568 20256
rect 7564 20247 7616 20256
rect 7564 20213 7573 20247
rect 7573 20213 7607 20247
rect 7607 20213 7616 20247
rect 7564 20204 7616 20213
rect 9496 20204 9548 20256
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 12440 20408 12492 20417
rect 12900 20408 12952 20460
rect 12256 20383 12308 20392
rect 12256 20349 12265 20383
rect 12265 20349 12299 20383
rect 12299 20349 12308 20383
rect 12256 20340 12308 20349
rect 14740 20408 14792 20460
rect 14924 20408 14976 20460
rect 13820 20340 13872 20392
rect 15016 20383 15068 20392
rect 15016 20349 15025 20383
rect 15025 20349 15059 20383
rect 15059 20349 15068 20383
rect 15016 20340 15068 20349
rect 15752 20408 15804 20460
rect 16028 20451 16080 20460
rect 15844 20417 15853 20444
rect 15853 20417 15887 20444
rect 15887 20417 15896 20444
rect 15844 20392 15896 20417
rect 16028 20417 16042 20451
rect 16042 20417 16076 20451
rect 16076 20417 16080 20451
rect 16028 20408 16080 20417
rect 17408 20408 17460 20460
rect 17868 20408 17920 20460
rect 20536 20476 20588 20528
rect 23480 20544 23532 20596
rect 24492 20544 24544 20596
rect 24952 20544 25004 20596
rect 27252 20544 27304 20596
rect 22192 20451 22244 20460
rect 19156 20383 19208 20392
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 22192 20417 22201 20451
rect 22201 20417 22235 20451
rect 22235 20417 22244 20451
rect 22192 20408 22244 20417
rect 23112 20519 23164 20528
rect 23112 20485 23121 20519
rect 23121 20485 23155 20519
rect 23155 20485 23164 20519
rect 23112 20476 23164 20485
rect 22560 20340 22612 20392
rect 12348 20272 12400 20324
rect 12532 20204 12584 20256
rect 12716 20204 12768 20256
rect 15752 20272 15804 20324
rect 16488 20272 16540 20324
rect 17684 20247 17736 20256
rect 17684 20213 17693 20247
rect 17693 20213 17727 20247
rect 17727 20213 17736 20247
rect 19432 20272 19484 20324
rect 23020 20451 23072 20460
rect 23020 20417 23029 20451
rect 23029 20417 23063 20451
rect 23063 20417 23072 20451
rect 23296 20451 23348 20460
rect 23020 20408 23072 20417
rect 23296 20417 23299 20451
rect 23299 20417 23348 20451
rect 23296 20408 23348 20417
rect 23756 20451 23808 20460
rect 23756 20417 23765 20451
rect 23765 20417 23799 20451
rect 23799 20417 23808 20451
rect 23756 20408 23808 20417
rect 23848 20451 23900 20460
rect 23848 20417 23857 20451
rect 23857 20417 23891 20451
rect 23891 20417 23900 20451
rect 26792 20476 26844 20528
rect 23848 20408 23900 20417
rect 25044 20408 25096 20460
rect 25596 20408 25648 20460
rect 26424 20408 26476 20460
rect 26516 20451 26568 20460
rect 26516 20417 26525 20451
rect 26525 20417 26559 20451
rect 26559 20417 26568 20451
rect 26516 20408 26568 20417
rect 23204 20272 23256 20324
rect 23388 20315 23440 20324
rect 23388 20281 23397 20315
rect 23397 20281 23431 20315
rect 23431 20281 23440 20315
rect 23388 20272 23440 20281
rect 24584 20272 24636 20324
rect 17684 20204 17736 20213
rect 21364 20204 21416 20256
rect 21456 20204 21508 20256
rect 22376 20247 22428 20256
rect 22376 20213 22385 20247
rect 22385 20213 22419 20247
rect 22419 20213 22428 20247
rect 22376 20204 22428 20213
rect 23112 20204 23164 20256
rect 23848 20204 23900 20256
rect 25320 20340 25372 20392
rect 27068 20408 27120 20460
rect 25596 20272 25648 20324
rect 26056 20272 26108 20324
rect 26884 20204 26936 20256
rect 5688 20102 5740 20154
rect 5752 20102 5804 20154
rect 5816 20102 5868 20154
rect 5880 20102 5932 20154
rect 5944 20102 5996 20154
rect 15163 20102 15215 20154
rect 15227 20102 15279 20154
rect 15291 20102 15343 20154
rect 15355 20102 15407 20154
rect 15419 20102 15471 20154
rect 24639 20102 24691 20154
rect 24703 20102 24755 20154
rect 24767 20102 24819 20154
rect 24831 20102 24883 20154
rect 24895 20102 24947 20154
rect 6552 20000 6604 20052
rect 9772 20000 9824 20052
rect 10968 20000 11020 20052
rect 13728 20043 13780 20052
rect 13728 20009 13737 20043
rect 13737 20009 13771 20043
rect 13771 20009 13780 20043
rect 13728 20000 13780 20009
rect 16028 20000 16080 20052
rect 17684 20043 17736 20052
rect 17684 20009 17693 20043
rect 17693 20009 17727 20043
rect 17727 20009 17736 20043
rect 17684 20000 17736 20009
rect 19156 20000 19208 20052
rect 19248 20000 19300 20052
rect 11060 19932 11112 19984
rect 8208 19907 8260 19916
rect 8208 19873 8217 19907
rect 8217 19873 8251 19907
rect 8251 19873 8260 19907
rect 8208 19864 8260 19873
rect 8576 19864 8628 19916
rect 8944 19864 8996 19916
rect 11336 19864 11388 19916
rect 13544 19864 13596 19916
rect 15752 19864 15804 19916
rect 20260 19932 20312 19984
rect 17868 19864 17920 19916
rect 4620 19839 4672 19848
rect 4620 19805 4629 19839
rect 4629 19805 4663 19839
rect 4663 19805 4672 19839
rect 4620 19796 4672 19805
rect 8760 19839 8812 19848
rect 8760 19805 8769 19839
rect 8769 19805 8803 19839
rect 8803 19805 8812 19839
rect 8760 19796 8812 19805
rect 12348 19839 12400 19848
rect 12348 19805 12357 19839
rect 12357 19805 12391 19839
rect 12391 19805 12400 19839
rect 12348 19796 12400 19805
rect 4988 19728 5040 19780
rect 6000 19703 6052 19712
rect 6000 19669 6009 19703
rect 6009 19669 6043 19703
rect 6043 19669 6052 19703
rect 6000 19660 6052 19669
rect 10048 19728 10100 19780
rect 11704 19728 11756 19780
rect 12716 19796 12768 19848
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 14924 19839 14976 19848
rect 14924 19805 14933 19839
rect 14933 19805 14967 19839
rect 14967 19805 14976 19839
rect 14924 19796 14976 19805
rect 15016 19796 15068 19848
rect 15476 19839 15528 19848
rect 10784 19660 10836 19712
rect 11060 19660 11112 19712
rect 11888 19660 11940 19712
rect 12624 19728 12676 19780
rect 13820 19728 13872 19780
rect 15476 19805 15485 19839
rect 15485 19805 15519 19839
rect 15519 19805 15528 19839
rect 15476 19796 15528 19805
rect 15568 19839 15620 19848
rect 15568 19805 15582 19839
rect 15582 19805 15616 19839
rect 15616 19805 15620 19839
rect 15568 19796 15620 19805
rect 15844 19796 15896 19848
rect 16212 19796 16264 19848
rect 16672 19796 16724 19848
rect 16856 19728 16908 19780
rect 15568 19660 15620 19712
rect 15752 19703 15804 19712
rect 15752 19669 15769 19703
rect 15769 19669 15803 19703
rect 15803 19669 15804 19703
rect 15752 19660 15804 19669
rect 17132 19660 17184 19712
rect 18144 19839 18196 19848
rect 18144 19805 18158 19839
rect 18158 19805 18192 19839
rect 18192 19805 18196 19839
rect 18144 19796 18196 19805
rect 17960 19771 18012 19780
rect 17960 19737 17969 19771
rect 17969 19737 18003 19771
rect 18003 19737 18012 19771
rect 17960 19728 18012 19737
rect 18788 19796 18840 19848
rect 19800 19796 19852 19848
rect 18604 19728 18656 19780
rect 20720 19864 20772 19916
rect 21180 20000 21232 20052
rect 23020 20000 23072 20052
rect 25320 20043 25372 20052
rect 25320 20009 25329 20043
rect 25329 20009 25363 20043
rect 25363 20009 25372 20043
rect 25320 20000 25372 20009
rect 25596 20043 25648 20052
rect 25596 20009 25605 20043
rect 25605 20009 25639 20043
rect 25639 20009 25648 20043
rect 25596 20000 25648 20009
rect 26332 20043 26384 20052
rect 26332 20009 26341 20043
rect 26341 20009 26375 20043
rect 26375 20009 26384 20043
rect 26332 20000 26384 20009
rect 23388 19932 23440 19984
rect 23296 19864 23348 19916
rect 20352 19839 20404 19848
rect 20352 19805 20355 19839
rect 20355 19805 20404 19839
rect 20352 19796 20404 19805
rect 21456 19839 21508 19848
rect 21456 19805 21465 19839
rect 21465 19805 21499 19839
rect 21499 19805 21508 19839
rect 21456 19796 21508 19805
rect 22192 19796 22244 19848
rect 22744 19796 22796 19848
rect 25044 19839 25096 19848
rect 25044 19805 25053 19839
rect 25053 19805 25087 19839
rect 25087 19805 25096 19839
rect 25044 19796 25096 19805
rect 26240 19864 26292 19916
rect 26884 19907 26936 19916
rect 26884 19873 26893 19907
rect 26893 19873 26927 19907
rect 26927 19873 26936 19907
rect 26884 19864 26936 19873
rect 20720 19728 20772 19780
rect 22100 19728 22152 19780
rect 22468 19728 22520 19780
rect 28172 19796 28224 19848
rect 27620 19728 27672 19780
rect 18696 19660 18748 19712
rect 21548 19660 21600 19712
rect 21824 19660 21876 19712
rect 22008 19660 22060 19712
rect 22284 19660 22336 19712
rect 25136 19660 25188 19712
rect 26976 19660 27028 19712
rect 28540 19703 28592 19712
rect 28540 19669 28549 19703
rect 28549 19669 28583 19703
rect 28583 19669 28592 19703
rect 28540 19660 28592 19669
rect 10425 19558 10477 19610
rect 10489 19558 10541 19610
rect 10553 19558 10605 19610
rect 10617 19558 10669 19610
rect 10681 19558 10733 19610
rect 19901 19558 19953 19610
rect 19965 19558 20017 19610
rect 20029 19558 20081 19610
rect 20093 19558 20145 19610
rect 20157 19558 20209 19610
rect 2964 19456 3016 19508
rect 4528 19456 4580 19508
rect 4988 19499 5040 19508
rect 4988 19465 4997 19499
rect 4997 19465 5031 19499
rect 5031 19465 5040 19499
rect 4988 19456 5040 19465
rect 6000 19456 6052 19508
rect 7288 19456 7340 19508
rect 7748 19499 7800 19508
rect 4068 19320 4120 19372
rect 6552 19388 6604 19440
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 5264 19320 5316 19329
rect 7012 19320 7064 19372
rect 7748 19465 7757 19499
rect 7757 19465 7791 19499
rect 7791 19465 7800 19499
rect 7748 19456 7800 19465
rect 7932 19431 7984 19440
rect 7932 19397 7941 19431
rect 7941 19397 7975 19431
rect 7975 19397 7984 19431
rect 7932 19388 7984 19397
rect 9588 19456 9640 19508
rect 10048 19456 10100 19508
rect 12900 19499 12952 19508
rect 12900 19465 12909 19499
rect 12909 19465 12943 19499
rect 12943 19465 12952 19499
rect 12900 19456 12952 19465
rect 13268 19456 13320 19508
rect 14924 19456 14976 19508
rect 16028 19456 16080 19508
rect 7564 19363 7616 19372
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 4160 19295 4212 19304
rect 4160 19261 4169 19295
rect 4169 19261 4203 19295
rect 4203 19261 4212 19295
rect 4160 19252 4212 19261
rect 5540 19295 5592 19304
rect 3884 19184 3936 19236
rect 5540 19261 5549 19295
rect 5549 19261 5583 19295
rect 5583 19261 5592 19295
rect 5540 19252 5592 19261
rect 7564 19329 7573 19363
rect 7573 19329 7607 19363
rect 7607 19329 7616 19363
rect 7564 19320 7616 19329
rect 9496 19320 9548 19372
rect 9680 19320 9732 19372
rect 9956 19320 10008 19372
rect 6552 19184 6604 19236
rect 9772 19252 9824 19304
rect 10140 19320 10192 19372
rect 10784 19388 10836 19440
rect 11980 19388 12032 19440
rect 12164 19388 12216 19440
rect 16856 19431 16908 19440
rect 16856 19397 16865 19431
rect 16865 19397 16899 19431
rect 16899 19397 16908 19431
rect 16856 19388 16908 19397
rect 11520 19184 11572 19236
rect 11704 19320 11756 19372
rect 11888 19320 11940 19372
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 12348 19320 12400 19372
rect 12624 19320 12676 19372
rect 13360 19363 13412 19372
rect 13360 19329 13369 19363
rect 13369 19329 13403 19363
rect 13403 19329 13412 19363
rect 13360 19320 13412 19329
rect 14372 19320 14424 19372
rect 15936 19320 15988 19372
rect 16672 19363 16724 19372
rect 13452 19252 13504 19304
rect 14280 19295 14332 19304
rect 14280 19261 14289 19295
rect 14289 19261 14323 19295
rect 14323 19261 14332 19295
rect 14280 19252 14332 19261
rect 16028 19295 16080 19304
rect 16028 19261 16037 19295
rect 16037 19261 16071 19295
rect 16071 19261 16080 19295
rect 16028 19252 16080 19261
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 18144 19456 18196 19508
rect 18052 19388 18104 19440
rect 18512 19456 18564 19508
rect 20720 19456 20772 19508
rect 18604 19431 18656 19440
rect 17684 19363 17736 19372
rect 17684 19329 17693 19363
rect 17693 19329 17727 19363
rect 17727 19329 17736 19363
rect 17684 19320 17736 19329
rect 18604 19397 18613 19431
rect 18613 19397 18647 19431
rect 18647 19397 18656 19431
rect 18604 19388 18656 19397
rect 22100 19456 22152 19508
rect 21732 19388 21784 19440
rect 18788 19363 18840 19372
rect 14556 19227 14608 19236
rect 14556 19193 14565 19227
rect 14565 19193 14599 19227
rect 14599 19193 14608 19227
rect 14556 19184 14608 19193
rect 14740 19227 14792 19236
rect 14740 19193 14749 19227
rect 14749 19193 14783 19227
rect 14783 19193 14792 19227
rect 14740 19184 14792 19193
rect 17132 19252 17184 19304
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 18788 19320 18840 19329
rect 20720 19320 20772 19372
rect 21364 19363 21416 19372
rect 21364 19329 21373 19363
rect 21373 19329 21407 19363
rect 21407 19329 21416 19363
rect 21364 19320 21416 19329
rect 21456 19363 21508 19372
rect 21456 19329 21465 19363
rect 21465 19329 21499 19363
rect 21499 19329 21508 19363
rect 21456 19320 21508 19329
rect 22008 19320 22060 19372
rect 22100 19320 22152 19372
rect 23480 19456 23532 19508
rect 22284 19388 22336 19440
rect 26424 19456 26476 19508
rect 27620 19499 27672 19508
rect 25228 19388 25280 19440
rect 20628 19295 20680 19304
rect 17776 19184 17828 19236
rect 3516 19159 3568 19168
rect 3516 19125 3525 19159
rect 3525 19125 3559 19159
rect 3559 19125 3568 19159
rect 3516 19116 3568 19125
rect 5540 19116 5592 19168
rect 6368 19159 6420 19168
rect 6368 19125 6377 19159
rect 6377 19125 6411 19159
rect 6411 19125 6420 19159
rect 6368 19116 6420 19125
rect 13268 19159 13320 19168
rect 13268 19125 13277 19159
rect 13277 19125 13311 19159
rect 13311 19125 13320 19159
rect 13268 19116 13320 19125
rect 13728 19116 13780 19168
rect 17500 19159 17552 19168
rect 17500 19125 17509 19159
rect 17509 19125 17543 19159
rect 17543 19125 17552 19159
rect 17500 19116 17552 19125
rect 18420 19116 18472 19168
rect 20628 19261 20637 19295
rect 20637 19261 20671 19295
rect 20671 19261 20680 19295
rect 20628 19252 20680 19261
rect 22744 19320 22796 19372
rect 22928 19320 22980 19372
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 23664 19320 23716 19372
rect 24308 19363 24360 19372
rect 24308 19329 24317 19363
rect 24317 19329 24351 19363
rect 24351 19329 24360 19363
rect 24308 19320 24360 19329
rect 26332 19320 26384 19372
rect 27620 19465 27629 19499
rect 27629 19465 27663 19499
rect 27663 19465 27672 19499
rect 27620 19456 27672 19465
rect 28540 19320 28592 19372
rect 22560 19184 22612 19236
rect 19064 19116 19116 19168
rect 21088 19116 21140 19168
rect 21456 19116 21508 19168
rect 22376 19116 22428 19168
rect 23388 19116 23440 19168
rect 23480 19159 23532 19168
rect 23480 19125 23489 19159
rect 23489 19125 23523 19159
rect 23523 19125 23532 19159
rect 23480 19116 23532 19125
rect 23664 19116 23716 19168
rect 24032 19116 24084 19168
rect 25780 19116 25832 19168
rect 26424 19116 26476 19168
rect 28356 19116 28408 19168
rect 5688 19014 5740 19066
rect 5752 19014 5804 19066
rect 5816 19014 5868 19066
rect 5880 19014 5932 19066
rect 5944 19014 5996 19066
rect 15163 19014 15215 19066
rect 15227 19014 15279 19066
rect 15291 19014 15343 19066
rect 15355 19014 15407 19066
rect 15419 19014 15471 19066
rect 24639 19014 24691 19066
rect 24703 19014 24755 19066
rect 24767 19014 24819 19066
rect 24831 19014 24883 19066
rect 24895 19014 24947 19066
rect 3516 18912 3568 18964
rect 6460 18912 6512 18964
rect 25228 18955 25280 18964
rect 9220 18776 9272 18828
rect 12348 18776 12400 18828
rect 12992 18844 13044 18896
rect 13268 18887 13320 18896
rect 13268 18853 13277 18887
rect 13277 18853 13311 18887
rect 13311 18853 13320 18887
rect 13268 18844 13320 18853
rect 15844 18844 15896 18896
rect 21548 18887 21600 18896
rect 21548 18853 21557 18887
rect 21557 18853 21591 18887
rect 21591 18853 21600 18887
rect 21548 18844 21600 18853
rect 23388 18844 23440 18896
rect 25228 18921 25237 18955
rect 25237 18921 25271 18955
rect 25271 18921 25280 18955
rect 25228 18912 25280 18921
rect 26332 18844 26384 18896
rect 12624 18776 12676 18828
rect 12716 18776 12768 18828
rect 13728 18776 13780 18828
rect 14280 18776 14332 18828
rect 14832 18776 14884 18828
rect 16120 18776 16172 18828
rect 18052 18819 18104 18828
rect 18052 18785 18061 18819
rect 18061 18785 18095 18819
rect 18095 18785 18104 18819
rect 18052 18776 18104 18785
rect 18328 18819 18380 18828
rect 18328 18785 18337 18819
rect 18337 18785 18371 18819
rect 18371 18785 18380 18819
rect 18328 18776 18380 18785
rect 24308 18776 24360 18828
rect 3700 18708 3752 18760
rect 4068 18751 4120 18760
rect 4068 18717 4077 18751
rect 4077 18717 4111 18751
rect 4111 18717 4120 18751
rect 4068 18708 4120 18717
rect 4160 18751 4212 18760
rect 4160 18717 4169 18751
rect 4169 18717 4203 18751
rect 4203 18717 4212 18751
rect 4160 18708 4212 18717
rect 4620 18708 4672 18760
rect 4896 18751 4948 18760
rect 4896 18717 4905 18751
rect 4905 18717 4939 18751
rect 4939 18717 4948 18751
rect 4896 18708 4948 18717
rect 7472 18751 7524 18760
rect 7472 18717 7481 18751
rect 7481 18717 7515 18751
rect 7515 18717 7524 18751
rect 7472 18708 7524 18717
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 10784 18751 10836 18760
rect 10784 18717 10793 18751
rect 10793 18717 10827 18751
rect 10827 18717 10836 18751
rect 10784 18708 10836 18717
rect 11060 18751 11112 18760
rect 11060 18717 11069 18751
rect 11069 18717 11103 18751
rect 11103 18717 11112 18751
rect 11060 18708 11112 18717
rect 11244 18708 11296 18760
rect 11520 18751 11572 18760
rect 3976 18640 4028 18692
rect 5264 18640 5316 18692
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 11888 18708 11940 18760
rect 12256 18751 12308 18760
rect 12256 18717 12265 18751
rect 12265 18717 12299 18751
rect 12299 18717 12308 18751
rect 12808 18751 12860 18760
rect 12256 18708 12308 18717
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 12992 18751 13044 18760
rect 12992 18717 13001 18751
rect 13001 18717 13035 18751
rect 13035 18717 13044 18751
rect 12992 18708 13044 18717
rect 12072 18640 12124 18692
rect 12900 18640 12952 18692
rect 13360 18708 13412 18760
rect 15660 18751 15712 18760
rect 15660 18717 15669 18751
rect 15669 18717 15703 18751
rect 15703 18717 15712 18751
rect 15660 18708 15712 18717
rect 16028 18708 16080 18760
rect 15016 18640 15068 18692
rect 17500 18640 17552 18692
rect 4344 18615 4396 18624
rect 4344 18581 4353 18615
rect 4353 18581 4387 18615
rect 4387 18581 4396 18615
rect 4344 18572 4396 18581
rect 6460 18572 6512 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 9956 18572 10008 18624
rect 12348 18572 12400 18624
rect 13268 18572 13320 18624
rect 13544 18572 13596 18624
rect 16304 18572 16356 18624
rect 17132 18572 17184 18624
rect 17408 18572 17460 18624
rect 20260 18751 20312 18760
rect 20260 18717 20294 18751
rect 20294 18717 20312 18751
rect 20260 18708 20312 18717
rect 21732 18751 21784 18760
rect 21732 18717 21741 18751
rect 21741 18717 21775 18751
rect 21775 18717 21784 18751
rect 21732 18708 21784 18717
rect 23664 18708 23716 18760
rect 24492 18708 24544 18760
rect 25136 18776 25188 18828
rect 26240 18776 26292 18828
rect 22376 18683 22428 18692
rect 22376 18649 22385 18683
rect 22385 18649 22419 18683
rect 22419 18649 22428 18683
rect 22376 18640 22428 18649
rect 23388 18640 23440 18692
rect 24400 18640 24452 18692
rect 18972 18615 19024 18624
rect 18972 18581 18981 18615
rect 18981 18581 19015 18615
rect 19015 18581 19024 18615
rect 18972 18572 19024 18581
rect 20720 18572 20772 18624
rect 21364 18615 21416 18624
rect 21364 18581 21373 18615
rect 21373 18581 21407 18615
rect 21407 18581 21416 18615
rect 21364 18572 21416 18581
rect 23756 18572 23808 18624
rect 26424 18751 26476 18760
rect 26424 18717 26433 18751
rect 26433 18717 26467 18751
rect 26467 18717 26476 18751
rect 26424 18708 26476 18717
rect 27712 18640 27764 18692
rect 28356 18640 28408 18692
rect 26240 18615 26292 18624
rect 26240 18581 26249 18615
rect 26249 18581 26283 18615
rect 26283 18581 26292 18615
rect 26240 18572 26292 18581
rect 27804 18572 27856 18624
rect 10425 18470 10477 18522
rect 10489 18470 10541 18522
rect 10553 18470 10605 18522
rect 10617 18470 10669 18522
rect 10681 18470 10733 18522
rect 19901 18470 19953 18522
rect 19965 18470 20017 18522
rect 20029 18470 20081 18522
rect 20093 18470 20145 18522
rect 20157 18470 20209 18522
rect 3516 18368 3568 18420
rect 4160 18368 4212 18420
rect 5080 18368 5132 18420
rect 5264 18411 5316 18420
rect 5264 18377 5273 18411
rect 5273 18377 5307 18411
rect 5307 18377 5316 18411
rect 5264 18368 5316 18377
rect 11152 18368 11204 18420
rect 12440 18368 12492 18420
rect 12532 18368 12584 18420
rect 15752 18411 15804 18420
rect 15752 18377 15761 18411
rect 15761 18377 15795 18411
rect 15795 18377 15804 18411
rect 15752 18368 15804 18377
rect 17684 18368 17736 18420
rect 17776 18368 17828 18420
rect 1400 18300 1452 18352
rect 4896 18300 4948 18352
rect 4344 18232 4396 18284
rect 4712 18275 4764 18284
rect 4712 18241 4721 18275
rect 4721 18241 4755 18275
rect 4755 18241 4764 18275
rect 4712 18232 4764 18241
rect 6460 18300 6512 18352
rect 7656 18300 7708 18352
rect 9220 18343 9272 18352
rect 9220 18309 9229 18343
rect 9229 18309 9263 18343
rect 9263 18309 9272 18343
rect 9220 18300 9272 18309
rect 9956 18300 10008 18352
rect 12808 18300 12860 18352
rect 13176 18300 13228 18352
rect 14372 18343 14424 18352
rect 14372 18309 14381 18343
rect 14381 18309 14415 18343
rect 14415 18309 14424 18343
rect 14372 18300 14424 18309
rect 18328 18300 18380 18352
rect 18420 18343 18472 18352
rect 18420 18309 18429 18343
rect 18429 18309 18463 18343
rect 18463 18309 18472 18343
rect 18420 18300 18472 18309
rect 18972 18300 19024 18352
rect 5080 18164 5132 18216
rect 6368 18232 6420 18284
rect 6644 18207 6696 18216
rect 6644 18173 6653 18207
rect 6653 18173 6687 18207
rect 6687 18173 6696 18207
rect 6644 18164 6696 18173
rect 6920 18207 6972 18216
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 8944 18207 8996 18216
rect 8944 18173 8953 18207
rect 8953 18173 8987 18207
rect 8987 18173 8996 18207
rect 8944 18164 8996 18173
rect 11980 18232 12032 18284
rect 12716 18232 12768 18284
rect 14280 18232 14332 18284
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 17408 18275 17460 18284
rect 17408 18241 17417 18275
rect 17417 18241 17451 18275
rect 17451 18241 17460 18275
rect 17408 18232 17460 18241
rect 18144 18275 18196 18284
rect 18144 18241 18153 18275
rect 18153 18241 18187 18275
rect 18187 18241 18196 18275
rect 18144 18232 18196 18241
rect 20720 18275 20772 18284
rect 20720 18241 20729 18275
rect 20729 18241 20763 18275
rect 20763 18241 20772 18275
rect 20720 18232 20772 18241
rect 21088 18275 21140 18284
rect 21088 18241 21097 18275
rect 21097 18241 21131 18275
rect 21131 18241 21140 18275
rect 21088 18232 21140 18241
rect 23388 18411 23440 18420
rect 23388 18377 23397 18411
rect 23397 18377 23431 18411
rect 23431 18377 23440 18411
rect 23388 18368 23440 18377
rect 24308 18368 24360 18420
rect 24032 18300 24084 18352
rect 15844 18207 15896 18216
rect 5540 18096 5592 18148
rect 15844 18173 15853 18207
rect 15853 18173 15887 18207
rect 15887 18173 15896 18207
rect 15844 18164 15896 18173
rect 16120 18164 16172 18216
rect 23756 18232 23808 18284
rect 23480 18164 23532 18216
rect 24492 18275 24544 18284
rect 26240 18300 26292 18352
rect 27252 18300 27304 18352
rect 24492 18241 24506 18275
rect 24506 18241 24540 18275
rect 24540 18241 24544 18275
rect 24492 18232 24544 18241
rect 26608 18232 26660 18284
rect 27344 18275 27396 18284
rect 27344 18241 27353 18275
rect 27353 18241 27387 18275
rect 27387 18241 27396 18275
rect 27344 18232 27396 18241
rect 3608 18028 3660 18080
rect 8300 18028 8352 18080
rect 10784 18028 10836 18080
rect 11980 18071 12032 18080
rect 11980 18037 11989 18071
rect 11989 18037 12023 18071
rect 12023 18037 12032 18071
rect 11980 18028 12032 18037
rect 13544 18096 13596 18148
rect 12900 18028 12952 18080
rect 14832 18071 14884 18080
rect 14832 18037 14841 18071
rect 14841 18037 14875 18071
rect 14875 18037 14884 18071
rect 14832 18028 14884 18037
rect 18236 18028 18288 18080
rect 19064 18028 19116 18080
rect 20352 18028 20404 18080
rect 20628 18071 20680 18080
rect 20628 18037 20637 18071
rect 20637 18037 20671 18071
rect 20671 18037 20680 18071
rect 20628 18028 20680 18037
rect 27068 18164 27120 18216
rect 27712 18139 27764 18148
rect 27712 18105 27721 18139
rect 27721 18105 27755 18139
rect 27755 18105 27764 18139
rect 27712 18096 27764 18105
rect 25044 18028 25096 18080
rect 27804 18028 27856 18080
rect 5688 17926 5740 17978
rect 5752 17926 5804 17978
rect 5816 17926 5868 17978
rect 5880 17926 5932 17978
rect 5944 17926 5996 17978
rect 15163 17926 15215 17978
rect 15227 17926 15279 17978
rect 15291 17926 15343 17978
rect 15355 17926 15407 17978
rect 15419 17926 15471 17978
rect 24639 17926 24691 17978
rect 24703 17926 24755 17978
rect 24767 17926 24819 17978
rect 24831 17926 24883 17978
rect 24895 17926 24947 17978
rect 3424 17824 3476 17876
rect 3884 17824 3936 17876
rect 4068 17824 4120 17876
rect 4252 17867 4304 17876
rect 4252 17833 4261 17867
rect 4261 17833 4295 17867
rect 4295 17833 4304 17867
rect 4252 17824 4304 17833
rect 6920 17824 6972 17876
rect 7472 17867 7524 17876
rect 7472 17833 7481 17867
rect 7481 17833 7515 17867
rect 7515 17833 7524 17867
rect 7472 17824 7524 17833
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 11060 17824 11112 17876
rect 12440 17824 12492 17876
rect 24492 17824 24544 17876
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 3240 17663 3292 17672
rect 3240 17629 3249 17663
rect 3249 17629 3283 17663
rect 3283 17629 3292 17663
rect 3240 17620 3292 17629
rect 6460 17731 6512 17740
rect 6460 17697 6469 17731
rect 6469 17697 6503 17731
rect 6503 17697 6512 17731
rect 6460 17688 6512 17697
rect 6552 17731 6604 17740
rect 6552 17697 6561 17731
rect 6561 17697 6595 17731
rect 6595 17697 6604 17731
rect 12532 17756 12584 17808
rect 19708 17756 19760 17808
rect 6552 17688 6604 17697
rect 3608 17663 3660 17672
rect 3608 17629 3617 17663
rect 3617 17629 3651 17663
rect 3651 17629 3660 17663
rect 3608 17620 3660 17629
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 4712 17620 4764 17672
rect 11796 17688 11848 17740
rect 14556 17688 14608 17740
rect 15660 17688 15712 17740
rect 18144 17688 18196 17740
rect 19616 17688 19668 17740
rect 20168 17688 20220 17740
rect 7564 17620 7616 17672
rect 9588 17620 9640 17672
rect 8300 17595 8352 17604
rect 8300 17561 8309 17595
rect 8309 17561 8343 17595
rect 8343 17561 8352 17595
rect 8300 17552 8352 17561
rect 8392 17595 8444 17604
rect 8392 17561 8401 17595
rect 8401 17561 8435 17595
rect 8435 17561 8444 17595
rect 12440 17629 12449 17650
rect 12449 17629 12483 17650
rect 12483 17629 12492 17650
rect 12440 17598 12492 17629
rect 12532 17619 12584 17671
rect 12992 17663 13044 17672
rect 12992 17629 13001 17663
rect 13001 17629 13035 17663
rect 13035 17629 13044 17663
rect 12992 17620 13044 17629
rect 13176 17620 13228 17672
rect 13544 17620 13596 17672
rect 14004 17620 14056 17672
rect 8392 17552 8444 17561
rect 12716 17552 12768 17604
rect 13728 17552 13780 17604
rect 14924 17620 14976 17672
rect 18236 17620 18288 17672
rect 21272 17756 21324 17808
rect 23572 17756 23624 17808
rect 27344 17799 27396 17808
rect 27344 17765 27353 17799
rect 27353 17765 27387 17799
rect 27387 17765 27396 17799
rect 27344 17756 27396 17765
rect 20720 17620 20772 17672
rect 20904 17620 20956 17672
rect 22836 17688 22888 17740
rect 23664 17688 23716 17740
rect 26424 17688 26476 17740
rect 23388 17663 23440 17672
rect 14556 17552 14608 17604
rect 15292 17552 15344 17604
rect 6092 17484 6144 17536
rect 9772 17527 9824 17536
rect 9772 17493 9781 17527
rect 9781 17493 9815 17527
rect 9815 17493 9824 17527
rect 9772 17484 9824 17493
rect 12164 17484 12216 17536
rect 14004 17484 14056 17536
rect 14188 17527 14240 17536
rect 14188 17493 14197 17527
rect 14197 17493 14231 17527
rect 14231 17493 14240 17527
rect 14188 17484 14240 17493
rect 14648 17484 14700 17536
rect 16672 17484 16724 17536
rect 17960 17527 18012 17536
rect 17960 17493 17969 17527
rect 17969 17493 18003 17527
rect 18003 17493 18012 17527
rect 17960 17484 18012 17493
rect 18236 17484 18288 17536
rect 22376 17595 22428 17604
rect 20260 17484 20312 17536
rect 22376 17561 22385 17595
rect 22385 17561 22419 17595
rect 22419 17561 22428 17595
rect 22376 17552 22428 17561
rect 23388 17629 23397 17663
rect 23397 17629 23431 17663
rect 23431 17629 23440 17663
rect 23388 17620 23440 17629
rect 24400 17620 24452 17672
rect 20628 17484 20680 17536
rect 20904 17527 20956 17536
rect 20904 17493 20913 17527
rect 20913 17493 20947 17527
rect 20947 17493 20956 17527
rect 20904 17484 20956 17493
rect 22100 17527 22152 17536
rect 22100 17493 22109 17527
rect 22109 17493 22143 17527
rect 22143 17493 22152 17527
rect 23480 17552 23532 17604
rect 23296 17527 23348 17536
rect 22100 17484 22152 17493
rect 23296 17493 23305 17527
rect 23305 17493 23339 17527
rect 23339 17493 23348 17527
rect 23296 17484 23348 17493
rect 26608 17620 26660 17672
rect 27436 17688 27488 17740
rect 27252 17663 27304 17672
rect 27252 17629 27255 17663
rect 27255 17629 27304 17663
rect 27252 17620 27304 17629
rect 25044 17527 25096 17536
rect 25044 17493 25053 17527
rect 25053 17493 25087 17527
rect 25087 17493 25096 17527
rect 25044 17484 25096 17493
rect 25228 17484 25280 17536
rect 10425 17382 10477 17434
rect 10489 17382 10541 17434
rect 10553 17382 10605 17434
rect 10617 17382 10669 17434
rect 10681 17382 10733 17434
rect 19901 17382 19953 17434
rect 19965 17382 20017 17434
rect 20029 17382 20081 17434
rect 20093 17382 20145 17434
rect 20157 17382 20209 17434
rect 4528 17144 4580 17196
rect 4896 17212 4948 17264
rect 6644 17212 6696 17264
rect 5356 17144 5408 17196
rect 7564 17144 7616 17196
rect 12992 17280 13044 17332
rect 13084 17280 13136 17332
rect 9956 17212 10008 17264
rect 8944 17144 8996 17196
rect 12072 17144 12124 17196
rect 12716 17144 12768 17196
rect 10968 17076 11020 17128
rect 12164 17119 12216 17128
rect 12164 17085 12173 17119
rect 12173 17085 12207 17119
rect 12207 17085 12216 17119
rect 12164 17076 12216 17085
rect 12992 17144 13044 17196
rect 14280 17212 14332 17264
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 13084 17119 13136 17128
rect 13084 17085 13093 17119
rect 13093 17085 13127 17119
rect 13127 17085 13136 17119
rect 13084 17076 13136 17085
rect 4344 16940 4396 16992
rect 6460 16940 6512 16992
rect 8300 16940 8352 16992
rect 10324 16940 10376 16992
rect 11152 16940 11204 16992
rect 11796 16940 11848 16992
rect 13636 17008 13688 17060
rect 14648 17076 14700 17128
rect 15936 17280 15988 17332
rect 16672 17323 16724 17332
rect 16672 17289 16681 17323
rect 16681 17289 16715 17323
rect 16715 17289 16724 17323
rect 16672 17280 16724 17289
rect 18328 17280 18380 17332
rect 15016 17144 15068 17196
rect 15476 17144 15528 17196
rect 15660 17144 15712 17196
rect 17960 17212 18012 17264
rect 19248 17212 19300 17264
rect 19708 17255 19760 17264
rect 19708 17221 19717 17255
rect 19717 17221 19751 17255
rect 19751 17221 19760 17255
rect 19708 17212 19760 17221
rect 19800 17212 19852 17264
rect 16212 17187 16264 17196
rect 16212 17153 16221 17187
rect 16221 17153 16255 17187
rect 16255 17153 16264 17187
rect 20628 17280 20680 17332
rect 21916 17280 21968 17332
rect 22652 17280 22704 17332
rect 21640 17212 21692 17264
rect 24492 17323 24544 17332
rect 24492 17289 24501 17323
rect 24501 17289 24535 17323
rect 24535 17289 24544 17323
rect 24492 17280 24544 17289
rect 23296 17212 23348 17264
rect 16212 17144 16264 17153
rect 15292 17119 15344 17128
rect 15292 17085 15301 17119
rect 15301 17085 15335 17119
rect 15335 17085 15344 17119
rect 15292 17076 15344 17085
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 19340 17076 19392 17128
rect 19616 17076 19668 17128
rect 14832 17008 14884 17060
rect 15568 17008 15620 17060
rect 20720 17187 20772 17196
rect 20720 17153 20729 17187
rect 20729 17153 20763 17187
rect 20763 17153 20772 17187
rect 20720 17144 20772 17153
rect 20996 17187 21048 17196
rect 20996 17153 21005 17187
rect 21005 17153 21039 17187
rect 21039 17153 21048 17187
rect 20996 17144 21048 17153
rect 21272 17144 21324 17196
rect 25228 17212 25280 17264
rect 27344 17212 27396 17264
rect 27988 17212 28040 17264
rect 23572 17119 23624 17128
rect 23572 17085 23581 17119
rect 23581 17085 23615 17119
rect 23615 17085 23624 17119
rect 23572 17076 23624 17085
rect 25964 17119 26016 17128
rect 14648 16940 14700 16992
rect 18144 16940 18196 16992
rect 20536 16940 20588 16992
rect 21548 16940 21600 16992
rect 22100 16983 22152 16992
rect 22100 16949 22109 16983
rect 22109 16949 22143 16983
rect 22143 16949 22152 16983
rect 22100 16940 22152 16949
rect 22560 16940 22612 16992
rect 25964 17085 25973 17119
rect 25973 17085 26007 17119
rect 26007 17085 26016 17119
rect 25964 17076 26016 17085
rect 26240 17119 26292 17128
rect 26240 17085 26249 17119
rect 26249 17085 26283 17119
rect 26283 17085 26292 17119
rect 26240 17076 26292 17085
rect 24400 16940 24452 16992
rect 26332 16940 26384 16992
rect 5688 16838 5740 16890
rect 5752 16838 5804 16890
rect 5816 16838 5868 16890
rect 5880 16838 5932 16890
rect 5944 16838 5996 16890
rect 15163 16838 15215 16890
rect 15227 16838 15279 16890
rect 15291 16838 15343 16890
rect 15355 16838 15407 16890
rect 15419 16838 15471 16890
rect 24639 16838 24691 16890
rect 24703 16838 24755 16890
rect 24767 16838 24819 16890
rect 24831 16838 24883 16890
rect 24895 16838 24947 16890
rect 4528 16736 4580 16788
rect 5356 16779 5408 16788
rect 5356 16745 5365 16779
rect 5365 16745 5399 16779
rect 5399 16745 5408 16779
rect 5356 16736 5408 16745
rect 5540 16736 5592 16788
rect 6644 16736 6696 16788
rect 9956 16779 10008 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 3240 16532 3292 16584
rect 3700 16532 3752 16584
rect 4160 16532 4212 16584
rect 4344 16575 4396 16584
rect 4344 16541 4353 16575
rect 4353 16541 4387 16575
rect 4387 16541 4396 16575
rect 4344 16532 4396 16541
rect 6092 16600 6144 16652
rect 6460 16643 6512 16652
rect 6460 16609 6469 16643
rect 6469 16609 6503 16643
rect 6503 16609 6512 16643
rect 6460 16600 6512 16609
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 9956 16745 9965 16779
rect 9965 16745 9999 16779
rect 9999 16745 10008 16779
rect 9956 16736 10008 16745
rect 11980 16736 12032 16788
rect 12072 16779 12124 16788
rect 12072 16745 12081 16779
rect 12081 16745 12115 16779
rect 12115 16745 12124 16779
rect 12072 16736 12124 16745
rect 9864 16668 9916 16720
rect 19340 16736 19392 16788
rect 21732 16736 21784 16788
rect 12532 16668 12584 16720
rect 13360 16668 13412 16720
rect 18328 16668 18380 16720
rect 19248 16711 19300 16720
rect 6552 16600 6604 16609
rect 10968 16643 11020 16652
rect 10968 16609 10977 16643
rect 10977 16609 11011 16643
rect 11011 16609 11020 16643
rect 10968 16600 11020 16609
rect 12440 16600 12492 16652
rect 12716 16600 12768 16652
rect 16764 16600 16816 16652
rect 2320 16464 2372 16516
rect 2780 16439 2832 16448
rect 2780 16405 2789 16439
rect 2789 16405 2823 16439
rect 2823 16405 2832 16439
rect 3976 16464 4028 16516
rect 4252 16507 4304 16516
rect 4252 16473 4261 16507
rect 4261 16473 4295 16507
rect 4295 16473 4304 16507
rect 4252 16464 4304 16473
rect 4620 16464 4672 16516
rect 5080 16464 5132 16516
rect 8300 16532 8352 16584
rect 9772 16575 9824 16584
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 10784 16532 10836 16584
rect 11152 16575 11204 16584
rect 7196 16507 7248 16516
rect 2780 16396 2832 16405
rect 5356 16396 5408 16448
rect 7196 16473 7205 16507
rect 7205 16473 7239 16507
rect 7239 16473 7248 16507
rect 7196 16464 7248 16473
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 11336 16575 11388 16584
rect 11336 16541 11345 16575
rect 11345 16541 11379 16575
rect 11379 16541 11388 16575
rect 11336 16532 11388 16541
rect 11520 16575 11572 16584
rect 11520 16541 11529 16575
rect 11529 16541 11563 16575
rect 11563 16541 11572 16575
rect 11520 16532 11572 16541
rect 11888 16532 11940 16584
rect 11980 16532 12032 16584
rect 13820 16532 13872 16584
rect 16580 16532 16632 16584
rect 17776 16532 17828 16584
rect 19248 16677 19257 16711
rect 19257 16677 19291 16711
rect 19291 16677 19300 16711
rect 19248 16668 19300 16677
rect 24492 16668 24544 16720
rect 25964 16736 26016 16788
rect 27988 16736 28040 16788
rect 25504 16668 25556 16720
rect 21548 16643 21600 16652
rect 21548 16609 21557 16643
rect 21557 16609 21591 16643
rect 21591 16609 21600 16643
rect 21548 16600 21600 16609
rect 22652 16600 22704 16652
rect 11244 16464 11296 16516
rect 8484 16396 8536 16448
rect 12348 16464 12400 16516
rect 15292 16464 15344 16516
rect 12624 16396 12676 16448
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 12716 16396 12768 16405
rect 13176 16396 13228 16448
rect 15200 16396 15252 16448
rect 16856 16439 16908 16448
rect 16856 16405 16865 16439
rect 16865 16405 16899 16439
rect 16899 16405 16908 16439
rect 16856 16396 16908 16405
rect 17040 16396 17092 16448
rect 18512 16396 18564 16448
rect 23756 16532 23808 16584
rect 24492 16575 24544 16584
rect 24492 16541 24501 16575
rect 24501 16541 24535 16575
rect 24535 16541 24544 16575
rect 24492 16532 24544 16541
rect 25320 16532 25372 16584
rect 27160 16575 27212 16584
rect 20536 16464 20588 16516
rect 26424 16464 26476 16516
rect 20904 16396 20956 16448
rect 23940 16396 23992 16448
rect 24032 16396 24084 16448
rect 27160 16541 27169 16575
rect 27169 16541 27203 16575
rect 27203 16541 27212 16575
rect 27160 16532 27212 16541
rect 27528 16575 27580 16584
rect 27528 16541 27542 16575
rect 27542 16541 27576 16575
rect 27576 16541 27580 16575
rect 27528 16532 27580 16541
rect 27068 16464 27120 16516
rect 27436 16507 27488 16516
rect 27436 16473 27445 16507
rect 27445 16473 27479 16507
rect 27479 16473 27488 16507
rect 27436 16464 27488 16473
rect 27712 16439 27764 16448
rect 27712 16405 27729 16439
rect 27729 16405 27763 16439
rect 27763 16405 27764 16439
rect 27712 16396 27764 16405
rect 10425 16294 10477 16346
rect 10489 16294 10541 16346
rect 10553 16294 10605 16346
rect 10617 16294 10669 16346
rect 10681 16294 10733 16346
rect 19901 16294 19953 16346
rect 19965 16294 20017 16346
rect 20029 16294 20081 16346
rect 20093 16294 20145 16346
rect 20157 16294 20209 16346
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 4068 16192 4120 16244
rect 5080 16235 5132 16244
rect 2320 16167 2372 16176
rect 2320 16133 2329 16167
rect 2329 16133 2363 16167
rect 2363 16133 2372 16167
rect 2320 16124 2372 16133
rect 3700 16167 3752 16176
rect 3700 16133 3709 16167
rect 3709 16133 3743 16167
rect 3743 16133 3752 16167
rect 3700 16124 3752 16133
rect 2780 16099 2832 16108
rect 2780 16065 2803 16099
rect 2803 16065 2832 16099
rect 2780 16056 2832 16065
rect 3976 16099 4028 16108
rect 3148 15988 3200 16040
rect 3332 15988 3384 16040
rect 3976 16065 3985 16099
rect 3985 16065 4019 16099
rect 4019 16065 4028 16099
rect 3976 16056 4028 16065
rect 4712 16124 4764 16176
rect 5080 16201 5089 16235
rect 5089 16201 5123 16235
rect 5123 16201 5132 16235
rect 5080 16192 5132 16201
rect 7196 16192 7248 16244
rect 8484 16235 8536 16244
rect 8484 16201 8493 16235
rect 8493 16201 8527 16235
rect 8527 16201 8536 16235
rect 8484 16192 8536 16201
rect 10968 16192 11020 16244
rect 11336 16192 11388 16244
rect 12900 16192 12952 16244
rect 14188 16192 14240 16244
rect 4620 16099 4672 16108
rect 4620 16065 4629 16099
rect 4629 16065 4663 16099
rect 4663 16065 4672 16099
rect 4620 16056 4672 16065
rect 4896 16099 4948 16108
rect 4896 16065 4905 16099
rect 4905 16065 4939 16099
rect 4939 16065 4948 16099
rect 4896 16056 4948 16065
rect 3608 15920 3660 15972
rect 8392 16056 8444 16108
rect 9128 16056 9180 16108
rect 8484 16031 8536 16040
rect 8484 15997 8493 16031
rect 8493 15997 8527 16031
rect 8527 15997 8536 16031
rect 8484 15988 8536 15997
rect 9220 16031 9272 16040
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 3056 15852 3108 15904
rect 4620 15852 4672 15904
rect 11888 16124 11940 16176
rect 10232 16056 10284 16108
rect 10324 15988 10376 16040
rect 11060 16056 11112 16108
rect 12716 16124 12768 16176
rect 12072 16099 12124 16108
rect 12072 16065 12095 16099
rect 12095 16065 12124 16099
rect 12072 16056 12124 16065
rect 12348 16056 12400 16108
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 12532 16031 12584 16040
rect 12532 15997 12541 16031
rect 12541 15997 12575 16031
rect 12575 15997 12584 16031
rect 12532 15988 12584 15997
rect 5540 15852 5592 15904
rect 8116 15852 8168 15904
rect 10784 15852 10836 15904
rect 10968 15852 11020 15904
rect 12440 15920 12492 15972
rect 13452 16056 13504 16108
rect 14280 16056 14332 16108
rect 14372 16056 14424 16108
rect 16028 16192 16080 16244
rect 16764 16192 16816 16244
rect 16948 16235 17000 16244
rect 16948 16201 16957 16235
rect 16957 16201 16991 16235
rect 16991 16201 17000 16235
rect 16948 16192 17000 16201
rect 15292 16099 15344 16108
rect 15292 16065 15301 16099
rect 15301 16065 15335 16099
rect 15335 16065 15344 16099
rect 15292 16056 15344 16065
rect 16120 16124 16172 16176
rect 19248 16192 19300 16244
rect 19524 16192 19576 16244
rect 17684 16124 17736 16176
rect 18328 16124 18380 16176
rect 18880 16124 18932 16176
rect 15936 16056 15988 16108
rect 16396 16056 16448 16108
rect 16672 16099 16724 16108
rect 16672 16065 16681 16099
rect 16681 16065 16715 16099
rect 16715 16065 16724 16099
rect 16672 16056 16724 16065
rect 16764 16056 16816 16108
rect 17040 16099 17092 16108
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 22192 16192 22244 16244
rect 22652 16192 22704 16244
rect 23940 16124 23992 16176
rect 21180 16056 21232 16108
rect 15200 16031 15252 16040
rect 12900 15920 12952 15972
rect 14556 15920 14608 15972
rect 14832 15920 14884 15972
rect 15200 15997 15209 16031
rect 15209 15997 15243 16031
rect 15243 15997 15252 16031
rect 15200 15988 15252 15997
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 17592 16031 17644 16040
rect 15936 15963 15988 15972
rect 15936 15929 15945 15963
rect 15945 15929 15979 15963
rect 15979 15929 15988 15963
rect 15936 15920 15988 15929
rect 13544 15852 13596 15904
rect 15660 15895 15712 15904
rect 15660 15861 15669 15895
rect 15669 15861 15703 15895
rect 15703 15861 15712 15895
rect 15660 15852 15712 15861
rect 16672 15852 16724 15904
rect 17592 15997 17601 16031
rect 17601 15997 17635 16031
rect 17635 15997 17644 16031
rect 17592 15988 17644 15997
rect 17776 15852 17828 15904
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 21088 15852 21140 15904
rect 22284 16099 22336 16108
rect 22284 16065 22298 16099
rect 22298 16065 22332 16099
rect 22332 16065 22336 16099
rect 22652 16099 22704 16108
rect 22284 16056 22336 16065
rect 22652 16065 22661 16099
rect 22661 16065 22695 16099
rect 22695 16065 22704 16099
rect 22652 16056 22704 16065
rect 24308 16056 24360 16108
rect 26240 16192 26292 16244
rect 26608 16124 26660 16176
rect 24952 16099 25004 16108
rect 24952 16065 24961 16099
rect 24961 16065 24995 16099
rect 24995 16065 25004 16099
rect 24952 16056 25004 16065
rect 27712 16124 27764 16176
rect 28632 16124 28684 16176
rect 24400 16031 24452 16040
rect 24400 15997 24409 16031
rect 24409 15997 24443 16031
rect 24443 15997 24452 16031
rect 24400 15988 24452 15997
rect 25228 16031 25280 16040
rect 25228 15997 25237 16031
rect 25237 15997 25271 16031
rect 25271 15997 25280 16031
rect 25228 15988 25280 15997
rect 25320 15852 25372 15904
rect 25412 15852 25464 15904
rect 27344 15852 27396 15904
rect 5688 15750 5740 15802
rect 5752 15750 5804 15802
rect 5816 15750 5868 15802
rect 5880 15750 5932 15802
rect 5944 15750 5996 15802
rect 15163 15750 15215 15802
rect 15227 15750 15279 15802
rect 15291 15750 15343 15802
rect 15355 15750 15407 15802
rect 15419 15750 15471 15802
rect 24639 15750 24691 15802
rect 24703 15750 24755 15802
rect 24767 15750 24819 15802
rect 24831 15750 24883 15802
rect 24895 15750 24947 15802
rect 3976 15648 4028 15700
rect 3884 15580 3936 15632
rect 3056 15555 3108 15564
rect 3056 15521 3065 15555
rect 3065 15521 3099 15555
rect 3099 15521 3108 15555
rect 3056 15512 3108 15521
rect 3240 15512 3292 15564
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 3148 15487 3200 15496
rect 3148 15453 3157 15487
rect 3157 15453 3191 15487
rect 3191 15453 3200 15487
rect 4252 15512 4304 15564
rect 8484 15648 8536 15700
rect 14372 15691 14424 15700
rect 14372 15657 14381 15691
rect 14381 15657 14415 15691
rect 14415 15657 14424 15691
rect 14372 15648 14424 15657
rect 16304 15648 16356 15700
rect 17592 15648 17644 15700
rect 18328 15648 18380 15700
rect 19524 15648 19576 15700
rect 3148 15444 3200 15453
rect 4528 15487 4580 15530
rect 4528 15478 4537 15487
rect 4537 15478 4571 15487
rect 4571 15478 4580 15487
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 5080 15444 5132 15496
rect 5356 15487 5408 15496
rect 5356 15453 5365 15487
rect 5365 15453 5399 15487
rect 5399 15453 5408 15487
rect 5356 15444 5408 15453
rect 5540 15487 5592 15496
rect 5540 15453 5554 15487
rect 5554 15453 5588 15487
rect 5588 15453 5592 15487
rect 5540 15444 5592 15453
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 8116 15487 8168 15496
rect 8116 15453 8125 15487
rect 8125 15453 8159 15487
rect 8159 15453 8168 15487
rect 8116 15444 8168 15453
rect 16212 15580 16264 15632
rect 21548 15648 21600 15700
rect 22652 15648 22704 15700
rect 23756 15691 23808 15700
rect 10968 15512 11020 15564
rect 9680 15487 9732 15496
rect 2044 15308 2096 15360
rect 3884 15308 3936 15360
rect 5448 15419 5500 15428
rect 5448 15385 5462 15419
rect 5462 15385 5496 15419
rect 5496 15385 5500 15419
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 11060 15444 11112 15496
rect 12716 15512 12768 15564
rect 13820 15444 13872 15496
rect 15844 15512 15896 15564
rect 16672 15512 16724 15564
rect 5448 15376 5500 15385
rect 4896 15351 4948 15360
rect 4896 15317 4905 15351
rect 4905 15317 4939 15351
rect 4939 15317 4948 15351
rect 4896 15308 4948 15317
rect 12348 15376 12400 15428
rect 13636 15376 13688 15428
rect 14096 15419 14148 15428
rect 14096 15385 14105 15419
rect 14105 15385 14139 15419
rect 14139 15385 14148 15419
rect 14096 15376 14148 15385
rect 16396 15444 16448 15496
rect 16580 15444 16632 15496
rect 16948 15444 17000 15496
rect 17684 15512 17736 15564
rect 19064 15512 19116 15564
rect 19248 15512 19300 15564
rect 22836 15512 22888 15564
rect 23756 15657 23765 15691
rect 23765 15657 23799 15691
rect 23799 15657 23808 15691
rect 23756 15648 23808 15657
rect 25228 15648 25280 15700
rect 25688 15648 25740 15700
rect 26608 15691 26660 15700
rect 25412 15580 25464 15632
rect 26608 15657 26617 15691
rect 26617 15657 26651 15691
rect 26651 15657 26660 15691
rect 26608 15648 26660 15657
rect 28632 15691 28684 15700
rect 28632 15657 28641 15691
rect 28641 15657 28675 15691
rect 28675 15657 28684 15691
rect 28632 15648 28684 15657
rect 27620 15580 27672 15632
rect 15016 15376 15068 15428
rect 15568 15376 15620 15428
rect 18788 15444 18840 15496
rect 18972 15487 19024 15496
rect 18972 15453 18981 15487
rect 18981 15453 19015 15487
rect 19015 15453 19024 15487
rect 18972 15444 19024 15453
rect 19708 15444 19760 15496
rect 23388 15487 23440 15496
rect 20812 15419 20864 15428
rect 7748 15308 7800 15360
rect 9312 15351 9364 15360
rect 9312 15317 9321 15351
rect 9321 15317 9355 15351
rect 9355 15317 9364 15351
rect 9312 15308 9364 15317
rect 9772 15308 9824 15360
rect 10324 15308 10376 15360
rect 10968 15308 11020 15360
rect 12716 15308 12768 15360
rect 13544 15308 13596 15360
rect 16028 15308 16080 15360
rect 18512 15351 18564 15360
rect 18512 15317 18521 15351
rect 18521 15317 18555 15351
rect 18555 15317 18564 15351
rect 18512 15308 18564 15317
rect 20812 15385 20821 15419
rect 20821 15385 20855 15419
rect 20855 15385 20864 15419
rect 20812 15376 20864 15385
rect 20536 15308 20588 15360
rect 23388 15453 23397 15487
rect 23397 15453 23431 15487
rect 23431 15453 23440 15487
rect 23388 15444 23440 15453
rect 23572 15487 23624 15496
rect 23572 15453 23581 15487
rect 23581 15453 23615 15487
rect 23615 15453 23624 15487
rect 23572 15444 23624 15453
rect 24032 15444 24084 15496
rect 24400 15444 24452 15496
rect 25320 15487 25372 15496
rect 25320 15453 25324 15487
rect 25324 15453 25358 15487
rect 25358 15453 25372 15487
rect 25320 15444 25372 15453
rect 26332 15487 26384 15496
rect 22836 15419 22888 15428
rect 22836 15385 22845 15419
rect 22845 15385 22879 15419
rect 22879 15385 22888 15419
rect 22836 15376 22888 15385
rect 22928 15376 22980 15428
rect 24308 15376 24360 15428
rect 25412 15419 25464 15428
rect 25412 15385 25421 15419
rect 25421 15385 25455 15419
rect 25455 15385 25464 15419
rect 25412 15376 25464 15385
rect 25504 15419 25556 15428
rect 25504 15385 25513 15419
rect 25513 15385 25547 15419
rect 25547 15385 25556 15419
rect 26332 15453 26341 15487
rect 26341 15453 26375 15487
rect 26375 15453 26384 15487
rect 26332 15444 26384 15453
rect 26884 15444 26936 15496
rect 27160 15487 27212 15496
rect 27160 15453 27169 15487
rect 27169 15453 27203 15487
rect 27203 15453 27212 15487
rect 27160 15444 27212 15453
rect 27528 15487 27580 15496
rect 27528 15453 27542 15487
rect 27542 15453 27576 15487
rect 27576 15453 27580 15487
rect 27528 15444 27580 15453
rect 25504 15376 25556 15385
rect 24492 15308 24544 15360
rect 26700 15376 26752 15428
rect 27436 15419 27488 15428
rect 27436 15385 27445 15419
rect 27445 15385 27479 15419
rect 27479 15385 27488 15419
rect 27436 15376 27488 15385
rect 27528 15308 27580 15360
rect 10425 15206 10477 15258
rect 10489 15206 10541 15258
rect 10553 15206 10605 15258
rect 10617 15206 10669 15258
rect 10681 15206 10733 15258
rect 19901 15206 19953 15258
rect 19965 15206 20017 15258
rect 20029 15206 20081 15258
rect 20093 15206 20145 15258
rect 20157 15206 20209 15258
rect 2964 15104 3016 15156
rect 4160 15104 4212 15156
rect 2780 15036 2832 15088
rect 1952 14968 2004 15020
rect 3240 15011 3292 15020
rect 3240 14977 3249 15011
rect 3249 14977 3283 15011
rect 3283 14977 3292 15011
rect 3240 14968 3292 14977
rect 3332 15011 3384 15020
rect 3332 14977 3341 15011
rect 3341 14977 3375 15011
rect 3375 14977 3384 15011
rect 4620 15036 4672 15088
rect 3332 14968 3384 14977
rect 3884 15011 3936 15020
rect 3148 14832 3200 14884
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 3792 14900 3844 14952
rect 4436 14900 4488 14952
rect 5448 15079 5500 15088
rect 5448 15045 5457 15079
rect 5457 15045 5491 15079
rect 5491 15045 5500 15079
rect 5448 15036 5500 15045
rect 4896 15011 4948 15020
rect 4896 14977 4905 15011
rect 4905 14977 4939 15011
rect 4939 14977 4948 15011
rect 4896 14968 4948 14977
rect 10232 15104 10284 15156
rect 7748 15079 7800 15088
rect 7748 15045 7757 15079
rect 7757 15045 7791 15079
rect 7791 15045 7800 15079
rect 7748 15036 7800 15045
rect 9312 15036 9364 15088
rect 11060 15104 11112 15156
rect 11888 15104 11940 15156
rect 12532 15036 12584 15088
rect 16120 15104 16172 15156
rect 17776 15104 17828 15156
rect 19800 15104 19852 15156
rect 20536 15104 20588 15156
rect 21180 15104 21232 15156
rect 21548 15147 21600 15156
rect 21548 15113 21557 15147
rect 21557 15113 21591 15147
rect 21591 15113 21600 15147
rect 21548 15104 21600 15113
rect 4528 14832 4580 14884
rect 3976 14764 4028 14816
rect 5356 14764 5408 14816
rect 6184 14968 6236 15020
rect 9772 14968 9824 15020
rect 10048 14968 10100 15020
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 6644 14900 6696 14952
rect 7380 14900 7432 14952
rect 12716 14968 12768 15020
rect 13268 14968 13320 15020
rect 13544 15036 13596 15088
rect 18788 15079 18840 15088
rect 14280 15011 14332 15020
rect 12348 14832 12400 14884
rect 12532 14875 12584 14884
rect 12532 14841 12541 14875
rect 12541 14841 12575 14875
rect 12575 14841 12584 14875
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 18788 15045 18797 15079
rect 18797 15045 18831 15079
rect 18831 15045 18840 15079
rect 18788 15036 18840 15045
rect 19524 15036 19576 15088
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 15016 15011 15068 15020
rect 12532 14832 12584 14841
rect 14096 14832 14148 14884
rect 15016 14977 15025 15011
rect 15025 14977 15059 15011
rect 15059 14977 15068 15011
rect 15016 14968 15068 14977
rect 14924 14900 14976 14952
rect 15568 15011 15620 15020
rect 15568 14977 15577 15011
rect 15577 14977 15611 15011
rect 15611 14977 15620 15011
rect 15568 14968 15620 14977
rect 16028 15011 16080 15020
rect 16028 14977 16037 15011
rect 16037 14977 16071 15011
rect 16071 14977 16080 15011
rect 16028 14968 16080 14977
rect 15292 14900 15344 14952
rect 16764 14968 16816 15020
rect 18972 15011 19024 15020
rect 18972 14977 18981 15011
rect 18981 14977 19015 15011
rect 19015 14977 19024 15011
rect 18972 14968 19024 14977
rect 16488 14832 16540 14884
rect 17224 14900 17276 14952
rect 17592 14832 17644 14884
rect 19800 14968 19852 15020
rect 19708 14832 19760 14884
rect 9220 14807 9272 14816
rect 9220 14773 9229 14807
rect 9229 14773 9263 14807
rect 9263 14773 9272 14807
rect 9220 14764 9272 14773
rect 9956 14764 10008 14816
rect 12164 14764 12216 14816
rect 12808 14764 12860 14816
rect 13268 14764 13320 14816
rect 13360 14764 13412 14816
rect 14832 14764 14884 14816
rect 16212 14764 16264 14816
rect 16396 14764 16448 14816
rect 20720 15011 20772 15020
rect 20720 14977 20723 15011
rect 20723 14977 20772 15011
rect 21088 15011 21140 15020
rect 20720 14968 20772 14977
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 21916 14968 21968 15020
rect 23388 15104 23440 15156
rect 24400 15147 24452 15156
rect 24400 15113 24409 15147
rect 24409 15113 24443 15147
rect 24443 15113 24452 15147
rect 24400 15104 24452 15113
rect 26332 15147 26384 15156
rect 26332 15113 26341 15147
rect 26341 15113 26375 15147
rect 26375 15113 26384 15147
rect 26332 15104 26384 15113
rect 27528 15104 27580 15156
rect 22284 15011 22336 15020
rect 22284 14977 22287 15011
rect 22287 14977 22336 15011
rect 22284 14968 22336 14977
rect 22560 15011 22612 15020
rect 22560 14977 22569 15011
rect 22569 14977 22603 15011
rect 22603 14977 22612 15011
rect 22560 14968 22612 14977
rect 23572 14968 23624 15020
rect 24308 15011 24360 15020
rect 24308 14977 24317 15011
rect 24317 14977 24351 15011
rect 24351 14977 24360 15011
rect 24308 14968 24360 14977
rect 20812 14875 20864 14884
rect 20812 14841 20821 14875
rect 20821 14841 20855 14875
rect 20855 14841 20864 14875
rect 20812 14832 20864 14841
rect 23480 14900 23532 14952
rect 26608 14968 26660 15020
rect 22284 14832 22336 14884
rect 22836 14832 22888 14884
rect 24492 14832 24544 14884
rect 21180 14764 21232 14816
rect 21364 14764 21416 14816
rect 23940 14764 23992 14816
rect 25228 14764 25280 14816
rect 26792 14764 26844 14816
rect 5688 14662 5740 14714
rect 5752 14662 5804 14714
rect 5816 14662 5868 14714
rect 5880 14662 5932 14714
rect 5944 14662 5996 14714
rect 15163 14662 15215 14714
rect 15227 14662 15279 14714
rect 15291 14662 15343 14714
rect 15355 14662 15407 14714
rect 15419 14662 15471 14714
rect 24639 14662 24691 14714
rect 24703 14662 24755 14714
rect 24767 14662 24819 14714
rect 24831 14662 24883 14714
rect 24895 14662 24947 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 3240 14603 3292 14612
rect 3240 14569 3249 14603
rect 3249 14569 3283 14603
rect 3283 14569 3292 14603
rect 3240 14560 3292 14569
rect 3792 14603 3844 14612
rect 3792 14569 3801 14603
rect 3801 14569 3835 14603
rect 3835 14569 3844 14603
rect 3792 14560 3844 14569
rect 12992 14603 13044 14612
rect 12992 14569 13001 14603
rect 13001 14569 13035 14603
rect 13035 14569 13044 14603
rect 12992 14560 13044 14569
rect 13176 14560 13228 14612
rect 14096 14560 14148 14612
rect 15016 14560 15068 14612
rect 15568 14603 15620 14612
rect 15568 14569 15577 14603
rect 15577 14569 15611 14603
rect 15611 14569 15620 14603
rect 15568 14560 15620 14569
rect 16764 14603 16816 14612
rect 16764 14569 16773 14603
rect 16773 14569 16807 14603
rect 16807 14569 16816 14603
rect 16764 14560 16816 14569
rect 19616 14560 19668 14612
rect 20720 14560 20772 14612
rect 22284 14560 22336 14612
rect 25780 14560 25832 14612
rect 9772 14424 9824 14476
rect 2044 14399 2096 14408
rect 2044 14365 2053 14399
rect 2053 14365 2087 14399
rect 2087 14365 2096 14399
rect 2044 14356 2096 14365
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 4252 14356 4304 14408
rect 5080 14356 5132 14408
rect 8484 14399 8536 14408
rect 4344 14288 4396 14340
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 8484 14356 8536 14365
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 12256 14424 12308 14476
rect 13268 14492 13320 14544
rect 14464 14492 14516 14544
rect 14004 14424 14056 14476
rect 16396 14492 16448 14544
rect 12716 14399 12768 14408
rect 8852 14288 8904 14340
rect 9128 14288 9180 14340
rect 5632 14220 5684 14272
rect 10140 14263 10192 14272
rect 10140 14229 10149 14263
rect 10149 14229 10183 14263
rect 10183 14229 10192 14263
rect 10140 14220 10192 14229
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 12808 14356 12860 14365
rect 14372 14399 14424 14408
rect 14372 14365 14381 14399
rect 14381 14365 14415 14399
rect 14415 14365 14424 14399
rect 14372 14356 14424 14365
rect 14648 14356 14700 14408
rect 15568 14424 15620 14476
rect 22192 14492 22244 14544
rect 23756 14492 23808 14544
rect 23848 14492 23900 14544
rect 25044 14492 25096 14544
rect 15660 14356 15712 14408
rect 15844 14356 15896 14408
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 16488 14356 16540 14408
rect 24492 14424 24544 14476
rect 17684 14356 17736 14408
rect 17960 14356 18012 14408
rect 19524 14356 19576 14408
rect 21364 14399 21416 14408
rect 12900 14288 12952 14340
rect 13452 14288 13504 14340
rect 15568 14288 15620 14340
rect 13360 14220 13412 14272
rect 16672 14288 16724 14340
rect 17040 14288 17092 14340
rect 17592 14331 17644 14340
rect 17592 14297 17601 14331
rect 17601 14297 17635 14331
rect 17635 14297 17644 14331
rect 17592 14288 17644 14297
rect 21364 14365 21373 14399
rect 21373 14365 21407 14399
rect 21407 14365 21416 14399
rect 21364 14356 21416 14365
rect 23296 14356 23348 14408
rect 23572 14399 23624 14408
rect 23572 14365 23581 14399
rect 23581 14365 23615 14399
rect 23615 14365 23624 14399
rect 23572 14356 23624 14365
rect 16212 14263 16264 14272
rect 16212 14229 16221 14263
rect 16221 14229 16255 14263
rect 16255 14229 16264 14263
rect 16212 14220 16264 14229
rect 16396 14220 16448 14272
rect 17500 14220 17552 14272
rect 20260 14288 20312 14340
rect 23940 14399 23992 14408
rect 23940 14365 23954 14399
rect 23954 14365 23988 14399
rect 23988 14365 23992 14399
rect 23940 14356 23992 14365
rect 25228 14399 25280 14408
rect 25228 14365 25231 14399
rect 25231 14365 25280 14399
rect 25228 14356 25280 14365
rect 27528 14356 27580 14408
rect 21548 14263 21600 14272
rect 21548 14229 21557 14263
rect 21557 14229 21591 14263
rect 21591 14229 21600 14263
rect 21548 14220 21600 14229
rect 22652 14220 22704 14272
rect 23756 14331 23808 14340
rect 23756 14297 23765 14331
rect 23765 14297 23799 14331
rect 23799 14297 23808 14331
rect 24492 14331 24544 14340
rect 23756 14288 23808 14297
rect 24492 14297 24501 14331
rect 24501 14297 24535 14331
rect 24535 14297 24544 14331
rect 24492 14288 24544 14297
rect 24952 14331 25004 14340
rect 24952 14297 24961 14331
rect 24961 14297 24995 14331
rect 24995 14297 25004 14331
rect 24952 14288 25004 14297
rect 24400 14220 24452 14272
rect 26792 14288 26844 14340
rect 27528 14220 27580 14272
rect 28632 14220 28684 14272
rect 10425 14118 10477 14170
rect 10489 14118 10541 14170
rect 10553 14118 10605 14170
rect 10617 14118 10669 14170
rect 10681 14118 10733 14170
rect 19901 14118 19953 14170
rect 19965 14118 20017 14170
rect 20029 14118 20081 14170
rect 20093 14118 20145 14170
rect 20157 14118 20209 14170
rect 3424 14016 3476 14068
rect 4896 14016 4948 14068
rect 5080 14059 5132 14068
rect 5080 14025 5089 14059
rect 5089 14025 5123 14059
rect 5123 14025 5132 14059
rect 5080 14016 5132 14025
rect 4436 13948 4488 14000
rect 2872 13880 2924 13932
rect 3700 13923 3752 13932
rect 3700 13889 3709 13923
rect 3709 13889 3743 13923
rect 3743 13889 3752 13923
rect 3700 13880 3752 13889
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 4344 13923 4396 13932
rect 4344 13889 4353 13923
rect 4353 13889 4387 13923
rect 4387 13889 4396 13923
rect 4344 13880 4396 13889
rect 4712 13948 4764 14000
rect 5540 13948 5592 14000
rect 8484 14016 8536 14068
rect 9128 14016 9180 14068
rect 12716 14016 12768 14068
rect 4804 13923 4856 13932
rect 4804 13889 4813 13923
rect 4813 13889 4847 13923
rect 4847 13889 4856 13923
rect 4804 13880 4856 13889
rect 4988 13880 5040 13932
rect 5448 13880 5500 13932
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 9680 13948 9732 14000
rect 10140 13948 10192 14000
rect 4252 13812 4304 13864
rect 5632 13855 5684 13864
rect 5632 13821 5641 13855
rect 5641 13821 5675 13855
rect 5675 13821 5684 13855
rect 5632 13812 5684 13821
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 9772 13812 9824 13864
rect 11980 13880 12032 13932
rect 12348 13948 12400 14000
rect 14372 14016 14424 14068
rect 15752 14016 15804 14068
rect 15936 14016 15988 14068
rect 12440 13880 12492 13932
rect 11336 13812 11388 13864
rect 11704 13812 11756 13864
rect 15016 13991 15068 14000
rect 15016 13957 15025 13991
rect 15025 13957 15059 13991
rect 15059 13957 15068 13991
rect 15016 13948 15068 13957
rect 16304 13991 16356 14000
rect 16304 13957 16313 13991
rect 16313 13957 16347 13991
rect 16347 13957 16356 13991
rect 16304 13948 16356 13957
rect 16396 13948 16448 14000
rect 17224 14016 17276 14068
rect 19524 14059 19576 14068
rect 19524 14025 19533 14059
rect 19533 14025 19567 14059
rect 19567 14025 19576 14059
rect 19524 14016 19576 14025
rect 20720 14016 20772 14068
rect 21180 14016 21232 14068
rect 16948 13948 17000 14000
rect 18696 13948 18748 14000
rect 14004 13880 14056 13932
rect 13636 13812 13688 13864
rect 14740 13880 14792 13932
rect 15660 13880 15712 13932
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 16764 13880 16816 13932
rect 17040 13923 17092 13932
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 17224 13923 17276 13932
rect 17224 13889 17233 13923
rect 17233 13889 17267 13923
rect 17267 13889 17276 13923
rect 17224 13880 17276 13889
rect 17500 13923 17552 13932
rect 17500 13889 17503 13923
rect 17503 13889 17552 13923
rect 17500 13880 17552 13889
rect 17776 13923 17828 13932
rect 17776 13889 17785 13923
rect 17785 13889 17819 13923
rect 17819 13889 17828 13923
rect 17776 13880 17828 13889
rect 20260 13880 20312 13932
rect 22376 14016 22428 14068
rect 23756 14016 23808 14068
rect 24952 14016 25004 14068
rect 25780 14016 25832 14068
rect 26608 14059 26660 14068
rect 26608 14025 26617 14059
rect 26617 14025 26651 14059
rect 26651 14025 26660 14059
rect 26608 14016 26660 14025
rect 27436 14016 27488 14068
rect 29092 14059 29144 14068
rect 29092 14025 29101 14059
rect 29101 14025 29135 14059
rect 29135 14025 29144 14059
rect 29092 14016 29144 14025
rect 27620 13991 27672 14000
rect 27620 13957 27629 13991
rect 27629 13957 27663 13991
rect 27663 13957 27672 13991
rect 27620 13948 27672 13957
rect 28632 13948 28684 14000
rect 20720 13923 20772 13932
rect 20720 13889 20729 13923
rect 20729 13889 20763 13923
rect 20763 13889 20772 13923
rect 20720 13880 20772 13889
rect 24400 13923 24452 13932
rect 4896 13744 4948 13796
rect 6092 13744 6144 13796
rect 12808 13787 12860 13796
rect 12808 13753 12817 13787
rect 12817 13753 12851 13787
rect 12851 13753 12860 13787
rect 12808 13744 12860 13753
rect 3884 13676 3936 13728
rect 5264 13676 5316 13728
rect 9036 13719 9088 13728
rect 9036 13685 9045 13719
rect 9045 13685 9079 13719
rect 9079 13685 9088 13719
rect 9036 13676 9088 13685
rect 16396 13812 16448 13864
rect 15016 13744 15068 13796
rect 16488 13744 16540 13796
rect 24400 13889 24409 13923
rect 24409 13889 24443 13923
rect 24443 13889 24452 13923
rect 24400 13880 24452 13889
rect 26332 13880 26384 13932
rect 20720 13744 20772 13796
rect 22284 13812 22336 13864
rect 22652 13812 22704 13864
rect 23848 13855 23900 13864
rect 23848 13821 23857 13855
rect 23857 13821 23891 13855
rect 23891 13821 23900 13855
rect 23848 13812 23900 13821
rect 25044 13812 25096 13864
rect 14464 13676 14516 13728
rect 20812 13676 20864 13728
rect 5688 13574 5740 13626
rect 5752 13574 5804 13626
rect 5816 13574 5868 13626
rect 5880 13574 5932 13626
rect 5944 13574 5996 13626
rect 15163 13574 15215 13626
rect 15227 13574 15279 13626
rect 15291 13574 15343 13626
rect 15355 13574 15407 13626
rect 15419 13574 15471 13626
rect 24639 13574 24691 13626
rect 24703 13574 24755 13626
rect 24767 13574 24819 13626
rect 24831 13574 24883 13626
rect 24895 13574 24947 13626
rect 4988 13472 5040 13524
rect 3424 13404 3476 13456
rect 5264 13404 5316 13456
rect 5540 13404 5592 13456
rect 8392 13404 8444 13456
rect 2780 13268 2832 13320
rect 4160 13336 4212 13388
rect 2412 13200 2464 13252
rect 4344 13268 4396 13320
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 6092 13336 6144 13388
rect 8852 13472 8904 13524
rect 11796 13472 11848 13524
rect 12440 13472 12492 13524
rect 16396 13472 16448 13524
rect 18696 13515 18748 13524
rect 14464 13404 14516 13456
rect 17132 13404 17184 13456
rect 15660 13336 15712 13388
rect 16580 13336 16632 13388
rect 17500 13336 17552 13388
rect 5540 13268 5592 13320
rect 6644 13311 6696 13320
rect 5264 13200 5316 13252
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 9036 13268 9088 13320
rect 11888 13311 11940 13320
rect 1768 13132 1820 13184
rect 2688 13132 2740 13184
rect 3700 13132 3752 13184
rect 4712 13132 4764 13184
rect 5100 13132 5152 13184
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 11888 13277 11897 13311
rect 11897 13277 11931 13311
rect 11931 13277 11940 13311
rect 11888 13268 11940 13277
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 13452 13268 13504 13320
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15568 13268 15620 13277
rect 18696 13481 18705 13515
rect 18705 13481 18739 13515
rect 18739 13481 18748 13515
rect 18696 13472 18748 13481
rect 22284 13515 22336 13524
rect 22284 13481 22293 13515
rect 22293 13481 22327 13515
rect 22327 13481 22336 13515
rect 22284 13472 22336 13481
rect 23848 13472 23900 13524
rect 24492 13472 24544 13524
rect 20536 13379 20588 13388
rect 20536 13345 20545 13379
rect 20545 13345 20579 13379
rect 20579 13345 20588 13379
rect 20536 13336 20588 13345
rect 20812 13379 20864 13388
rect 20812 13345 20821 13379
rect 20821 13345 20855 13379
rect 20855 13345 20864 13379
rect 20812 13336 20864 13345
rect 17960 13311 18012 13320
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 15660 13200 15712 13252
rect 6184 13132 6236 13141
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 13820 13175 13872 13184
rect 13820 13141 13829 13175
rect 13829 13141 13863 13175
rect 13863 13141 13872 13175
rect 13820 13132 13872 13141
rect 15016 13132 15068 13184
rect 16948 13175 17000 13184
rect 16948 13141 16957 13175
rect 16957 13141 16991 13175
rect 16991 13141 17000 13175
rect 16948 13132 17000 13141
rect 23480 13311 23532 13320
rect 23480 13277 23489 13311
rect 23489 13277 23523 13311
rect 23523 13277 23532 13311
rect 23480 13268 23532 13277
rect 23572 13311 23624 13320
rect 23572 13277 23581 13311
rect 23581 13277 23615 13311
rect 23615 13277 23624 13311
rect 23756 13311 23808 13320
rect 23572 13268 23624 13277
rect 23756 13277 23765 13311
rect 23765 13277 23799 13311
rect 23799 13277 23808 13311
rect 23756 13268 23808 13277
rect 21548 13200 21600 13252
rect 22744 13175 22796 13184
rect 22744 13141 22753 13175
rect 22753 13141 22787 13175
rect 22787 13141 22796 13175
rect 22744 13132 22796 13141
rect 23296 13175 23348 13184
rect 23296 13141 23305 13175
rect 23305 13141 23339 13175
rect 23339 13141 23348 13175
rect 23296 13132 23348 13141
rect 25228 13404 25280 13456
rect 23940 13311 23992 13320
rect 23940 13277 23954 13311
rect 23954 13277 23988 13311
rect 23988 13277 23992 13311
rect 23940 13268 23992 13277
rect 25044 13336 25096 13388
rect 24952 13243 25004 13252
rect 24952 13209 24961 13243
rect 24961 13209 24995 13243
rect 24995 13209 25004 13243
rect 24952 13200 25004 13209
rect 24400 13132 24452 13184
rect 26516 13200 26568 13252
rect 27160 13132 27212 13184
rect 10425 13030 10477 13082
rect 10489 13030 10541 13082
rect 10553 13030 10605 13082
rect 10617 13030 10669 13082
rect 10681 13030 10733 13082
rect 19901 13030 19953 13082
rect 19965 13030 20017 13082
rect 20029 13030 20081 13082
rect 20093 13030 20145 13082
rect 20157 13030 20209 13082
rect 2872 12928 2924 12980
rect 3424 12928 3476 12980
rect 2412 12903 2464 12912
rect 2412 12869 2421 12903
rect 2421 12869 2455 12903
rect 2455 12869 2464 12903
rect 2412 12860 2464 12869
rect 2688 12860 2740 12912
rect 4068 12928 4120 12980
rect 4436 12928 4488 12980
rect 4804 12928 4856 12980
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 5448 12971 5500 12980
rect 5448 12937 5457 12971
rect 5457 12937 5491 12971
rect 5491 12937 5500 12971
rect 5448 12928 5500 12937
rect 1768 12792 1820 12844
rect 5080 12860 5132 12912
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 5172 12792 5224 12844
rect 5356 12835 5408 12844
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 4528 12724 4580 12776
rect 5448 12724 5500 12776
rect 6920 12792 6972 12844
rect 9680 12792 9732 12844
rect 10876 12860 10928 12912
rect 9956 12792 10008 12844
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 13544 12928 13596 12980
rect 14372 12928 14424 12980
rect 12808 12903 12860 12912
rect 12808 12869 12817 12903
rect 12817 12869 12851 12903
rect 12851 12869 12860 12903
rect 12808 12860 12860 12869
rect 13820 12860 13872 12912
rect 16764 12860 16816 12912
rect 15016 12835 15068 12844
rect 15016 12801 15025 12835
rect 15025 12801 15059 12835
rect 15059 12801 15068 12835
rect 15016 12792 15068 12801
rect 16672 12792 16724 12844
rect 20536 12860 20588 12912
rect 25044 12928 25096 12980
rect 25228 12928 25280 12980
rect 26516 12971 26568 12980
rect 24400 12903 24452 12912
rect 20444 12792 20496 12844
rect 22376 12835 22428 12844
rect 22376 12801 22385 12835
rect 22385 12801 22419 12835
rect 22419 12801 22428 12835
rect 22376 12792 22428 12801
rect 24400 12869 24409 12903
rect 24409 12869 24443 12903
rect 24443 12869 24452 12903
rect 24400 12860 24452 12869
rect 25412 12860 25464 12912
rect 26516 12937 26525 12971
rect 26525 12937 26559 12971
rect 26559 12937 26568 12971
rect 26516 12928 26568 12937
rect 27068 12860 27120 12912
rect 2780 12656 2832 12708
rect 6644 12656 6696 12708
rect 12072 12724 12124 12776
rect 13544 12724 13596 12776
rect 23296 12724 23348 12776
rect 24492 12724 24544 12776
rect 12532 12656 12584 12708
rect 5540 12588 5592 12640
rect 9312 12588 9364 12640
rect 13360 12588 13412 12640
rect 18236 12588 18288 12640
rect 19248 12588 19300 12640
rect 20720 12588 20772 12640
rect 21180 12588 21232 12640
rect 22468 12631 22520 12640
rect 22468 12597 22477 12631
rect 22477 12597 22511 12631
rect 22511 12597 22520 12631
rect 22468 12588 22520 12597
rect 5688 12486 5740 12538
rect 5752 12486 5804 12538
rect 5816 12486 5868 12538
rect 5880 12486 5932 12538
rect 5944 12486 5996 12538
rect 15163 12486 15215 12538
rect 15227 12486 15279 12538
rect 15291 12486 15343 12538
rect 15355 12486 15407 12538
rect 15419 12486 15471 12538
rect 24639 12486 24691 12538
rect 24703 12486 24755 12538
rect 24767 12486 24819 12538
rect 24831 12486 24883 12538
rect 24895 12486 24947 12538
rect 4436 12384 4488 12436
rect 5080 12384 5132 12436
rect 14280 12427 14332 12436
rect 4988 12316 5040 12368
rect 4804 12248 4856 12300
rect 5540 12291 5592 12300
rect 5540 12257 5549 12291
rect 5549 12257 5583 12291
rect 5583 12257 5592 12291
rect 5540 12248 5592 12257
rect 2780 12180 2832 12232
rect 4528 12180 4580 12232
rect 4068 12112 4120 12164
rect 3884 12044 3936 12096
rect 5540 12112 5592 12164
rect 6092 12180 6144 12232
rect 8300 12316 8352 12368
rect 8944 12316 8996 12368
rect 9588 12316 9640 12368
rect 9956 12316 10008 12368
rect 10784 12359 10836 12368
rect 10784 12325 10793 12359
rect 10793 12325 10827 12359
rect 10827 12325 10836 12359
rect 10784 12316 10836 12325
rect 11520 12316 11572 12368
rect 8484 12248 8536 12300
rect 6368 12180 6420 12232
rect 6644 12180 6696 12232
rect 8392 12180 8444 12232
rect 7656 12112 7708 12164
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 8760 12044 8812 12096
rect 8852 12044 8904 12096
rect 10324 12248 10376 12300
rect 11888 12248 11940 12300
rect 10784 12180 10836 12232
rect 11612 12180 11664 12232
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 12900 12316 12952 12368
rect 14280 12393 14289 12427
rect 14289 12393 14323 12427
rect 14323 12393 14332 12427
rect 14280 12384 14332 12393
rect 14464 12384 14516 12436
rect 14832 12384 14884 12436
rect 16672 12384 16724 12436
rect 19248 12384 19300 12436
rect 22376 12427 22428 12436
rect 22376 12393 22385 12427
rect 22385 12393 22419 12427
rect 22419 12393 22428 12427
rect 22376 12384 22428 12393
rect 25412 12384 25464 12436
rect 12624 12180 12676 12232
rect 13820 12180 13872 12232
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 15476 12248 15528 12300
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 19340 12248 19392 12300
rect 22744 12316 22796 12368
rect 20444 12291 20496 12300
rect 11060 12112 11112 12164
rect 13728 12112 13780 12164
rect 15660 12180 15712 12232
rect 16396 12180 16448 12232
rect 16764 12180 16816 12232
rect 18236 12180 18288 12232
rect 19156 12180 19208 12232
rect 20444 12257 20453 12291
rect 20453 12257 20487 12291
rect 20487 12257 20496 12291
rect 20444 12248 20496 12257
rect 14648 12112 14700 12164
rect 15292 12112 15344 12164
rect 11336 12044 11388 12096
rect 11796 12044 11848 12096
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 12072 12044 12124 12096
rect 13544 12044 13596 12096
rect 16580 12087 16632 12096
rect 16580 12053 16589 12087
rect 16589 12053 16623 12087
rect 16623 12053 16632 12087
rect 16580 12044 16632 12053
rect 19524 12112 19576 12164
rect 19708 12155 19760 12164
rect 19708 12121 19717 12155
rect 19717 12121 19751 12155
rect 19751 12121 19760 12155
rect 19708 12112 19760 12121
rect 20260 12180 20312 12232
rect 21272 12248 21324 12300
rect 20720 12180 20772 12232
rect 21180 12223 21232 12232
rect 21180 12189 21189 12223
rect 21189 12189 21223 12223
rect 21223 12189 21232 12223
rect 21180 12180 21232 12189
rect 21640 12223 21692 12232
rect 21640 12189 21649 12223
rect 21649 12189 21683 12223
rect 21683 12189 21692 12223
rect 21640 12180 21692 12189
rect 21456 12112 21508 12164
rect 22192 12180 22244 12232
rect 22468 12180 22520 12232
rect 25044 12248 25096 12300
rect 24492 12180 24544 12232
rect 10425 11942 10477 11994
rect 10489 11942 10541 11994
rect 10553 11942 10605 11994
rect 10617 11942 10669 11994
rect 10681 11942 10733 11994
rect 19901 11942 19953 11994
rect 19965 11942 20017 11994
rect 20029 11942 20081 11994
rect 20093 11942 20145 11994
rect 20157 11942 20209 11994
rect 3792 11883 3844 11892
rect 3792 11849 3801 11883
rect 3801 11849 3835 11883
rect 3835 11849 3844 11883
rect 3792 11840 3844 11849
rect 3424 11815 3476 11824
rect 3424 11781 3433 11815
rect 3433 11781 3467 11815
rect 3467 11781 3476 11815
rect 3424 11772 3476 11781
rect 3884 11772 3936 11824
rect 5172 11840 5224 11892
rect 4436 11704 4488 11756
rect 4896 11704 4948 11756
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 7564 11840 7616 11892
rect 8392 11883 8444 11892
rect 6000 11772 6052 11824
rect 8392 11849 8401 11883
rect 8401 11849 8435 11883
rect 8435 11849 8444 11883
rect 8392 11840 8444 11849
rect 10784 11840 10836 11892
rect 11336 11840 11388 11892
rect 3884 11679 3936 11688
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 4712 11679 4764 11688
rect 4712 11645 4721 11679
rect 4721 11645 4755 11679
rect 4755 11645 4764 11679
rect 4712 11636 4764 11645
rect 5908 11747 5960 11756
rect 5908 11713 5922 11747
rect 5922 11713 5956 11747
rect 5956 11713 5960 11747
rect 5908 11704 5960 11713
rect 6092 11704 6144 11756
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 4252 11568 4304 11620
rect 3976 11500 4028 11552
rect 6276 11636 6328 11688
rect 6920 11704 6972 11756
rect 9864 11772 9916 11824
rect 6184 11568 6236 11620
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 8944 11747 8996 11756
rect 8944 11713 8953 11747
rect 8953 11713 8987 11747
rect 8987 11713 8996 11747
rect 8944 11704 8996 11713
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 9956 11747 10008 11756
rect 7932 11611 7984 11620
rect 7932 11577 7941 11611
rect 7941 11577 7975 11611
rect 7975 11577 7984 11611
rect 7932 11568 7984 11577
rect 6736 11500 6788 11552
rect 8208 11500 8260 11552
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 13084 11840 13136 11892
rect 15292 11883 15344 11892
rect 15292 11849 15301 11883
rect 15301 11849 15335 11883
rect 15335 11849 15344 11883
rect 15292 11840 15344 11849
rect 15844 11840 15896 11892
rect 16948 11840 17000 11892
rect 19800 11883 19852 11892
rect 19800 11849 19809 11883
rect 19809 11849 19843 11883
rect 19843 11849 19852 11883
rect 21456 11883 21508 11892
rect 19800 11840 19852 11849
rect 16580 11772 16632 11824
rect 12164 11747 12216 11756
rect 12164 11713 12173 11747
rect 12173 11713 12207 11747
rect 12207 11713 12216 11747
rect 12164 11704 12216 11713
rect 11520 11636 11572 11688
rect 11796 11636 11848 11688
rect 13728 11636 13780 11688
rect 15568 11704 15620 11756
rect 19248 11704 19300 11756
rect 20720 11772 20772 11824
rect 21456 11849 21465 11883
rect 21465 11849 21499 11883
rect 21499 11849 21508 11883
rect 21456 11840 21508 11849
rect 21640 11840 21692 11892
rect 21180 11772 21232 11824
rect 15844 11636 15896 11688
rect 10784 11568 10836 11620
rect 10968 11568 11020 11620
rect 12256 11611 12308 11620
rect 9864 11500 9916 11552
rect 11152 11500 11204 11552
rect 11612 11500 11664 11552
rect 12256 11577 12265 11611
rect 12265 11577 12299 11611
rect 12299 11577 12308 11611
rect 12256 11568 12308 11577
rect 15292 11568 15344 11620
rect 15752 11568 15804 11620
rect 12532 11543 12584 11552
rect 12532 11509 12541 11543
rect 12541 11509 12575 11543
rect 12575 11509 12584 11543
rect 12532 11500 12584 11509
rect 20720 11636 20772 11688
rect 20260 11611 20312 11620
rect 20260 11577 20269 11611
rect 20269 11577 20303 11611
rect 20303 11577 20312 11611
rect 20260 11568 20312 11577
rect 20812 11568 20864 11620
rect 19340 11500 19392 11552
rect 19616 11500 19668 11552
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 22284 11747 22336 11756
rect 22284 11713 22293 11747
rect 22293 11713 22327 11747
rect 22327 11713 22336 11747
rect 22560 11747 22612 11756
rect 22284 11704 22336 11713
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 27252 11747 27304 11756
rect 27252 11713 27286 11747
rect 27286 11713 27304 11747
rect 27252 11704 27304 11713
rect 25044 11636 25096 11688
rect 22284 11568 22336 11620
rect 21180 11543 21232 11552
rect 21180 11509 21189 11543
rect 21189 11509 21223 11543
rect 21223 11509 21232 11543
rect 21180 11500 21232 11509
rect 23020 11543 23072 11552
rect 23020 11509 23029 11543
rect 23029 11509 23063 11543
rect 23063 11509 23072 11543
rect 23020 11500 23072 11509
rect 28356 11543 28408 11552
rect 28356 11509 28365 11543
rect 28365 11509 28399 11543
rect 28399 11509 28408 11543
rect 28356 11500 28408 11509
rect 5688 11398 5740 11450
rect 5752 11398 5804 11450
rect 5816 11398 5868 11450
rect 5880 11398 5932 11450
rect 5944 11398 5996 11450
rect 15163 11398 15215 11450
rect 15227 11398 15279 11450
rect 15291 11398 15343 11450
rect 15355 11398 15407 11450
rect 15419 11398 15471 11450
rect 24639 11398 24691 11450
rect 24703 11398 24755 11450
rect 24767 11398 24819 11450
rect 24831 11398 24883 11450
rect 24895 11398 24947 11450
rect 3792 11296 3844 11348
rect 1952 11271 2004 11280
rect 1952 11237 1961 11271
rect 1961 11237 1995 11271
rect 1995 11237 2004 11271
rect 1952 11228 2004 11237
rect 4160 11160 4212 11212
rect 4712 11160 4764 11212
rect 6092 11228 6144 11280
rect 6736 11296 6788 11348
rect 8944 11296 8996 11348
rect 9128 11296 9180 11348
rect 10140 11296 10192 11348
rect 11336 11296 11388 11348
rect 11612 11296 11664 11348
rect 12164 11296 12216 11348
rect 13728 11296 13780 11348
rect 14648 11339 14700 11348
rect 7012 11228 7064 11280
rect 7656 11271 7708 11280
rect 7656 11237 7665 11271
rect 7665 11237 7699 11271
rect 7699 11237 7708 11271
rect 7656 11228 7708 11237
rect 10968 11228 11020 11280
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 4252 11092 4304 11144
rect 5540 11092 5592 11144
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 6184 11135 6236 11144
rect 6184 11101 6198 11135
rect 6198 11101 6232 11135
rect 6232 11101 6236 11135
rect 6184 11092 6236 11101
rect 7472 11092 7524 11144
rect 9220 11160 9272 11212
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8300 11135 8352 11144
rect 8116 11092 8168 11101
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 10140 11203 10192 11212
rect 10140 11169 10149 11203
rect 10149 11169 10183 11203
rect 10183 11169 10192 11203
rect 10140 11160 10192 11169
rect 10324 11135 10376 11144
rect 1492 10956 1544 11008
rect 5264 10999 5316 11008
rect 5264 10965 5273 10999
rect 5273 10965 5307 10999
rect 5307 10965 5316 10999
rect 5264 10956 5316 10965
rect 9036 11024 9088 11076
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 11152 11092 11204 11144
rect 11704 11203 11756 11212
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 11796 11203 11848 11212
rect 11796 11169 11805 11203
rect 11805 11169 11839 11203
rect 11839 11169 11848 11203
rect 11796 11160 11848 11169
rect 12532 11160 12584 11212
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 14648 11305 14657 11339
rect 14657 11305 14691 11339
rect 14691 11305 14700 11339
rect 14648 11296 14700 11305
rect 14740 11296 14792 11348
rect 15568 11339 15620 11348
rect 15568 11305 15577 11339
rect 15577 11305 15611 11339
rect 15611 11305 15620 11339
rect 15568 11296 15620 11305
rect 18144 11296 18196 11348
rect 19248 11296 19300 11348
rect 19524 11296 19576 11348
rect 15384 11160 15436 11212
rect 11520 11135 11572 11144
rect 10232 11024 10284 11076
rect 10968 11024 11020 11076
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 12256 11092 12308 11144
rect 13544 11092 13596 11144
rect 13912 11092 13964 11144
rect 14648 11135 14700 11144
rect 14648 11101 14657 11135
rect 14657 11101 14691 11135
rect 14691 11101 14700 11135
rect 14648 11092 14700 11101
rect 15752 11135 15804 11144
rect 11796 11024 11848 11076
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 19800 11160 19852 11212
rect 16672 11092 16724 11144
rect 19340 11092 19392 11144
rect 15568 11024 15620 11076
rect 15844 11024 15896 11076
rect 6276 10956 6328 11008
rect 7196 10999 7248 11008
rect 7196 10965 7205 10999
rect 7205 10965 7239 10999
rect 7239 10965 7248 10999
rect 7196 10956 7248 10965
rect 10876 10956 10928 11008
rect 11888 10956 11940 11008
rect 15108 10956 15160 11008
rect 15292 10956 15344 11008
rect 18052 11024 18104 11076
rect 19616 11135 19668 11144
rect 19616 11101 19625 11135
rect 19625 11101 19659 11135
rect 19659 11101 19668 11135
rect 19616 11092 19668 11101
rect 20812 11296 20864 11348
rect 22284 11296 22336 11348
rect 27252 11339 27304 11348
rect 27252 11305 27261 11339
rect 27261 11305 27295 11339
rect 27295 11305 27304 11339
rect 27252 11296 27304 11305
rect 21272 11160 21324 11212
rect 20720 11092 20772 11144
rect 20996 11092 21048 11144
rect 21364 11092 21416 11144
rect 23112 11092 23164 11144
rect 23848 11135 23900 11144
rect 23848 11101 23857 11135
rect 23857 11101 23891 11135
rect 23891 11101 23900 11135
rect 23848 11092 23900 11101
rect 24032 11135 24084 11144
rect 24032 11101 24041 11135
rect 24041 11101 24075 11135
rect 24075 11101 24084 11135
rect 24032 11092 24084 11101
rect 21456 11024 21508 11076
rect 22376 11024 22428 11076
rect 25044 11092 25096 11144
rect 26976 11135 27028 11144
rect 26976 11101 26985 11135
rect 26985 11101 27019 11135
rect 27019 11101 27028 11135
rect 26976 11092 27028 11101
rect 28448 11160 28500 11212
rect 24492 11024 24544 11076
rect 26056 11067 26108 11076
rect 26056 11033 26065 11067
rect 26065 11033 26099 11067
rect 26099 11033 26108 11067
rect 26056 11024 26108 11033
rect 26424 11067 26476 11076
rect 21364 10999 21416 11008
rect 21364 10965 21373 10999
rect 21373 10965 21407 10999
rect 21407 10965 21416 10999
rect 21364 10956 21416 10965
rect 22744 10956 22796 11008
rect 24768 10956 24820 11008
rect 26424 11033 26433 11067
rect 26433 11033 26467 11067
rect 26467 11033 26476 11067
rect 26424 11024 26476 11033
rect 27988 11092 28040 11144
rect 26332 10956 26384 11008
rect 27712 10999 27764 11008
rect 27712 10965 27721 10999
rect 27721 10965 27755 10999
rect 27755 10965 27764 10999
rect 27712 10956 27764 10965
rect 27896 10956 27948 11008
rect 10425 10854 10477 10906
rect 10489 10854 10541 10906
rect 10553 10854 10605 10906
rect 10617 10854 10669 10906
rect 10681 10854 10733 10906
rect 19901 10854 19953 10906
rect 19965 10854 20017 10906
rect 20029 10854 20081 10906
rect 20093 10854 20145 10906
rect 20157 10854 20209 10906
rect 4160 10795 4212 10804
rect 4160 10761 4169 10795
rect 4169 10761 4203 10795
rect 4203 10761 4212 10795
rect 4160 10752 4212 10761
rect 7472 10752 7524 10804
rect 8300 10752 8352 10804
rect 9680 10752 9732 10804
rect 10048 10752 10100 10804
rect 10324 10752 10376 10804
rect 11060 10752 11112 10804
rect 11612 10752 11664 10804
rect 13084 10795 13136 10804
rect 13084 10761 13093 10795
rect 13093 10761 13127 10795
rect 13127 10761 13136 10795
rect 13084 10752 13136 10761
rect 14648 10752 14700 10804
rect 15292 10752 15344 10804
rect 16488 10752 16540 10804
rect 16948 10752 17000 10804
rect 17316 10752 17368 10804
rect 18052 10752 18104 10804
rect 5816 10684 5868 10736
rect 8392 10684 8444 10736
rect 9956 10727 10008 10736
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 1860 10616 1912 10668
rect 3148 10616 3200 10668
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 5540 10616 5592 10668
rect 1676 10548 1728 10600
rect 7748 10616 7800 10668
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 9956 10693 9965 10727
rect 9965 10693 9999 10727
rect 9999 10693 10008 10727
rect 9956 10684 10008 10693
rect 10140 10727 10192 10736
rect 10140 10693 10149 10727
rect 10149 10693 10183 10727
rect 10183 10693 10192 10727
rect 10140 10684 10192 10693
rect 10232 10684 10284 10736
rect 19340 10727 19392 10736
rect 8116 10548 8168 10600
rect 2136 10412 2188 10464
rect 3240 10412 3292 10464
rect 4068 10412 4120 10464
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 9220 10455 9272 10464
rect 9220 10421 9229 10455
rect 9229 10421 9263 10455
rect 9263 10421 9272 10455
rect 9220 10412 9272 10421
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 10048 10616 10100 10668
rect 10508 10616 10560 10668
rect 10876 10616 10928 10668
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12072 10616 12124 10668
rect 10968 10591 11020 10600
rect 10416 10480 10468 10532
rect 10692 10412 10744 10464
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 11060 10548 11112 10600
rect 19340 10693 19349 10727
rect 19349 10693 19383 10727
rect 19383 10693 19392 10727
rect 19340 10684 19392 10693
rect 19708 10684 19760 10736
rect 13728 10616 13780 10668
rect 14832 10659 14884 10668
rect 14832 10625 14841 10659
rect 14841 10625 14875 10659
rect 14875 10625 14884 10659
rect 14832 10616 14884 10625
rect 15200 10659 15252 10668
rect 15200 10625 15209 10659
rect 15209 10625 15243 10659
rect 15243 10625 15252 10659
rect 15200 10616 15252 10625
rect 15384 10659 15436 10668
rect 15384 10625 15393 10659
rect 15393 10625 15427 10659
rect 15427 10625 15436 10659
rect 15384 10616 15436 10625
rect 18144 10659 18196 10668
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 18144 10625 18153 10659
rect 18153 10625 18187 10659
rect 18187 10625 18196 10659
rect 18144 10616 18196 10625
rect 18328 10616 18380 10668
rect 10876 10480 10928 10532
rect 15660 10480 15712 10532
rect 17408 10480 17460 10532
rect 18420 10548 18472 10600
rect 20444 10616 20496 10668
rect 21180 10616 21232 10668
rect 21456 10616 21508 10668
rect 22376 10616 22428 10668
rect 23112 10752 23164 10804
rect 24492 10752 24544 10804
rect 24768 10795 24820 10804
rect 24768 10761 24777 10795
rect 24777 10761 24811 10795
rect 24811 10761 24820 10795
rect 24768 10752 24820 10761
rect 27712 10795 27764 10804
rect 27712 10761 27721 10795
rect 27721 10761 27755 10795
rect 27755 10761 27764 10795
rect 27712 10752 27764 10761
rect 15752 10412 15804 10464
rect 21272 10480 21324 10532
rect 24492 10616 24544 10668
rect 26056 10616 26108 10668
rect 26424 10684 26476 10736
rect 26976 10727 27028 10736
rect 26700 10659 26752 10668
rect 23388 10548 23440 10600
rect 26332 10548 26384 10600
rect 26700 10625 26709 10659
rect 26709 10625 26743 10659
rect 26743 10625 26752 10659
rect 26700 10616 26752 10625
rect 26976 10693 26985 10727
rect 26985 10693 27019 10727
rect 27019 10693 27028 10727
rect 26976 10684 27028 10693
rect 28356 10684 28408 10736
rect 27896 10659 27948 10668
rect 27896 10625 27905 10659
rect 27905 10625 27939 10659
rect 27939 10625 27948 10659
rect 27896 10616 27948 10625
rect 25504 10480 25556 10532
rect 26700 10480 26752 10532
rect 26792 10480 26844 10532
rect 21548 10455 21600 10464
rect 21548 10421 21557 10455
rect 21557 10421 21591 10455
rect 21591 10421 21600 10455
rect 21548 10412 21600 10421
rect 21640 10412 21692 10464
rect 27528 10412 27580 10464
rect 5688 10310 5740 10362
rect 5752 10310 5804 10362
rect 5816 10310 5868 10362
rect 5880 10310 5932 10362
rect 5944 10310 5996 10362
rect 15163 10310 15215 10362
rect 15227 10310 15279 10362
rect 15291 10310 15343 10362
rect 15355 10310 15407 10362
rect 15419 10310 15471 10362
rect 24639 10310 24691 10362
rect 24703 10310 24755 10362
rect 24767 10310 24819 10362
rect 24831 10310 24883 10362
rect 24895 10310 24947 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 4528 10208 4580 10260
rect 7748 10208 7800 10260
rect 10324 10251 10376 10260
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 14832 10208 14884 10260
rect 16580 10208 16632 10260
rect 17684 10208 17736 10260
rect 24032 10208 24084 10260
rect 26332 10208 26384 10260
rect 1952 10072 2004 10124
rect 2136 10004 2188 10056
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 3976 10140 4028 10192
rect 4436 10115 4488 10124
rect 2412 10072 2464 10081
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 6000 10115 6052 10124
rect 6000 10081 6009 10115
rect 6009 10081 6043 10115
rect 6043 10081 6052 10115
rect 6000 10072 6052 10081
rect 10048 10140 10100 10192
rect 12716 10183 12768 10192
rect 12716 10149 12725 10183
rect 12725 10149 12759 10183
rect 12759 10149 12768 10183
rect 12716 10140 12768 10149
rect 3608 9979 3660 9988
rect 3608 9945 3617 9979
rect 3617 9945 3651 9979
rect 3651 9945 3660 9979
rect 3608 9936 3660 9945
rect 4160 10004 4212 10056
rect 6092 10004 6144 10056
rect 6368 10004 6420 10056
rect 8852 10072 8904 10124
rect 10416 10072 10468 10124
rect 10876 10115 10928 10124
rect 4344 9936 4396 9988
rect 4620 9936 4672 9988
rect 5264 9936 5316 9988
rect 8484 10004 8536 10056
rect 8944 10047 8996 10056
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 9220 10047 9272 10056
rect 9220 10013 9254 10047
rect 9254 10013 9272 10047
rect 9220 10004 9272 10013
rect 10876 10081 10885 10115
rect 10885 10081 10919 10115
rect 10919 10081 10928 10115
rect 10876 10072 10928 10081
rect 10968 10072 11020 10124
rect 21640 10140 21692 10192
rect 10968 9936 11020 9988
rect 4068 9868 4120 9920
rect 4252 9911 4304 9920
rect 4252 9877 4261 9911
rect 4261 9877 4295 9911
rect 4295 9877 4304 9911
rect 4988 9911 5040 9920
rect 4252 9868 4304 9877
rect 4988 9877 4997 9911
rect 4997 9877 5031 9911
rect 5031 9877 5040 9911
rect 4988 9868 5040 9877
rect 5448 9911 5500 9920
rect 5448 9877 5457 9911
rect 5457 9877 5491 9911
rect 5491 9877 5500 9911
rect 5448 9868 5500 9877
rect 7104 9868 7156 9920
rect 11244 10004 11296 10056
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 13820 10004 13872 10056
rect 17316 10072 17368 10124
rect 18328 10115 18380 10124
rect 18328 10081 18337 10115
rect 18337 10081 18371 10115
rect 18371 10081 18380 10115
rect 18328 10072 18380 10081
rect 19708 10072 19760 10124
rect 16672 10004 16724 10056
rect 11244 9868 11296 9920
rect 11796 9868 11848 9920
rect 16028 9936 16080 9988
rect 18144 10004 18196 10056
rect 16304 9911 16356 9920
rect 16304 9877 16313 9911
rect 16313 9877 16347 9911
rect 16347 9877 16356 9911
rect 16304 9868 16356 9877
rect 16580 9868 16632 9920
rect 19800 10047 19852 10056
rect 19800 10013 19809 10047
rect 19809 10013 19843 10047
rect 19843 10013 19852 10047
rect 19800 10004 19852 10013
rect 20444 10004 20496 10056
rect 21364 10047 21416 10056
rect 21364 10013 21373 10047
rect 21373 10013 21407 10047
rect 21407 10013 21416 10047
rect 21364 10004 21416 10013
rect 21548 10072 21600 10124
rect 22376 10115 22428 10124
rect 22376 10081 22385 10115
rect 22385 10081 22419 10115
rect 22419 10081 22428 10115
rect 22376 10072 22428 10081
rect 23020 10072 23072 10124
rect 26516 10072 26568 10124
rect 27988 10072 28040 10124
rect 22744 10047 22796 10056
rect 22744 10013 22753 10047
rect 22753 10013 22787 10047
rect 22787 10013 22796 10047
rect 22744 10004 22796 10013
rect 24492 10004 24544 10056
rect 24860 10047 24912 10056
rect 24860 10013 24869 10047
rect 24869 10013 24903 10047
rect 24903 10013 24912 10047
rect 24860 10004 24912 10013
rect 26700 10047 26752 10056
rect 26700 10013 26709 10047
rect 26709 10013 26743 10047
rect 26743 10013 26752 10047
rect 26700 10004 26752 10013
rect 26976 9979 27028 9988
rect 19064 9911 19116 9920
rect 19064 9877 19073 9911
rect 19073 9877 19107 9911
rect 19107 9877 19116 9911
rect 19064 9868 19116 9877
rect 19616 9868 19668 9920
rect 26976 9945 26985 9979
rect 26985 9945 27019 9979
rect 27019 9945 27028 9979
rect 26976 9936 27028 9945
rect 27620 9936 27672 9988
rect 22284 9868 22336 9920
rect 26792 9868 26844 9920
rect 28356 9868 28408 9920
rect 10425 9766 10477 9818
rect 10489 9766 10541 9818
rect 10553 9766 10605 9818
rect 10617 9766 10669 9818
rect 10681 9766 10733 9818
rect 19901 9766 19953 9818
rect 19965 9766 20017 9818
rect 20029 9766 20081 9818
rect 20093 9766 20145 9818
rect 20157 9766 20209 9818
rect 2412 9664 2464 9716
rect 4804 9664 4856 9716
rect 6000 9664 6052 9716
rect 10324 9664 10376 9716
rect 1676 9596 1728 9648
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 3424 9528 3476 9580
rect 6368 9596 6420 9648
rect 7932 9596 7984 9648
rect 8944 9596 8996 9648
rect 9588 9596 9640 9648
rect 5448 9528 5500 9580
rect 8116 9528 8168 9580
rect 10784 9596 10836 9648
rect 13912 9639 13964 9648
rect 13912 9605 13921 9639
rect 13921 9605 13955 9639
rect 13955 9605 13964 9639
rect 13912 9596 13964 9605
rect 14556 9596 14608 9648
rect 24860 9664 24912 9716
rect 15660 9596 15712 9648
rect 17224 9639 17276 9648
rect 11060 9528 11112 9580
rect 11980 9528 12032 9580
rect 12072 9528 12124 9580
rect 12716 9571 12768 9580
rect 12716 9537 12725 9571
rect 12725 9537 12759 9571
rect 12759 9537 12768 9571
rect 12716 9528 12768 9537
rect 14924 9528 14976 9580
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 2780 9392 2832 9444
rect 3608 9392 3660 9444
rect 6368 9392 6420 9444
rect 6552 9435 6604 9444
rect 6552 9401 6561 9435
rect 6561 9401 6595 9435
rect 6595 9401 6604 9435
rect 6552 9392 6604 9401
rect 7012 9435 7064 9444
rect 7012 9401 7021 9435
rect 7021 9401 7055 9435
rect 7055 9401 7064 9435
rect 7012 9392 7064 9401
rect 11336 9435 11388 9444
rect 11336 9401 11345 9435
rect 11345 9401 11379 9435
rect 11379 9401 11388 9435
rect 11336 9392 11388 9401
rect 1400 9324 1452 9376
rect 3792 9367 3844 9376
rect 3792 9333 3801 9367
rect 3801 9333 3835 9367
rect 3835 9333 3844 9367
rect 3792 9324 3844 9333
rect 6092 9367 6144 9376
rect 6092 9333 6101 9367
rect 6101 9333 6135 9367
rect 6135 9333 6144 9367
rect 6092 9324 6144 9333
rect 11152 9324 11204 9376
rect 11244 9324 11296 9376
rect 13084 9460 13136 9512
rect 12256 9392 12308 9444
rect 15476 9460 15528 9512
rect 15752 9503 15804 9512
rect 15752 9469 15761 9503
rect 15761 9469 15795 9503
rect 15795 9469 15804 9503
rect 15752 9460 15804 9469
rect 17224 9605 17233 9639
rect 17233 9605 17267 9639
rect 17267 9605 17276 9639
rect 17224 9596 17276 9605
rect 16212 9528 16264 9580
rect 16488 9528 16540 9580
rect 17132 9528 17184 9580
rect 19156 9596 19208 9648
rect 19800 9639 19852 9648
rect 19800 9605 19809 9639
rect 19809 9605 19843 9639
rect 19843 9605 19852 9639
rect 19800 9596 19852 9605
rect 19984 9596 20036 9648
rect 20260 9596 20312 9648
rect 17776 9571 17828 9580
rect 17776 9537 17785 9571
rect 17785 9537 17819 9571
rect 17819 9537 17828 9571
rect 17776 9528 17828 9537
rect 18512 9528 18564 9580
rect 19064 9571 19116 9580
rect 19064 9537 19073 9571
rect 19073 9537 19107 9571
rect 19107 9537 19116 9571
rect 19064 9528 19116 9537
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 15844 9392 15896 9444
rect 17316 9392 17368 9444
rect 17592 9392 17644 9444
rect 11704 9324 11756 9376
rect 14924 9324 14976 9376
rect 15660 9324 15712 9376
rect 16120 9324 16172 9376
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 20536 9528 20588 9580
rect 20720 9596 20772 9648
rect 22284 9639 22336 9648
rect 20812 9528 20864 9580
rect 20720 9503 20772 9512
rect 20720 9469 20729 9503
rect 20729 9469 20763 9503
rect 20763 9469 20772 9503
rect 20720 9460 20772 9469
rect 18420 9324 18472 9376
rect 20168 9324 20220 9376
rect 22284 9605 22293 9639
rect 22293 9605 22327 9639
rect 22327 9605 22336 9639
rect 22284 9596 22336 9605
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 22560 9528 22612 9580
rect 23112 9528 23164 9580
rect 27896 9596 27948 9648
rect 25964 9571 26016 9580
rect 25964 9537 25973 9571
rect 25973 9537 26007 9571
rect 26007 9537 26016 9571
rect 25964 9528 26016 9537
rect 26240 9571 26292 9580
rect 26240 9537 26249 9571
rect 26249 9537 26283 9571
rect 26283 9537 26292 9571
rect 26516 9571 26568 9580
rect 26240 9528 26292 9537
rect 26516 9537 26525 9571
rect 26525 9537 26559 9571
rect 26559 9537 26568 9571
rect 26516 9528 26568 9537
rect 22008 9460 22060 9512
rect 21916 9392 21968 9444
rect 26056 9460 26108 9512
rect 26976 9528 27028 9580
rect 27988 9571 28040 9580
rect 27988 9537 28022 9571
rect 28022 9537 28040 9571
rect 24860 9392 24912 9444
rect 25780 9392 25832 9444
rect 26976 9392 27028 9444
rect 22744 9324 22796 9376
rect 23756 9324 23808 9376
rect 26148 9367 26200 9376
rect 26148 9333 26157 9367
rect 26157 9333 26191 9367
rect 26191 9333 26200 9367
rect 26148 9324 26200 9333
rect 27160 9324 27212 9376
rect 27988 9528 28040 9537
rect 27712 9503 27764 9512
rect 27712 9469 27721 9503
rect 27721 9469 27755 9503
rect 27755 9469 27764 9503
rect 27712 9460 27764 9469
rect 5688 9222 5740 9274
rect 5752 9222 5804 9274
rect 5816 9222 5868 9274
rect 5880 9222 5932 9274
rect 5944 9222 5996 9274
rect 15163 9222 15215 9274
rect 15227 9222 15279 9274
rect 15291 9222 15343 9274
rect 15355 9222 15407 9274
rect 15419 9222 15471 9274
rect 24639 9222 24691 9274
rect 24703 9222 24755 9274
rect 24767 9222 24819 9274
rect 24831 9222 24883 9274
rect 24895 9222 24947 9274
rect 3608 9120 3660 9172
rect 7564 9120 7616 9172
rect 12900 9120 12952 9172
rect 14924 9120 14976 9172
rect 15568 9120 15620 9172
rect 16396 9120 16448 9172
rect 3424 9052 3476 9104
rect 3700 9052 3752 9104
rect 7840 9052 7892 9104
rect 16304 9095 16356 9104
rect 16304 9061 16313 9095
rect 16313 9061 16347 9095
rect 16347 9061 16356 9095
rect 16304 9052 16356 9061
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 3792 8984 3844 9036
rect 10324 8984 10376 9036
rect 11060 8984 11112 9036
rect 11520 8984 11572 9036
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 1952 8891 2004 8900
rect 1952 8857 1986 8891
rect 1986 8857 2004 8891
rect 3608 8891 3660 8900
rect 1952 8848 2004 8857
rect 3608 8857 3617 8891
rect 3617 8857 3651 8891
rect 3651 8857 3660 8891
rect 3608 8848 3660 8857
rect 7472 8916 7524 8968
rect 10876 8916 10928 8968
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 11612 8959 11664 8968
rect 4436 8891 4488 8900
rect 4436 8857 4445 8891
rect 4445 8857 4479 8891
rect 4479 8857 4488 8891
rect 4436 8848 4488 8857
rect 5080 8848 5132 8900
rect 7104 8848 7156 8900
rect 8024 8848 8076 8900
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 11704 8959 11756 8968
rect 11704 8925 11713 8959
rect 11713 8925 11747 8959
rect 11747 8925 11756 8959
rect 12256 8959 12308 8968
rect 11704 8916 11756 8925
rect 12256 8925 12290 8959
rect 12290 8925 12308 8959
rect 12256 8916 12308 8925
rect 15016 8916 15068 8968
rect 16672 8984 16724 9036
rect 15660 8959 15712 8968
rect 15660 8925 15669 8959
rect 15669 8925 15703 8959
rect 15703 8925 15712 8959
rect 15660 8916 15712 8925
rect 15936 8959 15988 8968
rect 15936 8925 15945 8959
rect 15945 8925 15979 8959
rect 15979 8925 15988 8959
rect 15936 8916 15988 8925
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 16488 8959 16540 8968
rect 16488 8925 16497 8959
rect 16497 8925 16531 8959
rect 16531 8925 16540 8959
rect 16488 8916 16540 8925
rect 16580 8959 16632 8968
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 17224 9120 17276 9172
rect 17316 9120 17368 9172
rect 17868 9120 17920 9172
rect 18144 9052 18196 9104
rect 16580 8916 16632 8925
rect 17592 9027 17644 9036
rect 17592 8993 17601 9027
rect 17601 8993 17635 9027
rect 17635 8993 17644 9027
rect 17592 8984 17644 8993
rect 18144 8959 18196 8968
rect 18144 8925 18153 8959
rect 18153 8925 18187 8959
rect 18187 8925 18196 8959
rect 18144 8916 18196 8925
rect 19340 9120 19392 9172
rect 19524 9120 19576 9172
rect 20720 9163 20772 9172
rect 12164 8848 12216 8900
rect 2228 8780 2280 8832
rect 10048 8780 10100 8832
rect 10876 8780 10928 8832
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 23112 9163 23164 9172
rect 23112 9129 23121 9163
rect 23121 9129 23155 9163
rect 23155 9129 23164 9163
rect 23112 9120 23164 9129
rect 27620 9163 27672 9172
rect 27620 9129 27629 9163
rect 27629 9129 27663 9163
rect 27663 9129 27672 9163
rect 27620 9120 27672 9129
rect 27988 9120 28040 9172
rect 21548 9095 21600 9104
rect 21548 9061 21557 9095
rect 21557 9061 21591 9095
rect 21591 9061 21600 9095
rect 21548 9052 21600 9061
rect 23388 9052 23440 9104
rect 19616 8984 19668 9036
rect 21916 8984 21968 9036
rect 22744 9027 22796 9036
rect 22744 8993 22753 9027
rect 22753 8993 22787 9027
rect 22787 8993 22796 9027
rect 22744 8984 22796 8993
rect 23112 8984 23164 9036
rect 23756 9027 23808 9036
rect 23756 8993 23765 9027
rect 23765 8993 23799 9027
rect 23799 8993 23808 9027
rect 23756 8984 23808 8993
rect 26240 9052 26292 9104
rect 18604 8959 18656 8968
rect 18604 8925 18613 8959
rect 18613 8925 18647 8959
rect 18647 8925 18656 8959
rect 18604 8916 18656 8925
rect 19064 8959 19116 8968
rect 19064 8925 19073 8959
rect 19073 8925 19107 8959
rect 19107 8925 19116 8959
rect 19064 8916 19116 8925
rect 22376 8959 22428 8968
rect 22376 8925 22385 8959
rect 22385 8925 22419 8959
rect 22419 8925 22428 8959
rect 22376 8916 22428 8925
rect 20720 8848 20772 8900
rect 17224 8780 17276 8832
rect 17500 8823 17552 8832
rect 17500 8789 17509 8823
rect 17509 8789 17543 8823
rect 17543 8789 17552 8823
rect 17500 8780 17552 8789
rect 19248 8780 19300 8832
rect 19708 8823 19760 8832
rect 19708 8789 19717 8823
rect 19717 8789 19751 8823
rect 19751 8789 19760 8823
rect 21824 8848 21876 8900
rect 21088 8823 21140 8832
rect 19708 8780 19760 8789
rect 21088 8789 21097 8823
rect 21097 8789 21131 8823
rect 21131 8789 21140 8823
rect 21088 8780 21140 8789
rect 22192 8848 22244 8900
rect 22560 8823 22612 8832
rect 22560 8789 22569 8823
rect 22569 8789 22603 8823
rect 22603 8789 22612 8823
rect 22560 8780 22612 8789
rect 23388 8780 23440 8832
rect 23664 8823 23716 8832
rect 23664 8789 23673 8823
rect 23673 8789 23707 8823
rect 23707 8789 23716 8823
rect 23664 8780 23716 8789
rect 24952 8916 25004 8968
rect 27712 8984 27764 9036
rect 28356 9027 28408 9036
rect 28356 8993 28365 9027
rect 28365 8993 28399 9027
rect 28399 8993 28408 9027
rect 28356 8984 28408 8993
rect 28448 9027 28500 9036
rect 28448 8993 28457 9027
rect 28457 8993 28491 9027
rect 28491 8993 28500 9027
rect 28448 8984 28500 8993
rect 26056 8916 26108 8968
rect 26516 8916 26568 8968
rect 26976 8959 27028 8968
rect 26976 8925 26985 8959
rect 26985 8925 27019 8959
rect 27019 8925 27028 8959
rect 26976 8916 27028 8925
rect 27160 8959 27212 8968
rect 27160 8925 27169 8959
rect 27169 8925 27203 8959
rect 27203 8925 27212 8959
rect 27160 8916 27212 8925
rect 25320 8848 25372 8900
rect 25872 8780 25924 8832
rect 27620 8916 27672 8968
rect 27620 8780 27672 8832
rect 10425 8678 10477 8730
rect 10489 8678 10541 8730
rect 10553 8678 10605 8730
rect 10617 8678 10669 8730
rect 10681 8678 10733 8730
rect 19901 8678 19953 8730
rect 19965 8678 20017 8730
rect 20029 8678 20081 8730
rect 20093 8678 20145 8730
rect 20157 8678 20209 8730
rect 1952 8576 2004 8628
rect 2228 8619 2280 8628
rect 2228 8585 2237 8619
rect 2237 8585 2271 8619
rect 2271 8585 2280 8619
rect 2228 8576 2280 8585
rect 2780 8576 2832 8628
rect 5264 8576 5316 8628
rect 3424 8508 3476 8560
rect 4252 8508 4304 8560
rect 5540 8508 5592 8560
rect 6092 8508 6144 8560
rect 9588 8576 9640 8628
rect 3608 8440 3660 8492
rect 4160 8483 4212 8492
rect 2412 8415 2464 8424
rect 2412 8381 2421 8415
rect 2421 8381 2455 8415
rect 2455 8381 2464 8415
rect 2412 8372 2464 8381
rect 3240 8372 3292 8424
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4488 8483
rect 4436 8440 4488 8449
rect 6552 8508 6604 8560
rect 8300 8508 8352 8560
rect 6644 8483 6696 8492
rect 6644 8449 6678 8483
rect 6678 8449 6696 8483
rect 5264 8372 5316 8424
rect 5448 8415 5500 8424
rect 5448 8381 5457 8415
rect 5457 8381 5491 8415
rect 5491 8381 5500 8415
rect 5448 8372 5500 8381
rect 6644 8440 6696 8449
rect 4896 8304 4948 8356
rect 4620 8236 4672 8288
rect 5080 8236 5132 8288
rect 6092 8372 6144 8424
rect 7840 8304 7892 8356
rect 11060 8576 11112 8628
rect 12072 8619 12124 8628
rect 12072 8585 12081 8619
rect 12081 8585 12115 8619
rect 12115 8585 12124 8619
rect 12072 8576 12124 8585
rect 15752 8576 15804 8628
rect 16212 8619 16264 8628
rect 16212 8585 16221 8619
rect 16221 8585 16255 8619
rect 16255 8585 16264 8619
rect 16212 8576 16264 8585
rect 10048 8508 10100 8560
rect 9956 8440 10008 8492
rect 11704 8508 11756 8560
rect 10048 8415 10100 8424
rect 10048 8381 10057 8415
rect 10057 8381 10091 8415
rect 10091 8381 10100 8415
rect 10048 8372 10100 8381
rect 10324 8372 10376 8424
rect 9772 8304 9824 8356
rect 10876 8483 10928 8492
rect 10876 8449 10885 8483
rect 10885 8449 10919 8483
rect 10919 8449 10928 8483
rect 10876 8440 10928 8449
rect 11060 8483 11112 8492
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 12164 8440 12216 8492
rect 15936 8508 15988 8560
rect 17500 8551 17552 8560
rect 11336 8304 11388 8356
rect 12716 8440 12768 8492
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 17132 8466 17184 8518
rect 17500 8517 17509 8551
rect 17509 8517 17543 8551
rect 17543 8517 17552 8551
rect 17500 8508 17552 8517
rect 17776 8576 17828 8628
rect 18144 8576 18196 8628
rect 19340 8576 19392 8628
rect 20352 8619 20404 8628
rect 20352 8585 20361 8619
rect 20361 8585 20395 8619
rect 20395 8585 20404 8619
rect 20352 8576 20404 8585
rect 20536 8619 20588 8628
rect 20536 8585 20545 8619
rect 20545 8585 20579 8619
rect 20579 8585 20588 8619
rect 20536 8576 20588 8585
rect 22376 8576 22428 8628
rect 25320 8619 25372 8628
rect 15752 8415 15804 8424
rect 15752 8381 15761 8415
rect 15761 8381 15795 8415
rect 15795 8381 15804 8415
rect 15752 8372 15804 8381
rect 16396 8372 16448 8424
rect 16028 8304 16080 8356
rect 6736 8236 6788 8288
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 16488 8304 16540 8356
rect 16764 8236 16816 8288
rect 17132 8236 17184 8288
rect 18236 8440 18288 8492
rect 19248 8440 19300 8492
rect 17776 8372 17828 8424
rect 19708 8440 19760 8492
rect 20260 8440 20312 8492
rect 20812 8483 20864 8492
rect 20812 8449 20821 8483
rect 20821 8449 20855 8483
rect 20855 8449 20864 8483
rect 20812 8440 20864 8449
rect 21548 8440 21600 8492
rect 22560 8440 22612 8492
rect 19616 8415 19668 8424
rect 19616 8381 19625 8415
rect 19625 8381 19659 8415
rect 19659 8381 19668 8415
rect 22928 8440 22980 8492
rect 24952 8508 25004 8560
rect 25320 8585 25329 8619
rect 25329 8585 25363 8619
rect 25363 8585 25372 8619
rect 25320 8576 25372 8585
rect 26148 8576 26200 8628
rect 25780 8551 25832 8560
rect 23388 8440 23440 8492
rect 19616 8372 19668 8381
rect 18604 8304 18656 8356
rect 23112 8304 23164 8356
rect 25228 8304 25280 8356
rect 25780 8517 25789 8551
rect 25789 8517 25823 8551
rect 25823 8517 25832 8551
rect 25780 8508 25832 8517
rect 27896 8483 27948 8492
rect 27896 8449 27905 8483
rect 27905 8449 27939 8483
rect 27939 8449 27948 8483
rect 27896 8440 27948 8449
rect 28080 8483 28132 8492
rect 28080 8449 28089 8483
rect 28089 8449 28123 8483
rect 28123 8449 28132 8483
rect 28080 8440 28132 8449
rect 25872 8415 25924 8424
rect 25872 8381 25881 8415
rect 25881 8381 25915 8415
rect 25915 8381 25924 8415
rect 25872 8372 25924 8381
rect 28540 8372 28592 8424
rect 26516 8304 26568 8356
rect 18052 8236 18104 8288
rect 21088 8236 21140 8288
rect 21272 8236 21324 8288
rect 22836 8236 22888 8288
rect 28448 8279 28500 8288
rect 28448 8245 28457 8279
rect 28457 8245 28491 8279
rect 28491 8245 28500 8279
rect 28448 8236 28500 8245
rect 29092 8236 29144 8288
rect 5688 8134 5740 8186
rect 5752 8134 5804 8186
rect 5816 8134 5868 8186
rect 5880 8134 5932 8186
rect 5944 8134 5996 8186
rect 15163 8134 15215 8186
rect 15227 8134 15279 8186
rect 15291 8134 15343 8186
rect 15355 8134 15407 8186
rect 15419 8134 15471 8186
rect 24639 8134 24691 8186
rect 24703 8134 24755 8186
rect 24767 8134 24819 8186
rect 24831 8134 24883 8186
rect 24895 8134 24947 8186
rect 2780 8032 2832 8084
rect 4344 8032 4396 8084
rect 5448 8032 5500 8084
rect 6644 8032 6696 8084
rect 9956 8032 10008 8084
rect 17592 8075 17644 8084
rect 17592 8041 17601 8075
rect 17601 8041 17635 8075
rect 17635 8041 17644 8075
rect 17592 8032 17644 8041
rect 21824 8075 21876 8084
rect 21824 8041 21833 8075
rect 21833 8041 21867 8075
rect 21867 8041 21876 8075
rect 21824 8032 21876 8041
rect 22836 8032 22888 8084
rect 23664 8032 23716 8084
rect 4068 7964 4120 8016
rect 8576 7964 8628 8016
rect 2136 7896 2188 7948
rect 5540 7939 5592 7948
rect 5540 7905 5549 7939
rect 5549 7905 5583 7939
rect 5583 7905 5592 7939
rect 5540 7896 5592 7905
rect 6092 7896 6144 7948
rect 7196 7896 7248 7948
rect 7656 7896 7708 7948
rect 17408 7896 17460 7948
rect 21272 7896 21324 7948
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4620 7828 4672 7880
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5316 7871
rect 5264 7828 5316 7837
rect 6920 7828 6972 7880
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 10048 7828 10100 7880
rect 11336 7871 11388 7880
rect 11336 7837 11354 7871
rect 11354 7837 11388 7871
rect 11336 7828 11388 7837
rect 11520 7828 11572 7880
rect 17500 7828 17552 7880
rect 19064 7871 19116 7880
rect 19064 7837 19073 7871
rect 19073 7837 19107 7871
rect 19107 7837 19116 7871
rect 19064 7828 19116 7837
rect 21364 7828 21416 7880
rect 22744 7828 22796 7880
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 26884 7964 26936 8016
rect 25228 7896 25280 7948
rect 26700 7896 26752 7948
rect 27436 7896 27488 7948
rect 28448 7939 28500 7948
rect 28448 7905 28457 7939
rect 28457 7905 28491 7939
rect 28491 7905 28500 7939
rect 28448 7896 28500 7905
rect 28540 7939 28592 7948
rect 28540 7905 28549 7939
rect 28549 7905 28583 7939
rect 28583 7905 28592 7939
rect 28540 7896 28592 7905
rect 25136 7871 25188 7880
rect 25136 7837 25145 7871
rect 25145 7837 25179 7871
rect 25179 7837 25188 7871
rect 25136 7828 25188 7837
rect 26240 7871 26292 7880
rect 26240 7837 26249 7871
rect 26249 7837 26283 7871
rect 26283 7837 26292 7871
rect 26792 7871 26844 7880
rect 26240 7828 26292 7837
rect 26792 7837 26801 7871
rect 26801 7837 26835 7871
rect 26835 7837 26844 7871
rect 26792 7828 26844 7837
rect 26884 7828 26936 7880
rect 27620 7828 27672 7880
rect 27896 7828 27948 7880
rect 28080 7828 28132 7880
rect 29000 7871 29052 7880
rect 29000 7837 29009 7871
rect 29009 7837 29043 7871
rect 29043 7837 29052 7871
rect 29000 7828 29052 7837
rect 4344 7803 4396 7812
rect 4344 7769 4353 7803
rect 4353 7769 4387 7803
rect 4387 7769 4396 7803
rect 4344 7760 4396 7769
rect 4896 7760 4948 7812
rect 7104 7803 7156 7812
rect 7104 7769 7113 7803
rect 7113 7769 7147 7803
rect 7147 7769 7156 7803
rect 7104 7760 7156 7769
rect 3332 7692 3384 7744
rect 21180 7760 21232 7812
rect 27528 7803 27580 7812
rect 9772 7692 9824 7744
rect 11060 7692 11112 7744
rect 18236 7692 18288 7744
rect 18328 7692 18380 7744
rect 20812 7692 20864 7744
rect 27528 7769 27537 7803
rect 27537 7769 27571 7803
rect 27571 7769 27580 7803
rect 27528 7760 27580 7769
rect 23296 7735 23348 7744
rect 23296 7701 23305 7735
rect 23305 7701 23339 7735
rect 23339 7701 23348 7735
rect 23296 7692 23348 7701
rect 23388 7692 23440 7744
rect 27988 7735 28040 7744
rect 27988 7701 27997 7735
rect 27997 7701 28031 7735
rect 28031 7701 28040 7735
rect 27988 7692 28040 7701
rect 10425 7590 10477 7642
rect 10489 7590 10541 7642
rect 10553 7590 10605 7642
rect 10617 7590 10669 7642
rect 10681 7590 10733 7642
rect 19901 7590 19953 7642
rect 19965 7590 20017 7642
rect 20029 7590 20081 7642
rect 20093 7590 20145 7642
rect 20157 7590 20209 7642
rect 2136 7420 2188 7472
rect 2780 7463 2832 7472
rect 2780 7429 2789 7463
rect 2789 7429 2823 7463
rect 2823 7429 2832 7463
rect 6920 7463 6972 7472
rect 2780 7420 2832 7429
rect 6920 7429 6929 7463
rect 6929 7429 6963 7463
rect 6963 7429 6972 7463
rect 6920 7420 6972 7429
rect 3332 7395 3384 7404
rect 2412 7284 2464 7336
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 7748 7352 7800 7404
rect 8300 7352 8352 7404
rect 8760 7352 8812 7404
rect 15844 7488 15896 7540
rect 17500 7488 17552 7540
rect 18328 7531 18380 7540
rect 18328 7497 18337 7531
rect 18337 7497 18371 7531
rect 18371 7497 18380 7531
rect 18328 7488 18380 7497
rect 19524 7488 19576 7540
rect 20260 7488 20312 7540
rect 22744 7531 22796 7540
rect 15936 7420 15988 7472
rect 18236 7420 18288 7472
rect 16028 7395 16080 7404
rect 2136 7216 2188 7268
rect 15660 7327 15712 7336
rect 15660 7293 15669 7327
rect 15669 7293 15703 7327
rect 15703 7293 15712 7327
rect 16028 7361 16037 7395
rect 16037 7361 16071 7395
rect 16071 7361 16080 7395
rect 16028 7352 16080 7361
rect 16672 7352 16724 7404
rect 15660 7284 15712 7293
rect 15936 7284 15988 7336
rect 15752 7216 15804 7268
rect 16580 7216 16632 7268
rect 17500 7352 17552 7404
rect 18788 7395 18840 7404
rect 18788 7361 18797 7395
rect 18797 7361 18831 7395
rect 18831 7361 18840 7395
rect 18788 7352 18840 7361
rect 19524 7352 19576 7404
rect 20812 7420 20864 7472
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 20444 7395 20496 7404
rect 17316 7284 17368 7336
rect 18144 7284 18196 7336
rect 18328 7216 18380 7268
rect 19708 7284 19760 7336
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 22744 7497 22753 7531
rect 22753 7497 22787 7531
rect 22787 7497 22796 7531
rect 22744 7488 22796 7497
rect 23848 7488 23900 7540
rect 25228 7488 25280 7540
rect 27252 7531 27304 7540
rect 21364 7395 21416 7404
rect 21364 7361 21373 7395
rect 21373 7361 21407 7395
rect 21407 7361 21416 7395
rect 21364 7352 21416 7361
rect 21548 7395 21600 7404
rect 21548 7361 21557 7395
rect 21557 7361 21591 7395
rect 21591 7361 21600 7395
rect 21548 7352 21600 7361
rect 23388 7420 23440 7472
rect 22928 7395 22980 7404
rect 22928 7361 22937 7395
rect 22937 7361 22971 7395
rect 22971 7361 22980 7395
rect 22928 7352 22980 7361
rect 23020 7352 23072 7404
rect 25136 7420 25188 7472
rect 27252 7497 27261 7531
rect 27261 7497 27295 7531
rect 27295 7497 27304 7531
rect 27252 7488 27304 7497
rect 29000 7488 29052 7540
rect 26792 7420 26844 7472
rect 21088 7327 21140 7336
rect 19432 7259 19484 7268
rect 19432 7225 19441 7259
rect 19441 7225 19475 7259
rect 19475 7225 19484 7259
rect 19432 7216 19484 7225
rect 21088 7293 21097 7327
rect 21097 7293 21131 7327
rect 21131 7293 21140 7327
rect 21088 7284 21140 7293
rect 22836 7284 22888 7336
rect 21180 7259 21232 7268
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 2228 7148 2280 7200
rect 7104 7191 7156 7200
rect 7104 7157 7113 7191
rect 7113 7157 7147 7191
rect 7147 7157 7156 7191
rect 7104 7148 7156 7157
rect 9588 7191 9640 7200
rect 9588 7157 9597 7191
rect 9597 7157 9631 7191
rect 9631 7157 9640 7191
rect 9588 7148 9640 7157
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 16212 7148 16264 7157
rect 16764 7148 16816 7200
rect 17408 7148 17460 7200
rect 17684 7148 17736 7200
rect 21180 7225 21189 7259
rect 21189 7225 21223 7259
rect 21223 7225 21232 7259
rect 21180 7216 21232 7225
rect 25136 7327 25188 7336
rect 25136 7293 25145 7327
rect 25145 7293 25179 7327
rect 25179 7293 25188 7327
rect 25136 7284 25188 7293
rect 25228 7216 25280 7268
rect 26240 7352 26292 7404
rect 27436 7420 27488 7472
rect 27344 7352 27396 7404
rect 27160 7284 27212 7336
rect 27436 7284 27488 7336
rect 26332 7216 26384 7268
rect 27528 7216 27580 7268
rect 27896 7327 27948 7336
rect 27896 7293 27905 7327
rect 27905 7293 27939 7327
rect 27939 7293 27948 7327
rect 27896 7284 27948 7293
rect 21916 7148 21968 7200
rect 27620 7148 27672 7200
rect 28540 7148 28592 7200
rect 5688 7046 5740 7098
rect 5752 7046 5804 7098
rect 5816 7046 5868 7098
rect 5880 7046 5932 7098
rect 5944 7046 5996 7098
rect 15163 7046 15215 7098
rect 15227 7046 15279 7098
rect 15291 7046 15343 7098
rect 15355 7046 15407 7098
rect 15419 7046 15471 7098
rect 24639 7046 24691 7098
rect 24703 7046 24755 7098
rect 24767 7046 24819 7098
rect 24831 7046 24883 7098
rect 24895 7046 24947 7098
rect 2136 6944 2188 6996
rect 3792 6987 3844 6996
rect 3792 6953 3801 6987
rect 3801 6953 3835 6987
rect 3835 6953 3844 6987
rect 3792 6944 3844 6953
rect 6552 6944 6604 6996
rect 6920 6987 6972 6996
rect 6920 6953 6929 6987
rect 6929 6953 6963 6987
rect 6963 6953 6972 6987
rect 6920 6944 6972 6953
rect 7196 6944 7248 6996
rect 8760 6987 8812 6996
rect 8760 6953 8769 6987
rect 8769 6953 8803 6987
rect 8803 6953 8812 6987
rect 8760 6944 8812 6953
rect 15752 6987 15804 6996
rect 15752 6953 15761 6987
rect 15761 6953 15795 6987
rect 15795 6953 15804 6987
rect 15752 6944 15804 6953
rect 17500 6944 17552 6996
rect 18788 6944 18840 6996
rect 2136 6808 2188 6860
rect 2412 6808 2464 6860
rect 4160 6808 4212 6860
rect 6736 6876 6788 6928
rect 10232 6876 10284 6928
rect 17408 6876 17460 6928
rect 19708 6944 19760 6996
rect 19800 6944 19852 6996
rect 21088 6944 21140 6996
rect 23020 6944 23072 6996
rect 25320 6944 25372 6996
rect 19064 6919 19116 6928
rect 19064 6885 19073 6919
rect 19073 6885 19107 6919
rect 19107 6885 19116 6919
rect 19064 6876 19116 6885
rect 7196 6808 7248 6860
rect 7656 6808 7708 6860
rect 9588 6808 9640 6860
rect 9864 6808 9916 6860
rect 1860 6740 1912 6792
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 6184 6740 6236 6792
rect 7288 6783 7340 6792
rect 1676 6604 1728 6656
rect 2964 6672 3016 6724
rect 7288 6749 7297 6783
rect 7297 6749 7331 6783
rect 7331 6749 7340 6783
rect 7288 6740 7340 6749
rect 7104 6672 7156 6724
rect 8484 6740 8536 6792
rect 3332 6604 3384 6656
rect 6092 6604 6144 6656
rect 6736 6604 6788 6656
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 11428 6740 11480 6792
rect 16212 6740 16264 6792
rect 16580 6808 16632 6860
rect 16672 6808 16724 6860
rect 17316 6808 17368 6860
rect 17224 6740 17276 6792
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 21364 6808 21416 6860
rect 21824 6808 21876 6860
rect 23112 6808 23164 6860
rect 24492 6808 24544 6860
rect 26792 6876 26844 6928
rect 26700 6851 26752 6860
rect 26700 6817 26709 6851
rect 26709 6817 26743 6851
rect 26743 6817 26752 6851
rect 26700 6808 26752 6817
rect 27528 6944 27580 6996
rect 27252 6851 27304 6860
rect 27252 6817 27261 6851
rect 27261 6817 27295 6851
rect 27295 6817 27304 6851
rect 27252 6808 27304 6817
rect 27712 6851 27764 6860
rect 27712 6817 27721 6851
rect 27721 6817 27755 6851
rect 27755 6817 27764 6851
rect 27712 6808 27764 6817
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 21272 6783 21324 6792
rect 20904 6740 20956 6749
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 21548 6740 21600 6792
rect 22100 6740 22152 6792
rect 22468 6783 22520 6792
rect 22468 6749 22477 6783
rect 22477 6749 22511 6783
rect 22511 6749 22520 6783
rect 22468 6740 22520 6749
rect 23388 6740 23440 6792
rect 25228 6740 25280 6792
rect 26332 6783 26384 6792
rect 26332 6749 26341 6783
rect 26341 6749 26375 6783
rect 26375 6749 26384 6783
rect 26332 6740 26384 6749
rect 26884 6783 26936 6792
rect 26884 6749 26893 6783
rect 26893 6749 26927 6783
rect 26927 6749 26936 6783
rect 26884 6740 26936 6749
rect 27344 6740 27396 6792
rect 27988 6783 28040 6792
rect 27988 6749 28022 6783
rect 28022 6749 28040 6783
rect 27988 6740 28040 6749
rect 16028 6672 16080 6724
rect 10232 6604 10284 6656
rect 10324 6604 10376 6656
rect 16396 6672 16448 6724
rect 16764 6715 16816 6724
rect 16764 6681 16773 6715
rect 16773 6681 16807 6715
rect 16807 6681 16816 6715
rect 18696 6715 18748 6724
rect 16764 6672 16816 6681
rect 18696 6681 18705 6715
rect 18705 6681 18739 6715
rect 18739 6681 18748 6715
rect 18696 6672 18748 6681
rect 17776 6604 17828 6656
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 24400 6672 24452 6724
rect 23296 6604 23348 6656
rect 26148 6647 26200 6656
rect 26148 6613 26157 6647
rect 26157 6613 26191 6647
rect 26191 6613 26200 6647
rect 26148 6604 26200 6613
rect 27160 6647 27212 6656
rect 27160 6613 27169 6647
rect 27169 6613 27203 6647
rect 27203 6613 27212 6647
rect 27160 6604 27212 6613
rect 10425 6502 10477 6554
rect 10489 6502 10541 6554
rect 10553 6502 10605 6554
rect 10617 6502 10669 6554
rect 10681 6502 10733 6554
rect 19901 6502 19953 6554
rect 19965 6502 20017 6554
rect 20029 6502 20081 6554
rect 20093 6502 20145 6554
rect 20157 6502 20209 6554
rect 2780 6400 2832 6452
rect 2964 6375 3016 6384
rect 2964 6341 2973 6375
rect 2973 6341 3007 6375
rect 3007 6341 3016 6375
rect 2964 6332 3016 6341
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 4344 6400 4396 6452
rect 5908 6400 5960 6452
rect 7288 6400 7340 6452
rect 8300 6443 8352 6452
rect 8300 6409 8309 6443
rect 8309 6409 8343 6443
rect 8343 6409 8352 6443
rect 8300 6400 8352 6409
rect 18696 6400 18748 6452
rect 21732 6400 21784 6452
rect 25412 6400 25464 6452
rect 26884 6400 26936 6452
rect 6552 6375 6604 6384
rect 6552 6341 6561 6375
rect 6561 6341 6595 6375
rect 6595 6341 6604 6375
rect 6552 6332 6604 6341
rect 6920 6332 6972 6384
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 5356 6264 5408 6316
rect 6184 6264 6236 6316
rect 17500 6332 17552 6384
rect 18788 6332 18840 6384
rect 25136 6332 25188 6384
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 7564 6264 7616 6316
rect 8484 6264 8536 6316
rect 11060 6307 11112 6316
rect 11060 6273 11078 6307
rect 11078 6273 11112 6307
rect 11060 6264 11112 6273
rect 11520 6264 11572 6316
rect 12900 6264 12952 6316
rect 16396 6264 16448 6316
rect 17776 6307 17828 6316
rect 17776 6273 17785 6307
rect 17785 6273 17819 6307
rect 17819 6273 17828 6307
rect 17776 6264 17828 6273
rect 19524 6264 19576 6316
rect 21272 6264 21324 6316
rect 23572 6307 23624 6316
rect 23572 6273 23581 6307
rect 23581 6273 23615 6307
rect 23615 6273 23624 6307
rect 23572 6264 23624 6273
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 4160 6196 4212 6248
rect 7288 6239 7340 6248
rect 3792 6060 3844 6112
rect 7288 6205 7297 6239
rect 7297 6205 7331 6239
rect 7331 6205 7340 6239
rect 7288 6196 7340 6205
rect 24400 6264 24452 6316
rect 25872 6332 25924 6384
rect 25964 6264 26016 6316
rect 27160 6307 27212 6316
rect 27160 6273 27169 6307
rect 27169 6273 27203 6307
rect 27203 6273 27212 6307
rect 27160 6264 27212 6273
rect 25044 6196 25096 6248
rect 25320 6239 25372 6248
rect 25320 6205 25329 6239
rect 25329 6205 25363 6239
rect 25363 6205 25372 6239
rect 25320 6196 25372 6205
rect 6368 6171 6420 6180
rect 6368 6137 6377 6171
rect 6377 6137 6411 6171
rect 6411 6137 6420 6171
rect 6368 6128 6420 6137
rect 8392 6128 8444 6180
rect 23480 6171 23532 6180
rect 23480 6137 23489 6171
rect 23489 6137 23523 6171
rect 23523 6137 23532 6171
rect 23480 6128 23532 6137
rect 26424 6128 26476 6180
rect 6920 6060 6972 6112
rect 9956 6103 10008 6112
rect 9956 6069 9965 6103
rect 9965 6069 9999 6103
rect 9999 6069 10008 6103
rect 9956 6060 10008 6069
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 18696 6060 18748 6112
rect 22008 6103 22060 6112
rect 22008 6069 22017 6103
rect 22017 6069 22051 6103
rect 22051 6069 22060 6103
rect 22008 6060 22060 6069
rect 22468 6060 22520 6112
rect 5688 5958 5740 6010
rect 5752 5958 5804 6010
rect 5816 5958 5868 6010
rect 5880 5958 5932 6010
rect 5944 5958 5996 6010
rect 15163 5958 15215 6010
rect 15227 5958 15279 6010
rect 15291 5958 15343 6010
rect 15355 5958 15407 6010
rect 15419 5958 15471 6010
rect 24639 5958 24691 6010
rect 24703 5958 24755 6010
rect 24767 5958 24819 6010
rect 24831 5958 24883 6010
rect 24895 5958 24947 6010
rect 3332 5899 3384 5908
rect 3332 5865 3341 5899
rect 3341 5865 3375 5899
rect 3375 5865 3384 5899
rect 3332 5856 3384 5865
rect 3976 5856 4028 5908
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 4068 5788 4120 5840
rect 9864 5856 9916 5908
rect 10324 5856 10376 5908
rect 11060 5856 11112 5908
rect 11428 5899 11480 5908
rect 11428 5865 11437 5899
rect 11437 5865 11471 5899
rect 11471 5865 11480 5899
rect 11428 5856 11480 5865
rect 15844 5856 15896 5908
rect 3884 5720 3936 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 1676 5695 1728 5704
rect 1676 5661 1710 5695
rect 1710 5661 1728 5695
rect 3424 5695 3476 5704
rect 1676 5652 1728 5661
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4528 5720 4580 5772
rect 6092 5788 6144 5840
rect 20628 5856 20680 5908
rect 23112 5856 23164 5908
rect 23388 5856 23440 5908
rect 23572 5856 23624 5908
rect 7656 5720 7708 5772
rect 8944 5720 8996 5772
rect 10324 5763 10376 5772
rect 10324 5729 10333 5763
rect 10333 5729 10367 5763
rect 10367 5729 10376 5763
rect 10324 5720 10376 5729
rect 15568 5763 15620 5772
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 7564 5652 7616 5704
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 10876 5652 10928 5704
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 4344 5584 4396 5636
rect 7196 5584 7248 5636
rect 8852 5584 8904 5636
rect 10232 5584 10284 5636
rect 15660 5652 15712 5704
rect 15936 5652 15988 5704
rect 16764 5720 16816 5772
rect 16212 5584 16264 5636
rect 14924 5559 14976 5568
rect 14924 5525 14933 5559
rect 14933 5525 14967 5559
rect 14967 5525 14976 5559
rect 14924 5516 14976 5525
rect 16580 5652 16632 5704
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 19708 5831 19760 5840
rect 19708 5797 19717 5831
rect 19717 5797 19751 5831
rect 19751 5797 19760 5831
rect 19708 5788 19760 5797
rect 19892 5788 19944 5840
rect 20352 5788 20404 5840
rect 17776 5763 17828 5772
rect 17776 5729 17785 5763
rect 17785 5729 17819 5763
rect 17819 5729 17828 5763
rect 17776 5720 17828 5729
rect 18328 5720 18380 5772
rect 19340 5763 19392 5772
rect 16764 5584 16816 5636
rect 18236 5652 18288 5704
rect 18696 5695 18748 5704
rect 18696 5661 18705 5695
rect 18705 5661 18739 5695
rect 18739 5661 18748 5695
rect 18696 5652 18748 5661
rect 19340 5729 19349 5763
rect 19349 5729 19383 5763
rect 19383 5729 19392 5763
rect 19340 5720 19392 5729
rect 20536 5763 20588 5772
rect 19616 5652 19668 5704
rect 17132 5559 17184 5568
rect 17132 5525 17141 5559
rect 17141 5525 17175 5559
rect 17175 5525 17184 5559
rect 17132 5516 17184 5525
rect 18236 5516 18288 5568
rect 18788 5559 18840 5568
rect 18788 5525 18797 5559
rect 18797 5525 18831 5559
rect 18831 5525 18840 5559
rect 18788 5516 18840 5525
rect 19708 5584 19760 5636
rect 20536 5729 20545 5763
rect 20545 5729 20579 5763
rect 20579 5729 20588 5763
rect 20536 5720 20588 5729
rect 19984 5652 20036 5704
rect 20628 5652 20680 5704
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 20904 5652 20956 5661
rect 19800 5516 19852 5568
rect 20812 5584 20864 5636
rect 21180 5652 21232 5704
rect 21548 5652 21600 5704
rect 22100 5652 22152 5704
rect 23204 5652 23256 5704
rect 24400 5856 24452 5908
rect 25964 5899 26016 5908
rect 20444 5516 20496 5568
rect 22836 5584 22888 5636
rect 22928 5584 22980 5636
rect 24860 5652 24912 5704
rect 25964 5865 25973 5899
rect 25973 5865 26007 5899
rect 26007 5865 26016 5899
rect 25964 5856 26016 5865
rect 26424 5763 26476 5772
rect 26424 5729 26433 5763
rect 26433 5729 26467 5763
rect 26467 5729 26476 5763
rect 26424 5720 26476 5729
rect 27528 5720 27580 5772
rect 27160 5652 27212 5704
rect 21088 5559 21140 5568
rect 21088 5525 21097 5559
rect 21097 5525 21131 5559
rect 21131 5525 21140 5559
rect 21088 5516 21140 5525
rect 21364 5516 21416 5568
rect 21916 5516 21968 5568
rect 22376 5559 22428 5568
rect 22376 5525 22385 5559
rect 22385 5525 22419 5559
rect 22419 5525 22428 5559
rect 22376 5516 22428 5525
rect 24492 5559 24544 5568
rect 24492 5525 24501 5559
rect 24501 5525 24535 5559
rect 24535 5525 24544 5559
rect 24492 5516 24544 5525
rect 24768 5516 24820 5568
rect 10425 5414 10477 5466
rect 10489 5414 10541 5466
rect 10553 5414 10605 5466
rect 10617 5414 10669 5466
rect 10681 5414 10733 5466
rect 19901 5414 19953 5466
rect 19965 5414 20017 5466
rect 20029 5414 20081 5466
rect 20093 5414 20145 5466
rect 20157 5414 20209 5466
rect 3424 5312 3476 5364
rect 2228 5287 2280 5296
rect 2228 5253 2262 5287
rect 2262 5253 2280 5287
rect 2228 5244 2280 5253
rect 6368 5287 6420 5296
rect 6368 5253 6377 5287
rect 6377 5253 6411 5287
rect 6411 5253 6420 5287
rect 6368 5244 6420 5253
rect 8852 5355 8904 5364
rect 8852 5321 8861 5355
rect 8861 5321 8895 5355
rect 8895 5321 8904 5355
rect 8852 5312 8904 5321
rect 9220 5312 9272 5364
rect 10232 5355 10284 5364
rect 1400 5176 1452 5228
rect 4068 5176 4120 5228
rect 4436 5176 4488 5228
rect 4988 5219 5040 5228
rect 3792 4972 3844 5024
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 4988 5176 5040 5185
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 8208 5176 8260 5228
rect 9496 5176 9548 5228
rect 10232 5321 10241 5355
rect 10241 5321 10275 5355
rect 10275 5321 10284 5355
rect 10232 5312 10284 5321
rect 16120 5312 16172 5364
rect 16580 5312 16632 5364
rect 17132 5355 17184 5364
rect 17132 5321 17141 5355
rect 17141 5321 17175 5355
rect 17175 5321 17184 5355
rect 17132 5312 17184 5321
rect 17776 5312 17828 5364
rect 19248 5312 19300 5364
rect 20536 5312 20588 5364
rect 20904 5312 20956 5364
rect 22376 5312 22428 5364
rect 22836 5312 22888 5364
rect 23480 5355 23532 5364
rect 23480 5321 23489 5355
rect 23489 5321 23523 5355
rect 23523 5321 23532 5355
rect 23480 5312 23532 5321
rect 8392 5108 8444 5160
rect 8668 5108 8720 5160
rect 8944 5151 8996 5160
rect 8944 5117 8953 5151
rect 8953 5117 8987 5151
rect 8987 5117 8996 5151
rect 8944 5108 8996 5117
rect 10140 5176 10192 5228
rect 10876 5219 10928 5228
rect 10876 5185 10885 5219
rect 10885 5185 10919 5219
rect 10919 5185 10928 5219
rect 10876 5176 10928 5185
rect 11060 5219 11112 5228
rect 11060 5185 11069 5219
rect 11069 5185 11103 5219
rect 11103 5185 11112 5219
rect 11060 5176 11112 5185
rect 16212 5219 16264 5228
rect 16212 5185 16221 5219
rect 16221 5185 16255 5219
rect 16255 5185 16264 5219
rect 16212 5176 16264 5185
rect 16764 5176 16816 5228
rect 9956 5151 10008 5160
rect 9956 5117 9965 5151
rect 9965 5117 9999 5151
rect 9999 5117 10008 5151
rect 9956 5108 10008 5117
rect 10324 5108 10376 5160
rect 15568 5108 15620 5160
rect 17684 5176 17736 5228
rect 19432 5244 19484 5296
rect 19708 5244 19760 5296
rect 17408 5108 17460 5160
rect 20812 5219 20864 5228
rect 19432 5151 19484 5160
rect 7012 5040 7064 5092
rect 4896 4972 4948 5024
rect 6092 4972 6144 5024
rect 6920 5015 6972 5024
rect 6920 4981 6929 5015
rect 6929 4981 6963 5015
rect 6963 4981 6972 5015
rect 6920 4972 6972 4981
rect 8116 4972 8168 5024
rect 9404 5040 9456 5092
rect 17040 5040 17092 5092
rect 19432 5117 19441 5151
rect 19441 5117 19475 5151
rect 19475 5117 19484 5151
rect 19432 5108 19484 5117
rect 20444 5151 20496 5160
rect 9864 5015 9916 5024
rect 9864 4981 9873 5015
rect 9873 4981 9907 5015
rect 9907 4981 9916 5015
rect 9864 4972 9916 4981
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 15568 4972 15620 5024
rect 17500 4972 17552 5024
rect 18052 4972 18104 5024
rect 19064 4972 19116 5024
rect 20444 5117 20453 5151
rect 20453 5117 20487 5151
rect 20487 5117 20496 5151
rect 20444 5108 20496 5117
rect 20812 5185 20821 5219
rect 20821 5185 20855 5219
rect 20855 5185 20864 5219
rect 20812 5176 20864 5185
rect 21180 5176 21232 5228
rect 22100 5244 22152 5296
rect 24768 5244 24820 5296
rect 21364 5108 21416 5160
rect 23940 5176 23992 5228
rect 28172 5176 28224 5228
rect 21824 5108 21876 5160
rect 23388 5108 23440 5160
rect 22008 5040 22060 5092
rect 23940 5040 23992 5092
rect 25412 5040 25464 5092
rect 19800 5015 19852 5024
rect 19800 4981 19809 5015
rect 19809 4981 19843 5015
rect 19843 4981 19852 5015
rect 19800 4972 19852 4981
rect 25504 4972 25556 5024
rect 5688 4870 5740 4922
rect 5752 4870 5804 4922
rect 5816 4870 5868 4922
rect 5880 4870 5932 4922
rect 5944 4870 5996 4922
rect 15163 4870 15215 4922
rect 15227 4870 15279 4922
rect 15291 4870 15343 4922
rect 15355 4870 15407 4922
rect 15419 4870 15471 4922
rect 24639 4870 24691 4922
rect 24703 4870 24755 4922
rect 24767 4870 24819 4922
rect 24831 4870 24883 4922
rect 24895 4870 24947 4922
rect 4988 4768 5040 4820
rect 7288 4768 7340 4820
rect 8208 4811 8260 4820
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 9864 4768 9916 4820
rect 11060 4811 11112 4820
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 3884 4496 3936 4548
rect 4344 4539 4396 4548
rect 4344 4505 4378 4539
rect 4378 4505 4396 4539
rect 4344 4496 4396 4505
rect 4528 4428 4580 4480
rect 6092 4564 6144 4616
rect 6368 4632 6420 4684
rect 6552 4675 6604 4684
rect 6552 4641 6561 4675
rect 6561 4641 6595 4675
rect 6595 4641 6604 4675
rect 6552 4632 6604 4641
rect 9956 4700 10008 4752
rect 11060 4777 11069 4811
rect 11069 4777 11103 4811
rect 11103 4777 11112 4811
rect 11060 4768 11112 4777
rect 18052 4811 18104 4820
rect 18052 4777 18061 4811
rect 18061 4777 18095 4811
rect 18095 4777 18104 4811
rect 18052 4768 18104 4777
rect 21180 4811 21232 4820
rect 21180 4777 21189 4811
rect 21189 4777 21223 4811
rect 21223 4777 21232 4811
rect 21180 4768 21232 4777
rect 21548 4768 21600 4820
rect 10968 4700 11020 4752
rect 20352 4700 20404 4752
rect 27528 4768 27580 4820
rect 28172 4811 28224 4820
rect 28172 4777 28181 4811
rect 28181 4777 28215 4811
rect 28215 4777 28224 4811
rect 28172 4768 28224 4777
rect 6920 4564 6972 4616
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 9496 4632 9548 4684
rect 12900 4675 12952 4684
rect 12900 4641 12909 4675
rect 12909 4641 12943 4675
rect 12943 4641 12952 4675
rect 12900 4632 12952 4641
rect 22376 4675 22428 4684
rect 22376 4641 22385 4675
rect 22385 4641 22419 4675
rect 22419 4641 22428 4675
rect 22376 4632 22428 4641
rect 23388 4632 23440 4684
rect 25320 4632 25372 4684
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 10048 4564 10100 4616
rect 10876 4607 10928 4616
rect 6460 4539 6512 4548
rect 6460 4505 6469 4539
rect 6469 4505 6503 4539
rect 6503 4505 6512 4539
rect 6460 4496 6512 4505
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 11520 4564 11572 4616
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 18144 4607 18196 4616
rect 18144 4573 18153 4607
rect 18153 4573 18187 4607
rect 18187 4573 18196 4607
rect 18144 4564 18196 4573
rect 21364 4607 21416 4616
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 23940 4607 23992 4616
rect 23940 4573 23949 4607
rect 23949 4573 23983 4607
rect 23983 4573 23992 4607
rect 23940 4564 23992 4573
rect 24492 4564 24544 4616
rect 25412 4607 25464 4616
rect 25412 4573 25421 4607
rect 25421 4573 25455 4607
rect 25455 4573 25464 4607
rect 25412 4564 25464 4573
rect 25504 4607 25556 4616
rect 25504 4573 25513 4607
rect 25513 4573 25547 4607
rect 25547 4573 25556 4607
rect 25504 4564 25556 4573
rect 27252 4564 27304 4616
rect 10784 4496 10836 4548
rect 22652 4496 22704 4548
rect 23756 4539 23808 4548
rect 23756 4505 23765 4539
rect 23765 4505 23799 4539
rect 23799 4505 23808 4539
rect 23756 4496 23808 4505
rect 24584 4539 24636 4548
rect 9404 4428 9456 4480
rect 10232 4471 10284 4480
rect 10232 4437 10241 4471
rect 10241 4437 10275 4471
rect 10275 4437 10284 4471
rect 10232 4428 10284 4437
rect 10968 4428 11020 4480
rect 16028 4471 16080 4480
rect 16028 4437 16037 4471
rect 16037 4437 16071 4471
rect 16071 4437 16080 4471
rect 16028 4428 16080 4437
rect 22284 4471 22336 4480
rect 22284 4437 22293 4471
rect 22293 4437 22327 4471
rect 22327 4437 22336 4471
rect 22284 4428 22336 4437
rect 23848 4428 23900 4480
rect 24584 4505 24593 4539
rect 24593 4505 24627 4539
rect 24627 4505 24636 4539
rect 24584 4496 24636 4505
rect 10425 4326 10477 4378
rect 10489 4326 10541 4378
rect 10553 4326 10605 4378
rect 10617 4326 10669 4378
rect 10681 4326 10733 4378
rect 19901 4326 19953 4378
rect 19965 4326 20017 4378
rect 20029 4326 20081 4378
rect 20093 4326 20145 4378
rect 20157 4326 20209 4378
rect 4436 4267 4488 4276
rect 4436 4233 4445 4267
rect 4445 4233 4479 4267
rect 4479 4233 4488 4267
rect 4436 4224 4488 4233
rect 10876 4224 10928 4276
rect 15936 4224 15988 4276
rect 16764 4267 16816 4276
rect 8116 4156 8168 4208
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 6368 4131 6420 4140
rect 4528 4088 4580 4097
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 7472 4088 7524 4140
rect 4712 4063 4764 4072
rect 4712 4029 4721 4063
rect 4721 4029 4755 4063
rect 4755 4029 4764 4063
rect 4712 4020 4764 4029
rect 9220 4088 9272 4140
rect 10232 4088 10284 4140
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 12900 4088 12952 4140
rect 14924 4088 14976 4140
rect 16764 4233 16773 4267
rect 16773 4233 16807 4267
rect 16807 4233 16816 4267
rect 16764 4224 16816 4233
rect 18144 4224 18196 4276
rect 18788 4224 18840 4276
rect 21364 4224 21416 4276
rect 16672 4156 16724 4208
rect 18052 4156 18104 4208
rect 18512 4156 18564 4208
rect 19800 4156 19852 4208
rect 22100 4156 22152 4208
rect 16304 4088 16356 4140
rect 18328 4088 18380 4140
rect 22376 4156 22428 4208
rect 24584 4224 24636 4276
rect 9588 4020 9640 4072
rect 9956 4020 10008 4072
rect 11060 4063 11112 4072
rect 11060 4029 11069 4063
rect 11069 4029 11103 4063
rect 11103 4029 11112 4063
rect 11060 4020 11112 4029
rect 4344 3952 4396 4004
rect 848 3884 900 3936
rect 11244 3952 11296 4004
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 6920 3884 6972 3936
rect 8116 3884 8168 3936
rect 9680 3884 9732 3936
rect 14648 3884 14700 3936
rect 16948 4020 17000 4072
rect 17224 4063 17276 4072
rect 17224 4029 17233 4063
rect 17233 4029 17267 4063
rect 17267 4029 17276 4063
rect 17224 4020 17276 4029
rect 15936 3952 15988 4004
rect 17776 4020 17828 4072
rect 18144 4063 18196 4072
rect 18144 4029 18153 4063
rect 18153 4029 18187 4063
rect 18187 4029 18196 4063
rect 18144 4020 18196 4029
rect 17868 3952 17920 4004
rect 23756 4156 23808 4208
rect 23204 4131 23256 4140
rect 23204 4097 23213 4131
rect 23213 4097 23247 4131
rect 23247 4097 23256 4131
rect 23204 4088 23256 4097
rect 23480 4131 23532 4140
rect 23480 4097 23514 4131
rect 23514 4097 23532 4131
rect 23480 4088 23532 4097
rect 25504 4088 25556 4140
rect 26148 4088 26200 4140
rect 20812 3995 20864 4004
rect 16672 3884 16724 3936
rect 17776 3884 17828 3936
rect 18144 3884 18196 3936
rect 20812 3961 20821 3995
rect 20821 3961 20855 3995
rect 20855 3961 20864 3995
rect 20812 3952 20864 3961
rect 24400 3952 24452 4004
rect 20536 3884 20588 3936
rect 23940 3884 23992 3936
rect 5688 3782 5740 3834
rect 5752 3782 5804 3834
rect 5816 3782 5868 3834
rect 5880 3782 5932 3834
rect 5944 3782 5996 3834
rect 15163 3782 15215 3834
rect 15227 3782 15279 3834
rect 15291 3782 15343 3834
rect 15355 3782 15407 3834
rect 15419 3782 15471 3834
rect 24639 3782 24691 3834
rect 24703 3782 24755 3834
rect 24767 3782 24819 3834
rect 24831 3782 24883 3834
rect 24895 3782 24947 3834
rect 2504 3680 2556 3732
rect 4252 3680 4304 3732
rect 7840 3680 7892 3732
rect 9588 3680 9640 3732
rect 10968 3680 11020 3732
rect 11152 3680 11204 3732
rect 14648 3680 14700 3732
rect 17776 3723 17828 3732
rect 17776 3689 17785 3723
rect 17785 3689 17819 3723
rect 17819 3689 17828 3723
rect 17776 3680 17828 3689
rect 18880 3723 18932 3732
rect 4896 3544 4948 3596
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 6920 3612 6972 3664
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 5816 3476 5868 3528
rect 6368 3476 6420 3528
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 7012 3476 7064 3528
rect 10784 3612 10836 3664
rect 11244 3612 11296 3664
rect 11428 3612 11480 3664
rect 12716 3612 12768 3664
rect 16672 3612 16724 3664
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 11060 3544 11112 3596
rect 8024 3476 8076 3485
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 3884 3340 3936 3392
rect 5908 3340 5960 3392
rect 6000 3340 6052 3392
rect 6736 3340 6788 3392
rect 8208 3340 8260 3392
rect 8300 3340 8352 3392
rect 9220 3340 9272 3392
rect 9956 3408 10008 3460
rect 15936 3587 15988 3596
rect 15936 3553 15945 3587
rect 15945 3553 15979 3587
rect 15979 3553 15988 3587
rect 15936 3544 15988 3553
rect 16304 3544 16356 3596
rect 11336 3519 11388 3528
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 16028 3476 16080 3528
rect 16764 3476 16816 3528
rect 18880 3689 18889 3723
rect 18889 3689 18923 3723
rect 18923 3689 18932 3723
rect 18880 3680 18932 3689
rect 19432 3680 19484 3732
rect 18972 3612 19024 3664
rect 18788 3544 18840 3596
rect 10140 3340 10192 3392
rect 10784 3383 10836 3392
rect 10784 3349 10793 3383
rect 10793 3349 10827 3383
rect 10827 3349 10836 3383
rect 10784 3340 10836 3349
rect 10968 3340 11020 3392
rect 11980 3340 12032 3392
rect 16396 3340 16448 3392
rect 17040 3408 17092 3460
rect 18604 3476 18656 3528
rect 18696 3519 18748 3528
rect 18696 3485 18705 3519
rect 18705 3485 18739 3519
rect 18739 3485 18748 3519
rect 18696 3476 18748 3485
rect 22100 3680 22152 3732
rect 22284 3680 22336 3732
rect 23480 3723 23532 3732
rect 23480 3689 23489 3723
rect 23489 3689 23523 3723
rect 23523 3689 23532 3723
rect 23480 3680 23532 3689
rect 23388 3612 23440 3664
rect 20536 3587 20588 3596
rect 20536 3553 20545 3587
rect 20545 3553 20579 3587
rect 20579 3553 20588 3587
rect 20536 3544 20588 3553
rect 18052 3340 18104 3392
rect 18512 3408 18564 3460
rect 20260 3408 20312 3460
rect 18696 3340 18748 3392
rect 20444 3340 20496 3392
rect 21088 3476 21140 3528
rect 20628 3408 20680 3460
rect 23940 3587 23992 3596
rect 23940 3553 23949 3587
rect 23949 3553 23983 3587
rect 23983 3553 23992 3587
rect 23940 3544 23992 3553
rect 22376 3519 22428 3528
rect 22376 3485 22385 3519
rect 22385 3485 22419 3519
rect 22419 3485 22428 3519
rect 22376 3476 22428 3485
rect 22652 3519 22704 3528
rect 22652 3485 22661 3519
rect 22661 3485 22695 3519
rect 22695 3485 22704 3519
rect 22652 3476 22704 3485
rect 23848 3519 23900 3528
rect 22008 3340 22060 3392
rect 22192 3408 22244 3460
rect 23848 3485 23857 3519
rect 23857 3485 23891 3519
rect 23891 3485 23900 3519
rect 23848 3476 23900 3485
rect 29828 3476 29880 3528
rect 22744 3340 22796 3392
rect 10425 3238 10477 3290
rect 10489 3238 10541 3290
rect 10553 3238 10605 3290
rect 10617 3238 10669 3290
rect 10681 3238 10733 3290
rect 19901 3238 19953 3290
rect 19965 3238 20017 3290
rect 20029 3238 20081 3290
rect 20093 3238 20145 3290
rect 20157 3238 20209 3290
rect 4620 3136 4672 3188
rect 8024 3136 8076 3188
rect 8208 3136 8260 3188
rect 9772 3136 9824 3188
rect 9956 3179 10008 3188
rect 9956 3145 9965 3179
rect 9965 3145 9999 3179
rect 9999 3145 10008 3179
rect 9956 3136 10008 3145
rect 11888 3136 11940 3188
rect 16212 3136 16264 3188
rect 18236 3136 18288 3188
rect 18788 3136 18840 3188
rect 18880 3136 18932 3188
rect 19800 3136 19852 3188
rect 20260 3136 20312 3188
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 4068 2932 4120 2984
rect 4436 3043 4488 3052
rect 4436 3009 4470 3043
rect 4470 3009 4488 3043
rect 5908 3043 5960 3052
rect 4436 3000 4488 3009
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 8392 3068 8444 3120
rect 6000 3000 6052 3009
rect 6460 3000 6512 3052
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 7656 2932 7708 2984
rect 14464 3068 14516 3120
rect 8852 3043 8904 3052
rect 8852 3009 8886 3043
rect 8886 3009 8904 3043
rect 8852 3000 8904 3009
rect 10784 3000 10836 3052
rect 10140 2932 10192 2984
rect 12440 3000 12492 3052
rect 12900 3000 12952 3052
rect 15016 3043 15068 3052
rect 15016 3009 15025 3043
rect 15025 3009 15059 3043
rect 15059 3009 15068 3043
rect 15016 3000 15068 3009
rect 15568 3000 15620 3052
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17868 3068 17920 3120
rect 17500 3043 17552 3052
rect 17500 3009 17534 3043
rect 17534 3009 17552 3043
rect 17500 3000 17552 3009
rect 5816 2864 5868 2916
rect 7380 2864 7432 2916
rect 4804 2796 4856 2848
rect 6184 2839 6236 2848
rect 6184 2805 6193 2839
rect 6193 2805 6227 2839
rect 6227 2805 6236 2839
rect 6184 2796 6236 2805
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 11060 2864 11112 2916
rect 16948 2932 17000 2984
rect 18236 2932 18288 2984
rect 19708 3068 19760 3120
rect 20444 3111 20496 3120
rect 20444 3077 20453 3111
rect 20453 3077 20487 3111
rect 20487 3077 20496 3111
rect 20444 3068 20496 3077
rect 20812 3111 20864 3120
rect 20812 3077 20821 3111
rect 20821 3077 20855 3111
rect 20855 3077 20864 3111
rect 20812 3068 20864 3077
rect 22652 3136 22704 3188
rect 21824 3111 21876 3120
rect 21824 3077 21833 3111
rect 21833 3077 21867 3111
rect 21867 3077 21876 3111
rect 21824 3068 21876 3077
rect 22008 3111 22060 3120
rect 22008 3077 22017 3111
rect 22017 3077 22051 3111
rect 22051 3077 22060 3111
rect 22008 3068 22060 3077
rect 19064 3043 19116 3052
rect 19064 3009 19098 3043
rect 19098 3009 19116 3043
rect 19064 3000 19116 3009
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 22192 3043 22244 3052
rect 22192 3009 22201 3043
rect 22201 3009 22235 3043
rect 22235 3009 22244 3043
rect 22192 3000 22244 3009
rect 22008 2932 22060 2984
rect 22376 2932 22428 2984
rect 9312 2796 9364 2848
rect 10968 2796 11020 2848
rect 14464 2796 14516 2848
rect 21732 2864 21784 2916
rect 19800 2796 19852 2848
rect 21824 2796 21876 2848
rect 5688 2694 5740 2746
rect 5752 2694 5804 2746
rect 5816 2694 5868 2746
rect 5880 2694 5932 2746
rect 5944 2694 5996 2746
rect 15163 2694 15215 2746
rect 15227 2694 15279 2746
rect 15291 2694 15343 2746
rect 15355 2694 15407 2746
rect 15419 2694 15471 2746
rect 24639 2694 24691 2746
rect 24703 2694 24755 2746
rect 24767 2694 24819 2746
rect 24831 2694 24883 2746
rect 24895 2694 24947 2746
rect 4436 2592 4488 2644
rect 6460 2635 6512 2644
rect 6460 2601 6469 2635
rect 6469 2601 6503 2635
rect 6503 2601 6512 2635
rect 6460 2592 6512 2601
rect 8852 2592 8904 2644
rect 12440 2592 12492 2644
rect 18052 2592 18104 2644
rect 4712 2524 4764 2576
rect 4804 2499 4856 2508
rect 4804 2465 4813 2499
rect 4813 2465 4847 2499
rect 4847 2465 4856 2499
rect 4804 2456 4856 2465
rect 6184 2456 6236 2508
rect 8668 2524 8720 2576
rect 8484 2456 8536 2508
rect 11980 2499 12032 2508
rect 11980 2465 11989 2499
rect 11989 2465 12023 2499
rect 12023 2465 12032 2499
rect 11980 2456 12032 2465
rect 4620 2388 4672 2440
rect 6736 2388 6788 2440
rect 9220 2388 9272 2440
rect 11060 2388 11112 2440
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 3424 2320 3476 2372
rect 9128 2320 9180 2372
rect 10425 2150 10477 2202
rect 10489 2150 10541 2202
rect 10553 2150 10605 2202
rect 10617 2150 10669 2202
rect 10681 2150 10733 2202
rect 19901 2150 19953 2202
rect 19965 2150 20017 2202
rect 20029 2150 20081 2202
rect 20093 2150 20145 2202
rect 20157 2150 20209 2202
rect 3148 1300 3200 1352
rect 9036 1300 9088 1352
rect 16856 1300 16908 1352
rect 27528 1300 27580 1352
<< metal2 >>
rect 570 32056 626 32856
rect 1766 32056 1822 32856
rect 2962 32056 3018 32856
rect 3882 32192 3938 32201
rect 3882 32127 3938 32136
rect 584 28966 612 32056
rect 572 28960 624 28966
rect 572 28902 624 28908
rect 1308 28960 1360 28966
rect 1308 28902 1360 28908
rect 1320 16017 1348 28902
rect 1780 26234 1808 32056
rect 2976 29714 3004 32056
rect 3896 30666 3924 32127
rect 4250 32056 4306 32856
rect 5446 32056 5502 32856
rect 6642 32056 6698 32856
rect 7930 32056 7986 32856
rect 9126 32056 9182 32856
rect 10322 32056 10378 32856
rect 11610 32056 11666 32856
rect 12806 32056 12862 32856
rect 14002 32056 14058 32856
rect 15290 32056 15346 32856
rect 16486 32056 16542 32856
rect 17774 32056 17830 32856
rect 18970 32056 19026 32856
rect 20166 32056 20222 32856
rect 21454 32056 21510 32856
rect 22650 32056 22706 32856
rect 23846 32056 23902 32856
rect 25134 32056 25190 32856
rect 26330 32056 26386 32856
rect 27342 32056 27398 32065
rect 27526 32056 27582 32856
rect 28814 32056 28870 32856
rect 30010 32056 30066 32856
rect 4066 30832 4122 30841
rect 4066 30767 4122 30776
rect 3884 30660 3936 30666
rect 3884 30602 3936 30608
rect 4080 30394 4108 30767
rect 4068 30388 4120 30394
rect 4068 30330 4120 30336
rect 4068 30116 4120 30122
rect 4068 30058 4120 30064
rect 2964 29708 3016 29714
rect 2964 29650 3016 29656
rect 4080 29481 4108 30058
rect 4264 29714 4292 32056
rect 4252 29708 4304 29714
rect 4252 29650 4304 29656
rect 4066 29472 4122 29481
rect 4066 29407 4122 29416
rect 4068 28144 4120 28150
rect 4066 28112 4068 28121
rect 4120 28112 4122 28121
rect 4066 28047 4122 28056
rect 5172 28008 5224 28014
rect 5172 27950 5224 27956
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4080 26761 4108 27270
rect 4160 27056 4212 27062
rect 4160 26998 4212 27004
rect 4066 26752 4122 26761
rect 4066 26687 4122 26696
rect 1504 26206 1808 26234
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1412 23866 1440 24686
rect 1400 23860 1452 23866
rect 1400 23802 1452 23808
rect 1412 23662 1440 23802
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1412 22642 1440 23598
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 22098 1440 22578
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 1504 21418 1532 26206
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 4080 25401 4108 25434
rect 4066 25392 4122 25401
rect 4172 25362 4200 26998
rect 4620 26988 4672 26994
rect 4620 26930 4672 26936
rect 4632 26586 4660 26930
rect 4988 26784 5040 26790
rect 4988 26726 5040 26732
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 5000 26382 5028 26726
rect 5184 26382 5212 27950
rect 5356 27940 5408 27946
rect 5356 27882 5408 27888
rect 5368 26518 5396 27882
rect 5356 26512 5408 26518
rect 5356 26454 5408 26460
rect 4988 26376 5040 26382
rect 4988 26318 5040 26324
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4252 25696 4304 25702
rect 4252 25638 4304 25644
rect 4712 25696 4764 25702
rect 4712 25638 4764 25644
rect 4066 25327 4122 25336
rect 4160 25356 4212 25362
rect 4160 25298 4212 25304
rect 4172 24886 4200 25298
rect 2688 24880 2740 24886
rect 2688 24822 2740 24828
rect 4160 24880 4212 24886
rect 4160 24822 4212 24828
rect 2700 24410 2728 24822
rect 3700 24744 3752 24750
rect 3700 24686 3752 24692
rect 3976 24744 4028 24750
rect 3976 24686 4028 24692
rect 3712 24614 3740 24686
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 2688 24404 2740 24410
rect 2688 24346 2740 24352
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 2332 23118 2360 24142
rect 2872 23792 2924 23798
rect 2872 23734 2924 23740
rect 2884 23322 2912 23734
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3436 23526 3464 23666
rect 3424 23520 3476 23526
rect 3424 23462 3476 23468
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 1676 22568 1728 22574
rect 1676 22510 1728 22516
rect 1688 22234 1716 22510
rect 2240 22234 2268 23054
rect 2332 22574 2360 23054
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 2424 22710 2452 22918
rect 2412 22704 2464 22710
rect 2412 22646 2464 22652
rect 2320 22568 2372 22574
rect 2320 22510 2372 22516
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2332 22030 2360 22510
rect 3056 22432 3108 22438
rect 3056 22374 3108 22380
rect 2320 22024 2372 22030
rect 2320 21966 2372 21972
rect 3068 21894 3096 22374
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 1492 21412 1544 21418
rect 1492 21354 1544 21360
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 19310 1440 20878
rect 3068 20602 3096 21830
rect 3436 21690 3464 23462
rect 3608 23112 3660 23118
rect 3608 23054 3660 23060
rect 3620 21962 3648 23054
rect 3608 21956 3660 21962
rect 3608 21898 3660 21904
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3620 21486 3648 21898
rect 3148 21480 3200 21486
rect 3148 21422 3200 21428
rect 3240 21480 3292 21486
rect 3240 21422 3292 21428
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3056 20596 3108 20602
rect 3056 20538 3108 20544
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 2976 19514 3004 20334
rect 3160 20330 3188 21422
rect 3252 21078 3280 21422
rect 3516 21344 3568 21350
rect 3516 21286 3568 21292
rect 3240 21072 3292 21078
rect 3240 21014 3292 21020
rect 3252 20942 3280 21014
rect 3424 21004 3476 21010
rect 3424 20946 3476 20952
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 3344 20534 3372 20878
rect 3332 20528 3384 20534
rect 3332 20470 3384 20476
rect 3148 20324 3200 20330
rect 3148 20266 3200 20272
rect 3436 20244 3464 20946
rect 3528 20466 3556 21286
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 3620 20602 3648 20878
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3516 20256 3568 20262
rect 3436 20216 3516 20244
rect 3516 20198 3568 20204
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1412 18358 1440 19246
rect 3528 19174 3556 20198
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3528 18970 3556 19110
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3528 18426 3556 18906
rect 3712 18766 3740 24550
rect 3988 23662 4016 24686
rect 4068 24064 4120 24070
rect 4066 24032 4068 24041
rect 4120 24032 4122 24041
rect 4066 23967 4122 23976
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3988 23322 4016 23598
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 3974 22672 4030 22681
rect 3974 22607 4030 22616
rect 3988 22234 4016 22607
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 4160 21956 4212 21962
rect 4160 21898 4212 21904
rect 4172 21690 4200 21898
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 4066 21312 4122 21321
rect 4066 21247 4122 21256
rect 4080 21146 4108 21247
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 4068 20868 4120 20874
rect 4068 20810 4120 20816
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 3896 20330 3924 20742
rect 4080 20602 4108 20810
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 3884 20324 3936 20330
rect 3884 20266 3936 20272
rect 3896 19242 3924 20266
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 3884 19236 3936 19242
rect 3884 19178 3936 19184
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3790 18592 3846 18601
rect 3790 18527 3846 18536
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 1400 18352 1452 18358
rect 1400 18294 1452 18300
rect 1412 17746 1440 18294
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 1412 16658 1440 17682
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 3252 16590 3280 17614
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2332 16182 2360 16458
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2320 16176 2372 16182
rect 2320 16118 2372 16124
rect 2792 16114 2820 16390
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 1306 16008 1362 16017
rect 1306 15943 1362 15952
rect 2044 15360 2096 15366
rect 2044 15302 2096 15308
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 1964 14618 1992 14962
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2056 14414 2084 15302
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2792 13326 2820 15030
rect 2884 13938 2912 16186
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3068 15570 3096 15846
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 3160 15502 3188 15982
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 2976 15162 3004 15438
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 3252 15026 3280 15506
rect 3344 15026 3372 15982
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3148 14884 3200 14890
rect 3148 14826 3200 14832
rect 3160 14414 3188 14826
rect 3252 14618 3280 14962
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3436 14074 3464 17818
rect 3620 17678 3648 18022
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3620 15978 3648 17614
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3712 16182 3740 16526
rect 3700 16176 3752 16182
rect 3804 16153 3832 18527
rect 3896 17882 3924 19178
rect 4080 18766 4108 19314
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4172 18766 4200 19246
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 3976 18692 4028 18698
rect 3976 18634 4028 18640
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3988 17678 4016 18634
rect 4080 17882 4108 18702
rect 4172 18426 4200 18702
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4264 18034 4292 25638
rect 4724 25294 4752 25638
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4816 25226 4844 25842
rect 5184 25770 5212 26318
rect 5368 26042 5396 26454
rect 5460 26042 5488 32056
rect 5688 29948 5996 29968
rect 5688 29946 5694 29948
rect 5750 29946 5774 29948
rect 5830 29946 5854 29948
rect 5910 29946 5934 29948
rect 5990 29946 5996 29948
rect 5750 29894 5752 29946
rect 5932 29894 5934 29946
rect 5688 29892 5694 29894
rect 5750 29892 5774 29894
rect 5830 29892 5854 29894
rect 5910 29892 5934 29894
rect 5990 29892 5996 29894
rect 5688 29872 5996 29892
rect 6656 29714 6684 32056
rect 6644 29708 6696 29714
rect 6644 29650 6696 29656
rect 6368 29640 6420 29646
rect 6368 29582 6420 29588
rect 5688 28860 5996 28880
rect 5688 28858 5694 28860
rect 5750 28858 5774 28860
rect 5830 28858 5854 28860
rect 5910 28858 5934 28860
rect 5990 28858 5996 28860
rect 5750 28806 5752 28858
rect 5932 28806 5934 28858
rect 5688 28804 5694 28806
rect 5750 28804 5774 28806
rect 5830 28804 5854 28806
rect 5910 28804 5934 28806
rect 5990 28804 5996 28806
rect 5688 28784 5996 28804
rect 6380 28082 6408 29582
rect 7564 29028 7616 29034
rect 7564 28970 7616 28976
rect 6460 28960 6512 28966
rect 6460 28902 6512 28908
rect 5540 28076 5592 28082
rect 5540 28018 5592 28024
rect 5724 28076 5776 28082
rect 5724 28018 5776 28024
rect 6368 28076 6420 28082
rect 6368 28018 6420 28024
rect 5552 27674 5580 28018
rect 5736 27946 5764 28018
rect 5724 27940 5776 27946
rect 5724 27882 5776 27888
rect 6276 27872 6328 27878
rect 6276 27814 6328 27820
rect 5688 27772 5996 27792
rect 5688 27770 5694 27772
rect 5750 27770 5774 27772
rect 5830 27770 5854 27772
rect 5910 27770 5934 27772
rect 5990 27770 5996 27772
rect 5750 27718 5752 27770
rect 5932 27718 5934 27770
rect 5688 27716 5694 27718
rect 5750 27716 5774 27718
rect 5830 27716 5854 27718
rect 5910 27716 5934 27718
rect 5990 27716 5996 27718
rect 5688 27696 5996 27716
rect 5540 27668 5592 27674
rect 5540 27610 5592 27616
rect 6092 27124 6144 27130
rect 6092 27066 6144 27072
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 5552 26586 5580 26930
rect 5688 26684 5996 26704
rect 5688 26682 5694 26684
rect 5750 26682 5774 26684
rect 5830 26682 5854 26684
rect 5910 26682 5934 26684
rect 5990 26682 5996 26684
rect 5750 26630 5752 26682
rect 5932 26630 5934 26682
rect 5688 26628 5694 26630
rect 5750 26628 5774 26630
rect 5830 26628 5854 26630
rect 5910 26628 5934 26630
rect 5990 26628 5996 26630
rect 5688 26608 5996 26628
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 6104 26382 6132 27066
rect 6184 26512 6236 26518
rect 6184 26454 6236 26460
rect 5724 26376 5776 26382
rect 5724 26318 5776 26324
rect 6092 26376 6144 26382
rect 6092 26318 6144 26324
rect 5736 26246 5764 26318
rect 5724 26240 5776 26246
rect 5724 26182 5776 26188
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 5448 26036 5500 26042
rect 5448 25978 5500 25984
rect 5736 25906 5764 26182
rect 6196 26058 6224 26454
rect 6288 26246 6316 27814
rect 6380 27062 6408 28018
rect 6472 27674 6500 28902
rect 6460 27668 6512 27674
rect 6460 27610 6512 27616
rect 7472 27532 7524 27538
rect 7472 27474 7524 27480
rect 7104 27396 7156 27402
rect 7104 27338 7156 27344
rect 6736 27328 6788 27334
rect 6736 27270 6788 27276
rect 6368 27056 6420 27062
rect 6368 26998 6420 27004
rect 6380 26518 6408 26998
rect 6748 26994 6776 27270
rect 7116 27130 7144 27338
rect 7104 27124 7156 27130
rect 7104 27066 7156 27072
rect 7484 27062 7512 27474
rect 7472 27056 7524 27062
rect 7472 26998 7524 27004
rect 6736 26988 6788 26994
rect 6736 26930 6788 26936
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 6368 26512 6420 26518
rect 6368 26454 6420 26460
rect 6920 26444 6972 26450
rect 6920 26386 6972 26392
rect 6368 26376 6420 26382
rect 6368 26318 6420 26324
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6736 26376 6788 26382
rect 6736 26318 6788 26324
rect 6276 26240 6328 26246
rect 6276 26182 6328 26188
rect 6196 26030 6316 26058
rect 5724 25900 5776 25906
rect 5724 25842 5776 25848
rect 6092 25832 6144 25838
rect 6092 25774 6144 25780
rect 5172 25764 5224 25770
rect 5172 25706 5224 25712
rect 5184 25430 5212 25706
rect 5688 25596 5996 25616
rect 5688 25594 5694 25596
rect 5750 25594 5774 25596
rect 5830 25594 5854 25596
rect 5910 25594 5934 25596
rect 5990 25594 5996 25596
rect 5750 25542 5752 25594
rect 5932 25542 5934 25594
rect 5688 25540 5694 25542
rect 5750 25540 5774 25542
rect 5830 25540 5854 25542
rect 5910 25540 5934 25542
rect 5990 25540 5996 25542
rect 5688 25520 5996 25540
rect 5172 25424 5224 25430
rect 5172 25366 5224 25372
rect 4804 25220 4856 25226
rect 4804 25162 4856 25168
rect 4620 24880 4672 24886
rect 4620 24822 4672 24828
rect 4632 23866 4660 24822
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4632 23730 4660 23802
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4908 23322 4936 23666
rect 4896 23316 4948 23322
rect 4896 23258 4948 23264
rect 5184 23186 5212 25366
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5552 23254 5580 24754
rect 5688 24508 5996 24528
rect 5688 24506 5694 24508
rect 5750 24506 5774 24508
rect 5830 24506 5854 24508
rect 5910 24506 5934 24508
rect 5990 24506 5996 24508
rect 5750 24454 5752 24506
rect 5932 24454 5934 24506
rect 5688 24452 5694 24454
rect 5750 24452 5774 24454
rect 5830 24452 5854 24454
rect 5910 24452 5934 24454
rect 5990 24452 5996 24454
rect 5688 24432 5996 24452
rect 6104 24410 6132 25774
rect 6092 24404 6144 24410
rect 6144 24364 6224 24392
rect 6092 24346 6144 24352
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 5688 23420 5996 23440
rect 5688 23418 5694 23420
rect 5750 23418 5774 23420
rect 5830 23418 5854 23420
rect 5910 23418 5934 23420
rect 5990 23418 5996 23420
rect 5750 23366 5752 23418
rect 5932 23366 5934 23418
rect 5688 23364 5694 23366
rect 5750 23364 5774 23366
rect 5830 23364 5854 23366
rect 5910 23364 5934 23366
rect 5990 23364 5996 23366
rect 5688 23344 5996 23364
rect 6104 23322 6132 23802
rect 6092 23316 6144 23322
rect 6092 23258 6144 23264
rect 5540 23248 5592 23254
rect 6196 23202 6224 24364
rect 6288 24018 6316 26030
rect 6380 25838 6408 26318
rect 6472 26042 6500 26318
rect 6460 26036 6512 26042
rect 6460 25978 6512 25984
rect 6748 25906 6776 26318
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 6368 25832 6420 25838
rect 6368 25774 6420 25780
rect 6380 24410 6408 25774
rect 6748 25702 6776 25842
rect 6932 25770 6960 26386
rect 7104 25968 7156 25974
rect 7104 25910 7156 25916
rect 6920 25764 6972 25770
rect 6920 25706 6972 25712
rect 6736 25696 6788 25702
rect 6736 25638 6788 25644
rect 6828 25152 6880 25158
rect 6932 25140 6960 25706
rect 6880 25112 6960 25140
rect 6828 25094 6880 25100
rect 6644 24812 6696 24818
rect 6644 24754 6696 24760
rect 6656 24410 6684 24754
rect 6368 24404 6420 24410
rect 6368 24346 6420 24352
rect 6644 24404 6696 24410
rect 6644 24346 6696 24352
rect 6380 24138 6408 24346
rect 6840 24206 6868 25094
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6368 24132 6420 24138
rect 6368 24074 6420 24080
rect 6736 24132 6788 24138
rect 6736 24074 6788 24080
rect 6288 23990 6408 24018
rect 5540 23190 5592 23196
rect 5644 23186 6224 23202
rect 5172 23180 5224 23186
rect 5172 23122 5224 23128
rect 5632 23180 6224 23186
rect 5684 23174 6224 23180
rect 5632 23122 5684 23128
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5092 21690 5120 22510
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5184 21962 5212 22374
rect 5172 21956 5224 21962
rect 5172 21898 5224 21904
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 4528 21616 4580 21622
rect 4528 21558 4580 21564
rect 4540 19514 4568 21558
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 4632 20330 4660 20878
rect 5172 20800 5224 20806
rect 5172 20742 5224 20748
rect 5184 20466 5212 20742
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 4620 20324 4672 20330
rect 4620 20266 4672 20272
rect 4632 19854 4660 20266
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4632 18766 4660 19790
rect 4988 19780 5040 19786
rect 4988 19722 5040 19728
rect 5000 19514 5028 19722
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 5276 19378 5304 20470
rect 5264 19372 5316 19378
rect 5092 19332 5264 19360
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4356 18290 4384 18566
rect 4908 18358 4936 18702
rect 5092 18426 5120 19332
rect 5264 19314 5316 19320
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5276 18426 5304 18634
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 4896 18352 4948 18358
rect 4896 18294 4948 18300
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4712 18284 4764 18290
rect 4712 18226 4764 18232
rect 4172 18006 4292 18034
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 3976 17672 4028 17678
rect 3896 17632 3976 17660
rect 3700 16118 3752 16124
rect 3790 16144 3846 16153
rect 3790 16079 3846 16088
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3896 15638 3924 17632
rect 3976 17614 4028 17620
rect 4066 17232 4122 17241
rect 4172 17218 4200 18006
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4122 17190 4200 17218
rect 4066 17167 4122 17176
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 3988 16114 4016 16458
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3976 16108 4028 16114
rect 3976 16050 4028 16056
rect 3988 15706 4016 16050
rect 4080 15745 4108 16186
rect 4066 15736 4122 15745
rect 3976 15700 4028 15706
rect 4066 15671 4122 15680
rect 3976 15642 4028 15648
rect 3884 15632 3936 15638
rect 3884 15574 3936 15580
rect 3896 15450 3924 15574
rect 3804 15422 3924 15450
rect 3804 14958 3832 15422
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3896 15026 3924 15302
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3804 14618 3832 14894
rect 3988 14822 4016 15642
rect 4172 15162 4200 16526
rect 4264 16522 4292 17818
rect 4724 17678 4752 18226
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4356 16590 4384 16934
rect 4540 16794 4568 17138
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 4252 15564 4304 15570
rect 4356 15552 4384 16526
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4632 16114 4660 16458
rect 4724 16182 4752 17614
rect 4908 17270 4936 18294
rect 5092 18222 5120 18362
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5368 17354 5396 23054
rect 5724 23044 5776 23050
rect 5724 22986 5776 22992
rect 5736 22556 5764 22986
rect 5552 22528 5764 22556
rect 5552 20534 5580 22528
rect 6276 22500 6328 22506
rect 6276 22442 6328 22448
rect 5688 22332 5996 22352
rect 5688 22330 5694 22332
rect 5750 22330 5774 22332
rect 5830 22330 5854 22332
rect 5910 22330 5934 22332
rect 5990 22330 5996 22332
rect 5750 22278 5752 22330
rect 5932 22278 5934 22330
rect 5688 22276 5694 22278
rect 5750 22276 5774 22278
rect 5830 22276 5854 22278
rect 5910 22276 5934 22278
rect 5990 22276 5996 22278
rect 5688 22256 5996 22276
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 5644 21622 5672 21830
rect 5632 21616 5684 21622
rect 5632 21558 5684 21564
rect 6196 21486 6224 21830
rect 6184 21480 6236 21486
rect 6184 21422 6236 21428
rect 5688 21244 5996 21264
rect 5688 21242 5694 21244
rect 5750 21242 5774 21244
rect 5830 21242 5854 21244
rect 5910 21242 5934 21244
rect 5990 21242 5996 21244
rect 5750 21190 5752 21242
rect 5932 21190 5934 21242
rect 5688 21188 5694 21190
rect 5750 21188 5774 21190
rect 5830 21188 5854 21190
rect 5910 21188 5934 21190
rect 5990 21188 5996 21190
rect 5688 21168 5996 21188
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5644 20244 5672 20742
rect 5552 20216 5672 20244
rect 5552 19310 5580 20216
rect 5688 20156 5996 20176
rect 5688 20154 5694 20156
rect 5750 20154 5774 20156
rect 5830 20154 5854 20156
rect 5910 20154 5934 20156
rect 5990 20154 5996 20156
rect 5750 20102 5752 20154
rect 5932 20102 5934 20154
rect 5688 20100 5694 20102
rect 5750 20100 5774 20102
rect 5830 20100 5854 20102
rect 5910 20100 5934 20102
rect 5990 20100 5996 20102
rect 5688 20080 5996 20100
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 6012 19514 6040 19654
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5552 18154 5580 19110
rect 5688 19068 5996 19088
rect 5688 19066 5694 19068
rect 5750 19066 5774 19068
rect 5830 19066 5854 19068
rect 5910 19066 5934 19068
rect 5990 19066 5996 19068
rect 5750 19014 5752 19066
rect 5932 19014 5934 19066
rect 5688 19012 5694 19014
rect 5750 19012 5774 19014
rect 5830 19012 5854 19014
rect 5910 19012 5934 19014
rect 5990 19012 5996 19014
rect 5688 18992 5996 19012
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5276 17326 5396 17354
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 5092 16250 5120 16458
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4632 15910 4660 16050
rect 4724 15994 4752 16118
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4908 15994 4936 16050
rect 4724 15966 4936 15994
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4304 15536 4568 15552
rect 4304 15530 4580 15536
rect 4304 15524 4528 15530
rect 4252 15506 4304 15512
rect 4528 15472 4580 15478
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4632 15094 4660 15438
rect 4620 15088 4672 15094
rect 4066 15056 4122 15065
rect 4620 15030 4672 15036
rect 4066 14991 4122 15000
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 4080 14385 4108 14991
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4252 14408 4304 14414
rect 4066 14376 4122 14385
rect 4252 14350 4304 14356
rect 4066 14311 4122 14320
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1780 12850 1808 13126
rect 2424 12918 2452 13194
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12918 2728 13126
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2688 12912 2740 12918
rect 2688 12854 2740 12860
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10674 1532 10950
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1688 9654 1716 10542
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1412 8974 1440 9318
rect 1688 9042 1716 9590
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1780 6610 1808 12786
rect 2792 12714 2820 13262
rect 2884 12986 2912 13874
rect 3436 13462 3464 14010
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3712 13190 3740 13874
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3896 13025 3924 13670
rect 4172 13394 4200 13874
rect 4264 13870 4292 14350
rect 4344 14340 4396 14346
rect 4344 14282 4396 14288
rect 4356 13938 4384 14282
rect 4448 14006 4476 14894
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 3882 13016 3938 13025
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 3424 12980 3476 12986
rect 4172 13002 4200 13330
rect 4356 13326 4384 13874
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4080 12986 4200 13002
rect 3882 12951 3938 12960
rect 4068 12980 4200 12986
rect 3424 12922 3476 12928
rect 4120 12974 4200 12980
rect 4436 12980 4488 12986
rect 4068 12922 4120 12928
rect 4436 12922 4488 12928
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 12238 2820 12650
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 3436 11830 3464 12922
rect 4448 12442 4476 12922
rect 4540 12782 4568 14826
rect 4712 14000 4764 14006
rect 4712 13942 4764 13948
rect 4724 13326 4752 13942
rect 4816 13938 4844 15966
rect 5092 15502 5120 16186
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4908 15026 4936 15302
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 5092 14074 5120 14350
rect 4896 14068 4948 14074
rect 5080 14068 5132 14074
rect 4948 14028 5028 14056
rect 4896 14010 4948 14016
rect 5000 13938 5028 14028
rect 5080 14010 5132 14016
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4724 12866 4752 13126
rect 4816 12986 4844 13262
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4802 12880 4858 12889
rect 4724 12838 4802 12866
rect 4908 12850 4936 13738
rect 5000 13530 5028 13874
rect 5276 13734 5304 17326
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5368 16794 5396 17138
rect 5552 16794 5580 18090
rect 5688 17980 5996 18000
rect 5688 17978 5694 17980
rect 5750 17978 5774 17980
rect 5830 17978 5854 17980
rect 5910 17978 5934 17980
rect 5990 17978 5996 17980
rect 5750 17926 5752 17978
rect 5932 17926 5934 17978
rect 5688 17924 5694 17926
rect 5750 17924 5774 17926
rect 5830 17924 5854 17926
rect 5910 17924 5934 17926
rect 5990 17924 5996 17926
rect 5688 17904 5996 17924
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 5688 16892 5996 16912
rect 5688 16890 5694 16892
rect 5750 16890 5774 16892
rect 5830 16890 5854 16892
rect 5910 16890 5934 16892
rect 5990 16890 5996 16892
rect 5750 16838 5752 16890
rect 5932 16838 5934 16890
rect 5688 16836 5694 16838
rect 5750 16836 5774 16838
rect 5830 16836 5854 16838
rect 5910 16836 5934 16838
rect 5990 16836 5996 16838
rect 5688 16816 5996 16836
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 6104 16658 6132 17478
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5368 15502 5396 16390
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5552 15502 5580 15846
rect 5688 15804 5996 15824
rect 5688 15802 5694 15804
rect 5750 15802 5774 15804
rect 5830 15802 5854 15804
rect 5910 15802 5934 15804
rect 5990 15802 5996 15804
rect 5750 15750 5752 15802
rect 5932 15750 5934 15802
rect 5688 15748 5694 15750
rect 5750 15748 5774 15750
rect 5830 15748 5854 15750
rect 5910 15748 5934 15750
rect 5990 15748 5996 15750
rect 5688 15728 5996 15748
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 5460 15094 5488 15370
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5276 13258 5304 13398
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5100 13184 5152 13190
rect 5000 13144 5100 13172
rect 5000 12986 5028 13144
rect 5100 13126 5152 13132
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 4802 12815 4858 12824
rect 4896 12844 4948 12850
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3804 11354 3832 11834
rect 3896 11830 3924 12038
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 3884 11688 3936 11694
rect 3936 11648 4016 11676
rect 4080 11665 4108 12106
rect 4448 11762 4476 12378
rect 4816 12306 4844 12815
rect 4896 12786 4948 12792
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4540 11694 4568 12174
rect 4528 11688 4580 11694
rect 3884 11630 3936 11636
rect 3988 11558 4016 11648
rect 4066 11656 4122 11665
rect 4528 11630 4580 11636
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4066 11591 4122 11600
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1872 10266 1900 10610
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1964 10130 1992 11222
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 2148 10062 2176 10406
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2240 9586 2268 11086
rect 4172 10810 4200 11154
rect 4264 11150 4292 11562
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10266 3188 10610
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2424 9722 2452 10066
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2228 9580 2280 9586
rect 2148 9540 2228 9568
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1964 8634 1992 8842
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2148 7954 2176 9540
rect 2228 9522 2280 9528
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2240 8634 2268 8774
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2424 8430 2452 9658
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2792 8634 2820 9386
rect 3252 8974 3280 10406
rect 3974 10296 4030 10305
rect 3974 10231 4030 10240
rect 3988 10198 4016 10231
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 3608 9988 3660 9994
rect 3608 9930 3660 9936
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3436 9110 3464 9522
rect 3620 9450 3648 9930
rect 4080 9926 4108 10406
rect 4540 10266 4568 11630
rect 4724 11218 4752 11630
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3620 9178 3648 9386
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3436 8974 3464 9046
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3424 8968 3476 8974
rect 3712 8945 3740 9046
rect 3804 9042 3832 9318
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3424 8910 3476 8916
rect 3698 8936 3754 8945
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 3252 8430 3280 8910
rect 3436 8566 3464 8910
rect 3608 8900 3660 8906
rect 3698 8871 3754 8880
rect 3608 8842 3660 8848
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3620 8498 3648 8842
rect 4172 8498 4200 9998
rect 4344 9988 4396 9994
rect 4344 9930 4396 9936
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4264 8566 4292 9862
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2148 7478 2176 7890
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 2424 7342 2452 8366
rect 4356 8090 4384 9930
rect 4448 8906 4476 10066
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 2792 7478 2820 8026
rect 4068 8016 4120 8022
rect 4448 7970 4476 8434
rect 4632 8294 4660 9930
rect 4816 9722 4844 12242
rect 4908 11762 4936 12786
rect 5092 12442 5120 12854
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 5000 9926 5028 12310
rect 5184 11898 5212 12786
rect 5276 12617 5304 13194
rect 5368 12850 5396 14758
rect 5688 14716 5996 14736
rect 5688 14714 5694 14716
rect 5750 14714 5774 14716
rect 5830 14714 5854 14716
rect 5910 14714 5934 14716
rect 5990 14714 5996 14716
rect 5750 14662 5752 14714
rect 5932 14662 5934 14714
rect 5688 14660 5694 14662
rect 5750 14660 5774 14662
rect 5830 14660 5854 14662
rect 5910 14660 5934 14662
rect 5990 14660 5996 14662
rect 5688 14640 5996 14660
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5460 12986 5488 13874
rect 5552 13462 5580 13942
rect 5644 13870 5672 14214
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 5688 13628 5996 13648
rect 5688 13626 5694 13628
rect 5750 13626 5774 13628
rect 5830 13626 5854 13628
rect 5910 13626 5934 13628
rect 5990 13626 5996 13628
rect 5750 13574 5752 13626
rect 5932 13574 5934 13626
rect 5688 13572 5694 13574
rect 5750 13572 5774 13574
rect 5830 13572 5854 13574
rect 5910 13572 5934 13574
rect 5990 13572 5996 13574
rect 5688 13552 5996 13572
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 6104 13394 6132 13738
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 5540 13320 5592 13326
rect 6196 13274 6224 14962
rect 5540 13262 5592 13268
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5460 12889 5488 12922
rect 5446 12880 5502 12889
rect 5356 12844 5408 12850
rect 5446 12815 5502 12824
rect 5356 12786 5408 12792
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5262 12608 5318 12617
rect 5262 12543 5318 12552
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5460 11762 5488 12718
rect 5552 12646 5580 13262
rect 6104 13246 6224 13274
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12306 5580 12582
rect 5688 12540 5996 12560
rect 5688 12538 5694 12540
rect 5750 12538 5774 12540
rect 5830 12538 5854 12540
rect 5910 12538 5934 12540
rect 5990 12538 5996 12540
rect 5750 12486 5752 12538
rect 5932 12486 5934 12538
rect 5688 12484 5694 12486
rect 5750 12484 5774 12486
rect 5830 12484 5854 12486
rect 5910 12484 5934 12486
rect 5990 12484 5996 12486
rect 5688 12464 5996 12484
rect 5906 12336 5962 12345
rect 5540 12300 5592 12306
rect 5906 12271 5962 12280
rect 5540 12242 5592 12248
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5276 10674 5304 10950
rect 5264 10668 5316 10674
rect 5460 10656 5488 11698
rect 5552 11150 5580 12106
rect 5920 11762 5948 12271
rect 6104 12238 6132 13246
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11830 6040 12038
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 5688 11452 5996 11472
rect 5688 11450 5694 11452
rect 5750 11450 5774 11452
rect 5830 11450 5854 11452
rect 5910 11450 5934 11452
rect 5990 11450 5996 11452
rect 5750 11398 5752 11450
rect 5932 11398 5934 11450
rect 5688 11396 5694 11398
rect 5750 11396 5774 11398
rect 5830 11396 5854 11398
rect 5910 11396 5934 11398
rect 5990 11396 5996 11398
rect 5688 11376 5996 11396
rect 6104 11370 6132 11698
rect 6196 11626 6224 13126
rect 6288 12434 6316 22442
rect 6380 22094 6408 23990
rect 6460 23044 6512 23050
rect 6460 22986 6512 22992
rect 6472 22778 6500 22986
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 6460 22772 6512 22778
rect 6460 22714 6512 22720
rect 6656 22642 6684 22918
rect 6644 22636 6696 22642
rect 6748 22624 6776 24074
rect 6840 22778 6868 24142
rect 6932 24070 6960 24754
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6828 22636 6880 22642
rect 6748 22596 6828 22624
rect 6644 22578 6696 22584
rect 6828 22578 6880 22584
rect 6380 22066 6500 22094
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6380 18290 6408 19110
rect 6472 18970 6500 22066
rect 6552 22092 6604 22098
rect 6552 22034 6604 22040
rect 6564 20058 6592 22034
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6656 20942 6684 21966
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 6748 21010 6776 21286
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6644 20936 6696 20942
rect 6644 20878 6696 20884
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 6564 19446 6592 19994
rect 6552 19440 6604 19446
rect 6552 19382 6604 19388
rect 7024 19378 7052 21490
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6552 19236 6604 19242
rect 6552 19178 6604 19184
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6472 18358 6500 18566
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6472 17746 6500 18294
rect 6564 17746 6592 19178
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6472 16658 6500 16934
rect 6564 16658 6592 17682
rect 6656 17270 6684 18158
rect 6932 17882 6960 18158
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6656 16794 6684 17206
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6656 13870 6684 14894
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6656 13326 6684 13806
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6656 12714 6684 13262
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6644 12708 6696 12714
rect 6644 12650 6696 12656
rect 6288 12406 6500 12434
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6380 11762 6408 12174
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6104 11342 6224 11370
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5828 10742 5856 11086
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5540 10668 5592 10674
rect 5460 10628 5540 10656
rect 5264 10610 5316 10616
rect 5540 10610 5592 10616
rect 5276 9994 5304 10610
rect 5688 10364 5996 10384
rect 5688 10362 5694 10364
rect 5750 10362 5774 10364
rect 5830 10362 5854 10364
rect 5910 10362 5934 10364
rect 5990 10362 5996 10364
rect 5750 10310 5752 10362
rect 5932 10310 5934 10362
rect 5688 10308 5694 10310
rect 5750 10308 5774 10310
rect 5830 10308 5854 10310
rect 5910 10308 5934 10310
rect 5990 10308 5996 10310
rect 5688 10288 5996 10308
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 5000 8378 5028 9862
rect 5460 9586 5488 9862
rect 6012 9722 6040 10066
rect 6104 10062 6132 11222
rect 6196 11150 6224 11342
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6288 11014 6316 11630
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6380 9654 6408 9998
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 6380 9450 6408 9590
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 5688 9276 5996 9296
rect 5688 9274 5694 9276
rect 5750 9274 5774 9276
rect 5830 9274 5854 9276
rect 5910 9274 5934 9276
rect 5990 9274 5996 9276
rect 5750 9222 5752 9274
rect 5932 9222 5934 9274
rect 5688 9220 5694 9222
rect 5750 9220 5774 9222
rect 5830 9220 5854 9222
rect 5910 9220 5934 9222
rect 5990 9220 5996 9222
rect 5688 9200 5996 9220
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4908 8362 5028 8378
rect 4896 8356 5028 8362
rect 4948 8350 5028 8356
rect 4896 8298 4948 8304
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4068 7958 4120 7964
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1860 6792 1912 6798
rect 2056 6780 2084 7142
rect 2148 7002 2176 7210
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2148 6866 2176 6938
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 1912 6752 2084 6780
rect 1860 6734 1912 6740
rect 1688 5710 1716 6598
rect 1780 6582 1900 6610
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1412 5234 1440 5646
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1872 4146 1900 6582
rect 2240 5302 2268 7142
rect 2424 6866 2452 7278
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2792 6458 2820 7414
rect 3344 7410 3372 7686
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3804 7002 3832 7822
rect 4080 7585 4108 7958
rect 4356 7942 4476 7970
rect 4356 7818 4384 7942
rect 4632 7886 4660 8230
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4908 7818 4936 8298
rect 5092 8294 5120 8842
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5276 8430 5304 8570
rect 6104 8566 6132 9318
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5276 7886 5304 8366
rect 5460 8090 5488 8366
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5552 7954 5580 8502
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 5688 8188 5996 8208
rect 5688 8186 5694 8188
rect 5750 8186 5774 8188
rect 5830 8186 5854 8188
rect 5910 8186 5934 8188
rect 5990 8186 5996 8188
rect 5750 8134 5752 8186
rect 5932 8134 5934 8186
rect 5688 8132 5694 8134
rect 5750 8132 5774 8134
rect 5830 8132 5854 8134
rect 5910 8132 5934 8134
rect 5990 8132 5996 8134
rect 5688 8112 5996 8132
rect 6104 7954 6132 8366
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2976 6390 3004 6666
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3344 6322 3372 6598
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3344 5914 3372 6258
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3804 5710 3832 6054
rect 3896 5778 3924 6258
rect 4172 6254 4200 6802
rect 4356 6458 4384 7754
rect 5688 7100 5996 7120
rect 5688 7098 5694 7100
rect 5750 7098 5774 7100
rect 5830 7098 5854 7100
rect 5910 7098 5934 7100
rect 5990 7098 5996 7100
rect 5750 7046 5752 7098
rect 5932 7046 5934 7098
rect 5688 7044 5694 7046
rect 5750 7044 5774 7046
rect 5830 7044 5854 7046
rect 5910 7044 5934 7046
rect 5990 7044 5996 7046
rect 5688 7024 5996 7044
rect 6472 6882 6500 12406
rect 6656 12238 6684 12650
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6932 11762 6960 12786
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 11354 6776 11494
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7024 9450 7052 11222
rect 7116 9926 7144 25910
rect 7300 25906 7328 26522
rect 7380 26308 7432 26314
rect 7380 26250 7432 26256
rect 7392 26042 7420 26250
rect 7380 26036 7432 26042
rect 7380 25978 7432 25984
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7484 25362 7512 26998
rect 7576 25498 7604 28970
rect 7944 28558 7972 32056
rect 9036 30252 9088 30258
rect 9036 30194 9088 30200
rect 8024 29572 8076 29578
rect 8024 29514 8076 29520
rect 8036 29306 8064 29514
rect 9048 29510 9076 30194
rect 8300 29504 8352 29510
rect 8300 29446 8352 29452
rect 9036 29504 9088 29510
rect 9036 29446 9088 29452
rect 8024 29300 8076 29306
rect 8024 29242 8076 29248
rect 8312 29238 8340 29446
rect 8300 29232 8352 29238
rect 8300 29174 8352 29180
rect 7932 28552 7984 28558
rect 7932 28494 7984 28500
rect 7656 28212 7708 28218
rect 7656 28154 7708 28160
rect 7668 27538 7696 28154
rect 7656 27532 7708 27538
rect 7656 27474 7708 27480
rect 7748 27328 7800 27334
rect 7748 27270 7800 27276
rect 7760 26586 7788 27270
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7656 26308 7708 26314
rect 7656 26250 7708 26256
rect 7564 25492 7616 25498
rect 7564 25434 7616 25440
rect 7472 25356 7524 25362
rect 7472 25298 7524 25304
rect 7380 24064 7432 24070
rect 7380 24006 7432 24012
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7300 22982 7328 23666
rect 7288 22976 7340 22982
rect 7288 22918 7340 22924
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7300 19514 7328 20402
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7392 17218 7420 24006
rect 7484 23662 7512 25298
rect 7668 23866 7696 26250
rect 8312 26042 8340 29174
rect 8760 29096 8812 29102
rect 8760 29038 8812 29044
rect 8668 27872 8720 27878
rect 8772 27860 8800 29038
rect 8944 28076 8996 28082
rect 8944 28018 8996 28024
rect 8720 27832 8800 27860
rect 8668 27814 8720 27820
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 7944 25498 7972 25842
rect 8588 25838 8616 26862
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 7932 25492 7984 25498
rect 7932 25434 7984 25440
rect 8680 25226 8708 27814
rect 8956 27606 8984 28018
rect 8944 27600 8996 27606
rect 8944 27542 8996 27548
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 8864 27130 8892 27270
rect 8852 27124 8904 27130
rect 8852 27066 8904 27072
rect 9048 26382 9076 29446
rect 9140 28014 9168 32056
rect 10140 30252 10192 30258
rect 10140 30194 10192 30200
rect 9680 30184 9732 30190
rect 9680 30126 9732 30132
rect 9864 30184 9916 30190
rect 9864 30126 9916 30132
rect 9496 30048 9548 30054
rect 9496 29990 9548 29996
rect 9508 29578 9536 29990
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 9496 29572 9548 29578
rect 9496 29514 9548 29520
rect 9600 29102 9628 29582
rect 9588 29096 9640 29102
rect 9588 29038 9640 29044
rect 9692 28966 9720 30126
rect 9876 29238 9904 30126
rect 9864 29232 9916 29238
rect 9864 29174 9916 29180
rect 9772 29164 9824 29170
rect 9772 29106 9824 29112
rect 9956 29164 10008 29170
rect 9956 29106 10008 29112
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 9404 28076 9456 28082
rect 9404 28018 9456 28024
rect 9128 28008 9180 28014
rect 9128 27950 9180 27956
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 9140 27470 9168 27814
rect 9220 27668 9272 27674
rect 9220 27610 9272 27616
rect 9232 27470 9260 27610
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9140 27062 9168 27406
rect 9128 27056 9180 27062
rect 9128 26998 9180 27004
rect 9416 26994 9444 28018
rect 9692 27606 9720 28902
rect 9784 28490 9812 29106
rect 9968 28762 9996 29106
rect 10048 28960 10100 28966
rect 10048 28902 10100 28908
rect 10060 28762 10088 28902
rect 9956 28756 10008 28762
rect 9956 28698 10008 28704
rect 10048 28756 10100 28762
rect 10048 28698 10100 28704
rect 10060 28626 10088 28698
rect 10048 28620 10100 28626
rect 10048 28562 10100 28568
rect 9864 28552 9916 28558
rect 9862 28520 9864 28529
rect 9916 28520 9918 28529
rect 9772 28484 9824 28490
rect 9862 28455 9918 28464
rect 9772 28426 9824 28432
rect 9784 28218 9812 28426
rect 9864 28416 9916 28422
rect 9864 28358 9916 28364
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9680 27464 9732 27470
rect 9784 27452 9812 28154
rect 9876 27674 9904 28358
rect 10152 27878 10180 30194
rect 10232 29232 10284 29238
rect 10232 29174 10284 29180
rect 10244 28558 10272 29174
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10244 28422 10272 28494
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 10336 27985 10364 32056
rect 11624 30734 11652 32056
rect 11152 30728 11204 30734
rect 11152 30670 11204 30676
rect 11612 30728 11664 30734
rect 11612 30670 11664 30676
rect 10784 30592 10836 30598
rect 10784 30534 10836 30540
rect 10425 30492 10733 30512
rect 10425 30490 10431 30492
rect 10487 30490 10511 30492
rect 10567 30490 10591 30492
rect 10647 30490 10671 30492
rect 10727 30490 10733 30492
rect 10487 30438 10489 30490
rect 10669 30438 10671 30490
rect 10425 30436 10431 30438
rect 10487 30436 10511 30438
rect 10567 30436 10591 30438
rect 10647 30436 10671 30438
rect 10727 30436 10733 30438
rect 10425 30416 10733 30436
rect 10796 30326 10824 30534
rect 10784 30320 10836 30326
rect 10784 30262 10836 30268
rect 10425 29404 10733 29424
rect 10425 29402 10431 29404
rect 10487 29402 10511 29404
rect 10567 29402 10591 29404
rect 10647 29402 10671 29404
rect 10727 29402 10733 29404
rect 10487 29350 10489 29402
rect 10669 29350 10671 29402
rect 10425 29348 10431 29350
rect 10487 29348 10511 29350
rect 10567 29348 10591 29350
rect 10647 29348 10671 29350
rect 10727 29348 10733 29350
rect 10425 29328 10733 29348
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 11072 28694 11100 28902
rect 11060 28688 11112 28694
rect 11060 28630 11112 28636
rect 10784 28552 10836 28558
rect 10598 28520 10654 28529
rect 10598 28455 10600 28464
rect 10652 28455 10654 28464
rect 10782 28520 10784 28529
rect 10836 28520 10838 28529
rect 10782 28455 10838 28464
rect 10600 28426 10652 28432
rect 10425 28316 10733 28336
rect 10425 28314 10431 28316
rect 10487 28314 10511 28316
rect 10567 28314 10591 28316
rect 10647 28314 10671 28316
rect 10727 28314 10733 28316
rect 10487 28262 10489 28314
rect 10669 28262 10671 28314
rect 10425 28260 10431 28262
rect 10487 28260 10511 28262
rect 10567 28260 10591 28262
rect 10647 28260 10671 28262
rect 10727 28260 10733 28262
rect 10425 28240 10733 28260
rect 10322 27976 10378 27985
rect 10322 27911 10378 27920
rect 10140 27872 10192 27878
rect 10140 27814 10192 27820
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 9732 27424 9812 27452
rect 9864 27464 9916 27470
rect 9680 27406 9732 27412
rect 9864 27406 9916 27412
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 9036 26376 9088 26382
rect 9036 26318 9088 26324
rect 9128 25764 9180 25770
rect 9128 25706 9180 25712
rect 8944 25696 8996 25702
rect 8944 25638 8996 25644
rect 8668 25220 8720 25226
rect 8668 25162 8720 25168
rect 7748 25152 7800 25158
rect 7748 25094 7800 25100
rect 7760 24614 7788 25094
rect 8680 24750 8708 25162
rect 8668 24744 8720 24750
rect 8668 24686 8720 24692
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 7760 24274 7788 24550
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 7748 24268 7800 24274
rect 7748 24210 7800 24216
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 8036 23118 8064 23462
rect 8312 23186 8340 24346
rect 8864 24070 8892 24550
rect 8956 24206 8984 25638
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 9036 24197 9088 24203
rect 9036 24139 9088 24145
rect 8484 24064 8536 24070
rect 8484 24006 8536 24012
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 8496 23866 8524 24006
rect 9048 23866 9076 24139
rect 8484 23860 8536 23866
rect 8484 23802 8536 23808
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7576 20262 7604 21558
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7564 20256 7616 20262
rect 7564 20198 7616 20204
rect 7760 19514 7788 20402
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7484 17882 7512 18702
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7576 17678 7604 19314
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7668 18358 7696 18566
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7392 17190 7512 17218
rect 7576 17202 7604 17614
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 7208 16250 7236 16458
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7392 14958 7420 15438
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7484 12434 7512 17190
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7760 15094 7788 15302
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 7392 12406 7512 12434
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6564 8566 6592 9386
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6656 8090 6684 8434
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6748 7410 6776 8230
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6932 7478 6960 7822
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6564 7002 6592 7346
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6748 6934 6776 7346
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 5644 6854 6500 6882
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 5644 6746 5672 6854
rect 5552 6718 5672 6746
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 3976 6248 4028 6254
rect 4160 6248 4212 6254
rect 3976 6190 4028 6196
rect 4066 6216 4122 6225
rect 3988 5914 4016 6190
rect 4160 6190 4212 6196
rect 4066 6151 4122 6160
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4080 5846 4108 6151
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3436 5370 3464 5646
rect 4356 5642 4384 6394
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4540 5778 4568 6258
rect 5368 5914 5396 6258
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3804 4622 3832 4966
rect 3882 4856 3938 4865
rect 3882 4791 3938 4800
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3896 4554 3924 4791
rect 4080 4622 4108 5170
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 3884 4548 3936 4554
rect 3884 4490 3936 4496
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 848 3936 900 3942
rect 848 3878 900 3884
rect 860 800 888 3878
rect 1872 3505 1900 4082
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 2516 800 2544 3674
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3058 3924 3334
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 4080 2990 4108 4558
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4356 4010 4384 4490
rect 4448 4282 4476 5170
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4540 4146 4568 4422
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 3436 2145 3464 2314
rect 3422 2136 3478 2145
rect 3422 2071 3478 2080
rect 3148 1352 3200 1358
rect 3148 1294 3200 1300
rect 846 0 902 800
rect 2502 0 2558 800
rect 3160 785 3188 1294
rect 4264 800 4292 3674
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4632 3194 4660 3470
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4448 2650 4476 2994
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4632 2446 4660 3130
rect 4724 2582 4752 4014
rect 4908 3602 4936 4966
rect 5000 4826 5028 5170
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4816 2514 4844 2790
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 3146 776 3202 785
rect 3146 711 3202 720
rect 4250 0 4306 800
rect 5552 762 5580 6718
rect 5920 6458 5948 6734
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5688 6012 5996 6032
rect 5688 6010 5694 6012
rect 5750 6010 5774 6012
rect 5830 6010 5854 6012
rect 5910 6010 5934 6012
rect 5990 6010 5996 6012
rect 5750 5958 5752 6010
rect 5932 5958 5934 6010
rect 5688 5956 5694 5958
rect 5750 5956 5774 5958
rect 5830 5956 5854 5958
rect 5910 5956 5934 5958
rect 5990 5956 5996 5958
rect 5688 5936 5996 5956
rect 6104 5846 6132 6598
rect 6196 6322 6224 6734
rect 6748 6662 6776 6870
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6932 6390 6960 6938
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 6380 5302 6408 6122
rect 6564 5710 6592 6326
rect 6932 6118 6960 6326
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 5688 4924 5996 4944
rect 5688 4922 5694 4924
rect 5750 4922 5774 4924
rect 5830 4922 5854 4924
rect 5910 4922 5934 4924
rect 5990 4922 5996 4924
rect 5750 4870 5752 4922
rect 5932 4870 5934 4922
rect 5688 4868 5694 4870
rect 5750 4868 5774 4870
rect 5830 4868 5854 4870
rect 5910 4868 5934 4870
rect 5990 4868 5996 4870
rect 5688 4848 5996 4868
rect 6104 4622 6132 4966
rect 6380 4690 6408 5238
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6564 4690 6592 5170
rect 7024 5098 7052 9386
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7116 7818 7144 8842
rect 7208 7954 7236 10950
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7116 6730 7144 7142
rect 7208 7002 7236 7346
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7208 6322 7236 6802
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7300 6458 7328 6734
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5642 7236 6258
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 5688 3836 5996 3856
rect 5688 3834 5694 3836
rect 5750 3834 5774 3836
rect 5830 3834 5854 3836
rect 5910 3834 5934 3836
rect 5990 3834 5996 3836
rect 5750 3782 5752 3834
rect 5932 3782 5934 3834
rect 5688 3780 5694 3782
rect 5750 3780 5774 3782
rect 5830 3780 5854 3782
rect 5910 3780 5934 3782
rect 5990 3780 5996 3782
rect 5688 3760 5996 3780
rect 6104 3602 6132 4558
rect 6380 4146 6408 4626
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6472 4026 6500 4490
rect 6564 4146 6592 4626
rect 6932 4622 6960 4966
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6380 3998 6500 4026
rect 6380 3942 6408 3998
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6380 3534 6408 3878
rect 6932 3670 6960 3878
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 7024 3534 7052 5034
rect 7300 4826 7328 6190
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 5828 2922 5856 3470
rect 6748 3398 6776 3470
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 5920 3058 5948 3334
rect 6012 3058 6040 3334
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 5688 2748 5996 2768
rect 5688 2746 5694 2748
rect 5750 2746 5774 2748
rect 5830 2746 5854 2748
rect 5910 2746 5934 2748
rect 5990 2746 5996 2748
rect 5750 2694 5752 2746
rect 5932 2694 5934 2746
rect 5688 2692 5694 2694
rect 5750 2692 5774 2694
rect 5830 2692 5854 2694
rect 5910 2692 5934 2694
rect 5990 2692 5996 2694
rect 5688 2672 5996 2692
rect 6196 2514 6224 2790
rect 6472 2650 6500 2994
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6748 2446 6776 3334
rect 7392 2922 7420 12406
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7484 10810 7512 11086
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7484 8974 7512 10746
rect 7576 9178 7604 11834
rect 7668 11286 7696 12106
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7760 10266 7788 10610
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7576 6322 7604 9114
rect 7852 9110 7880 22918
rect 8220 22642 8248 22918
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 8220 19922 8248 22102
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 8300 21480 8352 21486
rect 8300 21422 8352 21428
rect 8312 21078 8340 21422
rect 8300 21072 8352 21078
rect 8300 21014 8352 21020
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 7932 19440 7984 19446
rect 7930 19408 7932 19417
rect 7984 19408 7986 19417
rect 7930 19343 7986 19352
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8312 17610 8340 18022
rect 8404 17610 8432 21558
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16590 8340 16934
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8404 16114 8432 17546
rect 8496 16538 8524 23802
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 8668 21888 8720 21894
rect 8668 21830 8720 21836
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8588 21146 8616 21422
rect 8680 21350 8708 21830
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8588 19922 8616 21082
rect 8956 21078 8984 21422
rect 9048 21350 9076 22374
rect 9140 21554 9168 25706
rect 9312 25152 9364 25158
rect 9312 25094 9364 25100
rect 9324 24274 9352 25094
rect 9220 24268 9272 24274
rect 9220 24210 9272 24216
rect 9312 24268 9364 24274
rect 9312 24210 9364 24216
rect 9232 23866 9260 24210
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 9324 23254 9352 24210
rect 9416 23730 9444 26930
rect 9600 26926 9628 27270
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 9600 26450 9628 26862
rect 9876 26790 9904 27406
rect 10048 26988 10100 26994
rect 10048 26930 10100 26936
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9864 26784 9916 26790
rect 9864 26726 9916 26732
rect 9588 26444 9640 26450
rect 9588 26386 9640 26392
rect 9692 26246 9720 26726
rect 9876 26382 9904 26726
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9680 26240 9732 26246
rect 9680 26182 9732 26188
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9692 25430 9720 26182
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9680 25424 9732 25430
rect 9680 25366 9732 25372
rect 9784 25242 9812 25774
rect 9876 25294 9904 26182
rect 9600 25226 9812 25242
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9588 25220 9812 25226
rect 9640 25214 9812 25220
rect 9588 25162 9640 25168
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9508 24410 9536 24754
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9600 24274 9628 25162
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 9956 25152 10008 25158
rect 9956 25094 10008 25100
rect 9876 24954 9904 25094
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 9680 24676 9732 24682
rect 9680 24618 9732 24624
rect 9588 24268 9640 24274
rect 9508 24228 9588 24256
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 9312 23248 9364 23254
rect 9312 23190 9364 23196
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9324 22778 9352 23054
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9312 22500 9364 22506
rect 9312 22442 9364 22448
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 8944 21072 8996 21078
rect 8944 21014 8996 21020
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8772 19854 8800 20266
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 8956 18222 8984 19858
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8956 17202 8984 18158
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9048 17082 9076 21286
rect 9140 21078 9168 21490
rect 9232 21350 9260 21898
rect 9220 21344 9272 21350
rect 9220 21286 9272 21292
rect 9128 21072 9180 21078
rect 9128 21014 9180 21020
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9140 20466 9168 20878
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 8956 17054 9076 17082
rect 8496 16510 8616 16538
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8496 16250 8524 16390
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8128 15502 8156 15846
rect 8496 15706 8524 15982
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8496 14074 8524 14350
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8404 13462 8432 13874
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8404 13326 8432 13398
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8312 11642 8340 12310
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11898 8432 12174
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 8128 11614 8340 11642
rect 7944 9654 7972 11562
rect 8128 11150 8156 11614
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8220 10674 8248 11494
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8312 10810 8340 11086
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8404 10742 8432 11834
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8128 10470 8156 10542
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 8128 9586 8156 10406
rect 8496 10062 8524 12242
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7668 6866 7696 7890
rect 7760 7410 7788 8230
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7484 4146 7512 6258
rect 7576 5710 7604 6258
rect 7668 5778 7696 6802
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7852 3738 7880 8298
rect 8036 7886 8064 8842
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8312 7410 8340 8502
rect 8588 8022 8616 16510
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8864 13938 8892 14282
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8864 13530 8892 13874
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8956 12374 8984 17054
rect 9140 16946 9168 20402
rect 9324 19961 9352 22442
rect 9416 22094 9444 23666
rect 9508 22778 9536 24228
rect 9588 24210 9640 24216
rect 9692 24206 9720 24618
rect 9772 24336 9824 24342
rect 9772 24278 9824 24284
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9784 23730 9812 24278
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9876 23594 9904 24890
rect 9968 23662 9996 25094
rect 10060 24410 10088 26930
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 10152 24188 10180 27814
rect 10796 27674 10824 28455
rect 10876 27872 10928 27878
rect 10876 27814 10928 27820
rect 10888 27674 10916 27814
rect 10784 27668 10836 27674
rect 10784 27610 10836 27616
rect 10876 27668 10928 27674
rect 10876 27610 10928 27616
rect 11072 27606 11100 28630
rect 11060 27600 11112 27606
rect 11060 27542 11112 27548
rect 10232 27532 10284 27538
rect 10232 27474 10284 27480
rect 10244 26790 10272 27474
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 10425 27228 10733 27248
rect 10425 27226 10431 27228
rect 10487 27226 10511 27228
rect 10567 27226 10591 27228
rect 10647 27226 10671 27228
rect 10727 27226 10733 27228
rect 10487 27174 10489 27226
rect 10669 27174 10671 27226
rect 10425 27172 10431 27174
rect 10487 27172 10511 27174
rect 10567 27172 10591 27174
rect 10647 27172 10671 27174
rect 10727 27172 10733 27174
rect 10425 27152 10733 27172
rect 10980 26994 11008 27406
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 10244 26586 10272 26726
rect 10232 26580 10284 26586
rect 10232 26522 10284 26528
rect 10425 26140 10733 26160
rect 10425 26138 10431 26140
rect 10487 26138 10511 26140
rect 10567 26138 10591 26140
rect 10647 26138 10671 26140
rect 10727 26138 10733 26140
rect 10487 26086 10489 26138
rect 10669 26086 10671 26138
rect 10425 26084 10431 26086
rect 10487 26084 10511 26086
rect 10567 26084 10591 26086
rect 10647 26084 10671 26086
rect 10727 26084 10733 26086
rect 10425 26064 10733 26084
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10612 25498 10640 25842
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10324 25288 10376 25294
rect 10324 25230 10376 25236
rect 10232 25152 10284 25158
rect 10232 25094 10284 25100
rect 10244 24682 10272 25094
rect 10336 24954 10364 25230
rect 10425 25052 10733 25072
rect 10425 25050 10431 25052
rect 10487 25050 10511 25052
rect 10567 25050 10591 25052
rect 10647 25050 10671 25052
rect 10727 25050 10733 25052
rect 10487 24998 10489 25050
rect 10669 24998 10671 25050
rect 10425 24996 10431 24998
rect 10487 24996 10511 24998
rect 10567 24996 10591 24998
rect 10647 24996 10671 24998
rect 10727 24996 10733 24998
rect 10425 24976 10733 24996
rect 10324 24948 10376 24954
rect 10324 24890 10376 24896
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10232 24676 10284 24682
rect 10232 24618 10284 24624
rect 10060 24160 10180 24188
rect 10060 23730 10088 24160
rect 10048 23724 10100 23730
rect 10048 23666 10100 23672
rect 9956 23656 10008 23662
rect 9956 23598 10008 23604
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9772 23588 9824 23594
rect 9772 23530 9824 23536
rect 9864 23588 9916 23594
rect 9864 23530 9916 23536
rect 9600 23186 9628 23530
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9588 23180 9640 23186
rect 9588 23122 9640 23128
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9600 22642 9628 22918
rect 9588 22636 9640 22642
rect 9588 22578 9640 22584
rect 9600 22506 9628 22578
rect 9692 22506 9720 23258
rect 9784 22642 9812 23530
rect 10060 23322 10088 23666
rect 10232 23588 10284 23594
rect 10232 23530 10284 23536
rect 10048 23316 10100 23322
rect 10048 23258 10100 23264
rect 9956 23180 10008 23186
rect 9956 23122 10008 23128
rect 9968 22778 9996 23122
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 10060 22642 10088 22986
rect 9772 22636 9824 22642
rect 10048 22636 10100 22642
rect 9824 22596 9996 22624
rect 9772 22578 9824 22584
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9680 22500 9732 22506
rect 9680 22442 9732 22448
rect 9692 22094 9720 22442
rect 9416 22066 9536 22094
rect 9692 22066 9904 22094
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9416 20874 9444 21490
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 9416 20602 9444 20810
rect 9508 20806 9536 22066
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9770 21992 9826 22001
rect 9600 21146 9628 21966
rect 9770 21927 9826 21936
rect 9784 21894 9812 21927
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9876 21554 9904 22066
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9968 21468 9996 22596
rect 10048 22578 10100 22584
rect 10060 22001 10088 22578
rect 10244 22574 10272 23530
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10046 21992 10102 22001
rect 10152 21962 10180 22374
rect 10046 21927 10102 21936
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 10244 21554 10272 22510
rect 10336 21622 10364 24754
rect 10600 24676 10652 24682
rect 10600 24618 10652 24624
rect 10612 24206 10640 24618
rect 10784 24404 10836 24410
rect 10836 24364 10916 24392
rect 10784 24346 10836 24352
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10784 24132 10836 24138
rect 10784 24074 10836 24080
rect 10425 23964 10733 23984
rect 10425 23962 10431 23964
rect 10487 23962 10511 23964
rect 10567 23962 10591 23964
rect 10647 23962 10671 23964
rect 10727 23962 10733 23964
rect 10487 23910 10489 23962
rect 10669 23910 10671 23962
rect 10425 23908 10431 23910
rect 10487 23908 10511 23910
rect 10567 23908 10591 23910
rect 10647 23908 10671 23910
rect 10727 23908 10733 23910
rect 10425 23888 10733 23908
rect 10796 23746 10824 24074
rect 10704 23718 10824 23746
rect 10704 23594 10732 23718
rect 10692 23588 10744 23594
rect 10692 23530 10744 23536
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10612 23118 10640 23462
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 10425 22876 10733 22896
rect 10425 22874 10431 22876
rect 10487 22874 10511 22876
rect 10567 22874 10591 22876
rect 10647 22874 10671 22876
rect 10727 22874 10733 22876
rect 10487 22822 10489 22874
rect 10669 22822 10671 22874
rect 10425 22820 10431 22822
rect 10487 22820 10511 22822
rect 10567 22820 10591 22822
rect 10647 22820 10671 22822
rect 10727 22820 10733 22822
rect 10425 22800 10733 22820
rect 10784 21956 10836 21962
rect 10784 21898 10836 21904
rect 10425 21788 10733 21808
rect 10425 21786 10431 21788
rect 10487 21786 10511 21788
rect 10567 21786 10591 21788
rect 10647 21786 10671 21788
rect 10727 21786 10733 21788
rect 10487 21734 10489 21786
rect 10669 21734 10671 21786
rect 10425 21732 10431 21734
rect 10487 21732 10511 21734
rect 10567 21732 10591 21734
rect 10647 21732 10671 21734
rect 10727 21732 10733 21734
rect 10425 21712 10733 21732
rect 10796 21690 10824 21898
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10324 21616 10376 21622
rect 10324 21558 10376 21564
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10140 21480 10192 21486
rect 9968 21440 10140 21468
rect 10140 21422 10192 21428
rect 9588 21140 9640 21146
rect 9588 21082 9640 21088
rect 10336 20942 10364 21558
rect 10508 21480 10560 21486
rect 10508 21422 10560 21428
rect 10520 20942 10548 21422
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9784 20398 9812 20878
rect 9864 20800 9916 20806
rect 9864 20742 9916 20748
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9496 20256 9548 20262
rect 9548 20216 9812 20244
rect 9496 20198 9548 20204
rect 9784 20058 9812 20216
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9310 19952 9366 19961
rect 9310 19887 9366 19896
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9496 19372 9548 19378
rect 9600 19360 9628 19450
rect 9680 19372 9732 19378
rect 9548 19332 9680 19360
rect 9496 19314 9548 19320
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9232 18358 9260 18770
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9600 17678 9628 19332
rect 9680 19314 9732 19320
rect 9784 19310 9812 19994
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9692 17882 9720 18702
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9048 16918 9168 16946
rect 9048 13734 9076 16918
rect 9784 16590 9812 17478
rect 9876 16726 9904 20742
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 10060 19514 10088 19722
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 10152 19378 10180 20538
rect 10244 19825 10272 20742
rect 10425 20700 10733 20720
rect 10425 20698 10431 20700
rect 10487 20698 10511 20700
rect 10567 20698 10591 20700
rect 10647 20698 10671 20700
rect 10727 20698 10733 20700
rect 10487 20646 10489 20698
rect 10669 20646 10671 20698
rect 10425 20644 10431 20646
rect 10487 20644 10511 20646
rect 10567 20644 10591 20646
rect 10647 20644 10671 20646
rect 10727 20644 10733 20646
rect 10425 20624 10733 20644
rect 10796 20534 10824 21014
rect 10784 20528 10836 20534
rect 10784 20470 10836 20476
rect 10230 19816 10286 19825
rect 10230 19751 10286 19760
rect 9956 19372 10008 19378
rect 10140 19372 10192 19378
rect 10008 19332 10088 19360
rect 9956 19314 10008 19320
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9968 18358 9996 18566
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 9968 16794 9996 17206
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9140 14346 9168 16050
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9232 14822 9260 15982
rect 9770 15600 9826 15609
rect 9770 15535 9826 15544
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9324 15094 9352 15302
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 13326 9076 13670
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8772 11762 8800 12038
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8864 10130 8892 12038
rect 9140 11762 9168 14010
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8956 11354 8984 11698
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9140 11234 9168 11290
rect 9048 11206 9168 11234
rect 9232 11218 9260 14758
rect 9692 14006 9720 15438
rect 9784 15366 9812 15535
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9784 15026 9812 15302
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12646 9352 13126
rect 9692 12850 9720 13942
rect 9784 13870 9812 14418
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9220 11212 9272 11218
rect 9048 11082 9076 11206
rect 9220 11154 9272 11160
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8956 9654 8984 9998
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8300 7404 8352 7410
rect 8760 7404 8812 7410
rect 8352 7364 8432 7392
rect 8300 7346 8352 7352
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6458 8340 6598
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8404 6186 8432 7364
rect 8760 7346 8812 7352
rect 8772 7002 8800 7346
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8496 6322 8524 6734
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 5030 8156 5646
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8128 4622 8156 4966
rect 8220 4826 8248 5170
rect 8404 5166 8432 6122
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8864 5370 8892 5578
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8956 5166 8984 5714
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8128 3942 8156 4150
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8128 3602 8156 3878
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 8036 3194 8064 3470
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8220 3194 8248 3334
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8312 3058 8340 3334
rect 8404 3126 8432 5102
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 5828 870 5948 898
rect 5828 762 5856 870
rect 5920 800 5948 870
rect 7668 800 7696 2926
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8496 2514 8524 2790
rect 8680 2582 8708 5102
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8864 2650 8892 2994
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 9048 1358 9076 11018
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 10062 9260 10406
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9324 7562 9352 12582
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9600 11098 9628 12310
rect 9876 11830 9904 16662
rect 10060 15026 10088 19332
rect 10140 19314 10192 19320
rect 10244 19258 10272 19751
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10425 19612 10733 19632
rect 10425 19610 10431 19612
rect 10487 19610 10511 19612
rect 10567 19610 10591 19612
rect 10647 19610 10671 19612
rect 10727 19610 10733 19612
rect 10487 19558 10489 19610
rect 10669 19558 10671 19610
rect 10425 19556 10431 19558
rect 10487 19556 10511 19558
rect 10567 19556 10591 19558
rect 10647 19556 10671 19558
rect 10727 19556 10733 19558
rect 10425 19536 10733 19556
rect 10796 19446 10824 19654
rect 10784 19440 10836 19446
rect 10784 19382 10836 19388
rect 10152 19230 10272 19258
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10152 14906 10180 19230
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10425 18524 10733 18544
rect 10425 18522 10431 18524
rect 10487 18522 10511 18524
rect 10567 18522 10591 18524
rect 10647 18522 10671 18524
rect 10727 18522 10733 18524
rect 10487 18470 10489 18522
rect 10669 18470 10671 18522
rect 10425 18468 10431 18470
rect 10487 18468 10511 18470
rect 10567 18468 10591 18470
rect 10647 18468 10671 18470
rect 10727 18468 10733 18470
rect 10425 18448 10733 18468
rect 10796 18086 10824 18702
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10425 17436 10733 17456
rect 10425 17434 10431 17436
rect 10487 17434 10511 17436
rect 10567 17434 10591 17436
rect 10647 17434 10671 17436
rect 10727 17434 10733 17436
rect 10487 17382 10489 17434
rect 10669 17382 10671 17434
rect 10425 17380 10431 17382
rect 10487 17380 10511 17382
rect 10567 17380 10591 17382
rect 10647 17380 10671 17382
rect 10727 17380 10733 17382
rect 10425 17360 10733 17380
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10244 15162 10272 16050
rect 10336 16046 10364 16934
rect 10796 16590 10824 18022
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10425 16348 10733 16368
rect 10425 16346 10431 16348
rect 10487 16346 10511 16348
rect 10567 16346 10591 16348
rect 10647 16346 10671 16348
rect 10727 16346 10733 16348
rect 10487 16294 10489 16346
rect 10669 16294 10671 16346
rect 10425 16292 10431 16294
rect 10487 16292 10511 16294
rect 10567 16292 10591 16294
rect 10647 16292 10671 16294
rect 10727 16292 10733 16294
rect 10425 16272 10733 16292
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10336 15366 10364 15982
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10425 15260 10733 15280
rect 10425 15258 10431 15260
rect 10487 15258 10511 15260
rect 10567 15258 10591 15260
rect 10647 15258 10671 15260
rect 10727 15258 10733 15260
rect 10487 15206 10489 15258
rect 10669 15206 10671 15258
rect 10425 15204 10431 15206
rect 10487 15204 10511 15206
rect 10567 15204 10591 15206
rect 10647 15204 10671 15206
rect 10727 15204 10733 15206
rect 10425 15184 10733 15204
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10796 15026 10824 15846
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10888 14906 10916 24364
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10980 23254 11008 23462
rect 10968 23248 11020 23254
rect 10968 23190 11020 23196
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 10980 20058 11008 20878
rect 11072 20602 11100 20878
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 11072 19990 11100 20334
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 18766 11100 19654
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11072 17882 11100 18702
rect 11164 18426 11192 30670
rect 11704 30252 11756 30258
rect 11704 30194 11756 30200
rect 12532 30252 12584 30258
rect 12532 30194 12584 30200
rect 11612 30048 11664 30054
rect 11612 29990 11664 29996
rect 11520 29640 11572 29646
rect 11520 29582 11572 29588
rect 11532 29102 11560 29582
rect 11624 29578 11652 29990
rect 11612 29572 11664 29578
rect 11612 29514 11664 29520
rect 11716 29510 11744 30194
rect 11980 30184 12032 30190
rect 11980 30126 12032 30132
rect 11992 29714 12020 30126
rect 11980 29708 12032 29714
rect 11980 29650 12032 29656
rect 11704 29504 11756 29510
rect 11704 29446 11756 29452
rect 11520 29096 11572 29102
rect 11520 29038 11572 29044
rect 11244 28484 11296 28490
rect 11244 28426 11296 28432
rect 11256 27606 11284 28426
rect 11532 28014 11560 29038
rect 11992 28150 12020 29650
rect 12164 29504 12216 29510
rect 12164 29446 12216 29452
rect 12072 28212 12124 28218
rect 12072 28154 12124 28160
rect 11980 28144 12032 28150
rect 11980 28086 12032 28092
rect 11520 28008 11572 28014
rect 11520 27950 11572 27956
rect 11992 27606 12020 28086
rect 11244 27600 11296 27606
rect 11244 27542 11296 27548
rect 11980 27600 12032 27606
rect 11980 27542 12032 27548
rect 12084 27130 12112 28154
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 12072 26920 12124 26926
rect 11978 26888 12034 26897
rect 12072 26862 12124 26868
rect 11978 26823 11980 26832
rect 12032 26823 12034 26832
rect 11980 26794 12032 26800
rect 12084 26450 12112 26862
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 12084 25838 12112 26386
rect 12176 25974 12204 29446
rect 12440 28756 12492 28762
rect 12440 28698 12492 28704
rect 12256 28416 12308 28422
rect 12256 28358 12308 28364
rect 12268 28150 12296 28358
rect 12256 28144 12308 28150
rect 12256 28086 12308 28092
rect 12452 27878 12480 28698
rect 12440 27872 12492 27878
rect 12440 27814 12492 27820
rect 12544 27470 12572 30194
rect 12624 29504 12676 29510
rect 12624 29446 12676 29452
rect 12636 29238 12664 29446
rect 12624 29232 12676 29238
rect 12624 29174 12676 29180
rect 12820 28626 12848 32056
rect 13912 30660 13964 30666
rect 13912 30602 13964 30608
rect 13268 30252 13320 30258
rect 13268 30194 13320 30200
rect 12900 30116 12952 30122
rect 12900 30058 12952 30064
rect 12912 29646 12940 30058
rect 13280 29646 13308 30194
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 13268 29640 13320 29646
rect 13268 29582 13320 29588
rect 12912 28762 12940 29582
rect 12900 28756 12952 28762
rect 12900 28698 12952 28704
rect 12808 28620 12860 28626
rect 12808 28562 12860 28568
rect 12624 28552 12676 28558
rect 12622 28520 12624 28529
rect 12676 28520 12678 28529
rect 12622 28455 12678 28464
rect 12992 27872 13044 27878
rect 12992 27814 13044 27820
rect 13176 27872 13228 27878
rect 13176 27814 13228 27820
rect 13004 27606 13032 27814
rect 12992 27600 13044 27606
rect 12992 27542 13044 27548
rect 13188 27470 13216 27814
rect 13280 27538 13308 29582
rect 13636 29572 13688 29578
rect 13636 29514 13688 29520
rect 13648 29306 13676 29514
rect 13924 29306 13952 30602
rect 13636 29300 13688 29306
rect 13636 29242 13688 29248
rect 13912 29300 13964 29306
rect 13912 29242 13964 29248
rect 13268 27532 13320 27538
rect 13268 27474 13320 27480
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12900 27464 12952 27470
rect 12900 27406 12952 27412
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 12912 27334 12940 27406
rect 12532 27328 12584 27334
rect 12532 27270 12584 27276
rect 12900 27328 12952 27334
rect 12900 27270 12952 27276
rect 12256 26988 12308 26994
rect 12256 26930 12308 26936
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12164 25968 12216 25974
rect 12164 25910 12216 25916
rect 12072 25832 12124 25838
rect 12072 25774 12124 25780
rect 11520 25696 11572 25702
rect 11520 25638 11572 25644
rect 11532 25362 11560 25638
rect 12268 25498 12296 26930
rect 12360 26518 12388 26930
rect 12544 26926 12572 27270
rect 12532 26920 12584 26926
rect 12532 26862 12584 26868
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 12348 26512 12400 26518
rect 12348 26454 12400 26460
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 11336 25356 11388 25362
rect 11336 25298 11388 25304
rect 11520 25356 11572 25362
rect 11520 25298 11572 25304
rect 11348 24750 11376 25298
rect 12256 24880 12308 24886
rect 12256 24822 12308 24828
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 12072 24744 12124 24750
rect 12072 24686 12124 24692
rect 11428 24676 11480 24682
rect 11428 24618 11480 24624
rect 11440 24410 11468 24618
rect 11428 24404 11480 24410
rect 11428 24346 11480 24352
rect 11440 23730 11468 24346
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 11256 23118 11284 23598
rect 11716 23526 11744 23666
rect 11808 23662 11836 23802
rect 12084 23746 12112 24686
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 12176 23866 12204 24074
rect 12268 24070 12296 24822
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12164 23860 12216 23866
rect 12164 23802 12216 23808
rect 11888 23724 11940 23730
rect 12084 23718 12204 23746
rect 12268 23730 12296 24006
rect 11888 23666 11940 23672
rect 11796 23656 11848 23662
rect 11796 23598 11848 23604
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 11704 23112 11756 23118
rect 11808 23100 11836 23598
rect 11900 23186 11928 23666
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 11756 23072 11836 23100
rect 11704 23054 11756 23060
rect 11336 21004 11388 21010
rect 11336 20946 11388 20952
rect 11348 20398 11376 20946
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 11348 19922 11376 20334
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10980 16658 11008 17070
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 11164 16590 11192 16934
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11256 16522 11284 18702
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11244 16516 11296 16522
rect 11244 16458 11296 16464
rect 11348 16250 11376 16526
rect 10968 16244 11020 16250
rect 11336 16244 11388 16250
rect 11020 16204 11100 16232
rect 10968 16186 11020 16192
rect 11072 16114 11100 16204
rect 11336 16186 11388 16192
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 10980 15570 11008 15846
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10060 14878 10180 14906
rect 10796 14878 10916 14906
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 14414 9996 14758
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9968 12374 9996 12786
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9600 11070 9812 11098
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9692 10674 9720 10746
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9600 8634 9628 9590
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9784 8362 9812 11070
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9876 8242 9904 11494
rect 9968 10742 9996 11698
rect 10060 10810 10088 14878
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10152 14006 10180 14214
rect 10425 14172 10733 14192
rect 10425 14170 10431 14172
rect 10487 14170 10511 14172
rect 10567 14170 10591 14172
rect 10647 14170 10671 14172
rect 10727 14170 10733 14172
rect 10487 14118 10489 14170
rect 10669 14118 10671 14170
rect 10425 14116 10431 14118
rect 10487 14116 10511 14118
rect 10567 14116 10591 14118
rect 10647 14116 10671 14118
rect 10727 14116 10733 14118
rect 10425 14096 10733 14116
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10425 13084 10733 13104
rect 10425 13082 10431 13084
rect 10487 13082 10511 13084
rect 10567 13082 10591 13084
rect 10647 13082 10671 13084
rect 10727 13082 10733 13084
rect 10487 13030 10489 13082
rect 10669 13030 10671 13082
rect 10425 13028 10431 13030
rect 10487 13028 10511 13030
rect 10567 13028 10591 13030
rect 10647 13028 10671 13030
rect 10727 13028 10733 13030
rect 10425 13008 10733 13028
rect 10796 12374 10824 14878
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10336 11762 10364 12242
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10425 11996 10733 12016
rect 10425 11994 10431 11996
rect 10487 11994 10511 11996
rect 10567 11994 10591 11996
rect 10647 11994 10671 11996
rect 10727 11994 10733 11996
rect 10487 11942 10489 11994
rect 10669 11942 10671 11994
rect 10425 11940 10431 11942
rect 10487 11940 10511 11942
rect 10567 11940 10591 11942
rect 10647 11940 10671 11942
rect 10727 11940 10733 11942
rect 10425 11920 10733 11940
rect 10796 11898 10824 12174
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10152 11354 10180 11698
rect 10888 11642 10916 12854
rect 10980 12322 11008 15302
rect 11072 15162 11100 15438
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 13870 11376 14350
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 10980 12294 11284 12322
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 10796 11626 10916 11642
rect 10784 11620 10916 11626
rect 10836 11614 10916 11620
rect 10968 11620 11020 11626
rect 10784 11562 10836 11568
rect 10968 11562 11020 11568
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10152 10742 10180 11154
rect 10324 11144 10376 11150
rect 10692 11144 10744 11150
rect 10324 11086 10376 11092
rect 10690 11112 10692 11121
rect 10744 11112 10746 11121
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 10244 10742 10272 11018
rect 10336 10810 10364 11086
rect 10690 11047 10746 11056
rect 10425 10908 10733 10928
rect 10425 10906 10431 10908
rect 10487 10906 10511 10908
rect 10567 10906 10591 10908
rect 10647 10906 10671 10908
rect 10727 10906 10733 10908
rect 10487 10854 10489 10906
rect 10669 10854 10671 10906
rect 10425 10852 10431 10854
rect 10487 10852 10511 10854
rect 10567 10852 10591 10854
rect 10647 10852 10671 10854
rect 10727 10852 10733 10854
rect 10425 10832 10733 10852
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10060 10198 10088 10610
rect 10336 10266 10364 10746
rect 10506 10704 10562 10713
rect 10506 10639 10508 10648
rect 10560 10639 10562 10648
rect 10508 10610 10560 10616
rect 10690 10568 10746 10577
rect 10416 10532 10468 10538
rect 10690 10503 10746 10512
rect 10416 10474 10468 10480
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 10428 10130 10456 10474
rect 10704 10470 10732 10503
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10416 10124 10468 10130
rect 10336 10084 10416 10112
rect 10336 9722 10364 10084
rect 10416 10066 10468 10072
rect 10425 9820 10733 9840
rect 10425 9818 10431 9820
rect 10487 9818 10511 9820
rect 10567 9818 10591 9820
rect 10647 9818 10671 9820
rect 10727 9818 10733 9820
rect 10487 9766 10489 9818
rect 10669 9766 10671 9818
rect 10425 9764 10431 9766
rect 10487 9764 10511 9766
rect 10567 9764 10591 9766
rect 10647 9764 10671 9766
rect 10727 9764 10733 9766
rect 10425 9744 10733 9764
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10336 9042 10364 9658
rect 10796 9654 10824 11562
rect 10980 11286 11008 11562
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10674 10916 10950
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10980 10606 11008 11018
rect 11072 10810 11100 12106
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11164 11150 11192 11494
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11164 10713 11192 11086
rect 11150 10704 11206 10713
rect 11150 10639 11206 10648
rect 10968 10600 11020 10606
rect 10874 10568 10930 10577
rect 10968 10542 11020 10548
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10874 10503 10876 10512
rect 10928 10503 10930 10512
rect 10876 10474 10928 10480
rect 10888 10130 10916 10474
rect 10980 10130 11008 10542
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10060 8566 10088 8774
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9784 8214 9904 8242
rect 9784 7750 9812 8214
rect 9968 8090 9996 8434
rect 10060 8430 10088 8502
rect 10336 8430 10364 8978
rect 10888 8974 10916 10066
rect 11072 10010 11100 10542
rect 11256 10062 11284 12294
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11348 11898 11376 12038
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 10980 9994 11100 10010
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 10968 9988 11100 9994
rect 11020 9982 11100 9988
rect 10968 9930 11020 9936
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11072 9042 11100 9522
rect 11256 9382 11284 9862
rect 11348 9450 11376 11290
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10425 8732 10733 8752
rect 10425 8730 10431 8732
rect 10487 8730 10511 8732
rect 10567 8730 10591 8732
rect 10647 8730 10671 8732
rect 10727 8730 10733 8732
rect 10487 8678 10489 8730
rect 10669 8678 10671 8730
rect 10425 8676 10431 8678
rect 10487 8676 10511 8678
rect 10567 8676 10591 8678
rect 10647 8676 10671 8678
rect 10727 8676 10733 8678
rect 10425 8656 10733 8676
rect 10888 8498 10916 8774
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11072 8498 11100 8570
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10060 7886 10088 8366
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 11072 7750 11100 8434
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 9140 7534 9352 7562
rect 9140 2378 9168 7534
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9600 6866 9628 7142
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9232 4622 9260 5306
rect 9508 5234 9536 5646
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9232 4146 9260 4558
rect 9416 4486 9444 5034
rect 9508 4690 9536 5170
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9600 3738 9628 4014
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9692 3534 9720 3878
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9232 3398 9260 3470
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9232 2446 9260 3334
rect 9784 3194 9812 7686
rect 10425 7644 10733 7664
rect 10425 7642 10431 7644
rect 10487 7642 10511 7644
rect 10567 7642 10591 7644
rect 10647 7642 10671 7644
rect 10727 7642 10733 7644
rect 10487 7590 10489 7642
rect 10669 7590 10671 7642
rect 10425 7588 10431 7590
rect 10487 7588 10511 7590
rect 10567 7588 10591 7590
rect 10647 7588 10671 7590
rect 10727 7588 10733 7590
rect 10425 7568 10733 7588
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9876 5914 9904 6802
rect 10244 6662 10272 6870
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9968 5710 9996 6054
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9968 5386 9996 5646
rect 10244 5642 10272 6598
rect 10336 5914 10364 6598
rect 10425 6556 10733 6576
rect 10425 6554 10431 6556
rect 10487 6554 10511 6556
rect 10567 6554 10591 6556
rect 10647 6554 10671 6556
rect 10727 6554 10733 6556
rect 10487 6502 10489 6554
rect 10669 6502 10671 6554
rect 10425 6500 10431 6502
rect 10487 6500 10511 6502
rect 10567 6500 10591 6502
rect 10647 6500 10671 6502
rect 10727 6500 10733 6502
rect 10425 6480 10733 6500
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11072 5914 11100 6258
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 9876 5358 9996 5386
rect 10244 5370 10272 5578
rect 10232 5364 10284 5370
rect 9876 5030 9904 5358
rect 10232 5306 10284 5312
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 4826 9904 4966
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9968 4758 9996 5102
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9968 3466 9996 4014
rect 10060 3534 10088 4558
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 9968 3194 9996 3402
rect 10152 3398 10180 5170
rect 10336 5166 10364 5714
rect 11164 5710 11192 9318
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10425 5468 10733 5488
rect 10425 5466 10431 5468
rect 10487 5466 10511 5468
rect 10567 5466 10591 5468
rect 10647 5466 10671 5468
rect 10727 5466 10733 5468
rect 10487 5414 10489 5466
rect 10669 5414 10671 5466
rect 10425 5412 10431 5414
rect 10487 5412 10511 5414
rect 10567 5412 10591 5414
rect 10647 5412 10671 5414
rect 10727 5412 10733 5414
rect 10425 5392 10733 5412
rect 10888 5234 10916 5646
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 11072 4826 11100 5170
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10244 4146 10272 4422
rect 10425 4380 10733 4400
rect 10425 4378 10431 4380
rect 10487 4378 10511 4380
rect 10567 4378 10591 4380
rect 10647 4378 10671 4380
rect 10727 4378 10733 4380
rect 10487 4326 10489 4378
rect 10669 4326 10671 4378
rect 10425 4324 10431 4326
rect 10487 4324 10511 4326
rect 10567 4324 10591 4326
rect 10647 4324 10671 4326
rect 10727 4324 10733 4326
rect 10425 4304 10733 4324
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10796 3670 10824 4490
rect 10888 4282 10916 4558
rect 10980 4486 11008 4694
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10980 4146 11008 4422
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10980 3738 11008 4082
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 11072 3602 11100 4014
rect 11256 4010 11284 9318
rect 11348 8974 11376 9386
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 7886 11376 8298
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11440 7698 11468 23054
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 11900 22710 11928 22918
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 11900 21554 11928 21830
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 12084 20874 12112 23122
rect 12176 22778 12204 23718
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12176 22166 12204 22714
rect 12164 22160 12216 22166
rect 12164 22102 12216 22108
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11716 19378 11744 19722
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11900 19378 11928 19654
rect 12176 19446 12204 22102
rect 12360 21894 12388 25842
rect 12440 23520 12492 23526
rect 12438 23488 12440 23497
rect 12492 23488 12494 23497
rect 12438 23423 12494 23432
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12452 22438 12480 23054
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 21894 12480 22374
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12544 21554 12572 26726
rect 13188 26450 13216 27406
rect 13268 27328 13320 27334
rect 13266 27296 13268 27305
rect 13360 27328 13412 27334
rect 13320 27296 13322 27305
rect 13360 27270 13412 27276
rect 13266 27231 13322 27240
rect 13372 26897 13400 27270
rect 13358 26888 13414 26897
rect 13358 26823 13414 26832
rect 13176 26444 13228 26450
rect 13176 26386 13228 26392
rect 12716 26308 12768 26314
rect 12716 26250 12768 26256
rect 12728 23322 12756 26250
rect 12808 25832 12860 25838
rect 12808 25774 12860 25780
rect 12820 25362 12848 25774
rect 13648 25362 13676 29242
rect 14016 28966 14044 32056
rect 15304 30666 15332 32056
rect 15292 30660 15344 30666
rect 15292 30602 15344 30608
rect 16028 30660 16080 30666
rect 16028 30602 16080 30608
rect 14464 30252 14516 30258
rect 14740 30252 14792 30258
rect 14516 30212 14596 30240
rect 14464 30194 14516 30200
rect 14280 29572 14332 29578
rect 14280 29514 14332 29520
rect 14292 29306 14320 29514
rect 14372 29504 14424 29510
rect 14372 29446 14424 29452
rect 14462 29472 14518 29481
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 14384 29170 14412 29446
rect 14462 29407 14518 29416
rect 14372 29164 14424 29170
rect 14372 29106 14424 29112
rect 14004 28960 14056 28966
rect 14004 28902 14056 28908
rect 14188 28144 14240 28150
rect 14188 28086 14240 28092
rect 13820 28076 13872 28082
rect 13820 28018 13872 28024
rect 13832 27606 13860 28018
rect 13820 27600 13872 27606
rect 13820 27542 13872 27548
rect 13728 27464 13780 27470
rect 13728 27406 13780 27412
rect 13740 26790 13768 27406
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 14004 26784 14056 26790
rect 14004 26726 14056 26732
rect 13740 26314 13768 26726
rect 13728 26308 13780 26314
rect 13728 26250 13780 26256
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13912 25696 13964 25702
rect 13912 25638 13964 25644
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 12716 23316 12768 23322
rect 12716 23258 12768 23264
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12360 20806 12388 21354
rect 12440 21140 12492 21146
rect 12544 21128 12572 21490
rect 12636 21418 12664 21490
rect 12624 21412 12676 21418
rect 12624 21354 12676 21360
rect 12820 21298 12848 25298
rect 13084 25152 13136 25158
rect 13084 25094 13136 25100
rect 13096 24954 13124 25094
rect 13084 24948 13136 24954
rect 13084 24890 13136 24896
rect 13452 24880 13504 24886
rect 13452 24822 13504 24828
rect 13464 24206 13492 24822
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 13544 24132 13596 24138
rect 13596 24092 13676 24120
rect 13544 24074 13596 24080
rect 13648 23730 13676 24092
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13648 23050 13676 23666
rect 13636 23044 13688 23050
rect 13636 22986 13688 22992
rect 13648 22778 13676 22986
rect 13636 22772 13688 22778
rect 13636 22714 13688 22720
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13556 22030 13584 22578
rect 13832 22030 13860 25638
rect 13924 24206 13952 25638
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 14016 23730 14044 26726
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14108 24070 14136 24142
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 14108 23526 14136 24006
rect 14200 23866 14228 28086
rect 14280 27532 14332 27538
rect 14280 27474 14332 27480
rect 14292 26926 14320 27474
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14280 25832 14332 25838
rect 14280 25774 14332 25780
rect 14292 25294 14320 25774
rect 14384 25362 14412 29106
rect 14476 27130 14504 29407
rect 14568 29238 14596 30212
rect 14740 30194 14792 30200
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 14556 29232 14608 29238
rect 14556 29174 14608 29180
rect 14752 29102 14780 30194
rect 14832 30184 14884 30190
rect 14832 30126 14884 30132
rect 14844 29850 14872 30126
rect 14832 29844 14884 29850
rect 14832 29786 14884 29792
rect 14740 29096 14792 29102
rect 14740 29038 14792 29044
rect 14648 29028 14700 29034
rect 14648 28970 14700 28976
rect 14660 28762 14688 28970
rect 14752 28762 14780 29038
rect 14844 29034 14872 29786
rect 15028 29034 15056 30194
rect 15163 29948 15471 29968
rect 15163 29946 15169 29948
rect 15225 29946 15249 29948
rect 15305 29946 15329 29948
rect 15385 29946 15409 29948
rect 15465 29946 15471 29948
rect 15225 29894 15227 29946
rect 15407 29894 15409 29946
rect 15163 29892 15169 29894
rect 15225 29892 15249 29894
rect 15305 29892 15329 29894
rect 15385 29892 15409 29894
rect 15465 29892 15471 29894
rect 15163 29872 15471 29892
rect 15660 29504 15712 29510
rect 15660 29446 15712 29452
rect 15672 29170 15700 29446
rect 15660 29164 15712 29170
rect 15660 29106 15712 29112
rect 14832 29028 14884 29034
rect 14832 28970 14884 28976
rect 15016 29028 15068 29034
rect 15016 28970 15068 28976
rect 14648 28756 14700 28762
rect 14648 28698 14700 28704
rect 14740 28756 14792 28762
rect 14740 28698 14792 28704
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 14556 28212 14608 28218
rect 14556 28154 14608 28160
rect 14568 27538 14596 28154
rect 14752 28082 14780 28494
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14648 27668 14700 27674
rect 14648 27610 14700 27616
rect 14556 27532 14608 27538
rect 14556 27474 14608 27480
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14660 25498 14688 27610
rect 14844 27606 14872 28358
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 14936 27674 14964 27814
rect 14924 27668 14976 27674
rect 14924 27610 14976 27616
rect 14832 27600 14884 27606
rect 14832 27542 14884 27548
rect 14740 27328 14792 27334
rect 14740 27270 14792 27276
rect 14648 25492 14700 25498
rect 14648 25434 14700 25440
rect 14372 25356 14424 25362
rect 14372 25298 14424 25304
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14096 23520 14148 23526
rect 14096 23462 14148 23468
rect 14108 23118 14136 23462
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 14108 22778 14136 23054
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14004 22636 14056 22642
rect 14004 22578 14056 22584
rect 14016 22098 14044 22578
rect 14004 22094 14056 22098
rect 14292 22094 14320 25230
rect 14660 24886 14688 25434
rect 14556 24880 14608 24886
rect 14556 24822 14608 24828
rect 14648 24880 14700 24886
rect 14648 24822 14700 24828
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14384 24410 14412 24618
rect 14372 24404 14424 24410
rect 14372 24346 14424 24352
rect 14464 24336 14516 24342
rect 14464 24278 14516 24284
rect 14004 22092 14136 22094
rect 14056 22066 14136 22092
rect 14292 22066 14412 22094
rect 14004 22034 14056 22040
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13556 21554 13584 21966
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 14016 21622 14044 21830
rect 14004 21616 14056 21622
rect 14004 21558 14056 21564
rect 14108 21554 14136 22066
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 12492 21100 12572 21128
rect 12636 21270 12848 21298
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12440 21082 12492 21088
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12452 20602 12480 20878
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 12164 19440 12216 19446
rect 12164 19382 12216 19388
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11520 19236 11572 19242
rect 11520 19178 11572 19184
rect 11532 18766 11560 19178
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11808 16998 11836 17682
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11532 12374 11560 16526
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11532 11694 11560 12310
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11624 11558 11652 12174
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11624 11150 11652 11290
rect 11716 11218 11744 13806
rect 11808 13530 11836 16934
rect 11900 16590 11928 18702
rect 11992 18290 12020 19382
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 12084 18698 12112 19314
rect 12268 18766 12296 20334
rect 12348 20324 12400 20330
rect 12348 20266 12400 20272
rect 12360 19854 12388 20266
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12360 19378 12388 19790
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12452 18850 12480 20402
rect 12532 20256 12584 20262
rect 12636 20244 12664 21270
rect 12912 20874 12940 21286
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12584 20216 12664 20244
rect 12716 20256 12768 20262
rect 12532 20198 12584 20204
rect 12716 20198 12768 20204
rect 12544 19768 12572 20198
rect 12728 19854 12756 20198
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12624 19780 12676 19786
rect 12544 19740 12624 19768
rect 12624 19722 12676 19728
rect 12912 19514 12940 20402
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12360 18834 12480 18850
rect 12636 18834 12664 19314
rect 13004 18902 13032 19790
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 12348 18828 12480 18834
rect 12400 18822 12480 18828
rect 12624 18828 12676 18834
rect 12348 18770 12400 18776
rect 12624 18770 12676 18776
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12256 18760 12308 18766
rect 12176 18720 12256 18748
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11992 16794 12020 18022
rect 12176 17542 12204 18720
rect 12256 18702 12308 18708
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 12084 16946 12112 17138
rect 12176 17134 12204 17478
rect 12164 17128 12216 17134
rect 12360 17082 12388 18566
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12452 17882 12480 18362
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12544 17814 12572 18362
rect 12728 18290 12756 18770
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 12820 18358 12848 18702
rect 12900 18692 12952 18698
rect 12900 18634 12952 18640
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12912 18086 12940 18634
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12532 17671 12584 17677
rect 12440 17650 12492 17656
rect 12532 17613 12584 17619
rect 12440 17592 12492 17598
rect 12164 17070 12216 17076
rect 12268 17054 12388 17082
rect 12084 16918 12204 16946
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 11992 16590 12020 16730
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11900 16436 11928 16526
rect 12084 16436 12112 16730
rect 11900 16408 12112 16436
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11900 15162 11928 16118
rect 12072 16108 12124 16114
rect 12176 16096 12204 16918
rect 12124 16068 12204 16096
rect 12072 16050 12124 16056
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 12176 14822 12204 16068
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12268 14482 12296 17054
rect 12452 16658 12480 17592
rect 12544 17513 12572 17613
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12530 17504 12586 17513
rect 12530 17439 12586 17448
rect 12728 17202 12756 17546
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12360 16114 12388 16458
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12544 16046 12572 16662
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12728 16454 12756 16594
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12636 16114 12664 16390
rect 12912 16250 12940 18022
rect 13004 17678 13032 18702
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13004 17338 13032 17614
rect 13096 17338 13124 21490
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13280 21010 13308 21286
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13280 20380 13308 20946
rect 14384 20874 14412 22066
rect 14476 22030 14504 24278
rect 14568 24070 14596 24822
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14752 23118 14780 27270
rect 14832 26920 14884 26926
rect 14832 26862 14884 26868
rect 14844 26450 14872 26862
rect 14832 26444 14884 26450
rect 14832 26386 14884 26392
rect 15028 26042 15056 28970
rect 15163 28860 15471 28880
rect 15163 28858 15169 28860
rect 15225 28858 15249 28860
rect 15305 28858 15329 28860
rect 15385 28858 15409 28860
rect 15465 28858 15471 28860
rect 15225 28806 15227 28858
rect 15407 28806 15409 28858
rect 15163 28804 15169 28806
rect 15225 28804 15249 28806
rect 15305 28804 15329 28806
rect 15385 28804 15409 28806
rect 15465 28804 15471 28806
rect 15163 28784 15471 28804
rect 15568 28416 15620 28422
rect 15568 28358 15620 28364
rect 15163 27772 15471 27792
rect 15163 27770 15169 27772
rect 15225 27770 15249 27772
rect 15305 27770 15329 27772
rect 15385 27770 15409 27772
rect 15465 27770 15471 27772
rect 15225 27718 15227 27770
rect 15407 27718 15409 27770
rect 15163 27716 15169 27718
rect 15225 27716 15249 27718
rect 15305 27716 15329 27718
rect 15385 27716 15409 27718
rect 15465 27716 15471 27718
rect 15163 27696 15471 27716
rect 15292 27600 15344 27606
rect 15292 27542 15344 27548
rect 15304 27452 15332 27542
rect 15384 27464 15436 27470
rect 15304 27432 15384 27452
rect 15436 27432 15438 27441
rect 15304 27424 15382 27432
rect 15382 27367 15438 27376
rect 15163 26684 15471 26704
rect 15163 26682 15169 26684
rect 15225 26682 15249 26684
rect 15305 26682 15329 26684
rect 15385 26682 15409 26684
rect 15465 26682 15471 26684
rect 15225 26630 15227 26682
rect 15407 26630 15409 26682
rect 15163 26628 15169 26630
rect 15225 26628 15249 26630
rect 15305 26628 15329 26630
rect 15385 26628 15409 26630
rect 15465 26628 15471 26630
rect 15163 26608 15471 26628
rect 15108 26444 15160 26450
rect 15108 26386 15160 26392
rect 15016 26036 15068 26042
rect 15016 25978 15068 25984
rect 15120 25838 15148 26386
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14844 25430 14872 25638
rect 15163 25596 15471 25616
rect 15163 25594 15169 25596
rect 15225 25594 15249 25596
rect 15305 25594 15329 25596
rect 15385 25594 15409 25596
rect 15465 25594 15471 25596
rect 15225 25542 15227 25594
rect 15407 25542 15409 25594
rect 15163 25540 15169 25542
rect 15225 25540 15249 25542
rect 15305 25540 15329 25542
rect 15385 25540 15409 25542
rect 15465 25540 15471 25542
rect 15163 25520 15471 25540
rect 14832 25424 14884 25430
rect 14832 25366 14884 25372
rect 15476 25220 15528 25226
rect 15476 25162 15528 25168
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14844 24206 14872 25094
rect 14924 24880 14976 24886
rect 14924 24822 14976 24828
rect 14936 24274 14964 24822
rect 15108 24812 15160 24818
rect 15028 24772 15108 24800
rect 15028 24614 15056 24772
rect 15108 24754 15160 24760
rect 15488 24682 15516 25162
rect 15476 24676 15528 24682
rect 15476 24618 15528 24624
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 14924 24268 14976 24274
rect 14924 24210 14976 24216
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14924 23588 14976 23594
rect 14924 23530 14976 23536
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14936 23050 14964 23530
rect 15028 23118 15056 24550
rect 15163 24508 15471 24528
rect 15163 24506 15169 24508
rect 15225 24506 15249 24508
rect 15305 24506 15329 24508
rect 15385 24506 15409 24508
rect 15465 24506 15471 24508
rect 15225 24454 15227 24506
rect 15407 24454 15409 24506
rect 15163 24452 15169 24454
rect 15225 24452 15249 24454
rect 15305 24452 15329 24454
rect 15385 24452 15409 24454
rect 15465 24452 15471 24454
rect 15163 24432 15471 24452
rect 15163 23420 15471 23440
rect 15163 23418 15169 23420
rect 15225 23418 15249 23420
rect 15305 23418 15329 23420
rect 15385 23418 15409 23420
rect 15465 23418 15471 23420
rect 15225 23366 15227 23418
rect 15407 23366 15409 23418
rect 15163 23364 15169 23366
rect 15225 23364 15249 23366
rect 15305 23364 15329 23366
rect 15385 23364 15409 23366
rect 15465 23364 15471 23366
rect 15163 23344 15471 23364
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 14924 23044 14976 23050
rect 14924 22986 14976 22992
rect 14832 22568 14884 22574
rect 14832 22510 14884 22516
rect 14844 22166 14872 22510
rect 14936 22506 14964 22986
rect 15028 22642 15056 23054
rect 15488 22642 15516 23054
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 14832 22160 14884 22166
rect 14832 22102 14884 22108
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13188 20352 13308 20380
rect 13188 18442 13216 20352
rect 13556 19922 13584 20470
rect 13832 20398 13860 20810
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13280 19174 13308 19450
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13268 18896 13320 18902
rect 13268 18838 13320 18844
rect 13280 18630 13308 18838
rect 13372 18766 13400 19314
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13188 18414 13400 18442
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 13188 17762 13216 18294
rect 13188 17734 13308 17762
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12360 14890 12388 15370
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12360 14006 12388 14826
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12452 13938 12480 15914
rect 12728 15570 12756 16118
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12532 15088 12584 15094
rect 12584 15036 12664 15042
rect 12532 15030 12664 15036
rect 12544 15014 12664 15030
rect 12728 15026 12756 15302
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11992 13326 12020 13874
rect 12452 13530 12480 13874
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11808 12238 11836 12786
rect 11900 12306 11928 13262
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11992 12102 12020 13262
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12084 12238 12112 12718
rect 12544 12714 12572 14826
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12636 12238 12664 15014
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 14414 12848 14758
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12728 14074 12756 14350
rect 12912 14346 12940 15914
rect 13004 14618 13032 17138
rect 13096 17134 13124 17274
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 13188 16454 13216 17614
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13280 15026 13308 17734
rect 13372 16726 13400 18414
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13464 16114 13492 19246
rect 13740 19174 13768 19994
rect 13832 19786 13860 20334
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13740 18834 13768 19110
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13556 18154 13584 18566
rect 13832 18442 13860 19722
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14292 18834 14320 19246
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 13648 18414 13860 18442
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 13544 17672 13596 17678
rect 13648 17660 13676 18414
rect 14384 18358 14412 19314
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 13596 17632 13676 17660
rect 14004 17672 14056 17678
rect 13544 17614 13596 17620
rect 14004 17614 14056 17620
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13740 17513 13768 17546
rect 14016 17542 14044 17614
rect 14004 17536 14056 17542
rect 13726 17504 13782 17513
rect 14004 17478 14056 17484
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 13726 17439 13782 17448
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13268 15020 13320 15026
rect 13188 14980 13268 15008
rect 13188 14618 13216 14980
rect 13268 14962 13320 14968
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13280 14550 13308 14758
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12912 13977 12940 14282
rect 13372 14278 13400 14758
rect 13464 14346 13492 16050
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15366 13584 15846
rect 13648 15434 13676 17002
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13556 15094 13584 15302
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 12898 13968 12954 13977
rect 12898 13903 12954 13912
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12820 12918 12848 13738
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12912 12374 12940 13903
rect 13648 13870 13676 15370
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13360 12640 13412 12646
rect 13464 12628 13492 13262
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13556 12782 13584 12922
rect 13544 12776 13596 12782
rect 13596 12736 13676 12764
rect 13544 12718 13596 12724
rect 13464 12600 13584 12628
rect 13360 12582 13412 12588
rect 13372 12434 13400 12582
rect 13372 12406 13492 12434
rect 12900 12368 12952 12374
rect 12900 12310 12952 12316
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11808 11694 11836 12038
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 11218 11836 11630
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11532 10826 11560 11086
rect 11532 10810 11652 10826
rect 11532 10804 11664 10810
rect 11532 10798 11612 10804
rect 11612 10746 11664 10752
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11532 7886 11560 8978
rect 11624 8974 11652 10746
rect 11716 10674 11744 11154
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11808 9926 11836 11018
rect 11900 11014 11928 11698
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10674 11928 10950
rect 12084 10674 12112 12038
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12176 11354 12204 11698
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12268 11150 12296 11562
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 11218 12572 11494
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 13096 10810 13124 11834
rect 13464 11132 13492 12406
rect 13556 12102 13584 12600
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13648 11218 13676 12736
rect 13740 12170 13768 17439
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13832 16590 13860 17138
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13832 15502 13860 16526
rect 14200 16250 14228 17478
rect 14292 17270 14320 18226
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 14108 14890 14136 15370
rect 14292 15026 14320 16050
rect 14384 15706 14412 16050
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14280 15020 14332 15026
rect 14476 15008 14504 21490
rect 14554 19680 14610 19689
rect 14554 19615 14610 19624
rect 14568 19242 14596 19615
rect 14556 19236 14608 19242
rect 14556 19178 14608 19184
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14568 17610 14596 17682
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14660 17542 14688 21830
rect 14752 21554 14780 22034
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14752 19242 14780 20402
rect 14844 19961 14872 20946
rect 14936 20942 14964 21286
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 15028 20602 15056 22578
rect 15163 22332 15471 22352
rect 15163 22330 15169 22332
rect 15225 22330 15249 22332
rect 15305 22330 15329 22332
rect 15385 22330 15409 22332
rect 15465 22330 15471 22332
rect 15225 22278 15227 22330
rect 15407 22278 15409 22330
rect 15163 22276 15169 22278
rect 15225 22276 15249 22278
rect 15305 22276 15329 22278
rect 15385 22276 15409 22278
rect 15465 22276 15471 22278
rect 15163 22256 15471 22276
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 15304 21690 15332 21966
rect 15382 21720 15438 21729
rect 15292 21684 15344 21690
rect 15382 21655 15438 21664
rect 15292 21626 15344 21632
rect 15396 21622 15424 21655
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15163 21244 15471 21264
rect 15163 21242 15169 21244
rect 15225 21242 15249 21244
rect 15305 21242 15329 21244
rect 15385 21242 15409 21244
rect 15465 21242 15471 21244
rect 15225 21190 15227 21242
rect 15407 21190 15409 21242
rect 15163 21188 15169 21190
rect 15225 21188 15249 21190
rect 15305 21188 15329 21190
rect 15385 21188 15409 21190
rect 15465 21188 15471 21190
rect 15163 21168 15471 21188
rect 15108 20936 15160 20942
rect 15108 20878 15160 20884
rect 15016 20596 15068 20602
rect 15016 20538 15068 20544
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 14830 19952 14886 19961
rect 14830 19887 14886 19896
rect 14936 19854 14964 20402
rect 15016 20392 15068 20398
rect 15014 20360 15016 20369
rect 15068 20360 15070 20369
rect 15014 20295 15070 20304
rect 15120 20244 15148 20878
rect 15028 20216 15148 20244
rect 15028 19854 15056 20216
rect 15163 20156 15471 20176
rect 15163 20154 15169 20156
rect 15225 20154 15249 20156
rect 15305 20154 15329 20156
rect 15385 20154 15409 20156
rect 15465 20154 15471 20156
rect 15225 20102 15227 20154
rect 15407 20102 15409 20154
rect 15163 20100 15169 20102
rect 15225 20100 15249 20102
rect 15305 20100 15329 20102
rect 15385 20100 15409 20102
rect 15465 20100 15471 20102
rect 15163 20080 15471 20100
rect 15474 19952 15530 19961
rect 15474 19887 15530 19896
rect 15488 19854 15516 19887
rect 15580 19854 15608 28358
rect 15672 26450 15700 29106
rect 15936 28416 15988 28422
rect 15936 28358 15988 28364
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 15764 27538 15792 27814
rect 15856 27606 15884 28018
rect 15844 27600 15896 27606
rect 15844 27542 15896 27548
rect 15752 27532 15804 27538
rect 15752 27474 15804 27480
rect 15764 27112 15792 27474
rect 15844 27124 15896 27130
rect 15764 27084 15844 27112
rect 15844 27066 15896 27072
rect 15948 27062 15976 28358
rect 15936 27056 15988 27062
rect 15936 26998 15988 27004
rect 15752 26784 15804 26790
rect 15752 26726 15804 26732
rect 15660 26444 15712 26450
rect 15660 26386 15712 26392
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15672 23118 15700 24754
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15672 21350 15700 22578
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15660 21072 15712 21078
rect 15660 21014 15712 21020
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 14936 19514 14964 19790
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 15163 19068 15471 19088
rect 15163 19066 15169 19068
rect 15225 19066 15249 19068
rect 15305 19066 15329 19068
rect 15385 19066 15409 19068
rect 15465 19066 15471 19068
rect 15225 19014 15227 19066
rect 15407 19014 15409 19066
rect 15163 19012 15169 19014
rect 15225 19012 15249 19014
rect 15305 19012 15329 19014
rect 15385 19012 15409 19014
rect 15465 19012 15471 19014
rect 15163 18992 15471 19012
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14660 17218 14688 17478
rect 14568 17190 14688 17218
rect 14568 15978 14596 17190
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14660 16998 14688 17070
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14556 15020 14608 15026
rect 14476 14980 14556 15008
rect 14280 14962 14332 14968
rect 14556 14962 14608 14968
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14108 14618 14136 14826
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 14016 13938 14044 14418
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12918 13860 13126
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 14292 12442 14320 14962
rect 14568 14634 14596 14962
rect 14476 14606 14596 14634
rect 14476 14550 14504 14606
rect 14464 14544 14516 14550
rect 14464 14486 14516 14492
rect 14660 14414 14688 16934
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14384 14074 14412 14350
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14384 12986 14412 14010
rect 14752 13938 14780 18226
rect 14844 18086 14872 18770
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14844 17066 14872 18022
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 14844 14822 14872 15914
rect 14936 14958 14964 17614
rect 15028 17202 15056 18634
rect 15580 18578 15608 19654
rect 15672 18766 15700 21014
rect 15764 20942 15792 26726
rect 16040 25702 16068 30602
rect 16500 30598 16528 32056
rect 16488 30592 16540 30598
rect 16488 30534 16540 30540
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 16120 30048 16172 30054
rect 16120 29990 16172 29996
rect 16132 29238 16160 29990
rect 16488 29572 16540 29578
rect 16488 29514 16540 29520
rect 16764 29572 16816 29578
rect 16764 29514 16816 29520
rect 16120 29232 16172 29238
rect 16120 29174 16172 29180
rect 16500 29102 16528 29514
rect 16776 29306 16804 29514
rect 16764 29300 16816 29306
rect 16764 29242 16816 29248
rect 16488 29096 16540 29102
rect 16488 29038 16540 29044
rect 16578 29064 16634 29073
rect 16120 28620 16172 28626
rect 16120 28562 16172 28568
rect 16132 26926 16160 28562
rect 16500 28150 16528 29038
rect 16578 28999 16580 29008
rect 16632 28999 16634 29008
rect 16580 28970 16632 28976
rect 16488 28144 16540 28150
rect 16488 28086 16540 28092
rect 16500 28014 16528 28086
rect 16960 28082 16988 30194
rect 17132 30116 17184 30122
rect 17132 30058 17184 30064
rect 17040 30048 17092 30054
rect 17040 29990 17092 29996
rect 17052 29850 17080 29990
rect 17040 29844 17092 29850
rect 17040 29786 17092 29792
rect 17052 29102 17080 29786
rect 17144 29102 17172 30058
rect 17604 29782 17632 30194
rect 17684 30048 17736 30054
rect 17684 29990 17736 29996
rect 17592 29776 17644 29782
rect 17592 29718 17644 29724
rect 17604 29481 17632 29718
rect 17696 29578 17724 29990
rect 17684 29572 17736 29578
rect 17684 29514 17736 29520
rect 17590 29472 17646 29481
rect 17590 29407 17646 29416
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 17224 29164 17276 29170
rect 17276 29124 17356 29152
rect 17224 29106 17276 29112
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 17132 29096 17184 29102
rect 17132 29038 17184 29044
rect 17328 29034 17356 29124
rect 17420 29073 17448 29242
rect 17406 29064 17462 29073
rect 17316 29028 17368 29034
rect 17406 28999 17462 29008
rect 17316 28970 17368 28976
rect 17788 28694 17816 32056
rect 18786 29064 18842 29073
rect 18786 28999 18842 29008
rect 17776 28688 17828 28694
rect 17776 28630 17828 28636
rect 17776 28552 17828 28558
rect 17776 28494 17828 28500
rect 17040 28416 17092 28422
rect 17040 28358 17092 28364
rect 17132 28416 17184 28422
rect 17132 28358 17184 28364
rect 16580 28076 16632 28082
rect 16580 28018 16632 28024
rect 16948 28076 17000 28082
rect 16948 28018 17000 28024
rect 16488 28008 16540 28014
rect 16210 27976 16266 27985
rect 16488 27950 16540 27956
rect 16210 27911 16266 27920
rect 16120 26920 16172 26926
rect 16120 26862 16172 26868
rect 16120 26240 16172 26246
rect 16120 26182 16172 26188
rect 16028 25696 16080 25702
rect 16028 25638 16080 25644
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15856 23118 15884 23802
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15856 22710 15884 22918
rect 15844 22704 15896 22710
rect 15844 22646 15896 22652
rect 16132 22642 16160 26182
rect 16224 24818 16252 27911
rect 16394 27432 16450 27441
rect 16394 27367 16396 27376
rect 16448 27367 16450 27376
rect 16396 27338 16448 27344
rect 16304 26988 16356 26994
rect 16304 26930 16356 26936
rect 16316 26314 16344 26930
rect 16408 26450 16436 27338
rect 16396 26444 16448 26450
rect 16396 26386 16448 26392
rect 16304 26308 16356 26314
rect 16304 26250 16356 26256
rect 16396 26308 16448 26314
rect 16396 26250 16448 26256
rect 16408 25906 16436 26250
rect 16396 25900 16448 25906
rect 16396 25842 16448 25848
rect 16500 25362 16528 27950
rect 16592 27470 16620 28018
rect 16856 28008 16908 28014
rect 16856 27950 16908 27956
rect 16868 27606 16896 27950
rect 16856 27600 16908 27606
rect 16856 27542 16908 27548
rect 16580 27464 16632 27470
rect 16580 27406 16632 27412
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16592 26382 16620 27406
rect 16684 26790 16712 27406
rect 16868 27010 16896 27542
rect 16960 27130 16988 28018
rect 17052 27470 17080 28358
rect 17144 28082 17172 28358
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 17236 27402 17264 28018
rect 17224 27396 17276 27402
rect 17224 27338 17276 27344
rect 16948 27124 17000 27130
rect 16948 27066 17000 27072
rect 16868 26982 16988 27010
rect 16856 26920 16908 26926
rect 16856 26862 16908 26868
rect 16672 26784 16724 26790
rect 16672 26726 16724 26732
rect 16868 26586 16896 26862
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 16960 26450 16988 26982
rect 17592 26784 17644 26790
rect 17592 26726 17644 26732
rect 17604 26586 17632 26726
rect 17592 26580 17644 26586
rect 17592 26522 17644 26528
rect 16948 26444 17000 26450
rect 16948 26386 17000 26392
rect 16580 26376 16632 26382
rect 16580 26318 16632 26324
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16776 25702 16804 26318
rect 16764 25696 16816 25702
rect 16764 25638 16816 25644
rect 17592 25696 17644 25702
rect 17592 25638 17644 25644
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 16212 24812 16264 24818
rect 16212 24754 16264 24760
rect 16500 23730 16528 25298
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 16592 24954 16620 25230
rect 17408 25220 17460 25226
rect 17408 25162 17460 25168
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16684 24410 16712 24754
rect 17420 24682 17448 25162
rect 17408 24676 17460 24682
rect 17408 24618 17460 24624
rect 16672 24404 16724 24410
rect 16672 24346 16724 24352
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 16684 23730 16712 24142
rect 16488 23724 16540 23730
rect 16488 23666 16540 23672
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 16224 23322 16252 23598
rect 16212 23316 16264 23322
rect 16212 23258 16264 23264
rect 16488 22704 16540 22710
rect 16488 22646 16540 22652
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16040 21962 16068 22374
rect 16028 21956 16080 21962
rect 16028 21898 16080 21904
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15856 21010 15884 21830
rect 16316 21729 16344 22374
rect 16302 21720 16358 21729
rect 16212 21684 16264 21690
rect 16302 21655 16358 21664
rect 16212 21626 16264 21632
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15764 20466 15792 20742
rect 15752 20460 15804 20466
rect 15856 20450 15884 20810
rect 15752 20402 15804 20408
rect 15844 20444 15896 20450
rect 15844 20386 15896 20392
rect 15752 20324 15804 20330
rect 15752 20266 15804 20272
rect 15764 19922 15792 20266
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15580 18550 15700 18578
rect 15163 17980 15471 18000
rect 15163 17978 15169 17980
rect 15225 17978 15249 17980
rect 15305 17978 15329 17980
rect 15385 17978 15409 17980
rect 15465 17978 15471 17980
rect 15225 17926 15227 17978
rect 15407 17926 15409 17978
rect 15163 17924 15169 17926
rect 15225 17924 15249 17926
rect 15305 17924 15329 17926
rect 15385 17924 15409 17926
rect 15465 17924 15471 17926
rect 15163 17904 15471 17924
rect 15672 17746 15700 18550
rect 15764 18426 15792 19654
rect 15856 18902 15884 19790
rect 15948 19378 15976 21490
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16040 20058 16068 20402
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 16040 19514 16068 19994
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15856 18306 15884 18838
rect 15764 18278 15884 18306
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15304 17134 15332 17546
rect 15764 17354 15792 18278
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15488 17326 15792 17354
rect 15488 17202 15516 17326
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15660 17196 15712 17202
rect 15712 17156 15792 17184
rect 15660 17138 15712 17144
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15163 16892 15471 16912
rect 15163 16890 15169 16892
rect 15225 16890 15249 16892
rect 15305 16890 15329 16892
rect 15385 16890 15409 16892
rect 15465 16890 15471 16892
rect 15225 16838 15227 16890
rect 15407 16838 15409 16890
rect 15163 16836 15169 16838
rect 15225 16836 15249 16838
rect 15305 16836 15329 16838
rect 15385 16836 15409 16838
rect 15465 16836 15471 16838
rect 15163 16816 15471 16836
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15212 16046 15240 16390
rect 15304 16114 15332 16458
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15163 15804 15471 15824
rect 15163 15802 15169 15804
rect 15225 15802 15249 15804
rect 15305 15802 15329 15804
rect 15385 15802 15409 15804
rect 15465 15802 15471 15804
rect 15225 15750 15227 15802
rect 15407 15750 15409 15802
rect 15163 15748 15169 15750
rect 15225 15748 15249 15750
rect 15305 15748 15329 15750
rect 15385 15748 15409 15750
rect 15465 15748 15471 15750
rect 15163 15728 15471 15748
rect 15580 15434 15608 17002
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15028 15026 15056 15370
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 14924 14952 14976 14958
rect 15292 14952 15344 14958
rect 14924 14894 14976 14900
rect 15028 14900 15292 14906
rect 15028 14894 15344 14900
rect 15028 14878 15332 14894
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 13462 14504 13670
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14476 12238 14504 12378
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 11354 13768 11630
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13544 11144 13596 11150
rect 13464 11104 13544 11132
rect 13544 11086 13596 11092
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 12084 9738 12112 10610
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 11992 9710 12112 9738
rect 11992 9586 12020 9710
rect 12728 9586 12756 10134
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11716 8974 11744 9318
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11716 8566 11744 8910
rect 12084 8634 12112 9522
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12268 8974 12296 9386
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 12176 8498 12204 8842
rect 12728 8498 12756 9522
rect 12912 9178 12940 9998
rect 13096 9518 13124 10746
rect 13740 10674 13768 11290
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13832 10062 13860 12174
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14660 11354 14688 12106
rect 14752 11354 14780 13874
rect 14844 12442 14872 14758
rect 15028 14618 15056 14878
rect 15163 14716 15471 14736
rect 15163 14714 15169 14716
rect 15225 14714 15249 14716
rect 15305 14714 15329 14716
rect 15385 14714 15409 14716
rect 15465 14714 15471 14716
rect 15225 14662 15227 14714
rect 15407 14662 15409 14714
rect 15163 14660 15169 14662
rect 15225 14660 15249 14662
rect 15305 14660 15329 14662
rect 15385 14660 15409 14662
rect 15465 14660 15471 14662
rect 15163 14640 15471 14660
rect 15580 14618 15608 14962
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15580 14482 15608 14554
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15672 14414 15700 15846
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 15028 13802 15056 13942
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 15163 13628 15471 13648
rect 15163 13626 15169 13628
rect 15225 13626 15249 13628
rect 15305 13626 15329 13628
rect 15385 13626 15409 13628
rect 15465 13626 15471 13628
rect 15225 13574 15227 13626
rect 15407 13574 15409 13626
rect 15163 13572 15169 13574
rect 15225 13572 15249 13574
rect 15305 13572 15329 13574
rect 15385 13572 15409 13574
rect 15465 13572 15471 13574
rect 15163 13552 15471 13572
rect 15580 13326 15608 14282
rect 15764 14074 15792 17156
rect 15856 15570 15884 18158
rect 15948 17338 15976 19314
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16040 18766 16068 19246
rect 16132 18834 16160 21422
rect 16224 19854 16252 21626
rect 16500 21146 16528 22646
rect 16684 22642 16712 23666
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16684 21690 16712 22578
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 17052 21962 17080 22374
rect 17236 22166 17264 22918
rect 17328 22710 17356 23122
rect 17316 22704 17368 22710
rect 17316 22646 17368 22652
rect 17420 22642 17448 24142
rect 17500 23656 17552 23662
rect 17500 23598 17552 23604
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 17420 22098 17448 22578
rect 17512 22574 17540 23598
rect 17500 22568 17552 22574
rect 17500 22510 17552 22516
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17040 21956 17092 21962
rect 17040 21898 17092 21904
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16500 20330 16528 20946
rect 16868 20874 16896 21286
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 17144 20602 17172 21490
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 16488 20324 16540 20330
rect 16488 20266 16540 20272
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16684 19378 16712 19790
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16868 19553 16896 19722
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 16854 19544 16910 19553
rect 16854 19479 16910 19488
rect 16868 19446 16896 19479
rect 16856 19440 16908 19446
rect 16856 19382 16908 19388
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 17144 19310 17172 19654
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16132 18222 16160 18770
rect 17144 18630 17172 19246
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 15948 16114 15976 17274
rect 16132 17218 16160 18158
rect 16040 17190 16160 17218
rect 16212 17196 16264 17202
rect 16040 16250 16068 17190
rect 16212 17138 16264 17144
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16132 16182 16160 17070
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 16120 16040 16172 16046
rect 15934 16008 15990 16017
rect 16120 15982 16172 15988
rect 15934 15943 15936 15952
rect 15988 15943 15990 15952
rect 15936 15914 15988 15920
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 15856 14414 15884 15506
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15948 14074 15976 15914
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 16040 15026 16068 15302
rect 16132 15162 16160 15982
rect 16224 15638 16252 17138
rect 16316 15706 16344 18566
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16684 17338 16712 17478
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16408 15502 16436 16050
rect 16592 15502 16620 16526
rect 16776 16250 16804 16594
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16684 15910 16712 16050
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 15570 16712 15846
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16224 14278 16252 14758
rect 16408 14550 16436 14758
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16500 14414 16528 14826
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15658 13968 15714 13977
rect 15948 13938 15976 14010
rect 16316 14006 16344 14350
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 14006 16436 14214
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 15936 13932 15988 13938
rect 15658 13903 15660 13912
rect 15712 13903 15714 13912
rect 15660 13874 15712 13880
rect 15856 13892 15936 13920
rect 15672 13394 15700 13874
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15028 12850 15056 13126
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15163 12540 15471 12560
rect 15163 12538 15169 12540
rect 15225 12538 15249 12540
rect 15305 12538 15329 12540
rect 15385 12538 15409 12540
rect 15465 12538 15471 12540
rect 15225 12486 15227 12538
rect 15407 12486 15409 12538
rect 15163 12484 15169 12486
rect 15225 12484 15249 12486
rect 15305 12484 15329 12486
rect 15385 12484 15409 12486
rect 15465 12484 15471 12486
rect 15163 12464 15471 12484
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15304 11898 15332 12106
rect 15488 12050 15516 12242
rect 15672 12238 15700 13194
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15488 12022 15700 12050
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15304 11626 15332 11834
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15163 11452 15471 11472
rect 15163 11450 15169 11452
rect 15225 11450 15249 11452
rect 15305 11450 15329 11452
rect 15385 11450 15409 11452
rect 15465 11450 15471 11452
rect 15225 11398 15227 11450
rect 15407 11398 15409 11450
rect 15163 11396 15169 11398
rect 15225 11396 15249 11398
rect 15305 11396 15329 11398
rect 15385 11396 15409 11398
rect 15465 11396 15471 11398
rect 15163 11376 15471 11396
rect 15580 11354 15608 11698
rect 14648 11348 14700 11354
rect 14568 11308 14648 11336
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13924 9654 13952 11086
rect 14568 9654 14596 11308
rect 14648 11290 14700 11296
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14660 10810 14688 11086
rect 15108 11008 15160 11014
rect 15292 11008 15344 11014
rect 15160 10956 15240 10962
rect 15108 10950 15240 10956
rect 15292 10950 15344 10956
rect 15120 10934 15240 10950
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 15212 10674 15240 10934
rect 15304 10810 15332 10950
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15396 10674 15424 11154
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 14844 10266 14872 10610
rect 15163 10364 15471 10384
rect 15163 10362 15169 10364
rect 15225 10362 15249 10364
rect 15305 10362 15329 10364
rect 15385 10362 15409 10364
rect 15465 10362 15471 10364
rect 15225 10310 15227 10362
rect 15407 10310 15409 10362
rect 15163 10308 15169 10310
rect 15225 10308 15249 10310
rect 15305 10308 15329 10310
rect 15385 10308 15409 10310
rect 15465 10308 15471 10310
rect 15163 10288 15471 10308
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 15580 9586 15608 11018
rect 15672 10538 15700 12022
rect 15856 11898 15884 13892
rect 15936 13874 15988 13880
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16408 13530 16436 13806
rect 16500 13802 16528 14350
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16408 12238 16436 13466
rect 16592 13394 16620 15438
rect 16776 15178 16804 16050
rect 16684 15150 16804 15178
rect 16684 14346 16712 15150
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16776 14618 16804 14962
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16776 13938 16804 14554
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16776 12918 16804 13874
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16684 12442 16712 12786
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16396 12232 16448 12238
rect 16764 12232 16816 12238
rect 16396 12174 16448 12180
rect 16684 12192 16764 12220
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 16592 11830 16620 12038
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 15764 11150 15792 11562
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15856 11082 15884 11630
rect 16684 11150 16712 12192
rect 16764 12174 16816 12180
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15672 9654 15700 10474
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 10010 15792 10406
rect 15764 9994 16068 10010
rect 15764 9988 16080 9994
rect 15764 9982 16028 9988
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 14936 9382 14964 9522
rect 15764 9518 15792 9982
rect 16028 9930 16080 9936
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 15844 9580 15896 9586
rect 16212 9580 16264 9586
rect 15896 9540 15976 9568
rect 15844 9522 15896 9528
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15948 9466 15976 9540
rect 16212 9522 16264 9528
rect 14924 9376 14976 9382
rect 15488 9364 15516 9454
rect 15660 9376 15712 9382
rect 15488 9336 15608 9364
rect 14924 9318 14976 9324
rect 14936 9178 14964 9318
rect 15163 9276 15471 9296
rect 15163 9274 15169 9276
rect 15225 9274 15249 9276
rect 15305 9274 15329 9276
rect 15385 9274 15409 9276
rect 15465 9274 15471 9276
rect 15225 9222 15227 9274
rect 15407 9222 15409 9274
rect 15163 9220 15169 9222
rect 15225 9220 15249 9222
rect 15305 9220 15329 9222
rect 15385 9220 15409 9222
rect 15465 9220 15471 9222
rect 15163 9200 15471 9220
rect 15580 9178 15608 9336
rect 15660 9318 15712 9324
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 12912 8498 12940 9114
rect 15672 8974 15700 9318
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11348 7670 11468 7698
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10152 2990 10180 3334
rect 10425 3292 10733 3312
rect 10425 3290 10431 3292
rect 10487 3290 10511 3292
rect 10567 3290 10591 3292
rect 10647 3290 10671 3292
rect 10727 3290 10733 3292
rect 10487 3238 10489 3290
rect 10669 3238 10671 3290
rect 10425 3236 10431 3238
rect 10487 3236 10511 3238
rect 10567 3236 10591 3238
rect 10647 3236 10671 3238
rect 10727 3236 10733 3238
rect 10425 3216 10733 3236
rect 10796 3058 10824 3334
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10980 2854 11008 3334
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 9324 800 9352 2790
rect 11072 2446 11100 2858
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 10425 2204 10733 2224
rect 10425 2202 10431 2204
rect 10487 2202 10511 2204
rect 10567 2202 10591 2204
rect 10647 2202 10671 2204
rect 10727 2202 10733 2204
rect 10487 2150 10489 2202
rect 10669 2150 10671 2202
rect 10425 2148 10431 2150
rect 10487 2148 10511 2150
rect 10567 2148 10591 2150
rect 10647 2148 10671 2150
rect 10727 2148 10733 2150
rect 10425 2128 10733 2148
rect 11164 1850 11192 3674
rect 11244 3664 11296 3670
rect 11348 3652 11376 7670
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11440 5914 11468 6734
rect 11532 6322 11560 7822
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4622 11560 4966
rect 12912 4690 12940 6258
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 12912 4146 12940 4626
rect 14936 4146 14964 5510
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 11428 3664 11480 3670
rect 11348 3624 11428 3652
rect 11244 3606 11296 3612
rect 11428 3606 11480 3612
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 11256 3482 11284 3606
rect 11336 3528 11388 3534
rect 11256 3476 11336 3482
rect 11256 3470 11388 3476
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11256 3454 11376 3470
rect 11900 3194 11928 3470
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11992 2514 12020 3334
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12452 2650 12480 2994
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11072 1822 11192 1850
rect 11072 800 11100 1822
rect 12728 800 12756 3606
rect 12912 3058 12940 4082
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14660 3738 14688 3878
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14462 3224 14518 3233
rect 14462 3159 14518 3168
rect 14476 3126 14504 3159
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 15028 3058 15056 8910
rect 15764 8634 15792 9454
rect 15844 9444 15896 9450
rect 15948 9438 16068 9466
rect 15844 9386 15896 9392
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15752 8424 15804 8430
rect 15750 8392 15752 8401
rect 15804 8392 15806 8401
rect 15750 8327 15806 8336
rect 15163 8188 15471 8208
rect 15163 8186 15169 8188
rect 15225 8186 15249 8188
rect 15305 8186 15329 8188
rect 15385 8186 15409 8188
rect 15465 8186 15471 8188
rect 15225 8134 15227 8186
rect 15407 8134 15409 8186
rect 15163 8132 15169 8134
rect 15225 8132 15249 8134
rect 15305 8132 15329 8134
rect 15385 8132 15409 8134
rect 15465 8132 15471 8134
rect 15163 8112 15471 8132
rect 15856 7546 15884 9386
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15948 8566 15976 8910
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15948 7478 15976 8502
rect 16040 8362 16068 9438
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 8974 16160 9318
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16224 8634 16252 9522
rect 16316 9110 16344 9862
rect 16500 9586 16528 10746
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16592 9926 16620 10202
rect 16684 10062 16712 11086
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16408 8430 16436 9114
rect 16684 9042 16712 9998
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16500 8362 16528 8910
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 15936 7472 15988 7478
rect 15936 7414 15988 7420
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15163 7100 15471 7120
rect 15163 7098 15169 7100
rect 15225 7098 15249 7100
rect 15305 7098 15329 7100
rect 15385 7098 15409 7100
rect 15465 7098 15471 7100
rect 15225 7046 15227 7098
rect 15407 7046 15409 7098
rect 15163 7044 15169 7046
rect 15225 7044 15249 7046
rect 15305 7044 15329 7046
rect 15385 7044 15409 7046
rect 15465 7044 15471 7046
rect 15163 7024 15471 7044
rect 15163 6012 15471 6032
rect 15163 6010 15169 6012
rect 15225 6010 15249 6012
rect 15305 6010 15329 6012
rect 15385 6010 15409 6012
rect 15465 6010 15471 6012
rect 15225 5958 15227 6010
rect 15407 5958 15409 6010
rect 15163 5956 15169 5958
rect 15225 5956 15249 5958
rect 15305 5956 15329 5958
rect 15385 5956 15409 5958
rect 15465 5956 15471 5958
rect 15163 5936 15471 5956
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15580 5166 15608 5714
rect 15672 5710 15700 7278
rect 15752 7268 15804 7274
rect 15752 7210 15804 7216
rect 15764 7002 15792 7210
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15856 5914 15884 6054
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15948 5710 15976 7278
rect 16040 6730 16068 7346
rect 16592 7274 16620 8910
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 6798 16252 7142
rect 16592 6866 16620 7210
rect 16684 6866 16712 7346
rect 16776 7206 16804 8230
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16408 6322 16436 6666
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 16132 5370 16160 5714
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16224 5234 16252 5578
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15163 4924 15471 4944
rect 15163 4922 15169 4924
rect 15225 4922 15249 4924
rect 15305 4922 15329 4924
rect 15385 4922 15409 4924
rect 15465 4922 15471 4924
rect 15225 4870 15227 4922
rect 15407 4870 15409 4922
rect 15163 4868 15169 4870
rect 15225 4868 15249 4870
rect 15305 4868 15329 4870
rect 15385 4868 15409 4870
rect 15465 4868 15471 4870
rect 15163 4848 15471 4868
rect 15163 3836 15471 3856
rect 15163 3834 15169 3836
rect 15225 3834 15249 3836
rect 15305 3834 15329 3836
rect 15385 3834 15409 3836
rect 15465 3834 15471 3836
rect 15225 3782 15227 3834
rect 15407 3782 15409 3834
rect 15163 3780 15169 3782
rect 15225 3780 15249 3782
rect 15305 3780 15329 3782
rect 15385 3780 15409 3782
rect 15465 3780 15471 3782
rect 15163 3760 15471 3780
rect 15580 3058 15608 4966
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15948 4282 15976 4558
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15948 3602 15976 3946
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 16040 3534 16068 4422
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16316 3602 16344 4082
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16408 3398 16436 6258
rect 16776 5778 16804 6666
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16592 5370 16620 5646
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16776 5234 16804 5578
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16776 4282 16804 5170
rect 16764 4276 16816 4282
rect 16764 4218 16816 4224
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 16684 4060 16712 4150
rect 16684 4032 16804 4060
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16684 3670 16712 3878
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14476 800 14504 2790
rect 15163 2748 15471 2768
rect 15163 2746 15169 2748
rect 15225 2746 15249 2748
rect 15305 2746 15329 2748
rect 15385 2746 15409 2748
rect 15465 2746 15471 2748
rect 15225 2694 15227 2746
rect 15407 2694 15409 2746
rect 15163 2692 15169 2694
rect 15225 2692 15249 2694
rect 15305 2692 15329 2694
rect 15385 2692 15409 2694
rect 15465 2692 15471 2694
rect 15163 2672 15471 2692
rect 16224 800 16252 3130
rect 16684 3058 16712 3606
rect 16776 3534 16804 4032
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16776 3369 16804 3470
rect 16762 3360 16818 3369
rect 16762 3295 16818 3304
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16868 1358 16896 16390
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 16960 15502 16988 16186
rect 17052 16114 17080 16390
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16960 14006 16988 15438
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16960 13190 16988 13942
rect 17052 13938 17080 14282
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17144 13818 17172 18566
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17236 14074 17264 14894
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17236 13938 17264 14010
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17052 13790 17172 13818
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16960 11898 16988 13126
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16960 4078 16988 10746
rect 17052 5098 17080 13790
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17144 12306 17172 13398
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17328 10810 17356 20946
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 17512 20534 17540 20742
rect 17500 20528 17552 20534
rect 17500 20470 17552 20476
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17420 18630 17448 20402
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17512 18698 17540 19110
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17420 18290 17448 18566
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17604 17218 17632 25638
rect 17684 24608 17736 24614
rect 17684 24550 17736 24556
rect 17696 24138 17724 24550
rect 17684 24132 17736 24138
rect 17684 24074 17736 24080
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17696 23050 17724 23462
rect 17684 23044 17736 23050
rect 17684 22986 17736 22992
rect 17684 22160 17736 22166
rect 17684 22102 17736 22108
rect 17696 21010 17724 22102
rect 17684 21004 17736 21010
rect 17684 20946 17736 20952
rect 17788 20602 17816 28494
rect 18800 27402 18828 28999
rect 18984 28994 19012 32056
rect 20180 30682 20208 32056
rect 20180 30654 20300 30682
rect 19901 30492 20209 30512
rect 19901 30490 19907 30492
rect 19963 30490 19987 30492
rect 20043 30490 20067 30492
rect 20123 30490 20147 30492
rect 20203 30490 20209 30492
rect 19963 30438 19965 30490
rect 20145 30438 20147 30490
rect 19901 30436 19907 30438
rect 19963 30436 19987 30438
rect 20043 30436 20067 30438
rect 20123 30436 20147 30438
rect 20203 30436 20209 30438
rect 19901 30416 20209 30436
rect 19901 29404 20209 29424
rect 19901 29402 19907 29404
rect 19963 29402 19987 29404
rect 20043 29402 20067 29404
rect 20123 29402 20147 29404
rect 20203 29402 20209 29404
rect 19963 29350 19965 29402
rect 20145 29350 20147 29402
rect 19901 29348 19907 29350
rect 19963 29348 19987 29350
rect 20043 29348 20067 29350
rect 20123 29348 20147 29350
rect 20203 29348 20209 29350
rect 19901 29328 20209 29348
rect 18984 28966 19288 28994
rect 18880 27872 18932 27878
rect 18880 27814 18932 27820
rect 18892 27470 18920 27814
rect 19260 27690 19288 28966
rect 19901 28316 20209 28336
rect 19901 28314 19907 28316
rect 19963 28314 19987 28316
rect 20043 28314 20067 28316
rect 20123 28314 20147 28316
rect 20203 28314 20209 28316
rect 19963 28262 19965 28314
rect 20145 28262 20147 28314
rect 19901 28260 19907 28262
rect 19963 28260 19987 28262
rect 20043 28260 20067 28262
rect 20123 28260 20147 28262
rect 20203 28260 20209 28262
rect 19901 28240 20209 28260
rect 19260 27662 19380 27690
rect 18880 27464 18932 27470
rect 18880 27406 18932 27412
rect 18788 27396 18840 27402
rect 18788 27338 18840 27344
rect 18892 26382 18920 27406
rect 19248 27396 19300 27402
rect 19248 27338 19300 27344
rect 18972 26852 19024 26858
rect 18972 26794 19024 26800
rect 18984 26450 19012 26794
rect 19260 26518 19288 27338
rect 19248 26512 19300 26518
rect 19248 26454 19300 26460
rect 18972 26444 19024 26450
rect 18972 26386 19024 26392
rect 18880 26376 18932 26382
rect 18880 26318 18932 26324
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 17972 25362 18000 26250
rect 19352 26042 19380 27662
rect 20272 27538 20300 30654
rect 21468 29510 21496 32056
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 20260 27532 20312 27538
rect 20260 27474 20312 27480
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 19901 27228 20209 27248
rect 19901 27226 19907 27228
rect 19963 27226 19987 27228
rect 20043 27226 20067 27228
rect 20123 27226 20147 27228
rect 20203 27226 20209 27228
rect 19963 27174 19965 27226
rect 20145 27174 20147 27226
rect 19901 27172 19907 27174
rect 19963 27172 19987 27174
rect 20043 27172 20067 27174
rect 20123 27172 20147 27174
rect 20203 27172 20209 27174
rect 19901 27152 20209 27172
rect 20456 27062 20484 27474
rect 20720 27396 20772 27402
rect 20720 27338 20772 27344
rect 20444 27056 20496 27062
rect 20444 26998 20496 27004
rect 20352 26988 20404 26994
rect 20352 26930 20404 26936
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20260 26784 20312 26790
rect 20260 26726 20312 26732
rect 19524 26308 19576 26314
rect 19524 26250 19576 26256
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 19352 25362 19380 25978
rect 19536 25770 19564 26250
rect 19901 26140 20209 26160
rect 19901 26138 19907 26140
rect 19963 26138 19987 26140
rect 20043 26138 20067 26140
rect 20123 26138 20147 26140
rect 20203 26138 20209 26140
rect 19963 26086 19965 26138
rect 20145 26086 20147 26138
rect 19901 26084 19907 26086
rect 19963 26084 19987 26086
rect 20043 26084 20067 26086
rect 20123 26084 20147 26086
rect 20203 26084 20209 26086
rect 19901 26064 20209 26084
rect 20076 25968 20128 25974
rect 20076 25910 20128 25916
rect 19524 25764 19576 25770
rect 19524 25706 19576 25712
rect 19536 25430 19564 25706
rect 20088 25498 20116 25910
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 19524 25424 19576 25430
rect 19524 25366 19576 25372
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 19340 25356 19392 25362
rect 19340 25298 19392 25304
rect 17972 24750 18000 25298
rect 19616 25288 19668 25294
rect 19614 25256 19616 25265
rect 19668 25256 19670 25265
rect 19614 25191 19670 25200
rect 19800 25220 19852 25226
rect 19800 25162 19852 25168
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 18064 24818 18092 25094
rect 19812 24954 19840 25162
rect 19901 25052 20209 25072
rect 19901 25050 19907 25052
rect 19963 25050 19987 25052
rect 20043 25050 20067 25052
rect 20123 25050 20147 25052
rect 20203 25050 20209 25052
rect 19963 24998 19965 25050
rect 20145 24998 20147 25050
rect 19901 24996 19907 24998
rect 19963 24996 19987 24998
rect 20043 24996 20067 24998
rect 20123 24996 20147 24998
rect 20203 24996 20209 24998
rect 19901 24976 20209 24996
rect 19800 24948 19852 24954
rect 19800 24890 19852 24896
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 19708 24812 19760 24818
rect 19708 24754 19760 24760
rect 17960 24744 18012 24750
rect 17960 24686 18012 24692
rect 17972 24256 18000 24686
rect 18248 24410 18276 24754
rect 19432 24676 19484 24682
rect 19432 24618 19484 24624
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 18236 24268 18288 24274
rect 17972 24228 18236 24256
rect 18236 24210 18288 24216
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 17880 23730 17908 24142
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 18156 23730 18184 24006
rect 18234 23760 18290 23769
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 18144 23724 18196 23730
rect 18234 23695 18236 23704
rect 18144 23666 18196 23672
rect 18288 23695 18290 23704
rect 18512 23724 18564 23730
rect 18236 23666 18288 23672
rect 18512 23666 18564 23672
rect 17880 22642 17908 23666
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18156 22642 18184 23054
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 18144 22636 18196 22642
rect 18144 22578 18196 22584
rect 17880 21690 17908 22578
rect 18156 22094 18184 22578
rect 18248 22098 18276 23666
rect 18524 23322 18552 23666
rect 18708 23497 18736 24142
rect 19260 23526 19288 24550
rect 19444 24206 19472 24618
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 19720 24070 19748 24754
rect 20272 24614 20300 26726
rect 20364 26518 20392 26930
rect 20548 26790 20576 26930
rect 20732 26858 20760 27338
rect 20824 27130 20852 28018
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 20812 27124 20864 27130
rect 20812 27066 20864 27072
rect 20812 26988 20864 26994
rect 20996 26988 21048 26994
rect 20864 26948 20996 26976
rect 20812 26930 20864 26936
rect 20720 26852 20772 26858
rect 20720 26794 20772 26800
rect 20536 26784 20588 26790
rect 20536 26726 20588 26732
rect 20352 26512 20404 26518
rect 20352 26454 20404 26460
rect 20812 25832 20864 25838
rect 20812 25774 20864 25780
rect 20824 25498 20852 25774
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 20916 24614 20944 26948
rect 20996 26930 21048 26936
rect 21100 26246 21128 27406
rect 22112 27402 22140 27814
rect 22664 27606 22692 32056
rect 22652 27600 22704 27606
rect 22652 27542 22704 27548
rect 21548 27396 21600 27402
rect 21548 27338 21600 27344
rect 22100 27396 22152 27402
rect 22100 27338 22152 27344
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 21456 26988 21508 26994
rect 21456 26930 21508 26936
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 21100 25838 21128 26182
rect 21088 25832 21140 25838
rect 21088 25774 21140 25780
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 19800 24132 19852 24138
rect 19800 24074 19852 24080
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19432 23792 19484 23798
rect 19338 23760 19394 23769
rect 19432 23734 19484 23740
rect 19338 23695 19340 23704
rect 19392 23695 19394 23704
rect 19340 23666 19392 23672
rect 19444 23526 19472 23734
rect 19248 23520 19300 23526
rect 18694 23488 18750 23497
rect 19248 23462 19300 23468
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 18694 23423 18750 23432
rect 18512 23316 18564 23322
rect 18512 23258 18564 23264
rect 17972 22066 18184 22094
rect 18236 22092 18288 22098
rect 17972 21894 18000 22066
rect 18236 22034 18288 22040
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17972 21078 18000 21830
rect 18144 21616 18196 21622
rect 18064 21576 18144 21604
rect 17960 21072 18012 21078
rect 17960 21014 18012 21020
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 17880 20466 17908 20742
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17684 20256 17736 20262
rect 17684 20198 17736 20204
rect 17696 20058 17724 20198
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17696 18426 17724 19314
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17788 18426 17816 19178
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17420 17190 17632 17218
rect 17420 12434 17448 17190
rect 17788 16590 17816 18362
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17604 15706 17632 15982
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17696 15570 17724 16118
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17604 14346 17632 14826
rect 17696 14414 17724 15506
rect 17788 15162 17816 15846
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17512 13938 17540 14214
rect 17788 13938 17816 15098
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17776 13932 17828 13938
rect 17776 13874 17828 13880
rect 17512 13394 17540 13874
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17420 12406 17540 12434
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17328 10130 17356 10542
rect 17408 10532 17460 10538
rect 17408 10474 17460 10480
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17144 8524 17172 9522
rect 17236 9178 17264 9590
rect 17328 9450 17356 10066
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17420 9382 17448 10474
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17236 8838 17264 9114
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17132 8518 17184 8524
rect 17132 8460 17184 8466
rect 17132 8288 17184 8294
rect 17130 8256 17132 8265
rect 17184 8256 17186 8265
rect 17130 8191 17186 8200
rect 17328 7562 17356 9114
rect 17420 7954 17448 9318
rect 17512 8945 17540 12406
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17592 9444 17644 9450
rect 17592 9386 17644 9392
rect 17604 9042 17632 9386
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17498 8936 17554 8945
rect 17696 8922 17724 10202
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17498 8871 17554 8880
rect 17604 8894 17724 8922
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17512 8566 17540 8774
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17236 7534 17356 7562
rect 17236 6798 17264 7534
rect 17420 7426 17448 7890
rect 17512 7886 17540 8502
rect 17604 8090 17632 8894
rect 17682 8800 17738 8809
rect 17682 8735 17738 8744
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17512 7546 17540 7822
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17604 7426 17632 8026
rect 17328 7398 17448 7426
rect 17512 7410 17632 7426
rect 17500 7404 17632 7410
rect 17328 7342 17356 7398
rect 17552 7398 17632 7404
rect 17500 7346 17552 7352
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17328 6866 17356 7278
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17420 6934 17448 7142
rect 17512 7002 17540 7346
rect 17696 7290 17724 8735
rect 17788 8634 17816 9522
rect 17880 9178 17908 19858
rect 17960 19780 18012 19786
rect 18064 19768 18092 21576
rect 18144 21558 18196 21564
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 18156 20942 18184 21422
rect 18328 21072 18380 21078
rect 18328 21014 18380 21020
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18234 19816 18290 19825
rect 18012 19740 18092 19768
rect 17960 19722 18012 19728
rect 18156 19514 18184 19790
rect 18234 19751 18290 19760
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 18064 18834 18092 19382
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18156 17746 18184 18226
rect 18248 18170 18276 19751
rect 18340 18834 18368 21014
rect 18708 20942 18736 23423
rect 19536 23322 19564 24006
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19720 23186 19748 24006
rect 19812 23866 19840 24074
rect 19901 23964 20209 23984
rect 19901 23962 19907 23964
rect 19963 23962 19987 23964
rect 20043 23962 20067 23964
rect 20123 23962 20147 23964
rect 20203 23962 20209 23964
rect 19963 23910 19965 23962
rect 20145 23910 20147 23962
rect 19901 23908 19907 23910
rect 19963 23908 19987 23910
rect 20043 23908 20067 23910
rect 20123 23908 20147 23910
rect 20203 23908 20209 23910
rect 19901 23888 20209 23908
rect 19800 23860 19852 23866
rect 19800 23802 19852 23808
rect 20272 23798 20300 24550
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20260 23792 20312 23798
rect 20260 23734 20312 23740
rect 20640 23730 20668 24006
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20180 23633 20208 23666
rect 20166 23624 20222 23633
rect 19984 23588 20036 23594
rect 20166 23559 20222 23568
rect 19984 23530 20036 23536
rect 19996 23497 20024 23530
rect 20444 23520 20496 23526
rect 19982 23488 20038 23497
rect 20444 23462 20496 23468
rect 19982 23423 20038 23432
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 19260 22710 19288 23122
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 19340 22976 19392 22982
rect 20180 22964 20208 23054
rect 20180 22936 20300 22964
rect 19340 22918 19392 22924
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 18880 22092 18932 22098
rect 18880 22034 18932 22040
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18892 20806 18920 22034
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18984 20942 19012 21286
rect 19248 21072 19300 21078
rect 19248 21014 19300 21020
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18880 20800 18932 20806
rect 18880 20742 18932 20748
rect 18708 20534 18736 20742
rect 19260 20534 19288 21014
rect 18696 20528 18748 20534
rect 18696 20470 18748 20476
rect 19248 20528 19300 20534
rect 19248 20470 19300 20476
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19168 20058 19196 20334
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18328 18828 18380 18834
rect 18328 18770 18380 18776
rect 18340 18358 18368 18770
rect 18432 18358 18460 19110
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18248 18142 18368 18170
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18144 17740 18196 17746
rect 18144 17682 18196 17688
rect 18248 17678 18276 18022
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 17960 17536 18012 17542
rect 18236 17536 18288 17542
rect 17960 17478 18012 17484
rect 18156 17496 18236 17524
rect 17972 17270 18000 17478
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 18156 16998 18184 17496
rect 18236 17478 18288 17484
rect 18340 17338 18368 18142
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17972 13326 18000 14350
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18156 12434 18184 16934
rect 18340 16726 18368 17274
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18524 16454 18552 19450
rect 18616 19446 18644 19722
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18708 19553 18736 19654
rect 18694 19544 18750 19553
rect 18694 19479 18750 19488
rect 18604 19440 18656 19446
rect 18604 19382 18656 19388
rect 18800 19378 18828 19790
rect 19260 19689 19288 19994
rect 19246 19680 19302 19689
rect 19246 19615 19302 19624
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 18984 18358 19012 18566
rect 18972 18352 19024 18358
rect 18972 18294 19024 18300
rect 19076 18086 19104 19110
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 19248 17264 19300 17270
rect 19248 17206 19300 17212
rect 19260 16726 19288 17206
rect 19352 17134 19380 22918
rect 19901 22876 20209 22896
rect 19901 22874 19907 22876
rect 19963 22874 19987 22876
rect 20043 22874 20067 22876
rect 20123 22874 20147 22876
rect 20203 22874 20209 22876
rect 19963 22822 19965 22874
rect 20145 22822 20147 22874
rect 19901 22820 19907 22822
rect 19963 22820 19987 22822
rect 20043 22820 20067 22822
rect 20123 22820 20147 22822
rect 20203 22820 20209 22822
rect 19901 22800 20209 22820
rect 20272 22778 20300 22936
rect 20260 22772 20312 22778
rect 20260 22714 20312 22720
rect 19708 22636 19760 22642
rect 19708 22578 19760 22584
rect 19720 22030 19748 22578
rect 20168 22500 20220 22506
rect 20168 22442 20220 22448
rect 19984 22432 20036 22438
rect 20180 22386 20208 22442
rect 20036 22380 20208 22386
rect 19984 22374 20208 22380
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 19996 22358 20208 22374
rect 19800 22092 19852 22098
rect 19996 22094 20024 22358
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 20088 22098 20116 22170
rect 19800 22034 19852 22040
rect 19904 22066 20024 22094
rect 20076 22092 20128 22098
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19444 20330 19472 20878
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19338 16960 19394 16969
rect 19338 16895 19394 16904
rect 19352 16794 19380 16895
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 18328 16176 18380 16182
rect 18328 16118 18380 16124
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18340 15706 18368 16118
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18510 15600 18566 15609
rect 18892 15586 18920 16118
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 18510 15535 18566 15544
rect 18800 15558 18920 15586
rect 18970 15600 19026 15609
rect 18524 15366 18552 15535
rect 18800 15502 18828 15558
rect 19076 15570 19104 15846
rect 19260 15570 19288 16186
rect 18970 15535 19026 15544
rect 19064 15564 19116 15570
rect 18984 15502 19012 15535
rect 19064 15506 19116 15512
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18800 15094 18828 15438
rect 18788 15088 18840 15094
rect 18788 15030 18840 15036
rect 18984 15026 19012 15438
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18708 13530 18736 13942
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 17972 12406 18184 12434
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17776 8424 17828 8430
rect 17774 8392 17776 8401
rect 17828 8392 17830 8401
rect 17774 8327 17830 8336
rect 17604 7262 17724 7290
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17408 6928 17460 6934
rect 17408 6870 17460 6876
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17144 5370 17172 5510
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17420 5166 17448 6870
rect 17500 6384 17552 6390
rect 17500 6326 17552 6332
rect 17512 5710 17540 6326
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17040 5092 17092 5098
rect 17040 5034 17092 5040
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17236 3777 17264 4014
rect 17222 3768 17278 3777
rect 17222 3703 17278 3712
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 17052 3058 17080 3402
rect 17512 3058 17540 4966
rect 17604 3505 17632 7262
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17696 5234 17724 7142
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 6322 17816 6598
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17788 5370 17816 5714
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17774 4176 17830 4185
rect 17774 4111 17830 4120
rect 17788 4078 17816 4111
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17788 3738 17816 3878
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17590 3496 17646 3505
rect 17590 3431 17646 3440
rect 17880 3126 17908 3946
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16960 2446 16988 2926
rect 17972 2774 18000 12406
rect 18248 12238 18276 12582
rect 19260 12442 19288 12582
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19352 12306 19380 16730
rect 19444 12434 19472 20266
rect 19536 19417 19564 20742
rect 19522 19408 19578 19417
rect 19522 19343 19578 19352
rect 19536 16250 19564 19343
rect 19628 17746 19656 21830
rect 19720 21690 19748 21966
rect 19708 21684 19760 21690
rect 19708 21626 19760 21632
rect 19812 21622 19840 22034
rect 19904 22030 19932 22066
rect 20076 22034 20128 22040
rect 20364 22030 20392 22374
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 19901 21788 20209 21808
rect 19901 21786 19907 21788
rect 19963 21786 19987 21788
rect 20043 21786 20067 21788
rect 20123 21786 20147 21788
rect 20203 21786 20209 21788
rect 19963 21734 19965 21786
rect 20145 21734 20147 21786
rect 19901 21732 19907 21734
rect 19963 21732 19987 21734
rect 20043 21732 20067 21734
rect 20123 21732 20147 21734
rect 20203 21732 20209 21734
rect 19901 21712 20209 21732
rect 19800 21616 19852 21622
rect 19800 21558 19852 21564
rect 20272 21554 20300 21898
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 19800 21412 19852 21418
rect 19800 21354 19852 21360
rect 19812 21146 19840 21354
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19812 20942 19840 21082
rect 20272 21026 20300 21490
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 20088 20998 20300 21026
rect 20088 20942 20116 20998
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 20076 20936 20128 20942
rect 20168 20936 20220 20942
rect 20076 20878 20128 20884
rect 20166 20904 20168 20913
rect 20220 20904 20222 20913
rect 20166 20839 20222 20848
rect 19901 20700 20209 20720
rect 19901 20698 19907 20700
rect 19963 20698 19987 20700
rect 20043 20698 20067 20700
rect 20123 20698 20147 20700
rect 20203 20698 20209 20700
rect 19963 20646 19965 20698
rect 20145 20646 20147 20698
rect 19901 20644 19907 20646
rect 19963 20644 19987 20646
rect 20043 20644 20067 20646
rect 20123 20644 20147 20646
rect 20203 20644 20209 20646
rect 19901 20624 20209 20644
rect 20272 20602 20300 20998
rect 20364 20942 20392 21422
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20364 20806 20392 20878
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 19812 19854 19840 20538
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19901 19612 20209 19632
rect 19901 19610 19907 19612
rect 19963 19610 19987 19612
rect 20043 19610 20067 19612
rect 20123 19610 20147 19612
rect 20203 19610 20209 19612
rect 19963 19558 19965 19610
rect 20145 19558 20147 19610
rect 19901 19556 19907 19558
rect 19963 19556 19987 19558
rect 20043 19556 20067 19558
rect 20123 19556 20147 19558
rect 20203 19556 20209 19558
rect 19901 19536 20209 19556
rect 20272 18766 20300 19926
rect 20364 19854 20392 20742
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 19901 18524 20209 18544
rect 19901 18522 19907 18524
rect 19963 18522 19987 18524
rect 20043 18522 20067 18524
rect 20123 18522 20147 18524
rect 20203 18522 20209 18524
rect 19963 18470 19965 18522
rect 20145 18470 20147 18522
rect 19901 18468 19907 18470
rect 19963 18468 19987 18470
rect 20043 18468 20067 18470
rect 20123 18468 20147 18470
rect 20203 18468 20209 18470
rect 19901 18448 20209 18468
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 19708 17808 19760 17814
rect 19708 17750 19760 17756
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19720 17270 19748 17750
rect 20168 17740 20220 17746
rect 20168 17682 20220 17688
rect 20180 17524 20208 17682
rect 20260 17536 20312 17542
rect 20180 17496 20260 17524
rect 20260 17478 20312 17484
rect 19901 17436 20209 17456
rect 19901 17434 19907 17436
rect 19963 17434 19987 17436
rect 20043 17434 20067 17436
rect 20123 17434 20147 17436
rect 20203 17434 20209 17436
rect 19963 17382 19965 17434
rect 20145 17382 20147 17434
rect 19901 17380 19907 17382
rect 19963 17380 19987 17382
rect 20043 17380 20067 17382
rect 20123 17380 20147 17382
rect 20203 17380 20209 17382
rect 19901 17360 20209 17380
rect 19708 17264 19760 17270
rect 19708 17206 19760 17212
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19522 16144 19578 16153
rect 19522 16079 19578 16088
rect 19536 15706 19564 16079
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19536 15094 19564 15642
rect 19524 15088 19576 15094
rect 19524 15030 19576 15036
rect 19628 14618 19656 17070
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19720 14890 19748 15438
rect 19812 15162 19840 17206
rect 19901 16348 20209 16368
rect 19901 16346 19907 16348
rect 19963 16346 19987 16348
rect 20043 16346 20067 16348
rect 20123 16346 20147 16348
rect 20203 16346 20209 16348
rect 19963 16294 19965 16346
rect 20145 16294 20147 16346
rect 19901 16292 19907 16294
rect 19963 16292 19987 16294
rect 20043 16292 20067 16294
rect 20123 16292 20147 16294
rect 20203 16292 20209 16294
rect 19901 16272 20209 16292
rect 19901 15260 20209 15280
rect 19901 15258 19907 15260
rect 19963 15258 19987 15260
rect 20043 15258 20067 15260
rect 20123 15258 20147 15260
rect 20203 15258 20209 15260
rect 19963 15206 19965 15258
rect 20145 15206 20147 15258
rect 19901 15204 19907 15206
rect 19963 15204 19987 15206
rect 20043 15204 20067 15206
rect 20123 15204 20147 15206
rect 20203 15204 20209 15206
rect 19901 15184 20209 15204
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19708 14884 19760 14890
rect 19708 14826 19760 14832
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19536 14074 19564 14350
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 19812 12434 19840 14962
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 19901 14172 20209 14192
rect 19901 14170 19907 14172
rect 19963 14170 19987 14172
rect 20043 14170 20067 14172
rect 20123 14170 20147 14172
rect 20203 14170 20209 14172
rect 19963 14118 19965 14170
rect 20145 14118 20147 14170
rect 19901 14116 19907 14118
rect 19963 14116 19987 14118
rect 20043 14116 20067 14118
rect 20123 14116 20147 14118
rect 20203 14116 20209 14118
rect 19901 14096 20209 14116
rect 20272 13938 20300 14282
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 19901 13084 20209 13104
rect 19901 13082 19907 13084
rect 19963 13082 19987 13084
rect 20043 13082 20067 13084
rect 20123 13082 20147 13084
rect 20203 13082 20209 13084
rect 19963 13030 19965 13082
rect 20145 13030 20147 13082
rect 19901 13028 19907 13030
rect 19963 13028 19987 13030
rect 20043 13028 20067 13030
rect 20123 13028 20147 13030
rect 20203 13028 20209 13030
rect 19901 13008 20209 13028
rect 19444 12406 19564 12434
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 18064 10810 18092 11018
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 18156 10674 18184 11290
rect 18144 10668 18196 10674
rect 18064 10628 18144 10656
rect 18064 8294 18092 10628
rect 18144 10610 18196 10616
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18340 10130 18368 10610
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18156 9110 18184 9998
rect 18432 9382 18460 10542
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 19076 9586 19104 9862
rect 19168 9654 19196 12174
rect 19536 12170 19564 12406
rect 19720 12406 19840 12434
rect 19720 12170 19748 12406
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 11354 19288 11698
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19352 11150 19380 11494
rect 19536 11354 19564 12106
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19628 11150 19656 11494
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19352 10742 19380 11086
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19628 10112 19656 11086
rect 19720 10742 19748 12106
rect 19901 11996 20209 12016
rect 19901 11994 19907 11996
rect 19963 11994 19987 11996
rect 20043 11994 20067 11996
rect 20123 11994 20147 11996
rect 20203 11994 20209 11996
rect 19963 11942 19965 11994
rect 20145 11942 20147 11994
rect 19901 11940 19907 11942
rect 19963 11940 19987 11942
rect 20043 11940 20067 11942
rect 20123 11940 20147 11942
rect 20203 11940 20209 11942
rect 19901 11920 20209 11940
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19812 11218 19840 11834
rect 20272 11626 20300 12174
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19901 10908 20209 10928
rect 19901 10906 19907 10908
rect 19963 10906 19987 10908
rect 20043 10906 20067 10908
rect 20123 10906 20147 10908
rect 20203 10906 20209 10908
rect 19963 10854 19965 10906
rect 20145 10854 20147 10906
rect 19901 10852 19907 10854
rect 19963 10852 19987 10854
rect 20043 10852 20067 10854
rect 20123 10852 20147 10854
rect 20203 10852 20209 10854
rect 19901 10832 20209 10852
rect 20364 10826 20392 18022
rect 20456 17218 20484 23462
rect 20812 23044 20864 23050
rect 20812 22986 20864 22992
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20536 22432 20588 22438
rect 20536 22374 20588 22380
rect 20548 22234 20576 22374
rect 20536 22228 20588 22234
rect 20536 22170 20588 22176
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20548 21486 20576 21966
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20536 21072 20588 21078
rect 20536 21014 20588 21020
rect 20548 20534 20576 21014
rect 20536 20528 20588 20534
rect 20536 20470 20588 20476
rect 20640 19310 20668 22918
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20732 21554 20760 22374
rect 20824 22234 20852 22986
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 20732 19922 20760 21490
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20732 19514 20760 19722
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20732 19378 20760 19450
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20640 18086 20668 19246
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20732 18290 20760 18566
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20626 17912 20682 17921
rect 20626 17847 20682 17856
rect 20640 17542 20668 17847
rect 20916 17678 20944 24550
rect 21100 23866 21128 25774
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 21100 23118 21128 23802
rect 21192 23594 21220 26930
rect 21468 26738 21496 26930
rect 21560 26858 21588 27338
rect 22664 27062 22692 27542
rect 22652 27056 22704 27062
rect 22652 26998 22704 27004
rect 21548 26852 21600 26858
rect 21548 26794 21600 26800
rect 21468 26710 21588 26738
rect 21560 26518 21588 26710
rect 23860 26586 23888 32056
rect 24639 29948 24947 29968
rect 24639 29946 24645 29948
rect 24701 29946 24725 29948
rect 24781 29946 24805 29948
rect 24861 29946 24885 29948
rect 24941 29946 24947 29948
rect 24701 29894 24703 29946
rect 24883 29894 24885 29946
rect 24639 29892 24645 29894
rect 24701 29892 24725 29894
rect 24781 29892 24805 29894
rect 24861 29892 24885 29894
rect 24941 29892 24947 29894
rect 24639 29872 24947 29892
rect 24639 28860 24947 28880
rect 24639 28858 24645 28860
rect 24701 28858 24725 28860
rect 24781 28858 24805 28860
rect 24861 28858 24885 28860
rect 24941 28858 24947 28860
rect 24701 28806 24703 28858
rect 24883 28806 24885 28858
rect 24639 28804 24645 28806
rect 24701 28804 24725 28806
rect 24781 28804 24805 28806
rect 24861 28804 24885 28806
rect 24941 28804 24947 28806
rect 24639 28784 24947 28804
rect 24639 27772 24947 27792
rect 24639 27770 24645 27772
rect 24701 27770 24725 27772
rect 24781 27770 24805 27772
rect 24861 27770 24885 27772
rect 24941 27770 24947 27772
rect 24701 27718 24703 27770
rect 24883 27718 24885 27770
rect 24639 27716 24645 27718
rect 24701 27716 24725 27718
rect 24781 27716 24805 27718
rect 24861 27716 24885 27718
rect 24941 27716 24947 27718
rect 24639 27696 24947 27716
rect 24639 26684 24947 26704
rect 24639 26682 24645 26684
rect 24701 26682 24725 26684
rect 24781 26682 24805 26684
rect 24861 26682 24885 26684
rect 24941 26682 24947 26684
rect 24701 26630 24703 26682
rect 24883 26630 24885 26682
rect 24639 26628 24645 26630
rect 24701 26628 24725 26630
rect 24781 26628 24805 26630
rect 24861 26628 24885 26630
rect 24941 26628 24947 26630
rect 24639 26608 24947 26628
rect 23848 26580 23900 26586
rect 23848 26522 23900 26528
rect 21548 26512 21600 26518
rect 21548 26454 21600 26460
rect 21456 24812 21508 24818
rect 21376 24772 21456 24800
rect 21272 24744 21324 24750
rect 21376 24732 21404 24772
rect 21456 24754 21508 24760
rect 21324 24704 21404 24732
rect 21272 24686 21324 24692
rect 21376 24206 21404 24704
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 21180 23588 21232 23594
rect 21180 23530 21232 23536
rect 21088 23112 21140 23118
rect 21088 23054 21140 23060
rect 21100 22098 21128 23054
rect 21088 22092 21140 22098
rect 21088 22034 21140 22040
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 21008 21418 21036 21898
rect 20996 21412 21048 21418
rect 20996 21354 21048 21360
rect 21088 21344 21140 21350
rect 21088 21286 21140 21292
rect 21100 20942 21128 21286
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21100 19938 21128 20878
rect 21180 20868 21232 20874
rect 21180 20810 21232 20816
rect 21192 20058 21220 20810
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 21100 19910 21220 19938
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21100 18290 21128 19110
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20640 17338 20668 17478
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20456 17190 20668 17218
rect 20732 17202 20760 17614
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20548 16522 20576 16934
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20548 15162 20576 15302
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20548 13394 20576 15098
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20548 12918 20576 13330
rect 20536 12912 20588 12918
rect 20536 12854 20588 12860
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20456 12306 20484 12786
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20640 10962 20668 17190
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20916 17184 20944 17478
rect 20996 17196 21048 17202
rect 20916 17156 20996 17184
rect 20916 16454 20944 17156
rect 20996 17138 21048 17144
rect 21192 17082 21220 19910
rect 21284 17814 21312 24006
rect 21376 20262 21404 24142
rect 21560 24070 21588 26454
rect 22100 26444 22152 26450
rect 22100 26386 22152 26392
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 21916 26308 21968 26314
rect 21916 26250 21968 26256
rect 21640 25900 21692 25906
rect 21640 25842 21692 25848
rect 21652 25362 21680 25842
rect 21928 25770 21956 26250
rect 22112 26042 22140 26386
rect 23020 26308 23072 26314
rect 23020 26250 23072 26256
rect 22100 26036 22152 26042
rect 22100 25978 22152 25984
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22744 25900 22796 25906
rect 22744 25842 22796 25848
rect 21916 25764 21968 25770
rect 21916 25706 21968 25712
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 21640 25356 21692 25362
rect 21640 25298 21692 25304
rect 21652 24682 21680 25298
rect 21916 25288 21968 25294
rect 22020 25242 22048 25638
rect 21968 25236 22048 25242
rect 21916 25230 22048 25236
rect 21928 25214 22048 25230
rect 22020 24682 22048 25214
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 21640 24676 21692 24682
rect 21640 24618 21692 24624
rect 21732 24676 21784 24682
rect 21732 24618 21784 24624
rect 22008 24676 22060 24682
rect 22008 24618 22060 24624
rect 21652 24070 21680 24618
rect 21744 24206 21772 24618
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21928 24410 21956 24550
rect 21916 24404 21968 24410
rect 21916 24346 21968 24352
rect 22008 24336 22060 24342
rect 22008 24278 22060 24284
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21548 24064 21600 24070
rect 21548 24006 21600 24012
rect 21640 24064 21692 24070
rect 21640 24006 21692 24012
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21546 20904 21602 20913
rect 21546 20839 21602 20848
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21468 19854 21496 20198
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21468 19378 21496 19790
rect 21560 19718 21588 20839
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21376 18630 21404 19314
rect 21468 19174 21496 19314
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 21560 18902 21588 19654
rect 21548 18896 21600 18902
rect 21548 18838 21600 18844
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21272 17808 21324 17814
rect 21272 17750 21324 17756
rect 21284 17202 21312 17750
rect 21652 17270 21680 22918
rect 21836 19718 21864 24074
rect 22020 23866 22048 24278
rect 22008 23860 22060 23866
rect 22008 23802 22060 23808
rect 22112 23254 22140 25094
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22204 23594 22232 24754
rect 22192 23588 22244 23594
rect 22192 23530 22244 23536
rect 22100 23248 22152 23254
rect 22100 23190 22152 23196
rect 22296 22778 22324 25842
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22572 25158 22600 25230
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22572 24886 22600 25094
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 22376 22976 22428 22982
rect 22376 22918 22428 22924
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22388 22710 22416 22918
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 21916 22432 21968 22438
rect 21916 22374 21968 22380
rect 21928 21962 21956 22374
rect 22112 22234 22140 22578
rect 22100 22228 22152 22234
rect 22100 22170 22152 22176
rect 21916 21956 21968 21962
rect 21916 21898 21968 21904
rect 22112 21690 22140 22170
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 22020 20602 22048 20946
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 22204 20466 22232 21082
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22572 20754 22600 22714
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22664 21690 22692 21830
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 22664 20874 22692 21286
rect 22652 20868 22704 20874
rect 22652 20810 22704 20816
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22204 19854 22232 20402
rect 22388 20262 22416 20742
rect 22572 20726 22692 20754
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 22468 19780 22520 19786
rect 22468 19722 22520 19728
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21744 18766 21772 19382
rect 22020 19378 22048 19654
rect 22112 19514 22140 19722
rect 22284 19712 22336 19718
rect 22284 19654 22336 19660
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22296 19446 22324 19654
rect 22284 19440 22336 19446
rect 22284 19382 22336 19388
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 22100 19372 22152 19378
rect 22152 19332 22232 19360
rect 22100 19314 22152 19320
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 21916 17332 21968 17338
rect 21916 17274 21968 17280
rect 21640 17264 21692 17270
rect 21640 17206 21692 17212
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21192 17054 21312 17082
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20732 14618 20760 14962
rect 20824 14890 20852 15370
rect 20812 14884 20864 14890
rect 20812 14826 20864 14832
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20732 14074 20760 14554
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20732 13802 20760 13874
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20732 12646 20760 13738
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20824 13394 20852 13670
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20732 11830 20760 12174
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20732 11150 20760 11630
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20824 11354 20852 11562
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20640 10934 20760 10962
rect 20364 10798 20668 10826
rect 19708 10736 19760 10742
rect 19708 10678 19760 10684
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 19708 10124 19760 10130
rect 19628 10084 19708 10112
rect 19708 10066 19760 10072
rect 20456 10062 20484 10610
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18144 9104 18196 9110
rect 18196 9064 18276 9092
rect 18144 9046 18196 9052
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18156 8634 18184 8910
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18248 8498 18276 9064
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18248 7478 18276 7686
rect 18340 7546 18368 7686
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18236 7472 18288 7478
rect 18524 7426 18552 9522
rect 19076 8974 19104 9522
rect 19536 9178 19564 9522
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 18616 8362 18644 8910
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19260 8498 19288 8774
rect 19352 8634 19380 9114
rect 19628 9042 19656 9862
rect 19812 9654 19840 9998
rect 19901 9820 20209 9840
rect 19901 9818 19907 9820
rect 19963 9818 19987 9820
rect 20043 9818 20067 9820
rect 20123 9818 20147 9820
rect 20203 9818 20209 9820
rect 19963 9766 19965 9818
rect 20145 9766 20147 9818
rect 19901 9764 19907 9766
rect 19963 9764 19987 9766
rect 20043 9764 20067 9766
rect 20123 9764 20147 9766
rect 20203 9764 20209 9766
rect 19901 9744 20209 9764
rect 19800 9648 19852 9654
rect 19984 9648 20036 9654
rect 19800 9590 19852 9596
rect 19904 9608 19984 9636
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19628 8430 19656 8978
rect 19904 8956 19932 9608
rect 19984 9590 20036 9596
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 20168 9376 20220 9382
rect 20272 9330 20300 9590
rect 20220 9324 20300 9330
rect 20168 9318 20300 9324
rect 20180 9302 20300 9318
rect 19812 8928 19932 8956
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19720 8498 19748 8774
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18616 8265 18644 8298
rect 18602 8256 18658 8265
rect 18602 8191 18658 8200
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18236 7414 18288 7420
rect 18340 7398 18552 7426
rect 18788 7404 18840 7410
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 6798 18184 7278
rect 18340 7274 18368 7398
rect 18788 7346 18840 7352
rect 18328 7268 18380 7274
rect 18328 7210 18380 7216
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18340 5778 18368 7210
rect 18800 7002 18828 7346
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 19076 6934 19104 7822
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19536 7410 19564 7482
rect 19628 7426 19656 8366
rect 19524 7404 19576 7410
rect 19628 7398 19748 7426
rect 19812 7410 19840 8928
rect 19901 8732 20209 8752
rect 19901 8730 19907 8732
rect 19963 8730 19987 8732
rect 20043 8730 20067 8732
rect 20123 8730 20147 8732
rect 20203 8730 20209 8732
rect 19963 8678 19965 8730
rect 20145 8678 20147 8730
rect 19901 8676 19907 8678
rect 19963 8676 19987 8678
rect 20043 8676 20067 8678
rect 20123 8676 20147 8678
rect 20203 8676 20209 8678
rect 19901 8656 20209 8676
rect 20272 8498 20300 9302
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 19901 7644 20209 7664
rect 19901 7642 19907 7644
rect 19963 7642 19987 7644
rect 20043 7642 20067 7644
rect 20123 7642 20147 7644
rect 20203 7642 20209 7644
rect 19963 7590 19965 7642
rect 20145 7590 20147 7642
rect 19901 7588 19907 7590
rect 19963 7588 19987 7590
rect 20043 7588 20067 7590
rect 20123 7588 20147 7590
rect 20203 7588 20209 7590
rect 19901 7568 20209 7588
rect 20272 7546 20300 8434
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 19524 7346 19576 7352
rect 19720 7342 19748 7398
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19432 7268 19484 7274
rect 19432 7210 19484 7216
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 18696 6724 18748 6730
rect 18696 6666 18748 6672
rect 18708 6458 18736 6666
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18708 5710 18736 6054
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18248 5574 18276 5646
rect 18800 5574 18828 6326
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18788 5568 18840 5574
rect 18788 5510 18840 5516
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4826 18092 4966
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18156 4282 18184 4558
rect 18800 4282 18828 5510
rect 19248 5364 19300 5370
rect 19352 5352 19380 5714
rect 19300 5324 19380 5352
rect 19248 5306 19300 5312
rect 19444 5302 19472 7210
rect 19720 7002 19748 7278
rect 19812 7002 19840 7346
rect 19708 6996 19760 7002
rect 19708 6938 19760 6944
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19901 6556 20209 6576
rect 19901 6554 19907 6556
rect 19963 6554 19987 6556
rect 20043 6554 20067 6556
rect 20123 6554 20147 6556
rect 20203 6554 20209 6556
rect 19963 6502 19965 6554
rect 20145 6502 20147 6554
rect 19901 6500 19907 6502
rect 19963 6500 19987 6502
rect 20043 6500 20067 6502
rect 20123 6500 20147 6502
rect 20203 6500 20209 6502
rect 19901 6480 20209 6500
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19536 5692 19564 6258
rect 19720 5902 20024 5930
rect 19720 5846 19748 5902
rect 19708 5840 19760 5846
rect 19892 5840 19944 5846
rect 19708 5782 19760 5788
rect 19812 5788 19892 5794
rect 19812 5782 19944 5788
rect 19812 5766 19932 5782
rect 19616 5704 19668 5710
rect 19536 5664 19616 5692
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19432 5160 19484 5166
rect 19536 5114 19564 5664
rect 19616 5646 19668 5652
rect 19708 5636 19760 5642
rect 19708 5578 19760 5584
rect 19720 5302 19748 5578
rect 19812 5574 19840 5766
rect 19996 5710 20024 5902
rect 20364 5846 20392 8570
rect 20456 7410 20484 9998
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20548 8634 20576 9522
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20640 7290 20668 10798
rect 20732 9654 20760 10934
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20732 9178 20760 9454
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20824 9058 20852 9522
rect 20732 9030 20852 9058
rect 20732 8906 20760 9030
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20456 7262 20668 7290
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 19984 5704 20036 5710
rect 20456 5692 20484 7262
rect 20732 6780 20760 8842
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20824 7750 20852 8434
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20824 7478 20852 7686
rect 20916 7562 20944 16390
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21100 15026 21128 15846
rect 21192 15162 21220 16050
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 21100 14929 21128 14962
rect 21086 14920 21142 14929
rect 21086 14855 21142 14864
rect 21192 14822 21220 15098
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21192 14074 21220 14758
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21192 12238 21220 12582
rect 21284 12306 21312 17054
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21560 16658 21588 16934
rect 21652 16776 21680 17206
rect 21732 16788 21784 16794
rect 21652 16748 21732 16776
rect 21732 16730 21784 16736
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21548 15700 21600 15706
rect 21548 15642 21600 15648
rect 21560 15162 21588 15642
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21928 15026 21956 17274
rect 22112 16998 22140 17478
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22112 15065 22140 16934
rect 22204 16250 22232 19332
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22388 18698 22416 19110
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 22480 18578 22508 19722
rect 22572 19242 22600 20334
rect 22664 19334 22692 20726
rect 22756 19854 22784 25842
rect 23032 25498 23060 26250
rect 23388 26240 23440 26246
rect 23388 26182 23440 26188
rect 23400 25906 23428 26182
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23492 25498 23520 26386
rect 24492 26376 24544 26382
rect 24492 26318 24544 26324
rect 24400 26240 24452 26246
rect 24400 26182 24452 26188
rect 24412 25974 24440 26182
rect 24400 25968 24452 25974
rect 24400 25910 24452 25916
rect 24504 25498 24532 26318
rect 25148 26234 25176 32056
rect 26344 28422 26372 32056
rect 27342 31991 27398 32000
rect 26882 30696 26938 30705
rect 26882 30631 26938 30640
rect 26332 28416 26384 28422
rect 26332 28358 26384 28364
rect 25148 26206 25452 26234
rect 24639 25596 24947 25616
rect 24639 25594 24645 25596
rect 24701 25594 24725 25596
rect 24781 25594 24805 25596
rect 24861 25594 24885 25596
rect 24941 25594 24947 25596
rect 24701 25542 24703 25594
rect 24883 25542 24885 25594
rect 24639 25540 24645 25542
rect 24701 25540 24725 25542
rect 24781 25540 24805 25542
rect 24861 25540 24885 25542
rect 24941 25540 24947 25542
rect 24639 25520 24947 25540
rect 23020 25492 23072 25498
rect 23020 25434 23072 25440
rect 23480 25492 23532 25498
rect 23480 25434 23532 25440
rect 24492 25492 24544 25498
rect 24492 25434 24544 25440
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24412 24818 24440 25230
rect 24400 24812 24452 24818
rect 24400 24754 24452 24760
rect 24492 24744 24544 24750
rect 24492 24686 24544 24692
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23664 24268 23716 24274
rect 23664 24210 23716 24216
rect 23676 23866 23704 24210
rect 23768 24206 23796 24550
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 24032 24132 24084 24138
rect 24032 24074 24084 24080
rect 23664 23860 23716 23866
rect 23664 23802 23716 23808
rect 23020 23724 23072 23730
rect 23020 23666 23072 23672
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22848 22030 22876 23598
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 23032 21962 23060 23666
rect 23676 23662 23704 23802
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 23664 23656 23716 23662
rect 23664 23598 23716 23604
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 23204 22568 23256 22574
rect 23204 22510 23256 22516
rect 23216 22030 23244 22510
rect 23308 22098 23336 22578
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23020 21956 23072 21962
rect 23020 21898 23072 21904
rect 23032 21622 23060 21898
rect 23020 21616 23072 21622
rect 23020 21558 23072 21564
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 22848 20602 22876 21490
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 23112 20528 23164 20534
rect 23112 20470 23164 20476
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 23032 20058 23060 20402
rect 23124 20262 23152 20470
rect 23216 20330 23244 21966
rect 23308 21146 23336 22034
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23308 20466 23336 21082
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23400 20330 23428 20810
rect 23492 20602 23520 23598
rect 23676 22642 23704 23598
rect 23664 22636 23716 22642
rect 23664 22578 23716 22584
rect 23940 22568 23992 22574
rect 23940 22510 23992 22516
rect 23952 22234 23980 22510
rect 24044 22438 24072 24074
rect 24504 23866 24532 24686
rect 25320 24608 25372 24614
rect 25320 24550 25372 24556
rect 24639 24508 24947 24528
rect 24639 24506 24645 24508
rect 24701 24506 24725 24508
rect 24781 24506 24805 24508
rect 24861 24506 24885 24508
rect 24941 24506 24947 24508
rect 24701 24454 24703 24506
rect 24883 24454 24885 24506
rect 24639 24452 24645 24454
rect 24701 24452 24725 24454
rect 24781 24452 24805 24454
rect 24861 24452 24885 24454
rect 24941 24452 24947 24454
rect 24639 24432 24947 24452
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 24492 23860 24544 23866
rect 24492 23802 24544 23808
rect 25240 23798 25268 24210
rect 25332 24138 25360 24550
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 24860 23792 24912 23798
rect 25228 23792 25280 23798
rect 24912 23740 25084 23746
rect 24860 23734 25084 23740
rect 25228 23734 25280 23740
rect 24124 23724 24176 23730
rect 24872 23718 25084 23734
rect 24124 23666 24176 23672
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23754 20904 23810 20913
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23676 20369 23704 20878
rect 23754 20839 23810 20848
rect 23768 20466 23796 20839
rect 23848 20800 23900 20806
rect 23848 20742 23900 20748
rect 23860 20466 23888 20742
rect 23756 20460 23808 20466
rect 23756 20402 23808 20408
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23662 20360 23718 20369
rect 23204 20324 23256 20330
rect 23204 20266 23256 20272
rect 23388 20324 23440 20330
rect 23662 20295 23718 20304
rect 23388 20266 23440 20272
rect 23860 20262 23888 20402
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22744 19372 22796 19378
rect 22664 19320 22744 19334
rect 22928 19372 22980 19378
rect 22664 19314 22796 19320
rect 22848 19320 22928 19334
rect 22848 19314 22980 19320
rect 22664 19306 22784 19314
rect 22848 19306 22968 19314
rect 22560 19236 22612 19242
rect 22560 19178 22612 19184
rect 22388 18550 22508 18578
rect 22388 17610 22416 18550
rect 22376 17604 22428 17610
rect 22376 17546 22428 17552
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22098 15056 22154 15065
rect 21916 15020 21968 15026
rect 22098 14991 22154 15000
rect 21916 14962 21968 14968
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21376 14414 21404 14758
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21560 13258 21588 14214
rect 21928 13433 21956 14962
rect 22204 14550 22232 16186
rect 22284 16108 22336 16114
rect 22284 16050 22336 16056
rect 22296 15026 22324 16050
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22296 14618 22324 14826
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22388 14074 22416 17546
rect 22664 17338 22692 19306
rect 22848 17746 22876 19306
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22560 16992 22612 16998
rect 22612 16940 22692 16946
rect 22560 16934 22692 16940
rect 22572 16918 22692 16934
rect 22664 16658 22692 16918
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22664 16250 22692 16594
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22664 16114 22692 16186
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 22664 15706 22692 16050
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22848 15570 22968 15586
rect 22836 15564 22968 15570
rect 22888 15558 22968 15564
rect 22836 15506 22888 15512
rect 22940 15434 22968 15558
rect 22836 15428 22888 15434
rect 22836 15370 22888 15376
rect 22928 15428 22980 15434
rect 22928 15370 22980 15376
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22572 14929 22600 14962
rect 22558 14920 22614 14929
rect 22848 14890 22876 15370
rect 22558 14855 22614 14864
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22664 13870 22692 14214
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22296 13530 22324 13806
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 21914 13424 21970 13433
rect 21914 13359 21970 13368
rect 21548 13252 21600 13258
rect 21548 13194 21600 13200
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22388 12442 22416 12786
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 21192 11830 21220 12174
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21468 11898 21496 12106
rect 21652 11898 21680 12174
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21180 11824 21232 11830
rect 21180 11766 21232 11772
rect 21192 11642 21220 11766
rect 22204 11762 22232 12174
rect 22388 11778 22416 12378
rect 22480 12238 22508 12582
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22388 11762 22600 11778
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22388 11756 22612 11762
rect 22388 11750 22560 11756
rect 21100 11614 21220 11642
rect 22296 11626 22324 11698
rect 22284 11620 22336 11626
rect 20996 11144 21048 11150
rect 21100 11132 21128 11614
rect 22284 11562 22336 11568
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 21048 11104 21128 11132
rect 21192 11336 21220 11494
rect 22296 11354 22324 11562
rect 22284 11348 22336 11354
rect 21192 11308 21404 11336
rect 20996 11086 21048 11092
rect 21192 10674 21220 11308
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 21284 10538 21312 11154
rect 21376 11150 21404 11308
rect 22284 11290 22336 11296
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 22388 11082 22416 11750
rect 22560 11698 22612 11704
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21376 10062 21404 10950
rect 21468 10674 21496 11018
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21560 10130 21588 10406
rect 21652 10198 21680 10406
rect 21640 10192 21692 10198
rect 21640 10134 21692 10140
rect 22388 10130 22416 10610
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22296 9654 22324 9862
rect 22284 9648 22336 9654
rect 22284 9590 22336 9596
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 21916 9444 21968 9450
rect 21836 9404 21916 9432
rect 21548 9104 21600 9110
rect 21548 9046 21600 9052
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21100 8294 21128 8774
rect 21560 8498 21588 9046
rect 21836 8906 21864 9404
rect 21916 9386 21968 9392
rect 22020 9330 22048 9454
rect 21928 9302 22048 9330
rect 21928 9042 21956 9302
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 21284 7954 21312 8230
rect 21836 8090 21864 8842
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21928 7970 21956 8978
rect 22204 8906 22232 9522
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22192 8900 22244 8906
rect 22192 8842 22244 8848
rect 22388 8634 22416 8910
rect 22572 8838 22600 9522
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22572 8498 22600 8774
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 21272 7948 21324 7954
rect 21272 7890 21324 7896
rect 21836 7942 21956 7970
rect 21284 7834 21312 7890
rect 21192 7818 21312 7834
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 21180 7812 21312 7818
rect 21232 7806 21312 7812
rect 21180 7754 21232 7760
rect 20916 7534 21036 7562
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20904 6792 20956 6798
rect 20732 6752 20904 6780
rect 20904 6734 20956 6740
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20640 5914 20668 6598
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 19984 5646 20036 5652
rect 20364 5664 20484 5692
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19901 5468 20209 5488
rect 19901 5466 19907 5468
rect 19963 5466 19987 5468
rect 20043 5466 20067 5468
rect 20123 5466 20147 5468
rect 20203 5466 20209 5468
rect 19963 5414 19965 5466
rect 20145 5414 20147 5466
rect 19901 5412 19907 5414
rect 19963 5412 19987 5414
rect 20043 5412 20067 5414
rect 20123 5412 20147 5414
rect 20203 5412 20209 5414
rect 19901 5392 20209 5412
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 19484 5108 19564 5114
rect 19432 5102 19564 5108
rect 19444 5086 19564 5102
rect 19706 5128 19762 5137
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18052 4208 18104 4214
rect 18512 4208 18564 4214
rect 18052 4150 18104 4156
rect 18326 4176 18382 4185
rect 18064 3398 18092 4150
rect 18512 4150 18564 4156
rect 18326 4111 18328 4120
rect 18380 4111 18382 4120
rect 18328 4082 18380 4088
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18156 3942 18184 4014
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18524 3466 18552 4150
rect 18878 3768 18934 3777
rect 18878 3703 18880 3712
rect 18932 3703 18934 3712
rect 18880 3674 18932 3680
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18788 3596 18840 3602
rect 18788 3538 18840 3544
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18512 3460 18564 3466
rect 18512 3402 18564 3408
rect 18052 3392 18104 3398
rect 18616 3346 18644 3470
rect 18708 3398 18736 3470
rect 18104 3340 18644 3346
rect 18052 3334 18644 3340
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 17880 2746 18000 2774
rect 18064 3318 18644 3334
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 17880 800 17908 2746
rect 18064 2650 18092 3318
rect 18800 3194 18828 3538
rect 18878 3360 18934 3369
rect 18878 3295 18934 3304
rect 18892 3194 18920 3295
rect 18984 3233 19012 3606
rect 18970 3224 19026 3233
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18880 3188 18932 3194
rect 18970 3159 19026 3168
rect 18880 3130 18932 3136
rect 18248 2990 18276 3130
rect 19076 3058 19104 4966
rect 19444 3738 19472 5086
rect 19706 5063 19762 5072
rect 19614 4040 19670 4049
rect 19614 3975 19670 3984
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 18236 2984 18288 2990
rect 18236 2926 18288 2932
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 19628 800 19656 3975
rect 19720 3126 19748 5063
rect 19800 5024 19852 5030
rect 19800 4966 19852 4972
rect 19812 4214 19840 4966
rect 20364 4758 20392 5664
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20456 5166 20484 5510
rect 20548 5370 20576 5714
rect 20640 5710 20668 5850
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20904 5704 20956 5710
rect 20904 5646 20956 5652
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20824 5234 20852 5578
rect 20916 5370 20944 5646
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20352 4752 20404 4758
rect 20352 4694 20404 4700
rect 19901 4380 20209 4400
rect 19901 4378 19907 4380
rect 19963 4378 19987 4380
rect 20043 4378 20067 4380
rect 20123 4378 20147 4380
rect 20203 4378 20209 4380
rect 19963 4326 19965 4378
rect 20145 4326 20147 4378
rect 19901 4324 19907 4326
rect 19963 4324 19987 4326
rect 20043 4324 20067 4326
rect 20123 4324 20147 4326
rect 20203 4324 20209 4326
rect 19901 4304 20209 4324
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20548 3602 20576 3878
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 20260 3460 20312 3466
rect 20260 3402 20312 3408
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 19901 3292 20209 3312
rect 19901 3290 19907 3292
rect 19963 3290 19987 3292
rect 20043 3290 20067 3292
rect 20123 3290 20147 3292
rect 20203 3290 20209 3292
rect 19963 3238 19965 3290
rect 20145 3238 20147 3290
rect 19901 3236 19907 3238
rect 19963 3236 19987 3238
rect 20043 3236 20067 3238
rect 20123 3236 20147 3238
rect 20203 3236 20209 3238
rect 19901 3216 20209 3236
rect 20272 3194 20300 3402
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 20260 3188 20312 3194
rect 20260 3130 20312 3136
rect 19708 3120 19760 3126
rect 19708 3062 19760 3068
rect 19812 2854 19840 3130
rect 20456 3126 20484 3334
rect 20444 3120 20496 3126
rect 20444 3062 20496 3068
rect 20640 3058 20668 3402
rect 20824 3126 20852 3946
rect 20812 3120 20864 3126
rect 20812 3062 20864 3068
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19901 2204 20209 2224
rect 19901 2202 19907 2204
rect 19963 2202 19987 2204
rect 20043 2202 20067 2204
rect 20123 2202 20147 2204
rect 20203 2202 20209 2204
rect 19963 2150 19965 2202
rect 20145 2150 20147 2202
rect 19901 2148 19907 2150
rect 19963 2148 19987 2150
rect 20043 2148 20067 2150
rect 20123 2148 20147 2150
rect 20203 2148 20209 2150
rect 19901 2128 20209 2148
rect 5552 734 5856 762
rect 5906 0 5962 800
rect 7654 0 7710 800
rect 9310 0 9366 800
rect 11058 0 11114 800
rect 12714 0 12770 800
rect 14462 0 14518 800
rect 16210 0 16266 800
rect 17866 0 17922 800
rect 19614 0 19670 800
rect 21008 762 21036 7534
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 21100 7002 21128 7278
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 21192 5710 21220 7210
rect 21284 6798 21312 7806
rect 21376 7410 21404 7822
rect 21364 7404 21416 7410
rect 21364 7346 21416 7352
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21376 6866 21404 7346
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21560 6798 21588 7346
rect 21836 6866 21864 7942
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 21928 6882 21956 7142
rect 22664 6914 22692 13806
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22756 12374 22784 13126
rect 23124 12434 23152 20198
rect 23388 19984 23440 19990
rect 23388 19926 23440 19932
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 23308 19825 23336 19858
rect 23294 19816 23350 19825
rect 23294 19751 23350 19760
rect 23308 19378 23336 19751
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23400 19258 23428 19926
rect 23480 19508 23532 19514
rect 23480 19450 23532 19456
rect 23308 19230 23428 19258
rect 23308 18306 23336 19230
rect 23492 19174 23520 19450
rect 23664 19372 23716 19378
rect 23716 19320 23796 19334
rect 23664 19314 23796 19320
rect 23676 19306 23796 19314
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23400 18902 23428 19110
rect 23388 18896 23440 18902
rect 23388 18838 23440 18844
rect 23676 18766 23704 19110
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23400 18426 23428 18634
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23308 18278 23428 18306
rect 23400 17678 23428 18278
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23308 17270 23336 17478
rect 23296 17264 23348 17270
rect 23296 17206 23348 17212
rect 23400 15586 23428 17614
rect 23492 17610 23520 18158
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23480 17604 23532 17610
rect 23480 17546 23532 17552
rect 23584 17134 23612 17750
rect 23676 17746 23704 18702
rect 23768 18630 23796 19306
rect 23756 18624 23808 18630
rect 23756 18566 23808 18572
rect 23768 18290 23796 18566
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 23860 17626 23888 20198
rect 24044 19174 24072 21830
rect 24136 21146 24164 23666
rect 24639 23420 24947 23440
rect 24639 23418 24645 23420
rect 24701 23418 24725 23420
rect 24781 23418 24805 23420
rect 24861 23418 24885 23420
rect 24941 23418 24947 23420
rect 24701 23366 24703 23418
rect 24883 23366 24885 23418
rect 24639 23364 24645 23366
rect 24701 23364 24725 23366
rect 24781 23364 24805 23366
rect 24861 23364 24885 23366
rect 24941 23364 24947 23366
rect 24639 23344 24947 23364
rect 24308 23248 24360 23254
rect 24308 23190 24360 23196
rect 24320 21894 24348 23190
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24504 22234 24532 23054
rect 25056 23050 25084 23718
rect 25044 23044 25096 23050
rect 25044 22986 25096 22992
rect 24676 22976 24728 22982
rect 24676 22918 24728 22924
rect 24688 22710 24716 22918
rect 24676 22704 24728 22710
rect 24676 22646 24728 22652
rect 25424 22574 25452 26206
rect 26698 24712 26754 24721
rect 26698 24647 26754 24656
rect 25872 24608 25924 24614
rect 25872 24550 25924 24556
rect 25596 24064 25648 24070
rect 25596 24006 25648 24012
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25516 22710 25544 22918
rect 25504 22704 25556 22710
rect 25504 22646 25556 22652
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 24639 22332 24947 22352
rect 24639 22330 24645 22332
rect 24701 22330 24725 22332
rect 24781 22330 24805 22332
rect 24861 22330 24885 22332
rect 24941 22330 24947 22332
rect 24701 22278 24703 22330
rect 24883 22278 24885 22330
rect 24639 22276 24645 22278
rect 24701 22276 24725 22278
rect 24781 22276 24805 22278
rect 24861 22276 24885 22278
rect 24941 22276 24947 22278
rect 24639 22256 24947 22276
rect 24492 22228 24544 22234
rect 24492 22170 24544 22176
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 24308 21888 24360 21894
rect 24308 21830 24360 21836
rect 24504 21554 24532 21966
rect 25424 21962 25452 22510
rect 25516 22166 25544 22646
rect 25608 22642 25636 24006
rect 25884 23798 25912 24550
rect 26148 24404 26200 24410
rect 26148 24346 26200 24352
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 25872 23792 25924 23798
rect 25872 23734 25924 23740
rect 25688 23248 25740 23254
rect 25688 23190 25740 23196
rect 25700 23050 25728 23190
rect 25688 23044 25740 23050
rect 25688 22986 25740 22992
rect 25700 22642 25728 22986
rect 26068 22642 26096 24142
rect 26160 24070 26188 24346
rect 26712 24206 26740 24647
rect 26896 24410 26924 30631
rect 27356 26234 27384 31991
rect 27540 30258 27568 32056
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 27434 29200 27490 29209
rect 27434 29135 27490 29144
rect 27448 27334 27476 29135
rect 28828 29034 28856 32056
rect 28816 29028 28868 29034
rect 28816 28970 28868 28976
rect 30024 28966 30052 32056
rect 30012 28960 30064 28966
rect 30012 28902 30064 28908
rect 27526 27704 27582 27713
rect 27526 27639 27582 27648
rect 27436 27328 27488 27334
rect 27436 27270 27488 27276
rect 27540 27130 27568 27639
rect 27528 27124 27580 27130
rect 27528 27066 27580 27072
rect 27356 26206 27476 26234
rect 27448 24410 27476 26206
rect 27526 26208 27582 26217
rect 27526 26143 27582 26152
rect 27540 26042 27568 26143
rect 27528 26036 27580 26042
rect 27528 25978 27580 25984
rect 26884 24404 26936 24410
rect 26884 24346 26936 24352
rect 27436 24404 27488 24410
rect 27436 24346 27488 24352
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 26160 22778 26188 24006
rect 26608 23724 26660 23730
rect 26608 23666 26660 23672
rect 26620 23118 26648 23666
rect 26712 23662 26740 24142
rect 26792 24132 26844 24138
rect 26792 24074 26844 24080
rect 26700 23656 26752 23662
rect 26700 23598 26752 23604
rect 26804 23526 26832 24074
rect 27068 24064 27120 24070
rect 26988 24024 27068 24052
rect 26988 23798 27016 24024
rect 27068 24006 27120 24012
rect 27356 23866 27384 24142
rect 27448 23866 27476 24346
rect 27620 24132 27672 24138
rect 27620 24074 27672 24080
rect 28632 24132 28684 24138
rect 28632 24074 28684 24080
rect 27344 23860 27396 23866
rect 27344 23802 27396 23808
rect 27436 23860 27488 23866
rect 27436 23802 27488 23808
rect 26976 23792 27028 23798
rect 26976 23734 27028 23740
rect 26792 23520 26844 23526
rect 26792 23462 26844 23468
rect 26988 23254 27016 23734
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 26976 23248 27028 23254
rect 26976 23190 27028 23196
rect 27172 23118 27200 23598
rect 27252 23520 27304 23526
rect 27252 23462 27304 23468
rect 26608 23112 26660 23118
rect 26608 23054 26660 23060
rect 27160 23112 27212 23118
rect 27160 23054 27212 23060
rect 27264 23066 27292 23462
rect 27356 23186 27384 23802
rect 27632 23594 27660 24074
rect 28644 23866 28672 24074
rect 28632 23860 28684 23866
rect 28632 23802 28684 23808
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 27620 23588 27672 23594
rect 27620 23530 27672 23536
rect 28184 23526 28212 23666
rect 28172 23520 28224 23526
rect 28172 23462 28224 23468
rect 27436 23316 27488 23322
rect 27436 23258 27488 23264
rect 27448 23225 27476 23258
rect 27434 23216 27490 23225
rect 27344 23180 27396 23186
rect 27434 23151 27490 23160
rect 27344 23122 27396 23128
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 25688 22636 25740 22642
rect 25688 22578 25740 22584
rect 26056 22636 26108 22642
rect 26056 22578 26108 22584
rect 26516 22636 26568 22642
rect 26516 22578 26568 22584
rect 25504 22160 25556 22166
rect 25504 22102 25556 22108
rect 25412 21956 25464 21962
rect 25412 21898 25464 21904
rect 25608 21622 25636 22578
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 24124 21140 24176 21146
rect 24124 21082 24176 21088
rect 24228 21078 24256 21490
rect 24308 21412 24360 21418
rect 24308 21354 24360 21360
rect 24216 21072 24268 21078
rect 24216 21014 24268 21020
rect 24320 21010 24348 21354
rect 24504 21350 24532 21490
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 25044 21344 25096 21350
rect 25044 21286 25096 21292
rect 24400 21140 24452 21146
rect 24400 21082 24452 21088
rect 24308 21004 24360 21010
rect 24308 20946 24360 20952
rect 24320 19378 24348 20946
rect 24412 20874 24440 21082
rect 24400 20868 24452 20874
rect 24400 20810 24452 20816
rect 24504 20602 24532 21286
rect 24639 21244 24947 21264
rect 24639 21242 24645 21244
rect 24701 21242 24725 21244
rect 24781 21242 24805 21244
rect 24861 21242 24885 21244
rect 24941 21242 24947 21244
rect 24701 21190 24703 21242
rect 24883 21190 24885 21242
rect 24639 21188 24645 21190
rect 24701 21188 24725 21190
rect 24781 21188 24805 21190
rect 24861 21188 24885 21190
rect 24941 21188 24947 21190
rect 24639 21168 24947 21188
rect 24952 20868 25004 20874
rect 24952 20810 25004 20816
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24492 20596 24544 20602
rect 24492 20538 24544 20544
rect 24596 20330 24624 20742
rect 24964 20602 24992 20810
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 25056 20466 25084 21286
rect 25608 20466 25636 21558
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 25596 20460 25648 20466
rect 25596 20402 25648 20408
rect 25320 20392 25372 20398
rect 25320 20334 25372 20340
rect 24584 20324 24636 20330
rect 24584 20266 24636 20272
rect 24639 20156 24947 20176
rect 24639 20154 24645 20156
rect 24701 20154 24725 20156
rect 24781 20154 24805 20156
rect 24861 20154 24885 20156
rect 24941 20154 24947 20156
rect 24701 20102 24703 20154
rect 24883 20102 24885 20154
rect 24639 20100 24645 20102
rect 24701 20100 24725 20102
rect 24781 20100 24805 20102
rect 24861 20100 24885 20102
rect 24941 20100 24947 20102
rect 24639 20080 24947 20100
rect 25332 20058 25360 20334
rect 25596 20324 25648 20330
rect 25596 20266 25648 20272
rect 25608 20058 25636 20266
rect 25320 20052 25372 20058
rect 25320 19994 25372 20000
rect 25596 20052 25648 20058
rect 25596 19994 25648 20000
rect 25044 19848 25096 19854
rect 25042 19816 25044 19825
rect 25096 19816 25098 19825
rect 25042 19751 25098 19760
rect 25136 19712 25188 19718
rect 25136 19654 25188 19660
rect 24308 19372 24360 19378
rect 24308 19314 24360 19320
rect 24032 19168 24084 19174
rect 24032 19110 24084 19116
rect 24044 18358 24072 19110
rect 24320 18834 24348 19314
rect 24639 19068 24947 19088
rect 24639 19066 24645 19068
rect 24701 19066 24725 19068
rect 24781 19066 24805 19068
rect 24861 19066 24885 19068
rect 24941 19066 24947 19068
rect 24701 19014 24703 19066
rect 24883 19014 24885 19066
rect 24639 19012 24645 19014
rect 24701 19012 24725 19014
rect 24781 19012 24805 19014
rect 24861 19012 24885 19014
rect 24941 19012 24947 19014
rect 24639 18992 24947 19012
rect 25148 18834 25176 19654
rect 25228 19440 25280 19446
rect 25228 19382 25280 19388
rect 25240 18970 25268 19382
rect 25228 18964 25280 18970
rect 25228 18906 25280 18912
rect 24308 18828 24360 18834
rect 24308 18770 24360 18776
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 24320 18426 24348 18770
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24400 18692 24452 18698
rect 24400 18634 24452 18640
rect 24308 18420 24360 18426
rect 24308 18362 24360 18368
rect 24032 18352 24084 18358
rect 24032 18294 24084 18300
rect 24412 17678 24440 18634
rect 24504 18290 24532 18702
rect 24492 18284 24544 18290
rect 24492 18226 24544 18232
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 24639 17980 24947 18000
rect 24639 17978 24645 17980
rect 24701 17978 24725 17980
rect 24781 17978 24805 17980
rect 24861 17978 24885 17980
rect 24941 17978 24947 17980
rect 24701 17926 24703 17978
rect 24883 17926 24885 17978
rect 24639 17924 24645 17926
rect 24701 17924 24725 17926
rect 24781 17924 24805 17926
rect 24861 17924 24885 17926
rect 24941 17924 24947 17926
rect 24639 17904 24947 17924
rect 24492 17876 24544 17882
rect 24492 17818 24544 17824
rect 23676 17598 23888 17626
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 23400 15558 23520 15586
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23400 15162 23428 15438
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23492 14958 23520 15558
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23584 15026 23612 15438
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23480 14952 23532 14958
rect 23480 14894 23532 14900
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 23308 13190 23336 14350
rect 23492 13326 23520 14894
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23584 13326 23612 14350
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23572 13320 23624 13326
rect 23572 13262 23624 13268
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12782 23336 13126
rect 23296 12776 23348 12782
rect 23296 12718 23348 12724
rect 23124 12406 23244 12434
rect 22744 12368 22796 12374
rect 22744 12310 22796 12316
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22756 10062 22784 10950
rect 23032 10130 23060 11494
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 23124 10810 23152 11086
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22756 9042 22784 9318
rect 23124 9178 23152 9522
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 22756 8242 22784 8978
rect 22928 8492 22980 8498
rect 22928 8434 22980 8440
rect 22836 8288 22888 8294
rect 22756 8236 22836 8242
rect 22756 8230 22888 8236
rect 22756 8214 22876 8230
rect 22848 8090 22876 8214
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22756 7546 22784 7822
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22848 7342 22876 8026
rect 22940 7410 22968 8434
rect 23124 8362 23152 8978
rect 23112 8356 23164 8362
rect 23112 8298 23164 8304
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 22664 6886 22784 6914
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 21928 6854 22140 6882
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21284 6322 21312 6734
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21560 5710 21588 6734
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21100 3534 21128 5510
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21192 4826 21220 5170
rect 21376 5166 21404 5510
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21560 4826 21588 5646
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21376 4282 21404 4558
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21744 2922 21772 6394
rect 21836 5166 21864 6802
rect 21928 5574 21956 6854
rect 22112 6798 22140 6854
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 22480 6118 22508 6734
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 21916 5568 21968 5574
rect 21916 5510 21968 5516
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 22020 5098 22048 6054
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 22112 5302 22140 5646
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22388 5370 22416 5510
rect 22376 5364 22428 5370
rect 22376 5306 22428 5312
rect 22100 5296 22152 5302
rect 22100 5238 22152 5244
rect 22008 5092 22060 5098
rect 22008 5034 22060 5040
rect 22376 4684 22428 4690
rect 22376 4626 22428 4632
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 22112 3738 22140 4150
rect 22296 3738 22324 4422
rect 22388 4214 22416 4626
rect 22652 4548 22704 4554
rect 22652 4490 22704 4496
rect 22376 4208 22428 4214
rect 22376 4150 22428 4156
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 22284 3732 22336 3738
rect 22284 3674 22336 3680
rect 22664 3534 22692 4490
rect 22376 3528 22428 3534
rect 22376 3470 22428 3476
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22020 3126 22048 3334
rect 21824 3120 21876 3126
rect 21824 3062 21876 3068
rect 22008 3120 22060 3126
rect 22008 3062 22060 3068
rect 21836 2972 21864 3062
rect 22204 3058 22232 3402
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22388 2990 22416 3470
rect 22664 3194 22692 3470
rect 22756 3398 22784 6886
rect 22940 5642 22968 7346
rect 23032 7002 23060 7346
rect 23020 6996 23072 7002
rect 23020 6938 23072 6944
rect 23124 6866 23152 8298
rect 23112 6860 23164 6866
rect 23112 6802 23164 6808
rect 23124 5914 23152 6802
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23216 5794 23244 12406
rect 23676 10962 23704 17598
rect 24504 17338 24532 17818
rect 25056 17542 25084 18022
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 23756 16584 23808 16590
rect 23756 16526 23808 16532
rect 23768 15706 23796 16526
rect 23940 16448 23992 16454
rect 23940 16390 23992 16396
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 23952 16182 23980 16390
rect 23940 16176 23992 16182
rect 23940 16118 23992 16124
rect 23756 15700 23808 15706
rect 23756 15642 23808 15648
rect 24044 15502 24072 16390
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24032 15496 24084 15502
rect 24032 15438 24084 15444
rect 24320 15434 24348 16050
rect 24412 16046 24440 16934
rect 24504 16726 24532 17274
rect 24639 16892 24947 16912
rect 24639 16890 24645 16892
rect 24701 16890 24725 16892
rect 24781 16890 24805 16892
rect 24861 16890 24885 16892
rect 24941 16890 24947 16892
rect 24701 16838 24703 16890
rect 24883 16838 24885 16890
rect 24639 16836 24645 16838
rect 24701 16836 24725 16838
rect 24781 16836 24805 16838
rect 24861 16836 24885 16838
rect 24941 16836 24947 16838
rect 24639 16816 24947 16836
rect 24492 16720 24544 16726
rect 24492 16662 24544 16668
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 25056 16538 25084 17478
rect 25240 17270 25268 17478
rect 25228 17264 25280 17270
rect 25228 17206 25280 17212
rect 25504 16720 25556 16726
rect 25504 16662 25556 16668
rect 25320 16584 25372 16590
rect 24400 16040 24452 16046
rect 24400 15982 24452 15988
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24308 15428 24360 15434
rect 24308 15370 24360 15376
rect 24320 15026 24348 15370
rect 24412 15162 24440 15438
rect 24504 15366 24532 16526
rect 25056 16510 25176 16538
rect 25320 16526 25372 16532
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24964 15994 24992 16050
rect 24964 15966 25084 15994
rect 24639 15804 24947 15824
rect 24639 15802 24645 15804
rect 24701 15802 24725 15804
rect 24781 15802 24805 15804
rect 24861 15802 24885 15804
rect 24941 15802 24947 15804
rect 24701 15750 24703 15802
rect 24883 15750 24885 15802
rect 24639 15748 24645 15750
rect 24701 15748 24725 15750
rect 24781 15748 24805 15750
rect 24861 15748 24885 15750
rect 24941 15748 24947 15750
rect 24639 15728 24947 15748
rect 24492 15360 24544 15366
rect 24492 15302 24544 15308
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24492 14884 24544 14890
rect 24492 14826 24544 14832
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23756 14544 23808 14550
rect 23756 14486 23808 14492
rect 23848 14544 23900 14550
rect 23848 14486 23900 14492
rect 23768 14346 23796 14486
rect 23756 14340 23808 14346
rect 23756 14282 23808 14288
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23768 13326 23796 14010
rect 23860 13870 23888 14486
rect 23952 14414 23980 14758
rect 24504 14482 24532 14826
rect 24639 14716 24947 14736
rect 24639 14714 24645 14716
rect 24701 14714 24725 14716
rect 24781 14714 24805 14716
rect 24861 14714 24885 14716
rect 24941 14714 24947 14716
rect 24701 14662 24703 14714
rect 24883 14662 24885 14714
rect 24639 14660 24645 14662
rect 24701 14660 24725 14662
rect 24781 14660 24805 14662
rect 24861 14660 24885 14662
rect 24941 14660 24947 14662
rect 24639 14640 24947 14660
rect 25056 14550 25084 15966
rect 25044 14544 25096 14550
rect 25044 14486 25096 14492
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23860 11150 23888 13466
rect 23952 13326 23980 14350
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24952 14340 25004 14346
rect 24952 14282 25004 14288
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24412 13938 24440 14214
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24504 13530 24532 14282
rect 24964 14074 24992 14282
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 25056 13870 25084 14486
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 24639 13628 24947 13648
rect 24639 13626 24645 13628
rect 24701 13626 24725 13628
rect 24781 13626 24805 13628
rect 24861 13626 24885 13628
rect 24941 13626 24947 13628
rect 24701 13574 24703 13626
rect 24883 13574 24885 13626
rect 24639 13572 24645 13574
rect 24701 13572 24725 13574
rect 24781 13572 24805 13574
rect 24861 13572 24885 13574
rect 24941 13572 24947 13574
rect 24639 13552 24947 13572
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24950 13424 25006 13433
rect 25056 13394 25084 13806
rect 24950 13359 25006 13368
rect 25044 13388 25096 13394
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 24964 13258 24992 13359
rect 25044 13330 25096 13336
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24412 12918 24440 13126
rect 25056 12986 25084 13330
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 24400 12912 24452 12918
rect 24400 12854 24452 12860
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24504 12238 24532 12718
rect 24639 12540 24947 12560
rect 24639 12538 24645 12540
rect 24701 12538 24725 12540
rect 24781 12538 24805 12540
rect 24861 12538 24885 12540
rect 24941 12538 24947 12540
rect 24701 12486 24703 12538
rect 24883 12486 24885 12538
rect 24639 12484 24645 12486
rect 24701 12484 24725 12486
rect 24781 12484 24805 12486
rect 24861 12484 24885 12486
rect 24941 12484 24947 12486
rect 24639 12464 24947 12484
rect 25056 12306 25084 12922
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 24492 12232 24544 12238
rect 25148 12220 25176 16510
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 25240 15706 25268 15982
rect 25332 15910 25360 16526
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 25228 15700 25280 15706
rect 25228 15642 25280 15648
rect 25332 15502 25360 15846
rect 25424 15638 25452 15846
rect 25412 15632 25464 15638
rect 25412 15574 25464 15580
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25424 15434 25452 15574
rect 25516 15434 25544 16662
rect 25700 15706 25728 22578
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25976 21486 26004 21830
rect 26068 21706 26096 22578
rect 26148 22432 26200 22438
rect 26148 22374 26200 22380
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 26160 22234 26188 22374
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 26344 21962 26372 22374
rect 26332 21956 26384 21962
rect 26332 21898 26384 21904
rect 26528 21894 26556 22578
rect 26516 21888 26568 21894
rect 26516 21830 26568 21836
rect 26068 21678 26280 21706
rect 25964 21480 26016 21486
rect 25964 21422 26016 21428
rect 26068 20330 26096 21678
rect 26252 21622 26280 21678
rect 26240 21616 26292 21622
rect 26240 21558 26292 21564
rect 26240 21480 26292 21486
rect 26240 21422 26292 21428
rect 26252 21010 26280 21422
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26240 21004 26292 21010
rect 26240 20946 26292 20952
rect 26344 20992 26372 21286
rect 26620 21146 26648 23054
rect 26792 23044 26844 23050
rect 26792 22986 26844 22992
rect 26608 21140 26660 21146
rect 26608 21082 26660 21088
rect 26424 21004 26476 21010
rect 26344 20964 26424 20992
rect 26056 20324 26108 20330
rect 26056 20266 26108 20272
rect 26252 19922 26280 20946
rect 26344 20058 26372 20964
rect 26424 20946 26476 20952
rect 26516 20936 26568 20942
rect 26516 20878 26568 20884
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 26436 20466 26464 20742
rect 26528 20466 26556 20878
rect 26424 20460 26476 20466
rect 26424 20402 26476 20408
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 26422 20224 26478 20233
rect 26422 20159 26478 20168
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26240 19916 26292 19922
rect 26240 19858 26292 19864
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25688 15700 25740 15706
rect 25688 15642 25740 15648
rect 25412 15428 25464 15434
rect 25412 15370 25464 15376
rect 25504 15428 25556 15434
rect 25504 15370 25556 15376
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25424 14770 25452 15370
rect 25240 14414 25268 14758
rect 25424 14742 25544 14770
rect 25228 14408 25280 14414
rect 25228 14350 25280 14356
rect 25228 13456 25280 13462
rect 25228 13398 25280 13404
rect 25240 12986 25268 13398
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25412 12912 25464 12918
rect 25412 12854 25464 12860
rect 25424 12442 25452 12854
rect 25412 12436 25464 12442
rect 25412 12378 25464 12384
rect 25148 12192 25452 12220
rect 24492 12174 24544 12180
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 24639 11452 24947 11472
rect 24639 11450 24645 11452
rect 24701 11450 24725 11452
rect 24781 11450 24805 11452
rect 24861 11450 24885 11452
rect 24941 11450 24947 11452
rect 24701 11398 24703 11450
rect 24883 11398 24885 11450
rect 24639 11396 24645 11398
rect 24701 11396 24725 11398
rect 24781 11396 24805 11398
rect 24861 11396 24885 11398
rect 24941 11396 24947 11398
rect 24639 11376 24947 11396
rect 25056 11150 25084 11630
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 23676 10934 23980 10962
rect 23388 10600 23440 10606
rect 23388 10542 23440 10548
rect 23400 9110 23428 10542
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23388 9104 23440 9110
rect 23388 9046 23440 9052
rect 23768 9042 23796 9318
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23400 8498 23428 8774
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23676 8090 23704 8774
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23308 6662 23336 7686
rect 23400 7478 23428 7686
rect 23860 7546 23888 7822
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23400 6798 23428 7414
rect 23952 6914 23980 10934
rect 24044 10266 24072 11086
rect 24492 11076 24544 11082
rect 24492 11018 24544 11024
rect 24504 10810 24532 11018
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24780 10810 24808 10950
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24492 10668 24544 10674
rect 24492 10610 24544 10616
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 24504 10062 24532 10610
rect 24639 10364 24947 10384
rect 24639 10362 24645 10364
rect 24701 10362 24725 10364
rect 24781 10362 24805 10364
rect 24861 10362 24885 10364
rect 24941 10362 24947 10364
rect 24701 10310 24703 10362
rect 24883 10310 24885 10362
rect 24639 10308 24645 10310
rect 24701 10308 24725 10310
rect 24781 10308 24805 10310
rect 24861 10308 24885 10310
rect 24941 10308 24947 10310
rect 24639 10288 24947 10308
rect 24492 10056 24544 10062
rect 24492 9998 24544 10004
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24872 9722 24900 9998
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24872 9450 24900 9658
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 24639 9276 24947 9296
rect 24639 9274 24645 9276
rect 24701 9274 24725 9276
rect 24781 9274 24805 9276
rect 24861 9274 24885 9276
rect 24941 9274 24947 9276
rect 24701 9222 24703 9274
rect 24883 9222 24885 9274
rect 24639 9220 24645 9222
rect 24701 9220 24725 9222
rect 24781 9220 24805 9222
rect 24861 9220 24885 9222
rect 24941 9220 24947 9222
rect 24639 9200 24947 9220
rect 24952 8968 25004 8974
rect 25056 8956 25084 11086
rect 25004 8928 25084 8956
rect 24952 8910 25004 8916
rect 24964 8566 24992 8910
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 25332 8634 25360 8842
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 24952 8560 25004 8566
rect 25004 8508 25084 8514
rect 24952 8502 25084 8508
rect 24964 8486 25084 8502
rect 24639 8188 24947 8208
rect 24639 8186 24645 8188
rect 24701 8186 24725 8188
rect 24781 8186 24805 8188
rect 24861 8186 24885 8188
rect 24941 8186 24947 8188
rect 24701 8134 24703 8186
rect 24883 8134 24885 8186
rect 24639 8132 24645 8134
rect 24701 8132 24725 8134
rect 24781 8132 24805 8134
rect 24861 8132 24885 8134
rect 24941 8132 24947 8134
rect 24639 8112 24947 8132
rect 24639 7100 24947 7120
rect 24639 7098 24645 7100
rect 24701 7098 24725 7100
rect 24781 7098 24805 7100
rect 24861 7098 24885 7100
rect 24941 7098 24947 7100
rect 24701 7046 24703 7098
rect 24883 7046 24885 7098
rect 24639 7044 24645 7046
rect 24701 7044 24725 7046
rect 24781 7044 24805 7046
rect 24861 7044 24885 7046
rect 24941 7044 24947 7046
rect 24639 7024 24947 7044
rect 23952 6886 24348 6914
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23480 6180 23532 6186
rect 23480 6122 23532 6128
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 23032 5766 23244 5794
rect 22836 5636 22888 5642
rect 22836 5578 22888 5584
rect 22928 5636 22980 5642
rect 22928 5578 22980 5584
rect 22848 5370 22876 5578
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22008 2984 22060 2990
rect 21836 2944 22008 2972
rect 21732 2916 21784 2922
rect 21732 2858 21784 2864
rect 21836 2854 21864 2944
rect 22008 2926 22060 2932
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21192 870 21312 898
rect 21192 762 21220 870
rect 21284 800 21312 870
rect 23032 800 23060 5766
rect 23204 5704 23256 5710
rect 23204 5646 23256 5652
rect 23216 4146 23244 5646
rect 23400 5166 23428 5850
rect 23492 5370 23520 6122
rect 23584 5914 23612 6258
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23400 4690 23428 5102
rect 23952 5098 23980 5170
rect 23940 5092 23992 5098
rect 23940 5034 23992 5040
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23400 3670 23428 4626
rect 23952 4622 23980 5034
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23756 4548 23808 4554
rect 23756 4490 23808 4496
rect 23768 4214 23796 4490
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23492 3738 23520 4082
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23388 3664 23440 3670
rect 23388 3606 23440 3612
rect 23860 3534 23888 4422
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23952 3602 23980 3878
rect 23940 3596 23992 3602
rect 23940 3538 23992 3544
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 21008 734 21220 762
rect 21270 0 21326 800
rect 23018 0 23074 800
rect 24320 762 24348 6886
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24400 6724 24452 6730
rect 24400 6666 24452 6672
rect 24412 6322 24440 6666
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 24412 5914 24440 6258
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24412 4010 24440 5850
rect 24504 5658 24532 6802
rect 25056 6254 25084 8486
rect 25228 8356 25280 8362
rect 25228 8298 25280 8304
rect 25240 7954 25268 8298
rect 25228 7948 25280 7954
rect 25228 7890 25280 7896
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25148 7478 25176 7822
rect 25240 7546 25268 7890
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 25240 7392 25268 7482
rect 25240 7364 25360 7392
rect 25136 7336 25188 7342
rect 25136 7278 25188 7284
rect 25148 6390 25176 7278
rect 25228 7268 25280 7274
rect 25228 7210 25280 7216
rect 25240 6798 25268 7210
rect 25332 7002 25360 7364
rect 25320 6996 25372 7002
rect 25320 6938 25372 6944
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25424 6458 25452 12192
rect 25516 10538 25544 14742
rect 25792 14618 25820 19110
rect 26252 18834 26280 19858
rect 26344 19378 26372 19994
rect 26436 19514 26464 20159
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26332 18896 26384 18902
rect 26332 18838 26384 18844
rect 26240 18828 26292 18834
rect 26240 18770 26292 18776
rect 26344 18737 26372 18838
rect 26436 18766 26464 19110
rect 26424 18760 26476 18766
rect 26330 18728 26386 18737
rect 26424 18702 26476 18708
rect 26330 18663 26386 18672
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26252 18358 26280 18566
rect 26240 18352 26292 18358
rect 26240 18294 26292 18300
rect 26620 18290 26648 21082
rect 26804 20534 26832 22986
rect 27172 22114 27200 23054
rect 27264 23038 27476 23066
rect 27172 22086 27292 22114
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 27172 21570 27200 21966
rect 27080 21542 27200 21570
rect 27080 21486 27108 21542
rect 27068 21480 27120 21486
rect 27068 21422 27120 21428
rect 27264 20602 27292 22086
rect 27344 21684 27396 21690
rect 27344 21626 27396 21632
rect 27252 20596 27304 20602
rect 27252 20538 27304 20544
rect 26792 20528 26844 20534
rect 26792 20470 26844 20476
rect 27068 20460 27120 20466
rect 27068 20402 27120 20408
rect 27080 20346 27108 20402
rect 26988 20318 27108 20346
rect 26884 20256 26936 20262
rect 26884 20198 26936 20204
rect 26896 19922 26924 20198
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26988 19718 27016 20318
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 26608 18284 26660 18290
rect 26608 18226 26660 18232
rect 26424 17740 26476 17746
rect 26424 17682 26476 17688
rect 26330 17232 26386 17241
rect 26330 17167 26386 17176
rect 25964 17128 26016 17134
rect 25964 17070 26016 17076
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 25976 16794 26004 17070
rect 25964 16788 26016 16794
rect 25964 16730 26016 16736
rect 26252 16250 26280 17070
rect 26344 16998 26372 17167
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26436 16522 26464 17682
rect 26620 17678 26648 18226
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26424 16516 26476 16522
rect 26424 16458 26476 16464
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26608 16176 26660 16182
rect 26608 16118 26660 16124
rect 26620 15706 26648 16118
rect 26608 15700 26660 15706
rect 26608 15642 26660 15648
rect 26332 15496 26384 15502
rect 26884 15496 26936 15502
rect 26332 15438 26384 15444
rect 26712 15444 26884 15450
rect 26712 15438 26936 15444
rect 26344 15162 26372 15438
rect 26712 15434 26924 15438
rect 26700 15428 26924 15434
rect 26752 15422 26924 15428
rect 26700 15370 26752 15376
rect 26332 15156 26384 15162
rect 26332 15098 26384 15104
rect 25780 14612 25832 14618
rect 25780 14554 25832 14560
rect 25792 14074 25820 14554
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 26344 13938 26372 15098
rect 26608 15020 26660 15026
rect 26608 14962 26660 14968
rect 26620 14074 26648 14962
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26804 14346 26832 14758
rect 26792 14340 26844 14346
rect 26792 14282 26844 14288
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26516 13252 26568 13258
rect 26516 13194 26568 13200
rect 26528 12986 26556 13194
rect 26516 12980 26568 12986
rect 26516 12922 26568 12928
rect 26988 12434 27016 19654
rect 27264 18358 27292 20538
rect 27252 18352 27304 18358
rect 27252 18294 27304 18300
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 27080 16522 27108 18158
rect 27264 17678 27292 18294
rect 27356 18290 27384 21626
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27344 17808 27396 17814
rect 27344 17750 27396 17756
rect 27252 17672 27304 17678
rect 27252 17614 27304 17620
rect 27356 17270 27384 17750
rect 27448 17746 27476 23038
rect 28184 22642 28212 23462
rect 28632 23044 28684 23050
rect 28632 22986 28684 22992
rect 28644 22778 28672 22986
rect 28632 22772 28684 22778
rect 28632 22714 28684 22720
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 27988 21616 28040 21622
rect 27988 21558 28040 21564
rect 28000 21146 28028 21558
rect 27988 21140 28040 21146
rect 27988 21082 28040 21088
rect 28184 19854 28212 22578
rect 28814 21720 28870 21729
rect 28814 21655 28816 21664
rect 28868 21655 28870 21664
rect 28816 21626 28868 21632
rect 28172 19848 28224 19854
rect 28172 19790 28224 19796
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 27632 19514 27660 19722
rect 28540 19712 28592 19718
rect 28540 19654 28592 19660
rect 27620 19508 27672 19514
rect 27620 19450 27672 19456
rect 28552 19378 28580 19654
rect 28540 19372 28592 19378
rect 28540 19314 28592 19320
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 28368 18698 28396 19110
rect 27712 18692 27764 18698
rect 27712 18634 27764 18640
rect 28356 18692 28408 18698
rect 28356 18634 28408 18640
rect 27724 18154 27752 18634
rect 27804 18624 27856 18630
rect 27804 18566 27856 18572
rect 27712 18148 27764 18154
rect 27712 18090 27764 18096
rect 27816 18086 27844 18566
rect 27804 18080 27856 18086
rect 27804 18022 27856 18028
rect 27436 17740 27488 17746
rect 27436 17682 27488 17688
rect 27344 17264 27396 17270
rect 27344 17206 27396 17212
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27528 16584 27580 16590
rect 27528 16526 27580 16532
rect 27068 16516 27120 16522
rect 27068 16458 27120 16464
rect 27172 15502 27200 16526
rect 27436 16516 27488 16522
rect 27436 16458 27488 16464
rect 27448 15994 27476 16458
rect 27356 15966 27476 15994
rect 27356 15910 27384 15966
rect 27344 15904 27396 15910
rect 27344 15846 27396 15852
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 27160 13184 27212 13190
rect 27160 13126 27212 13132
rect 27068 12912 27120 12918
rect 27068 12854 27120 12860
rect 26620 12406 27016 12434
rect 26056 11076 26108 11082
rect 26056 11018 26108 11024
rect 26424 11076 26476 11082
rect 26424 11018 26476 11024
rect 26068 10674 26096 11018
rect 26332 11008 26384 11014
rect 26332 10950 26384 10956
rect 26056 10668 26108 10674
rect 26056 10610 26108 10616
rect 25504 10532 25556 10538
rect 25504 10474 25556 10480
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 25792 8566 25820 9386
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25780 8560 25832 8566
rect 25780 8502 25832 8508
rect 25884 8430 25912 8774
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 25976 6914 26004 9522
rect 26068 9518 26096 10610
rect 26344 10606 26372 10950
rect 26436 10742 26464 11018
rect 26424 10736 26476 10742
rect 26424 10678 26476 10684
rect 26332 10600 26384 10606
rect 26332 10542 26384 10548
rect 26344 10266 26372 10542
rect 26332 10260 26384 10266
rect 26332 10202 26384 10208
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 26528 9586 26556 10066
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 26516 9580 26568 9586
rect 26516 9522 26568 9528
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 26068 8974 26096 9454
rect 26148 9376 26200 9382
rect 26148 9318 26200 9324
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 26160 8634 26188 9318
rect 26252 9110 26280 9522
rect 26240 9104 26292 9110
rect 26240 9046 26292 9052
rect 26528 8974 26556 9522
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 26516 8356 26568 8362
rect 26516 8298 26568 8304
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 26252 7410 26280 7822
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 26332 7268 26384 7274
rect 26332 7210 26384 7216
rect 25884 6886 26004 6914
rect 25412 6452 25464 6458
rect 25412 6394 25464 6400
rect 25884 6390 25912 6886
rect 26344 6798 26372 7210
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26148 6656 26200 6662
rect 26148 6598 26200 6604
rect 25136 6384 25188 6390
rect 25136 6326 25188 6332
rect 25872 6384 25924 6390
rect 25872 6326 25924 6332
rect 25964 6316 26016 6322
rect 25964 6258 26016 6264
rect 25044 6248 25096 6254
rect 25044 6190 25096 6196
rect 25320 6248 25372 6254
rect 25320 6190 25372 6196
rect 24639 6012 24947 6032
rect 24639 6010 24645 6012
rect 24701 6010 24725 6012
rect 24781 6010 24805 6012
rect 24861 6010 24885 6012
rect 24941 6010 24947 6012
rect 24701 5958 24703 6010
rect 24883 5958 24885 6010
rect 24639 5956 24645 5958
rect 24701 5956 24725 5958
rect 24781 5956 24805 5958
rect 24861 5956 24885 5958
rect 24941 5956 24947 5958
rect 24639 5936 24947 5956
rect 24860 5704 24912 5710
rect 24504 5652 24860 5658
rect 24504 5646 24912 5652
rect 24504 5630 24900 5646
rect 24780 5574 24808 5630
rect 24492 5568 24544 5574
rect 24492 5510 24544 5516
rect 24768 5568 24820 5574
rect 24768 5510 24820 5516
rect 24504 4622 24532 5510
rect 24780 5302 24808 5510
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24639 4924 24947 4944
rect 24639 4922 24645 4924
rect 24701 4922 24725 4924
rect 24781 4922 24805 4924
rect 24861 4922 24885 4924
rect 24941 4922 24947 4924
rect 24701 4870 24703 4922
rect 24883 4870 24885 4922
rect 24639 4868 24645 4870
rect 24701 4868 24725 4870
rect 24781 4868 24805 4870
rect 24861 4868 24885 4870
rect 24941 4868 24947 4870
rect 24639 4848 24947 4868
rect 25332 4690 25360 6190
rect 25976 5914 26004 6258
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 25412 5092 25464 5098
rect 25412 5034 25464 5040
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25424 4622 25452 5034
rect 25504 5024 25556 5030
rect 25504 4966 25556 4972
rect 25516 4622 25544 4966
rect 24492 4616 24544 4622
rect 24492 4558 24544 4564
rect 25412 4616 25464 4622
rect 25412 4558 25464 4564
rect 25504 4616 25556 4622
rect 25504 4558 25556 4564
rect 24584 4548 24636 4554
rect 24584 4490 24636 4496
rect 24596 4282 24624 4490
rect 24584 4276 24636 4282
rect 24584 4218 24636 4224
rect 25516 4146 25544 4558
rect 26160 4146 26188 6598
rect 26424 6180 26476 6186
rect 26424 6122 26476 6128
rect 26436 5778 26464 6122
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 26148 4140 26200 4146
rect 26148 4082 26200 4088
rect 24400 4004 24452 4010
rect 24400 3946 24452 3952
rect 24639 3836 24947 3856
rect 24639 3834 24645 3836
rect 24701 3834 24725 3836
rect 24781 3834 24805 3836
rect 24861 3834 24885 3836
rect 24941 3834 24947 3836
rect 24701 3782 24703 3834
rect 24883 3782 24885 3834
rect 24639 3780 24645 3782
rect 24701 3780 24725 3782
rect 24781 3780 24805 3782
rect 24861 3780 24885 3782
rect 24941 3780 24947 3782
rect 24639 3760 24947 3780
rect 26422 3496 26478 3505
rect 26422 3431 26478 3440
rect 24639 2748 24947 2768
rect 24639 2746 24645 2748
rect 24701 2746 24725 2748
rect 24781 2746 24805 2748
rect 24861 2746 24885 2748
rect 24941 2746 24947 2748
rect 24701 2694 24703 2746
rect 24883 2694 24885 2746
rect 24639 2692 24645 2694
rect 24701 2692 24725 2694
rect 24781 2692 24805 2694
rect 24861 2692 24885 2694
rect 24941 2692 24947 2694
rect 24639 2672 24947 2692
rect 24596 870 24716 898
rect 24596 762 24624 870
rect 24688 800 24716 870
rect 26436 800 26464 3431
rect 26528 2281 26556 8298
rect 26620 5137 26648 12406
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 26988 10742 27016 11086
rect 26976 10736 27028 10742
rect 26976 10678 27028 10684
rect 26700 10668 26752 10674
rect 26752 10628 26832 10656
rect 26700 10610 26752 10616
rect 26804 10538 26832 10628
rect 26700 10532 26752 10538
rect 26700 10474 26752 10480
rect 26792 10532 26844 10538
rect 26792 10474 26844 10480
rect 26712 10062 26740 10474
rect 26700 10056 26752 10062
rect 26700 9998 26752 10004
rect 26804 10010 26832 10474
rect 26804 9982 26924 10010
rect 26792 9920 26844 9926
rect 26792 9862 26844 9868
rect 26700 7948 26752 7954
rect 26700 7890 26752 7896
rect 26712 6866 26740 7890
rect 26804 7886 26832 9862
rect 26896 8022 26924 9982
rect 26976 9988 27028 9994
rect 26976 9930 27028 9936
rect 26988 9586 27016 9930
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 26976 9444 27028 9450
rect 26976 9386 27028 9392
rect 26988 8974 27016 9386
rect 26976 8968 27028 8974
rect 26976 8910 27028 8916
rect 26884 8016 26936 8022
rect 26884 7958 26936 7964
rect 26896 7886 26924 7958
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26884 7880 26936 7886
rect 26884 7822 26936 7828
rect 26804 7478 26832 7822
rect 26792 7472 26844 7478
rect 26792 7414 26844 7420
rect 26804 6934 26832 7414
rect 26792 6928 26844 6934
rect 26792 6870 26844 6876
rect 26700 6860 26752 6866
rect 26700 6802 26752 6808
rect 26884 6792 26936 6798
rect 26884 6734 26936 6740
rect 26896 6458 26924 6734
rect 26884 6452 26936 6458
rect 26884 6394 26936 6400
rect 26606 5128 26662 5137
rect 26606 5063 26662 5072
rect 27080 3777 27108 12854
rect 27172 11234 27200 13126
rect 27356 12753 27384 15846
rect 27540 15502 27568 16526
rect 27712 16448 27764 16454
rect 27712 16390 27764 16396
rect 27724 16182 27752 16390
rect 27712 16176 27764 16182
rect 27712 16118 27764 16124
rect 27620 15632 27672 15638
rect 27620 15574 27672 15580
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27436 15428 27488 15434
rect 27436 15370 27488 15376
rect 27448 14074 27476 15370
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27540 15162 27568 15302
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 27540 14414 27568 15098
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27528 14272 27580 14278
rect 27528 14214 27580 14220
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 27342 12744 27398 12753
rect 27342 12679 27398 12688
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27264 11354 27292 11698
rect 27252 11348 27304 11354
rect 27252 11290 27304 11296
rect 27540 11257 27568 14214
rect 27632 14006 27660 15574
rect 27620 14000 27672 14006
rect 27620 13942 27672 13948
rect 27526 11248 27582 11257
rect 27172 11206 27292 11234
rect 27160 9376 27212 9382
rect 27160 9318 27212 9324
rect 27172 8974 27200 9318
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 27264 8820 27292 11206
rect 27526 11183 27582 11192
rect 27712 11008 27764 11014
rect 27712 10950 27764 10956
rect 27724 10810 27752 10950
rect 27712 10804 27764 10810
rect 27712 10746 27764 10752
rect 27528 10464 27580 10470
rect 27528 10406 27580 10412
rect 27540 9761 27568 10406
rect 27620 9988 27672 9994
rect 27620 9930 27672 9936
rect 27526 9752 27582 9761
rect 27526 9687 27582 9696
rect 27632 9178 27660 9930
rect 27712 9512 27764 9518
rect 27712 9454 27764 9460
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 27632 8974 27660 9114
rect 27724 9042 27752 9454
rect 27712 9036 27764 9042
rect 27712 8978 27764 8984
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 27172 8792 27292 8820
rect 27620 8832 27672 8838
rect 27172 7342 27200 8792
rect 27620 8774 27672 8780
rect 27436 7948 27488 7954
rect 27436 7890 27488 7896
rect 27252 7540 27304 7546
rect 27252 7482 27304 7488
rect 27160 7336 27212 7342
rect 27160 7278 27212 7284
rect 27264 6866 27292 7482
rect 27448 7478 27476 7890
rect 27632 7886 27660 8774
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27528 7812 27580 7818
rect 27528 7754 27580 7760
rect 27436 7472 27488 7478
rect 27436 7414 27488 7420
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27252 6860 27304 6866
rect 27252 6802 27304 6808
rect 27160 6656 27212 6662
rect 27160 6598 27212 6604
rect 27172 6322 27200 6598
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 27172 5710 27200 6258
rect 27160 5704 27212 5710
rect 27160 5646 27212 5652
rect 27264 4622 27292 6802
rect 27356 6798 27384 7346
rect 27436 7336 27488 7342
rect 27436 7278 27488 7284
rect 27344 6792 27396 6798
rect 27448 6769 27476 7278
rect 27540 7274 27568 7754
rect 27528 7268 27580 7274
rect 27528 7210 27580 7216
rect 27540 7002 27568 7210
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 27344 6734 27396 6740
rect 27434 6760 27490 6769
rect 27434 6695 27490 6704
rect 27632 5794 27660 7142
rect 27724 6866 27752 8978
rect 27816 6914 27844 18022
rect 27988 17264 28040 17270
rect 27988 17206 28040 17212
rect 28000 16794 28028 17206
rect 27988 16788 28040 16794
rect 27988 16730 28040 16736
rect 28632 16176 28684 16182
rect 28632 16118 28684 16124
rect 28644 15706 28672 16118
rect 28632 15700 28684 15706
rect 28632 15642 28684 15648
rect 28632 14272 28684 14278
rect 28632 14214 28684 14220
rect 29090 14240 29146 14249
rect 28644 14006 28672 14214
rect 29090 14175 29146 14184
rect 29104 14074 29132 14175
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 28632 14000 28684 14006
rect 28632 13942 28684 13948
rect 28356 11552 28408 11558
rect 28356 11494 28408 11500
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 27896 11008 27948 11014
rect 27896 10950 27948 10956
rect 27908 10674 27936 10950
rect 27896 10668 27948 10674
rect 27896 10610 27948 10616
rect 28000 10130 28028 11086
rect 28368 10742 28396 11494
rect 28448 11212 28500 11218
rect 28448 11154 28500 11160
rect 28356 10736 28408 10742
rect 28356 10678 28408 10684
rect 27988 10124 28040 10130
rect 27988 10066 28040 10072
rect 28000 9874 28028 10066
rect 27908 9846 28028 9874
rect 28356 9920 28408 9926
rect 28356 9862 28408 9868
rect 27908 9654 27936 9846
rect 27896 9648 27948 9654
rect 27896 9590 27948 9596
rect 27908 8498 27936 9590
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 28000 9178 28028 9522
rect 27988 9172 28040 9178
rect 27988 9114 28040 9120
rect 28368 9042 28396 9862
rect 28460 9042 28488 11154
rect 28356 9036 28408 9042
rect 28356 8978 28408 8984
rect 28448 9036 28500 9042
rect 28448 8978 28500 8984
rect 28460 8616 28488 8978
rect 28460 8588 28580 8616
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 28080 8492 28132 8498
rect 28080 8434 28132 8440
rect 28092 7886 28120 8434
rect 28552 8430 28580 8588
rect 28540 8424 28592 8430
rect 28540 8366 28592 8372
rect 28448 8288 28500 8294
rect 28448 8230 28500 8236
rect 28460 7954 28488 8230
rect 28552 7954 28580 8366
rect 29092 8288 29144 8294
rect 29090 8256 29092 8265
rect 29144 8256 29146 8265
rect 29090 8191 29146 8200
rect 28448 7948 28500 7954
rect 28448 7890 28500 7896
rect 28540 7948 28592 7954
rect 28540 7890 28592 7896
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 27908 7342 27936 7822
rect 27988 7744 28040 7750
rect 27988 7686 28040 7692
rect 27896 7336 27948 7342
rect 27896 7278 27948 7284
rect 27816 6886 27936 6914
rect 27712 6860 27764 6866
rect 27712 6802 27764 6808
rect 27540 5778 27660 5794
rect 27528 5772 27660 5778
rect 27580 5766 27660 5772
rect 27528 5714 27580 5720
rect 27526 5264 27582 5273
rect 27526 5199 27582 5208
rect 27540 4826 27568 5199
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 27252 4616 27304 4622
rect 27252 4558 27304 4564
rect 27066 3768 27122 3777
rect 27066 3703 27122 3712
rect 27908 3482 27936 6886
rect 28000 6798 28028 7686
rect 28552 7206 28580 7890
rect 29000 7880 29052 7886
rect 29000 7822 29052 7828
rect 29012 7546 29040 7822
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 28184 4826 28212 5170
rect 28172 4820 28224 4826
rect 28172 4762 28224 4768
rect 29828 3528 29880 3534
rect 27908 3454 28120 3482
rect 29828 3470 29880 3476
rect 26514 2272 26570 2281
rect 26514 2207 26570 2216
rect 27528 1352 27580 1358
rect 27528 1294 27580 1300
rect 24320 734 24624 762
rect 24674 0 24730 800
rect 26422 0 26478 800
rect 27540 785 27568 1294
rect 28092 800 28120 3454
rect 29840 800 29868 3470
rect 27526 776 27582 785
rect 27526 711 27582 720
rect 28078 0 28134 800
rect 29826 0 29882 800
<< via2 >>
rect 3882 32136 3938 32192
rect 4066 30776 4122 30832
rect 4066 29416 4122 29472
rect 4066 28092 4068 28112
rect 4068 28092 4120 28112
rect 4120 28092 4122 28112
rect 4066 28056 4122 28092
rect 4066 26696 4122 26752
rect 4066 25336 4122 25392
rect 4066 24012 4068 24032
rect 4068 24012 4120 24032
rect 4120 24012 4122 24032
rect 4066 23976 4122 24012
rect 3974 22616 4030 22672
rect 4066 21256 4122 21312
rect 3790 18536 3846 18592
rect 1306 15952 1362 16008
rect 5694 29946 5750 29948
rect 5774 29946 5830 29948
rect 5854 29946 5910 29948
rect 5934 29946 5990 29948
rect 5694 29894 5740 29946
rect 5740 29894 5750 29946
rect 5774 29894 5804 29946
rect 5804 29894 5816 29946
rect 5816 29894 5830 29946
rect 5854 29894 5868 29946
rect 5868 29894 5880 29946
rect 5880 29894 5910 29946
rect 5934 29894 5944 29946
rect 5944 29894 5990 29946
rect 5694 29892 5750 29894
rect 5774 29892 5830 29894
rect 5854 29892 5910 29894
rect 5934 29892 5990 29894
rect 5694 28858 5750 28860
rect 5774 28858 5830 28860
rect 5854 28858 5910 28860
rect 5934 28858 5990 28860
rect 5694 28806 5740 28858
rect 5740 28806 5750 28858
rect 5774 28806 5804 28858
rect 5804 28806 5816 28858
rect 5816 28806 5830 28858
rect 5854 28806 5868 28858
rect 5868 28806 5880 28858
rect 5880 28806 5910 28858
rect 5934 28806 5944 28858
rect 5944 28806 5990 28858
rect 5694 28804 5750 28806
rect 5774 28804 5830 28806
rect 5854 28804 5910 28806
rect 5934 28804 5990 28806
rect 5694 27770 5750 27772
rect 5774 27770 5830 27772
rect 5854 27770 5910 27772
rect 5934 27770 5990 27772
rect 5694 27718 5740 27770
rect 5740 27718 5750 27770
rect 5774 27718 5804 27770
rect 5804 27718 5816 27770
rect 5816 27718 5830 27770
rect 5854 27718 5868 27770
rect 5868 27718 5880 27770
rect 5880 27718 5910 27770
rect 5934 27718 5944 27770
rect 5944 27718 5990 27770
rect 5694 27716 5750 27718
rect 5774 27716 5830 27718
rect 5854 27716 5910 27718
rect 5934 27716 5990 27718
rect 5694 26682 5750 26684
rect 5774 26682 5830 26684
rect 5854 26682 5910 26684
rect 5934 26682 5990 26684
rect 5694 26630 5740 26682
rect 5740 26630 5750 26682
rect 5774 26630 5804 26682
rect 5804 26630 5816 26682
rect 5816 26630 5830 26682
rect 5854 26630 5868 26682
rect 5868 26630 5880 26682
rect 5880 26630 5910 26682
rect 5934 26630 5944 26682
rect 5944 26630 5990 26682
rect 5694 26628 5750 26630
rect 5774 26628 5830 26630
rect 5854 26628 5910 26630
rect 5934 26628 5990 26630
rect 5694 25594 5750 25596
rect 5774 25594 5830 25596
rect 5854 25594 5910 25596
rect 5934 25594 5990 25596
rect 5694 25542 5740 25594
rect 5740 25542 5750 25594
rect 5774 25542 5804 25594
rect 5804 25542 5816 25594
rect 5816 25542 5830 25594
rect 5854 25542 5868 25594
rect 5868 25542 5880 25594
rect 5880 25542 5910 25594
rect 5934 25542 5944 25594
rect 5944 25542 5990 25594
rect 5694 25540 5750 25542
rect 5774 25540 5830 25542
rect 5854 25540 5910 25542
rect 5934 25540 5990 25542
rect 5694 24506 5750 24508
rect 5774 24506 5830 24508
rect 5854 24506 5910 24508
rect 5934 24506 5990 24508
rect 5694 24454 5740 24506
rect 5740 24454 5750 24506
rect 5774 24454 5804 24506
rect 5804 24454 5816 24506
rect 5816 24454 5830 24506
rect 5854 24454 5868 24506
rect 5868 24454 5880 24506
rect 5880 24454 5910 24506
rect 5934 24454 5944 24506
rect 5944 24454 5990 24506
rect 5694 24452 5750 24454
rect 5774 24452 5830 24454
rect 5854 24452 5910 24454
rect 5934 24452 5990 24454
rect 5694 23418 5750 23420
rect 5774 23418 5830 23420
rect 5854 23418 5910 23420
rect 5934 23418 5990 23420
rect 5694 23366 5740 23418
rect 5740 23366 5750 23418
rect 5774 23366 5804 23418
rect 5804 23366 5816 23418
rect 5816 23366 5830 23418
rect 5854 23366 5868 23418
rect 5868 23366 5880 23418
rect 5880 23366 5910 23418
rect 5934 23366 5944 23418
rect 5944 23366 5990 23418
rect 5694 23364 5750 23366
rect 5774 23364 5830 23366
rect 5854 23364 5910 23366
rect 5934 23364 5990 23366
rect 3790 16088 3846 16144
rect 4066 17176 4122 17232
rect 4066 15680 4122 15736
rect 5694 22330 5750 22332
rect 5774 22330 5830 22332
rect 5854 22330 5910 22332
rect 5934 22330 5990 22332
rect 5694 22278 5740 22330
rect 5740 22278 5750 22330
rect 5774 22278 5804 22330
rect 5804 22278 5816 22330
rect 5816 22278 5830 22330
rect 5854 22278 5868 22330
rect 5868 22278 5880 22330
rect 5880 22278 5910 22330
rect 5934 22278 5944 22330
rect 5944 22278 5990 22330
rect 5694 22276 5750 22278
rect 5774 22276 5830 22278
rect 5854 22276 5910 22278
rect 5934 22276 5990 22278
rect 5694 21242 5750 21244
rect 5774 21242 5830 21244
rect 5854 21242 5910 21244
rect 5934 21242 5990 21244
rect 5694 21190 5740 21242
rect 5740 21190 5750 21242
rect 5774 21190 5804 21242
rect 5804 21190 5816 21242
rect 5816 21190 5830 21242
rect 5854 21190 5868 21242
rect 5868 21190 5880 21242
rect 5880 21190 5910 21242
rect 5934 21190 5944 21242
rect 5944 21190 5990 21242
rect 5694 21188 5750 21190
rect 5774 21188 5830 21190
rect 5854 21188 5910 21190
rect 5934 21188 5990 21190
rect 5694 20154 5750 20156
rect 5774 20154 5830 20156
rect 5854 20154 5910 20156
rect 5934 20154 5990 20156
rect 5694 20102 5740 20154
rect 5740 20102 5750 20154
rect 5774 20102 5804 20154
rect 5804 20102 5816 20154
rect 5816 20102 5830 20154
rect 5854 20102 5868 20154
rect 5868 20102 5880 20154
rect 5880 20102 5910 20154
rect 5934 20102 5944 20154
rect 5944 20102 5990 20154
rect 5694 20100 5750 20102
rect 5774 20100 5830 20102
rect 5854 20100 5910 20102
rect 5934 20100 5990 20102
rect 5694 19066 5750 19068
rect 5774 19066 5830 19068
rect 5854 19066 5910 19068
rect 5934 19066 5990 19068
rect 5694 19014 5740 19066
rect 5740 19014 5750 19066
rect 5774 19014 5804 19066
rect 5804 19014 5816 19066
rect 5816 19014 5830 19066
rect 5854 19014 5868 19066
rect 5868 19014 5880 19066
rect 5880 19014 5910 19066
rect 5934 19014 5944 19066
rect 5944 19014 5990 19066
rect 5694 19012 5750 19014
rect 5774 19012 5830 19014
rect 5854 19012 5910 19014
rect 5934 19012 5990 19014
rect 4066 15000 4122 15056
rect 4066 14320 4122 14376
rect 3882 12960 3938 13016
rect 4802 12824 4858 12880
rect 5694 17978 5750 17980
rect 5774 17978 5830 17980
rect 5854 17978 5910 17980
rect 5934 17978 5990 17980
rect 5694 17926 5740 17978
rect 5740 17926 5750 17978
rect 5774 17926 5804 17978
rect 5804 17926 5816 17978
rect 5816 17926 5830 17978
rect 5854 17926 5868 17978
rect 5868 17926 5880 17978
rect 5880 17926 5910 17978
rect 5934 17926 5944 17978
rect 5944 17926 5990 17978
rect 5694 17924 5750 17926
rect 5774 17924 5830 17926
rect 5854 17924 5910 17926
rect 5934 17924 5990 17926
rect 5694 16890 5750 16892
rect 5774 16890 5830 16892
rect 5854 16890 5910 16892
rect 5934 16890 5990 16892
rect 5694 16838 5740 16890
rect 5740 16838 5750 16890
rect 5774 16838 5804 16890
rect 5804 16838 5816 16890
rect 5816 16838 5830 16890
rect 5854 16838 5868 16890
rect 5868 16838 5880 16890
rect 5880 16838 5910 16890
rect 5934 16838 5944 16890
rect 5944 16838 5990 16890
rect 5694 16836 5750 16838
rect 5774 16836 5830 16838
rect 5854 16836 5910 16838
rect 5934 16836 5990 16838
rect 5694 15802 5750 15804
rect 5774 15802 5830 15804
rect 5854 15802 5910 15804
rect 5934 15802 5990 15804
rect 5694 15750 5740 15802
rect 5740 15750 5750 15802
rect 5774 15750 5804 15802
rect 5804 15750 5816 15802
rect 5816 15750 5830 15802
rect 5854 15750 5868 15802
rect 5868 15750 5880 15802
rect 5880 15750 5910 15802
rect 5934 15750 5944 15802
rect 5944 15750 5990 15802
rect 5694 15748 5750 15750
rect 5774 15748 5830 15750
rect 5854 15748 5910 15750
rect 5934 15748 5990 15750
rect 4066 11600 4122 11656
rect 3974 10240 4030 10296
rect 3698 8880 3754 8936
rect 5694 14714 5750 14716
rect 5774 14714 5830 14716
rect 5854 14714 5910 14716
rect 5934 14714 5990 14716
rect 5694 14662 5740 14714
rect 5740 14662 5750 14714
rect 5774 14662 5804 14714
rect 5804 14662 5816 14714
rect 5816 14662 5830 14714
rect 5854 14662 5868 14714
rect 5868 14662 5880 14714
rect 5880 14662 5910 14714
rect 5934 14662 5944 14714
rect 5944 14662 5990 14714
rect 5694 14660 5750 14662
rect 5774 14660 5830 14662
rect 5854 14660 5910 14662
rect 5934 14660 5990 14662
rect 5694 13626 5750 13628
rect 5774 13626 5830 13628
rect 5854 13626 5910 13628
rect 5934 13626 5990 13628
rect 5694 13574 5740 13626
rect 5740 13574 5750 13626
rect 5774 13574 5804 13626
rect 5804 13574 5816 13626
rect 5816 13574 5830 13626
rect 5854 13574 5868 13626
rect 5868 13574 5880 13626
rect 5880 13574 5910 13626
rect 5934 13574 5944 13626
rect 5944 13574 5990 13626
rect 5694 13572 5750 13574
rect 5774 13572 5830 13574
rect 5854 13572 5910 13574
rect 5934 13572 5990 13574
rect 5446 12824 5502 12880
rect 5262 12552 5318 12608
rect 5694 12538 5750 12540
rect 5774 12538 5830 12540
rect 5854 12538 5910 12540
rect 5934 12538 5990 12540
rect 5694 12486 5740 12538
rect 5740 12486 5750 12538
rect 5774 12486 5804 12538
rect 5804 12486 5816 12538
rect 5816 12486 5830 12538
rect 5854 12486 5868 12538
rect 5868 12486 5880 12538
rect 5880 12486 5910 12538
rect 5934 12486 5944 12538
rect 5944 12486 5990 12538
rect 5694 12484 5750 12486
rect 5774 12484 5830 12486
rect 5854 12484 5910 12486
rect 5934 12484 5990 12486
rect 5906 12280 5962 12336
rect 5694 11450 5750 11452
rect 5774 11450 5830 11452
rect 5854 11450 5910 11452
rect 5934 11450 5990 11452
rect 5694 11398 5740 11450
rect 5740 11398 5750 11450
rect 5774 11398 5804 11450
rect 5804 11398 5816 11450
rect 5816 11398 5830 11450
rect 5854 11398 5868 11450
rect 5868 11398 5880 11450
rect 5880 11398 5910 11450
rect 5934 11398 5944 11450
rect 5944 11398 5990 11450
rect 5694 11396 5750 11398
rect 5774 11396 5830 11398
rect 5854 11396 5910 11398
rect 5934 11396 5990 11398
rect 5694 10362 5750 10364
rect 5774 10362 5830 10364
rect 5854 10362 5910 10364
rect 5934 10362 5990 10364
rect 5694 10310 5740 10362
rect 5740 10310 5750 10362
rect 5774 10310 5804 10362
rect 5804 10310 5816 10362
rect 5816 10310 5830 10362
rect 5854 10310 5868 10362
rect 5868 10310 5880 10362
rect 5880 10310 5910 10362
rect 5934 10310 5944 10362
rect 5944 10310 5990 10362
rect 5694 10308 5750 10310
rect 5774 10308 5830 10310
rect 5854 10308 5910 10310
rect 5934 10308 5990 10310
rect 5694 9274 5750 9276
rect 5774 9274 5830 9276
rect 5854 9274 5910 9276
rect 5934 9274 5990 9276
rect 5694 9222 5740 9274
rect 5740 9222 5750 9274
rect 5774 9222 5804 9274
rect 5804 9222 5816 9274
rect 5816 9222 5830 9274
rect 5854 9222 5868 9274
rect 5868 9222 5880 9274
rect 5880 9222 5910 9274
rect 5934 9222 5944 9274
rect 5944 9222 5990 9274
rect 5694 9220 5750 9222
rect 5774 9220 5830 9222
rect 5854 9220 5910 9222
rect 5934 9220 5990 9222
rect 5694 8186 5750 8188
rect 5774 8186 5830 8188
rect 5854 8186 5910 8188
rect 5934 8186 5990 8188
rect 5694 8134 5740 8186
rect 5740 8134 5750 8186
rect 5774 8134 5804 8186
rect 5804 8134 5816 8186
rect 5816 8134 5830 8186
rect 5854 8134 5868 8186
rect 5868 8134 5880 8186
rect 5880 8134 5910 8186
rect 5934 8134 5944 8186
rect 5944 8134 5990 8186
rect 5694 8132 5750 8134
rect 5774 8132 5830 8134
rect 5854 8132 5910 8134
rect 5934 8132 5990 8134
rect 4066 7520 4122 7576
rect 5694 7098 5750 7100
rect 5774 7098 5830 7100
rect 5854 7098 5910 7100
rect 5934 7098 5990 7100
rect 5694 7046 5740 7098
rect 5740 7046 5750 7098
rect 5774 7046 5804 7098
rect 5804 7046 5816 7098
rect 5816 7046 5830 7098
rect 5854 7046 5868 7098
rect 5868 7046 5880 7098
rect 5880 7046 5910 7098
rect 5934 7046 5944 7098
rect 5944 7046 5990 7098
rect 5694 7044 5750 7046
rect 5774 7044 5830 7046
rect 5854 7044 5910 7046
rect 5934 7044 5990 7046
rect 9862 28500 9864 28520
rect 9864 28500 9916 28520
rect 9916 28500 9918 28520
rect 9862 28464 9918 28500
rect 10431 30490 10487 30492
rect 10511 30490 10567 30492
rect 10591 30490 10647 30492
rect 10671 30490 10727 30492
rect 10431 30438 10477 30490
rect 10477 30438 10487 30490
rect 10511 30438 10541 30490
rect 10541 30438 10553 30490
rect 10553 30438 10567 30490
rect 10591 30438 10605 30490
rect 10605 30438 10617 30490
rect 10617 30438 10647 30490
rect 10671 30438 10681 30490
rect 10681 30438 10727 30490
rect 10431 30436 10487 30438
rect 10511 30436 10567 30438
rect 10591 30436 10647 30438
rect 10671 30436 10727 30438
rect 10431 29402 10487 29404
rect 10511 29402 10567 29404
rect 10591 29402 10647 29404
rect 10671 29402 10727 29404
rect 10431 29350 10477 29402
rect 10477 29350 10487 29402
rect 10511 29350 10541 29402
rect 10541 29350 10553 29402
rect 10553 29350 10567 29402
rect 10591 29350 10605 29402
rect 10605 29350 10617 29402
rect 10617 29350 10647 29402
rect 10671 29350 10681 29402
rect 10681 29350 10727 29402
rect 10431 29348 10487 29350
rect 10511 29348 10567 29350
rect 10591 29348 10647 29350
rect 10671 29348 10727 29350
rect 10598 28484 10654 28520
rect 10598 28464 10600 28484
rect 10600 28464 10652 28484
rect 10652 28464 10654 28484
rect 10782 28500 10784 28520
rect 10784 28500 10836 28520
rect 10836 28500 10838 28520
rect 10782 28464 10838 28500
rect 10431 28314 10487 28316
rect 10511 28314 10567 28316
rect 10591 28314 10647 28316
rect 10671 28314 10727 28316
rect 10431 28262 10477 28314
rect 10477 28262 10487 28314
rect 10511 28262 10541 28314
rect 10541 28262 10553 28314
rect 10553 28262 10567 28314
rect 10591 28262 10605 28314
rect 10605 28262 10617 28314
rect 10617 28262 10647 28314
rect 10671 28262 10681 28314
rect 10681 28262 10727 28314
rect 10431 28260 10487 28262
rect 10511 28260 10567 28262
rect 10591 28260 10647 28262
rect 10671 28260 10727 28262
rect 10322 27920 10378 27976
rect 4066 6160 4122 6216
rect 3882 4800 3938 4856
rect 1858 3440 1914 3496
rect 3422 2080 3478 2136
rect 3146 720 3202 776
rect 5694 6010 5750 6012
rect 5774 6010 5830 6012
rect 5854 6010 5910 6012
rect 5934 6010 5990 6012
rect 5694 5958 5740 6010
rect 5740 5958 5750 6010
rect 5774 5958 5804 6010
rect 5804 5958 5816 6010
rect 5816 5958 5830 6010
rect 5854 5958 5868 6010
rect 5868 5958 5880 6010
rect 5880 5958 5910 6010
rect 5934 5958 5944 6010
rect 5944 5958 5990 6010
rect 5694 5956 5750 5958
rect 5774 5956 5830 5958
rect 5854 5956 5910 5958
rect 5934 5956 5990 5958
rect 5694 4922 5750 4924
rect 5774 4922 5830 4924
rect 5854 4922 5910 4924
rect 5934 4922 5990 4924
rect 5694 4870 5740 4922
rect 5740 4870 5750 4922
rect 5774 4870 5804 4922
rect 5804 4870 5816 4922
rect 5816 4870 5830 4922
rect 5854 4870 5868 4922
rect 5868 4870 5880 4922
rect 5880 4870 5910 4922
rect 5934 4870 5944 4922
rect 5944 4870 5990 4922
rect 5694 4868 5750 4870
rect 5774 4868 5830 4870
rect 5854 4868 5910 4870
rect 5934 4868 5990 4870
rect 5694 3834 5750 3836
rect 5774 3834 5830 3836
rect 5854 3834 5910 3836
rect 5934 3834 5990 3836
rect 5694 3782 5740 3834
rect 5740 3782 5750 3834
rect 5774 3782 5804 3834
rect 5804 3782 5816 3834
rect 5816 3782 5830 3834
rect 5854 3782 5868 3834
rect 5868 3782 5880 3834
rect 5880 3782 5910 3834
rect 5934 3782 5944 3834
rect 5944 3782 5990 3834
rect 5694 3780 5750 3782
rect 5774 3780 5830 3782
rect 5854 3780 5910 3782
rect 5934 3780 5990 3782
rect 5694 2746 5750 2748
rect 5774 2746 5830 2748
rect 5854 2746 5910 2748
rect 5934 2746 5990 2748
rect 5694 2694 5740 2746
rect 5740 2694 5750 2746
rect 5774 2694 5804 2746
rect 5804 2694 5816 2746
rect 5816 2694 5830 2746
rect 5854 2694 5868 2746
rect 5868 2694 5880 2746
rect 5880 2694 5910 2746
rect 5934 2694 5944 2746
rect 5944 2694 5990 2746
rect 5694 2692 5750 2694
rect 5774 2692 5830 2694
rect 5854 2692 5910 2694
rect 5934 2692 5990 2694
rect 7930 19388 7932 19408
rect 7932 19388 7984 19408
rect 7984 19388 7986 19408
rect 7930 19352 7986 19388
rect 10431 27226 10487 27228
rect 10511 27226 10567 27228
rect 10591 27226 10647 27228
rect 10671 27226 10727 27228
rect 10431 27174 10477 27226
rect 10477 27174 10487 27226
rect 10511 27174 10541 27226
rect 10541 27174 10553 27226
rect 10553 27174 10567 27226
rect 10591 27174 10605 27226
rect 10605 27174 10617 27226
rect 10617 27174 10647 27226
rect 10671 27174 10681 27226
rect 10681 27174 10727 27226
rect 10431 27172 10487 27174
rect 10511 27172 10567 27174
rect 10591 27172 10647 27174
rect 10671 27172 10727 27174
rect 10431 26138 10487 26140
rect 10511 26138 10567 26140
rect 10591 26138 10647 26140
rect 10671 26138 10727 26140
rect 10431 26086 10477 26138
rect 10477 26086 10487 26138
rect 10511 26086 10541 26138
rect 10541 26086 10553 26138
rect 10553 26086 10567 26138
rect 10591 26086 10605 26138
rect 10605 26086 10617 26138
rect 10617 26086 10647 26138
rect 10671 26086 10681 26138
rect 10681 26086 10727 26138
rect 10431 26084 10487 26086
rect 10511 26084 10567 26086
rect 10591 26084 10647 26086
rect 10671 26084 10727 26086
rect 10431 25050 10487 25052
rect 10511 25050 10567 25052
rect 10591 25050 10647 25052
rect 10671 25050 10727 25052
rect 10431 24998 10477 25050
rect 10477 24998 10487 25050
rect 10511 24998 10541 25050
rect 10541 24998 10553 25050
rect 10553 24998 10567 25050
rect 10591 24998 10605 25050
rect 10605 24998 10617 25050
rect 10617 24998 10647 25050
rect 10671 24998 10681 25050
rect 10681 24998 10727 25050
rect 10431 24996 10487 24998
rect 10511 24996 10567 24998
rect 10591 24996 10647 24998
rect 10671 24996 10727 24998
rect 9770 21936 9826 21992
rect 10046 21936 10102 21992
rect 10431 23962 10487 23964
rect 10511 23962 10567 23964
rect 10591 23962 10647 23964
rect 10671 23962 10727 23964
rect 10431 23910 10477 23962
rect 10477 23910 10487 23962
rect 10511 23910 10541 23962
rect 10541 23910 10553 23962
rect 10553 23910 10567 23962
rect 10591 23910 10605 23962
rect 10605 23910 10617 23962
rect 10617 23910 10647 23962
rect 10671 23910 10681 23962
rect 10681 23910 10727 23962
rect 10431 23908 10487 23910
rect 10511 23908 10567 23910
rect 10591 23908 10647 23910
rect 10671 23908 10727 23910
rect 10431 22874 10487 22876
rect 10511 22874 10567 22876
rect 10591 22874 10647 22876
rect 10671 22874 10727 22876
rect 10431 22822 10477 22874
rect 10477 22822 10487 22874
rect 10511 22822 10541 22874
rect 10541 22822 10553 22874
rect 10553 22822 10567 22874
rect 10591 22822 10605 22874
rect 10605 22822 10617 22874
rect 10617 22822 10647 22874
rect 10671 22822 10681 22874
rect 10681 22822 10727 22874
rect 10431 22820 10487 22822
rect 10511 22820 10567 22822
rect 10591 22820 10647 22822
rect 10671 22820 10727 22822
rect 10431 21786 10487 21788
rect 10511 21786 10567 21788
rect 10591 21786 10647 21788
rect 10671 21786 10727 21788
rect 10431 21734 10477 21786
rect 10477 21734 10487 21786
rect 10511 21734 10541 21786
rect 10541 21734 10553 21786
rect 10553 21734 10567 21786
rect 10591 21734 10605 21786
rect 10605 21734 10617 21786
rect 10617 21734 10647 21786
rect 10671 21734 10681 21786
rect 10681 21734 10727 21786
rect 10431 21732 10487 21734
rect 10511 21732 10567 21734
rect 10591 21732 10647 21734
rect 10671 21732 10727 21734
rect 9310 19896 9366 19952
rect 10431 20698 10487 20700
rect 10511 20698 10567 20700
rect 10591 20698 10647 20700
rect 10671 20698 10727 20700
rect 10431 20646 10477 20698
rect 10477 20646 10487 20698
rect 10511 20646 10541 20698
rect 10541 20646 10553 20698
rect 10553 20646 10567 20698
rect 10591 20646 10605 20698
rect 10605 20646 10617 20698
rect 10617 20646 10647 20698
rect 10671 20646 10681 20698
rect 10681 20646 10727 20698
rect 10431 20644 10487 20646
rect 10511 20644 10567 20646
rect 10591 20644 10647 20646
rect 10671 20644 10727 20646
rect 10230 19760 10286 19816
rect 9770 15544 9826 15600
rect 10431 19610 10487 19612
rect 10511 19610 10567 19612
rect 10591 19610 10647 19612
rect 10671 19610 10727 19612
rect 10431 19558 10477 19610
rect 10477 19558 10487 19610
rect 10511 19558 10541 19610
rect 10541 19558 10553 19610
rect 10553 19558 10567 19610
rect 10591 19558 10605 19610
rect 10605 19558 10617 19610
rect 10617 19558 10647 19610
rect 10671 19558 10681 19610
rect 10681 19558 10727 19610
rect 10431 19556 10487 19558
rect 10511 19556 10567 19558
rect 10591 19556 10647 19558
rect 10671 19556 10727 19558
rect 10431 18522 10487 18524
rect 10511 18522 10567 18524
rect 10591 18522 10647 18524
rect 10671 18522 10727 18524
rect 10431 18470 10477 18522
rect 10477 18470 10487 18522
rect 10511 18470 10541 18522
rect 10541 18470 10553 18522
rect 10553 18470 10567 18522
rect 10591 18470 10605 18522
rect 10605 18470 10617 18522
rect 10617 18470 10647 18522
rect 10671 18470 10681 18522
rect 10681 18470 10727 18522
rect 10431 18468 10487 18470
rect 10511 18468 10567 18470
rect 10591 18468 10647 18470
rect 10671 18468 10727 18470
rect 10431 17434 10487 17436
rect 10511 17434 10567 17436
rect 10591 17434 10647 17436
rect 10671 17434 10727 17436
rect 10431 17382 10477 17434
rect 10477 17382 10487 17434
rect 10511 17382 10541 17434
rect 10541 17382 10553 17434
rect 10553 17382 10567 17434
rect 10591 17382 10605 17434
rect 10605 17382 10617 17434
rect 10617 17382 10647 17434
rect 10671 17382 10681 17434
rect 10681 17382 10727 17434
rect 10431 17380 10487 17382
rect 10511 17380 10567 17382
rect 10591 17380 10647 17382
rect 10671 17380 10727 17382
rect 10431 16346 10487 16348
rect 10511 16346 10567 16348
rect 10591 16346 10647 16348
rect 10671 16346 10727 16348
rect 10431 16294 10477 16346
rect 10477 16294 10487 16346
rect 10511 16294 10541 16346
rect 10541 16294 10553 16346
rect 10553 16294 10567 16346
rect 10591 16294 10605 16346
rect 10605 16294 10617 16346
rect 10617 16294 10647 16346
rect 10671 16294 10681 16346
rect 10681 16294 10727 16346
rect 10431 16292 10487 16294
rect 10511 16292 10567 16294
rect 10591 16292 10647 16294
rect 10671 16292 10727 16294
rect 10431 15258 10487 15260
rect 10511 15258 10567 15260
rect 10591 15258 10647 15260
rect 10671 15258 10727 15260
rect 10431 15206 10477 15258
rect 10477 15206 10487 15258
rect 10511 15206 10541 15258
rect 10541 15206 10553 15258
rect 10553 15206 10567 15258
rect 10591 15206 10605 15258
rect 10605 15206 10617 15258
rect 10617 15206 10647 15258
rect 10671 15206 10681 15258
rect 10681 15206 10727 15258
rect 10431 15204 10487 15206
rect 10511 15204 10567 15206
rect 10591 15204 10647 15206
rect 10671 15204 10727 15206
rect 11978 26852 12034 26888
rect 11978 26832 11980 26852
rect 11980 26832 12032 26852
rect 12032 26832 12034 26852
rect 12622 28500 12624 28520
rect 12624 28500 12676 28520
rect 12676 28500 12678 28520
rect 12622 28464 12678 28500
rect 10431 14170 10487 14172
rect 10511 14170 10567 14172
rect 10591 14170 10647 14172
rect 10671 14170 10727 14172
rect 10431 14118 10477 14170
rect 10477 14118 10487 14170
rect 10511 14118 10541 14170
rect 10541 14118 10553 14170
rect 10553 14118 10567 14170
rect 10591 14118 10605 14170
rect 10605 14118 10617 14170
rect 10617 14118 10647 14170
rect 10671 14118 10681 14170
rect 10681 14118 10727 14170
rect 10431 14116 10487 14118
rect 10511 14116 10567 14118
rect 10591 14116 10647 14118
rect 10671 14116 10727 14118
rect 10431 13082 10487 13084
rect 10511 13082 10567 13084
rect 10591 13082 10647 13084
rect 10671 13082 10727 13084
rect 10431 13030 10477 13082
rect 10477 13030 10487 13082
rect 10511 13030 10541 13082
rect 10541 13030 10553 13082
rect 10553 13030 10567 13082
rect 10591 13030 10605 13082
rect 10605 13030 10617 13082
rect 10617 13030 10647 13082
rect 10671 13030 10681 13082
rect 10681 13030 10727 13082
rect 10431 13028 10487 13030
rect 10511 13028 10567 13030
rect 10591 13028 10647 13030
rect 10671 13028 10727 13030
rect 10431 11994 10487 11996
rect 10511 11994 10567 11996
rect 10591 11994 10647 11996
rect 10671 11994 10727 11996
rect 10431 11942 10477 11994
rect 10477 11942 10487 11994
rect 10511 11942 10541 11994
rect 10541 11942 10553 11994
rect 10553 11942 10567 11994
rect 10591 11942 10605 11994
rect 10605 11942 10617 11994
rect 10617 11942 10647 11994
rect 10671 11942 10681 11994
rect 10681 11942 10727 11994
rect 10431 11940 10487 11942
rect 10511 11940 10567 11942
rect 10591 11940 10647 11942
rect 10671 11940 10727 11942
rect 10690 11092 10692 11112
rect 10692 11092 10744 11112
rect 10744 11092 10746 11112
rect 10690 11056 10746 11092
rect 10431 10906 10487 10908
rect 10511 10906 10567 10908
rect 10591 10906 10647 10908
rect 10671 10906 10727 10908
rect 10431 10854 10477 10906
rect 10477 10854 10487 10906
rect 10511 10854 10541 10906
rect 10541 10854 10553 10906
rect 10553 10854 10567 10906
rect 10591 10854 10605 10906
rect 10605 10854 10617 10906
rect 10617 10854 10647 10906
rect 10671 10854 10681 10906
rect 10681 10854 10727 10906
rect 10431 10852 10487 10854
rect 10511 10852 10567 10854
rect 10591 10852 10647 10854
rect 10671 10852 10727 10854
rect 10506 10668 10562 10704
rect 10506 10648 10508 10668
rect 10508 10648 10560 10668
rect 10560 10648 10562 10668
rect 10690 10512 10746 10568
rect 10431 9818 10487 9820
rect 10511 9818 10567 9820
rect 10591 9818 10647 9820
rect 10671 9818 10727 9820
rect 10431 9766 10477 9818
rect 10477 9766 10487 9818
rect 10511 9766 10541 9818
rect 10541 9766 10553 9818
rect 10553 9766 10567 9818
rect 10591 9766 10605 9818
rect 10605 9766 10617 9818
rect 10617 9766 10647 9818
rect 10671 9766 10681 9818
rect 10681 9766 10727 9818
rect 10431 9764 10487 9766
rect 10511 9764 10567 9766
rect 10591 9764 10647 9766
rect 10671 9764 10727 9766
rect 11150 10648 11206 10704
rect 10874 10532 10930 10568
rect 10874 10512 10876 10532
rect 10876 10512 10928 10532
rect 10928 10512 10930 10532
rect 10431 8730 10487 8732
rect 10511 8730 10567 8732
rect 10591 8730 10647 8732
rect 10671 8730 10727 8732
rect 10431 8678 10477 8730
rect 10477 8678 10487 8730
rect 10511 8678 10541 8730
rect 10541 8678 10553 8730
rect 10553 8678 10567 8730
rect 10591 8678 10605 8730
rect 10605 8678 10617 8730
rect 10617 8678 10647 8730
rect 10671 8678 10681 8730
rect 10681 8678 10727 8730
rect 10431 8676 10487 8678
rect 10511 8676 10567 8678
rect 10591 8676 10647 8678
rect 10671 8676 10727 8678
rect 10431 7642 10487 7644
rect 10511 7642 10567 7644
rect 10591 7642 10647 7644
rect 10671 7642 10727 7644
rect 10431 7590 10477 7642
rect 10477 7590 10487 7642
rect 10511 7590 10541 7642
rect 10541 7590 10553 7642
rect 10553 7590 10567 7642
rect 10591 7590 10605 7642
rect 10605 7590 10617 7642
rect 10617 7590 10647 7642
rect 10671 7590 10681 7642
rect 10681 7590 10727 7642
rect 10431 7588 10487 7590
rect 10511 7588 10567 7590
rect 10591 7588 10647 7590
rect 10671 7588 10727 7590
rect 10431 6554 10487 6556
rect 10511 6554 10567 6556
rect 10591 6554 10647 6556
rect 10671 6554 10727 6556
rect 10431 6502 10477 6554
rect 10477 6502 10487 6554
rect 10511 6502 10541 6554
rect 10541 6502 10553 6554
rect 10553 6502 10567 6554
rect 10591 6502 10605 6554
rect 10605 6502 10617 6554
rect 10617 6502 10647 6554
rect 10671 6502 10681 6554
rect 10681 6502 10727 6554
rect 10431 6500 10487 6502
rect 10511 6500 10567 6502
rect 10591 6500 10647 6502
rect 10671 6500 10727 6502
rect 10431 5466 10487 5468
rect 10511 5466 10567 5468
rect 10591 5466 10647 5468
rect 10671 5466 10727 5468
rect 10431 5414 10477 5466
rect 10477 5414 10487 5466
rect 10511 5414 10541 5466
rect 10541 5414 10553 5466
rect 10553 5414 10567 5466
rect 10591 5414 10605 5466
rect 10605 5414 10617 5466
rect 10617 5414 10647 5466
rect 10671 5414 10681 5466
rect 10681 5414 10727 5466
rect 10431 5412 10487 5414
rect 10511 5412 10567 5414
rect 10591 5412 10647 5414
rect 10671 5412 10727 5414
rect 10431 4378 10487 4380
rect 10511 4378 10567 4380
rect 10591 4378 10647 4380
rect 10671 4378 10727 4380
rect 10431 4326 10477 4378
rect 10477 4326 10487 4378
rect 10511 4326 10541 4378
rect 10541 4326 10553 4378
rect 10553 4326 10567 4378
rect 10591 4326 10605 4378
rect 10605 4326 10617 4378
rect 10617 4326 10647 4378
rect 10671 4326 10681 4378
rect 10681 4326 10727 4378
rect 10431 4324 10487 4326
rect 10511 4324 10567 4326
rect 10591 4324 10647 4326
rect 10671 4324 10727 4326
rect 12438 23468 12440 23488
rect 12440 23468 12492 23488
rect 12492 23468 12494 23488
rect 12438 23432 12494 23468
rect 13266 27276 13268 27296
rect 13268 27276 13320 27296
rect 13320 27276 13322 27296
rect 13266 27240 13322 27276
rect 13358 26832 13414 26888
rect 14462 29416 14518 29472
rect 15169 29946 15225 29948
rect 15249 29946 15305 29948
rect 15329 29946 15385 29948
rect 15409 29946 15465 29948
rect 15169 29894 15215 29946
rect 15215 29894 15225 29946
rect 15249 29894 15279 29946
rect 15279 29894 15291 29946
rect 15291 29894 15305 29946
rect 15329 29894 15343 29946
rect 15343 29894 15355 29946
rect 15355 29894 15385 29946
rect 15409 29894 15419 29946
rect 15419 29894 15465 29946
rect 15169 29892 15225 29894
rect 15249 29892 15305 29894
rect 15329 29892 15385 29894
rect 15409 29892 15465 29894
rect 12530 17448 12586 17504
rect 15169 28858 15225 28860
rect 15249 28858 15305 28860
rect 15329 28858 15385 28860
rect 15409 28858 15465 28860
rect 15169 28806 15215 28858
rect 15215 28806 15225 28858
rect 15249 28806 15279 28858
rect 15279 28806 15291 28858
rect 15291 28806 15305 28858
rect 15329 28806 15343 28858
rect 15343 28806 15355 28858
rect 15355 28806 15385 28858
rect 15409 28806 15419 28858
rect 15419 28806 15465 28858
rect 15169 28804 15225 28806
rect 15249 28804 15305 28806
rect 15329 28804 15385 28806
rect 15409 28804 15465 28806
rect 15169 27770 15225 27772
rect 15249 27770 15305 27772
rect 15329 27770 15385 27772
rect 15409 27770 15465 27772
rect 15169 27718 15215 27770
rect 15215 27718 15225 27770
rect 15249 27718 15279 27770
rect 15279 27718 15291 27770
rect 15291 27718 15305 27770
rect 15329 27718 15343 27770
rect 15343 27718 15355 27770
rect 15355 27718 15385 27770
rect 15409 27718 15419 27770
rect 15419 27718 15465 27770
rect 15169 27716 15225 27718
rect 15249 27716 15305 27718
rect 15329 27716 15385 27718
rect 15409 27716 15465 27718
rect 15382 27412 15384 27432
rect 15384 27412 15436 27432
rect 15436 27412 15438 27432
rect 15382 27376 15438 27412
rect 15169 26682 15225 26684
rect 15249 26682 15305 26684
rect 15329 26682 15385 26684
rect 15409 26682 15465 26684
rect 15169 26630 15215 26682
rect 15215 26630 15225 26682
rect 15249 26630 15279 26682
rect 15279 26630 15291 26682
rect 15291 26630 15305 26682
rect 15329 26630 15343 26682
rect 15343 26630 15355 26682
rect 15355 26630 15385 26682
rect 15409 26630 15419 26682
rect 15419 26630 15465 26682
rect 15169 26628 15225 26630
rect 15249 26628 15305 26630
rect 15329 26628 15385 26630
rect 15409 26628 15465 26630
rect 15169 25594 15225 25596
rect 15249 25594 15305 25596
rect 15329 25594 15385 25596
rect 15409 25594 15465 25596
rect 15169 25542 15215 25594
rect 15215 25542 15225 25594
rect 15249 25542 15279 25594
rect 15279 25542 15291 25594
rect 15291 25542 15305 25594
rect 15329 25542 15343 25594
rect 15343 25542 15355 25594
rect 15355 25542 15385 25594
rect 15409 25542 15419 25594
rect 15419 25542 15465 25594
rect 15169 25540 15225 25542
rect 15249 25540 15305 25542
rect 15329 25540 15385 25542
rect 15409 25540 15465 25542
rect 15169 24506 15225 24508
rect 15249 24506 15305 24508
rect 15329 24506 15385 24508
rect 15409 24506 15465 24508
rect 15169 24454 15215 24506
rect 15215 24454 15225 24506
rect 15249 24454 15279 24506
rect 15279 24454 15291 24506
rect 15291 24454 15305 24506
rect 15329 24454 15343 24506
rect 15343 24454 15355 24506
rect 15355 24454 15385 24506
rect 15409 24454 15419 24506
rect 15419 24454 15465 24506
rect 15169 24452 15225 24454
rect 15249 24452 15305 24454
rect 15329 24452 15385 24454
rect 15409 24452 15465 24454
rect 15169 23418 15225 23420
rect 15249 23418 15305 23420
rect 15329 23418 15385 23420
rect 15409 23418 15465 23420
rect 15169 23366 15215 23418
rect 15215 23366 15225 23418
rect 15249 23366 15279 23418
rect 15279 23366 15291 23418
rect 15291 23366 15305 23418
rect 15329 23366 15343 23418
rect 15343 23366 15355 23418
rect 15355 23366 15385 23418
rect 15409 23366 15419 23418
rect 15419 23366 15465 23418
rect 15169 23364 15225 23366
rect 15249 23364 15305 23366
rect 15329 23364 15385 23366
rect 15409 23364 15465 23366
rect 13726 17448 13782 17504
rect 12898 13912 12954 13968
rect 14554 19624 14610 19680
rect 15169 22330 15225 22332
rect 15249 22330 15305 22332
rect 15329 22330 15385 22332
rect 15409 22330 15465 22332
rect 15169 22278 15215 22330
rect 15215 22278 15225 22330
rect 15249 22278 15279 22330
rect 15279 22278 15291 22330
rect 15291 22278 15305 22330
rect 15329 22278 15343 22330
rect 15343 22278 15355 22330
rect 15355 22278 15385 22330
rect 15409 22278 15419 22330
rect 15419 22278 15465 22330
rect 15169 22276 15225 22278
rect 15249 22276 15305 22278
rect 15329 22276 15385 22278
rect 15409 22276 15465 22278
rect 15382 21664 15438 21720
rect 15169 21242 15225 21244
rect 15249 21242 15305 21244
rect 15329 21242 15385 21244
rect 15409 21242 15465 21244
rect 15169 21190 15215 21242
rect 15215 21190 15225 21242
rect 15249 21190 15279 21242
rect 15279 21190 15291 21242
rect 15291 21190 15305 21242
rect 15329 21190 15343 21242
rect 15343 21190 15355 21242
rect 15355 21190 15385 21242
rect 15409 21190 15419 21242
rect 15419 21190 15465 21242
rect 15169 21188 15225 21190
rect 15249 21188 15305 21190
rect 15329 21188 15385 21190
rect 15409 21188 15465 21190
rect 14830 19896 14886 19952
rect 15014 20340 15016 20360
rect 15016 20340 15068 20360
rect 15068 20340 15070 20360
rect 15014 20304 15070 20340
rect 15169 20154 15225 20156
rect 15249 20154 15305 20156
rect 15329 20154 15385 20156
rect 15409 20154 15465 20156
rect 15169 20102 15215 20154
rect 15215 20102 15225 20154
rect 15249 20102 15279 20154
rect 15279 20102 15291 20154
rect 15291 20102 15305 20154
rect 15329 20102 15343 20154
rect 15343 20102 15355 20154
rect 15355 20102 15385 20154
rect 15409 20102 15419 20154
rect 15419 20102 15465 20154
rect 15169 20100 15225 20102
rect 15249 20100 15305 20102
rect 15329 20100 15385 20102
rect 15409 20100 15465 20102
rect 15474 19896 15530 19952
rect 15169 19066 15225 19068
rect 15249 19066 15305 19068
rect 15329 19066 15385 19068
rect 15409 19066 15465 19068
rect 15169 19014 15215 19066
rect 15215 19014 15225 19066
rect 15249 19014 15279 19066
rect 15279 19014 15291 19066
rect 15291 19014 15305 19066
rect 15329 19014 15343 19066
rect 15343 19014 15355 19066
rect 15355 19014 15385 19066
rect 15409 19014 15419 19066
rect 15419 19014 15465 19066
rect 15169 19012 15225 19014
rect 15249 19012 15305 19014
rect 15329 19012 15385 19014
rect 15409 19012 15465 19014
rect 16578 29028 16634 29064
rect 16578 29008 16580 29028
rect 16580 29008 16632 29028
rect 16632 29008 16634 29028
rect 17590 29416 17646 29472
rect 17406 29008 17462 29064
rect 18786 29008 18842 29064
rect 16210 27920 16266 27976
rect 16394 27396 16450 27432
rect 16394 27376 16396 27396
rect 16396 27376 16448 27396
rect 16448 27376 16450 27396
rect 16302 21664 16358 21720
rect 15169 17978 15225 17980
rect 15249 17978 15305 17980
rect 15329 17978 15385 17980
rect 15409 17978 15465 17980
rect 15169 17926 15215 17978
rect 15215 17926 15225 17978
rect 15249 17926 15279 17978
rect 15279 17926 15291 17978
rect 15291 17926 15305 17978
rect 15329 17926 15343 17978
rect 15343 17926 15355 17978
rect 15355 17926 15385 17978
rect 15409 17926 15419 17978
rect 15419 17926 15465 17978
rect 15169 17924 15225 17926
rect 15249 17924 15305 17926
rect 15329 17924 15385 17926
rect 15409 17924 15465 17926
rect 15169 16890 15225 16892
rect 15249 16890 15305 16892
rect 15329 16890 15385 16892
rect 15409 16890 15465 16892
rect 15169 16838 15215 16890
rect 15215 16838 15225 16890
rect 15249 16838 15279 16890
rect 15279 16838 15291 16890
rect 15291 16838 15305 16890
rect 15329 16838 15343 16890
rect 15343 16838 15355 16890
rect 15355 16838 15385 16890
rect 15409 16838 15419 16890
rect 15419 16838 15465 16890
rect 15169 16836 15225 16838
rect 15249 16836 15305 16838
rect 15329 16836 15385 16838
rect 15409 16836 15465 16838
rect 15169 15802 15225 15804
rect 15249 15802 15305 15804
rect 15329 15802 15385 15804
rect 15409 15802 15465 15804
rect 15169 15750 15215 15802
rect 15215 15750 15225 15802
rect 15249 15750 15279 15802
rect 15279 15750 15291 15802
rect 15291 15750 15305 15802
rect 15329 15750 15343 15802
rect 15343 15750 15355 15802
rect 15355 15750 15385 15802
rect 15409 15750 15419 15802
rect 15419 15750 15465 15802
rect 15169 15748 15225 15750
rect 15249 15748 15305 15750
rect 15329 15748 15385 15750
rect 15409 15748 15465 15750
rect 15169 14714 15225 14716
rect 15249 14714 15305 14716
rect 15329 14714 15385 14716
rect 15409 14714 15465 14716
rect 15169 14662 15215 14714
rect 15215 14662 15225 14714
rect 15249 14662 15279 14714
rect 15279 14662 15291 14714
rect 15291 14662 15305 14714
rect 15329 14662 15343 14714
rect 15343 14662 15355 14714
rect 15355 14662 15385 14714
rect 15409 14662 15419 14714
rect 15419 14662 15465 14714
rect 15169 14660 15225 14662
rect 15249 14660 15305 14662
rect 15329 14660 15385 14662
rect 15409 14660 15465 14662
rect 15169 13626 15225 13628
rect 15249 13626 15305 13628
rect 15329 13626 15385 13628
rect 15409 13626 15465 13628
rect 15169 13574 15215 13626
rect 15215 13574 15225 13626
rect 15249 13574 15279 13626
rect 15279 13574 15291 13626
rect 15291 13574 15305 13626
rect 15329 13574 15343 13626
rect 15343 13574 15355 13626
rect 15355 13574 15385 13626
rect 15409 13574 15419 13626
rect 15419 13574 15465 13626
rect 15169 13572 15225 13574
rect 15249 13572 15305 13574
rect 15329 13572 15385 13574
rect 15409 13572 15465 13574
rect 16854 19488 16910 19544
rect 15934 15972 15990 16008
rect 15934 15952 15936 15972
rect 15936 15952 15988 15972
rect 15988 15952 15990 15972
rect 15658 13932 15714 13968
rect 15658 13912 15660 13932
rect 15660 13912 15712 13932
rect 15712 13912 15714 13932
rect 15169 12538 15225 12540
rect 15249 12538 15305 12540
rect 15329 12538 15385 12540
rect 15409 12538 15465 12540
rect 15169 12486 15215 12538
rect 15215 12486 15225 12538
rect 15249 12486 15279 12538
rect 15279 12486 15291 12538
rect 15291 12486 15305 12538
rect 15329 12486 15343 12538
rect 15343 12486 15355 12538
rect 15355 12486 15385 12538
rect 15409 12486 15419 12538
rect 15419 12486 15465 12538
rect 15169 12484 15225 12486
rect 15249 12484 15305 12486
rect 15329 12484 15385 12486
rect 15409 12484 15465 12486
rect 15169 11450 15225 11452
rect 15249 11450 15305 11452
rect 15329 11450 15385 11452
rect 15409 11450 15465 11452
rect 15169 11398 15215 11450
rect 15215 11398 15225 11450
rect 15249 11398 15279 11450
rect 15279 11398 15291 11450
rect 15291 11398 15305 11450
rect 15329 11398 15343 11450
rect 15343 11398 15355 11450
rect 15355 11398 15385 11450
rect 15409 11398 15419 11450
rect 15419 11398 15465 11450
rect 15169 11396 15225 11398
rect 15249 11396 15305 11398
rect 15329 11396 15385 11398
rect 15409 11396 15465 11398
rect 15169 10362 15225 10364
rect 15249 10362 15305 10364
rect 15329 10362 15385 10364
rect 15409 10362 15465 10364
rect 15169 10310 15215 10362
rect 15215 10310 15225 10362
rect 15249 10310 15279 10362
rect 15279 10310 15291 10362
rect 15291 10310 15305 10362
rect 15329 10310 15343 10362
rect 15343 10310 15355 10362
rect 15355 10310 15385 10362
rect 15409 10310 15419 10362
rect 15419 10310 15465 10362
rect 15169 10308 15225 10310
rect 15249 10308 15305 10310
rect 15329 10308 15385 10310
rect 15409 10308 15465 10310
rect 15169 9274 15225 9276
rect 15249 9274 15305 9276
rect 15329 9274 15385 9276
rect 15409 9274 15465 9276
rect 15169 9222 15215 9274
rect 15215 9222 15225 9274
rect 15249 9222 15279 9274
rect 15279 9222 15291 9274
rect 15291 9222 15305 9274
rect 15329 9222 15343 9274
rect 15343 9222 15355 9274
rect 15355 9222 15385 9274
rect 15409 9222 15419 9274
rect 15419 9222 15465 9274
rect 15169 9220 15225 9222
rect 15249 9220 15305 9222
rect 15329 9220 15385 9222
rect 15409 9220 15465 9222
rect 10431 3290 10487 3292
rect 10511 3290 10567 3292
rect 10591 3290 10647 3292
rect 10671 3290 10727 3292
rect 10431 3238 10477 3290
rect 10477 3238 10487 3290
rect 10511 3238 10541 3290
rect 10541 3238 10553 3290
rect 10553 3238 10567 3290
rect 10591 3238 10605 3290
rect 10605 3238 10617 3290
rect 10617 3238 10647 3290
rect 10671 3238 10681 3290
rect 10681 3238 10727 3290
rect 10431 3236 10487 3238
rect 10511 3236 10567 3238
rect 10591 3236 10647 3238
rect 10671 3236 10727 3238
rect 10431 2202 10487 2204
rect 10511 2202 10567 2204
rect 10591 2202 10647 2204
rect 10671 2202 10727 2204
rect 10431 2150 10477 2202
rect 10477 2150 10487 2202
rect 10511 2150 10541 2202
rect 10541 2150 10553 2202
rect 10553 2150 10567 2202
rect 10591 2150 10605 2202
rect 10605 2150 10617 2202
rect 10617 2150 10647 2202
rect 10671 2150 10681 2202
rect 10681 2150 10727 2202
rect 10431 2148 10487 2150
rect 10511 2148 10567 2150
rect 10591 2148 10647 2150
rect 10671 2148 10727 2150
rect 14462 3168 14518 3224
rect 15750 8372 15752 8392
rect 15752 8372 15804 8392
rect 15804 8372 15806 8392
rect 15750 8336 15806 8372
rect 15169 8186 15225 8188
rect 15249 8186 15305 8188
rect 15329 8186 15385 8188
rect 15409 8186 15465 8188
rect 15169 8134 15215 8186
rect 15215 8134 15225 8186
rect 15249 8134 15279 8186
rect 15279 8134 15291 8186
rect 15291 8134 15305 8186
rect 15329 8134 15343 8186
rect 15343 8134 15355 8186
rect 15355 8134 15385 8186
rect 15409 8134 15419 8186
rect 15419 8134 15465 8186
rect 15169 8132 15225 8134
rect 15249 8132 15305 8134
rect 15329 8132 15385 8134
rect 15409 8132 15465 8134
rect 15169 7098 15225 7100
rect 15249 7098 15305 7100
rect 15329 7098 15385 7100
rect 15409 7098 15465 7100
rect 15169 7046 15215 7098
rect 15215 7046 15225 7098
rect 15249 7046 15279 7098
rect 15279 7046 15291 7098
rect 15291 7046 15305 7098
rect 15329 7046 15343 7098
rect 15343 7046 15355 7098
rect 15355 7046 15385 7098
rect 15409 7046 15419 7098
rect 15419 7046 15465 7098
rect 15169 7044 15225 7046
rect 15249 7044 15305 7046
rect 15329 7044 15385 7046
rect 15409 7044 15465 7046
rect 15169 6010 15225 6012
rect 15249 6010 15305 6012
rect 15329 6010 15385 6012
rect 15409 6010 15465 6012
rect 15169 5958 15215 6010
rect 15215 5958 15225 6010
rect 15249 5958 15279 6010
rect 15279 5958 15291 6010
rect 15291 5958 15305 6010
rect 15329 5958 15343 6010
rect 15343 5958 15355 6010
rect 15355 5958 15385 6010
rect 15409 5958 15419 6010
rect 15419 5958 15465 6010
rect 15169 5956 15225 5958
rect 15249 5956 15305 5958
rect 15329 5956 15385 5958
rect 15409 5956 15465 5958
rect 15169 4922 15225 4924
rect 15249 4922 15305 4924
rect 15329 4922 15385 4924
rect 15409 4922 15465 4924
rect 15169 4870 15215 4922
rect 15215 4870 15225 4922
rect 15249 4870 15279 4922
rect 15279 4870 15291 4922
rect 15291 4870 15305 4922
rect 15329 4870 15343 4922
rect 15343 4870 15355 4922
rect 15355 4870 15385 4922
rect 15409 4870 15419 4922
rect 15419 4870 15465 4922
rect 15169 4868 15225 4870
rect 15249 4868 15305 4870
rect 15329 4868 15385 4870
rect 15409 4868 15465 4870
rect 15169 3834 15225 3836
rect 15249 3834 15305 3836
rect 15329 3834 15385 3836
rect 15409 3834 15465 3836
rect 15169 3782 15215 3834
rect 15215 3782 15225 3834
rect 15249 3782 15279 3834
rect 15279 3782 15291 3834
rect 15291 3782 15305 3834
rect 15329 3782 15343 3834
rect 15343 3782 15355 3834
rect 15355 3782 15385 3834
rect 15409 3782 15419 3834
rect 15419 3782 15465 3834
rect 15169 3780 15225 3782
rect 15249 3780 15305 3782
rect 15329 3780 15385 3782
rect 15409 3780 15465 3782
rect 15169 2746 15225 2748
rect 15249 2746 15305 2748
rect 15329 2746 15385 2748
rect 15409 2746 15465 2748
rect 15169 2694 15215 2746
rect 15215 2694 15225 2746
rect 15249 2694 15279 2746
rect 15279 2694 15291 2746
rect 15291 2694 15305 2746
rect 15329 2694 15343 2746
rect 15343 2694 15355 2746
rect 15355 2694 15385 2746
rect 15409 2694 15419 2746
rect 15419 2694 15465 2746
rect 15169 2692 15225 2694
rect 15249 2692 15305 2694
rect 15329 2692 15385 2694
rect 15409 2692 15465 2694
rect 16762 3304 16818 3360
rect 19907 30490 19963 30492
rect 19987 30490 20043 30492
rect 20067 30490 20123 30492
rect 20147 30490 20203 30492
rect 19907 30438 19953 30490
rect 19953 30438 19963 30490
rect 19987 30438 20017 30490
rect 20017 30438 20029 30490
rect 20029 30438 20043 30490
rect 20067 30438 20081 30490
rect 20081 30438 20093 30490
rect 20093 30438 20123 30490
rect 20147 30438 20157 30490
rect 20157 30438 20203 30490
rect 19907 30436 19963 30438
rect 19987 30436 20043 30438
rect 20067 30436 20123 30438
rect 20147 30436 20203 30438
rect 19907 29402 19963 29404
rect 19987 29402 20043 29404
rect 20067 29402 20123 29404
rect 20147 29402 20203 29404
rect 19907 29350 19953 29402
rect 19953 29350 19963 29402
rect 19987 29350 20017 29402
rect 20017 29350 20029 29402
rect 20029 29350 20043 29402
rect 20067 29350 20081 29402
rect 20081 29350 20093 29402
rect 20093 29350 20123 29402
rect 20147 29350 20157 29402
rect 20157 29350 20203 29402
rect 19907 29348 19963 29350
rect 19987 29348 20043 29350
rect 20067 29348 20123 29350
rect 20147 29348 20203 29350
rect 19907 28314 19963 28316
rect 19987 28314 20043 28316
rect 20067 28314 20123 28316
rect 20147 28314 20203 28316
rect 19907 28262 19953 28314
rect 19953 28262 19963 28314
rect 19987 28262 20017 28314
rect 20017 28262 20029 28314
rect 20029 28262 20043 28314
rect 20067 28262 20081 28314
rect 20081 28262 20093 28314
rect 20093 28262 20123 28314
rect 20147 28262 20157 28314
rect 20157 28262 20203 28314
rect 19907 28260 19963 28262
rect 19987 28260 20043 28262
rect 20067 28260 20123 28262
rect 20147 28260 20203 28262
rect 19907 27226 19963 27228
rect 19987 27226 20043 27228
rect 20067 27226 20123 27228
rect 20147 27226 20203 27228
rect 19907 27174 19953 27226
rect 19953 27174 19963 27226
rect 19987 27174 20017 27226
rect 20017 27174 20029 27226
rect 20029 27174 20043 27226
rect 20067 27174 20081 27226
rect 20081 27174 20093 27226
rect 20093 27174 20123 27226
rect 20147 27174 20157 27226
rect 20157 27174 20203 27226
rect 19907 27172 19963 27174
rect 19987 27172 20043 27174
rect 20067 27172 20123 27174
rect 20147 27172 20203 27174
rect 19907 26138 19963 26140
rect 19987 26138 20043 26140
rect 20067 26138 20123 26140
rect 20147 26138 20203 26140
rect 19907 26086 19953 26138
rect 19953 26086 19963 26138
rect 19987 26086 20017 26138
rect 20017 26086 20029 26138
rect 20029 26086 20043 26138
rect 20067 26086 20081 26138
rect 20081 26086 20093 26138
rect 20093 26086 20123 26138
rect 20147 26086 20157 26138
rect 20157 26086 20203 26138
rect 19907 26084 19963 26086
rect 19987 26084 20043 26086
rect 20067 26084 20123 26086
rect 20147 26084 20203 26086
rect 19614 25236 19616 25256
rect 19616 25236 19668 25256
rect 19668 25236 19670 25256
rect 19614 25200 19670 25236
rect 19907 25050 19963 25052
rect 19987 25050 20043 25052
rect 20067 25050 20123 25052
rect 20147 25050 20203 25052
rect 19907 24998 19953 25050
rect 19953 24998 19963 25050
rect 19987 24998 20017 25050
rect 20017 24998 20029 25050
rect 20029 24998 20043 25050
rect 20067 24998 20081 25050
rect 20081 24998 20093 25050
rect 20093 24998 20123 25050
rect 20147 24998 20157 25050
rect 20157 24998 20203 25050
rect 19907 24996 19963 24998
rect 19987 24996 20043 24998
rect 20067 24996 20123 24998
rect 20147 24996 20203 24998
rect 18234 23724 18290 23760
rect 18234 23704 18236 23724
rect 18236 23704 18288 23724
rect 18288 23704 18290 23724
rect 19338 23724 19394 23760
rect 19338 23704 19340 23724
rect 19340 23704 19392 23724
rect 19392 23704 19394 23724
rect 18694 23432 18750 23488
rect 17130 8236 17132 8256
rect 17132 8236 17184 8256
rect 17184 8236 17186 8256
rect 17130 8200 17186 8236
rect 17498 8880 17554 8936
rect 17682 8744 17738 8800
rect 18234 19760 18290 19816
rect 19907 23962 19963 23964
rect 19987 23962 20043 23964
rect 20067 23962 20123 23964
rect 20147 23962 20203 23964
rect 19907 23910 19953 23962
rect 19953 23910 19963 23962
rect 19987 23910 20017 23962
rect 20017 23910 20029 23962
rect 20029 23910 20043 23962
rect 20067 23910 20081 23962
rect 20081 23910 20093 23962
rect 20093 23910 20123 23962
rect 20147 23910 20157 23962
rect 20157 23910 20203 23962
rect 19907 23908 19963 23910
rect 19987 23908 20043 23910
rect 20067 23908 20123 23910
rect 20147 23908 20203 23910
rect 20166 23568 20222 23624
rect 19982 23432 20038 23488
rect 18694 19488 18750 19544
rect 19246 19624 19302 19680
rect 19907 22874 19963 22876
rect 19987 22874 20043 22876
rect 20067 22874 20123 22876
rect 20147 22874 20203 22876
rect 19907 22822 19953 22874
rect 19953 22822 19963 22874
rect 19987 22822 20017 22874
rect 20017 22822 20029 22874
rect 20029 22822 20043 22874
rect 20067 22822 20081 22874
rect 20081 22822 20093 22874
rect 20093 22822 20123 22874
rect 20147 22822 20157 22874
rect 20157 22822 20203 22874
rect 19907 22820 19963 22822
rect 19987 22820 20043 22822
rect 20067 22820 20123 22822
rect 20147 22820 20203 22822
rect 19338 16904 19394 16960
rect 18510 15544 18566 15600
rect 18970 15544 19026 15600
rect 17774 8372 17776 8392
rect 17776 8372 17828 8392
rect 17828 8372 17830 8392
rect 17774 8336 17830 8372
rect 17222 3712 17278 3768
rect 17774 4120 17830 4176
rect 17590 3440 17646 3496
rect 19522 19352 19578 19408
rect 19907 21786 19963 21788
rect 19987 21786 20043 21788
rect 20067 21786 20123 21788
rect 20147 21786 20203 21788
rect 19907 21734 19953 21786
rect 19953 21734 19963 21786
rect 19987 21734 20017 21786
rect 20017 21734 20029 21786
rect 20029 21734 20043 21786
rect 20067 21734 20081 21786
rect 20081 21734 20093 21786
rect 20093 21734 20123 21786
rect 20147 21734 20157 21786
rect 20157 21734 20203 21786
rect 19907 21732 19963 21734
rect 19987 21732 20043 21734
rect 20067 21732 20123 21734
rect 20147 21732 20203 21734
rect 20166 20884 20168 20904
rect 20168 20884 20220 20904
rect 20220 20884 20222 20904
rect 20166 20848 20222 20884
rect 19907 20698 19963 20700
rect 19987 20698 20043 20700
rect 20067 20698 20123 20700
rect 20147 20698 20203 20700
rect 19907 20646 19953 20698
rect 19953 20646 19963 20698
rect 19987 20646 20017 20698
rect 20017 20646 20029 20698
rect 20029 20646 20043 20698
rect 20067 20646 20081 20698
rect 20081 20646 20093 20698
rect 20093 20646 20123 20698
rect 20147 20646 20157 20698
rect 20157 20646 20203 20698
rect 19907 20644 19963 20646
rect 19987 20644 20043 20646
rect 20067 20644 20123 20646
rect 20147 20644 20203 20646
rect 19907 19610 19963 19612
rect 19987 19610 20043 19612
rect 20067 19610 20123 19612
rect 20147 19610 20203 19612
rect 19907 19558 19953 19610
rect 19953 19558 19963 19610
rect 19987 19558 20017 19610
rect 20017 19558 20029 19610
rect 20029 19558 20043 19610
rect 20067 19558 20081 19610
rect 20081 19558 20093 19610
rect 20093 19558 20123 19610
rect 20147 19558 20157 19610
rect 20157 19558 20203 19610
rect 19907 19556 19963 19558
rect 19987 19556 20043 19558
rect 20067 19556 20123 19558
rect 20147 19556 20203 19558
rect 19907 18522 19963 18524
rect 19987 18522 20043 18524
rect 20067 18522 20123 18524
rect 20147 18522 20203 18524
rect 19907 18470 19953 18522
rect 19953 18470 19963 18522
rect 19987 18470 20017 18522
rect 20017 18470 20029 18522
rect 20029 18470 20043 18522
rect 20067 18470 20081 18522
rect 20081 18470 20093 18522
rect 20093 18470 20123 18522
rect 20147 18470 20157 18522
rect 20157 18470 20203 18522
rect 19907 18468 19963 18470
rect 19987 18468 20043 18470
rect 20067 18468 20123 18470
rect 20147 18468 20203 18470
rect 19907 17434 19963 17436
rect 19987 17434 20043 17436
rect 20067 17434 20123 17436
rect 20147 17434 20203 17436
rect 19907 17382 19953 17434
rect 19953 17382 19963 17434
rect 19987 17382 20017 17434
rect 20017 17382 20029 17434
rect 20029 17382 20043 17434
rect 20067 17382 20081 17434
rect 20081 17382 20093 17434
rect 20093 17382 20123 17434
rect 20147 17382 20157 17434
rect 20157 17382 20203 17434
rect 19907 17380 19963 17382
rect 19987 17380 20043 17382
rect 20067 17380 20123 17382
rect 20147 17380 20203 17382
rect 19522 16088 19578 16144
rect 19907 16346 19963 16348
rect 19987 16346 20043 16348
rect 20067 16346 20123 16348
rect 20147 16346 20203 16348
rect 19907 16294 19953 16346
rect 19953 16294 19963 16346
rect 19987 16294 20017 16346
rect 20017 16294 20029 16346
rect 20029 16294 20043 16346
rect 20067 16294 20081 16346
rect 20081 16294 20093 16346
rect 20093 16294 20123 16346
rect 20147 16294 20157 16346
rect 20157 16294 20203 16346
rect 19907 16292 19963 16294
rect 19987 16292 20043 16294
rect 20067 16292 20123 16294
rect 20147 16292 20203 16294
rect 19907 15258 19963 15260
rect 19987 15258 20043 15260
rect 20067 15258 20123 15260
rect 20147 15258 20203 15260
rect 19907 15206 19953 15258
rect 19953 15206 19963 15258
rect 19987 15206 20017 15258
rect 20017 15206 20029 15258
rect 20029 15206 20043 15258
rect 20067 15206 20081 15258
rect 20081 15206 20093 15258
rect 20093 15206 20123 15258
rect 20147 15206 20157 15258
rect 20157 15206 20203 15258
rect 19907 15204 19963 15206
rect 19987 15204 20043 15206
rect 20067 15204 20123 15206
rect 20147 15204 20203 15206
rect 19907 14170 19963 14172
rect 19987 14170 20043 14172
rect 20067 14170 20123 14172
rect 20147 14170 20203 14172
rect 19907 14118 19953 14170
rect 19953 14118 19963 14170
rect 19987 14118 20017 14170
rect 20017 14118 20029 14170
rect 20029 14118 20043 14170
rect 20067 14118 20081 14170
rect 20081 14118 20093 14170
rect 20093 14118 20123 14170
rect 20147 14118 20157 14170
rect 20157 14118 20203 14170
rect 19907 14116 19963 14118
rect 19987 14116 20043 14118
rect 20067 14116 20123 14118
rect 20147 14116 20203 14118
rect 19907 13082 19963 13084
rect 19987 13082 20043 13084
rect 20067 13082 20123 13084
rect 20147 13082 20203 13084
rect 19907 13030 19953 13082
rect 19953 13030 19963 13082
rect 19987 13030 20017 13082
rect 20017 13030 20029 13082
rect 20029 13030 20043 13082
rect 20067 13030 20081 13082
rect 20081 13030 20093 13082
rect 20093 13030 20123 13082
rect 20147 13030 20157 13082
rect 20157 13030 20203 13082
rect 19907 13028 19963 13030
rect 19987 13028 20043 13030
rect 20067 13028 20123 13030
rect 20147 13028 20203 13030
rect 19907 11994 19963 11996
rect 19987 11994 20043 11996
rect 20067 11994 20123 11996
rect 20147 11994 20203 11996
rect 19907 11942 19953 11994
rect 19953 11942 19963 11994
rect 19987 11942 20017 11994
rect 20017 11942 20029 11994
rect 20029 11942 20043 11994
rect 20067 11942 20081 11994
rect 20081 11942 20093 11994
rect 20093 11942 20123 11994
rect 20147 11942 20157 11994
rect 20157 11942 20203 11994
rect 19907 11940 19963 11942
rect 19987 11940 20043 11942
rect 20067 11940 20123 11942
rect 20147 11940 20203 11942
rect 19907 10906 19963 10908
rect 19987 10906 20043 10908
rect 20067 10906 20123 10908
rect 20147 10906 20203 10908
rect 19907 10854 19953 10906
rect 19953 10854 19963 10906
rect 19987 10854 20017 10906
rect 20017 10854 20029 10906
rect 20029 10854 20043 10906
rect 20067 10854 20081 10906
rect 20081 10854 20093 10906
rect 20093 10854 20123 10906
rect 20147 10854 20157 10906
rect 20157 10854 20203 10906
rect 19907 10852 19963 10854
rect 19987 10852 20043 10854
rect 20067 10852 20123 10854
rect 20147 10852 20203 10854
rect 20626 17856 20682 17912
rect 24645 29946 24701 29948
rect 24725 29946 24781 29948
rect 24805 29946 24861 29948
rect 24885 29946 24941 29948
rect 24645 29894 24691 29946
rect 24691 29894 24701 29946
rect 24725 29894 24755 29946
rect 24755 29894 24767 29946
rect 24767 29894 24781 29946
rect 24805 29894 24819 29946
rect 24819 29894 24831 29946
rect 24831 29894 24861 29946
rect 24885 29894 24895 29946
rect 24895 29894 24941 29946
rect 24645 29892 24701 29894
rect 24725 29892 24781 29894
rect 24805 29892 24861 29894
rect 24885 29892 24941 29894
rect 24645 28858 24701 28860
rect 24725 28858 24781 28860
rect 24805 28858 24861 28860
rect 24885 28858 24941 28860
rect 24645 28806 24691 28858
rect 24691 28806 24701 28858
rect 24725 28806 24755 28858
rect 24755 28806 24767 28858
rect 24767 28806 24781 28858
rect 24805 28806 24819 28858
rect 24819 28806 24831 28858
rect 24831 28806 24861 28858
rect 24885 28806 24895 28858
rect 24895 28806 24941 28858
rect 24645 28804 24701 28806
rect 24725 28804 24781 28806
rect 24805 28804 24861 28806
rect 24885 28804 24941 28806
rect 24645 27770 24701 27772
rect 24725 27770 24781 27772
rect 24805 27770 24861 27772
rect 24885 27770 24941 27772
rect 24645 27718 24691 27770
rect 24691 27718 24701 27770
rect 24725 27718 24755 27770
rect 24755 27718 24767 27770
rect 24767 27718 24781 27770
rect 24805 27718 24819 27770
rect 24819 27718 24831 27770
rect 24831 27718 24861 27770
rect 24885 27718 24895 27770
rect 24895 27718 24941 27770
rect 24645 27716 24701 27718
rect 24725 27716 24781 27718
rect 24805 27716 24861 27718
rect 24885 27716 24941 27718
rect 24645 26682 24701 26684
rect 24725 26682 24781 26684
rect 24805 26682 24861 26684
rect 24885 26682 24941 26684
rect 24645 26630 24691 26682
rect 24691 26630 24701 26682
rect 24725 26630 24755 26682
rect 24755 26630 24767 26682
rect 24767 26630 24781 26682
rect 24805 26630 24819 26682
rect 24819 26630 24831 26682
rect 24831 26630 24861 26682
rect 24885 26630 24895 26682
rect 24895 26630 24941 26682
rect 24645 26628 24701 26630
rect 24725 26628 24781 26630
rect 24805 26628 24861 26630
rect 24885 26628 24941 26630
rect 21546 20848 21602 20904
rect 19907 9818 19963 9820
rect 19987 9818 20043 9820
rect 20067 9818 20123 9820
rect 20147 9818 20203 9820
rect 19907 9766 19953 9818
rect 19953 9766 19963 9818
rect 19987 9766 20017 9818
rect 20017 9766 20029 9818
rect 20029 9766 20043 9818
rect 20067 9766 20081 9818
rect 20081 9766 20093 9818
rect 20093 9766 20123 9818
rect 20147 9766 20157 9818
rect 20157 9766 20203 9818
rect 19907 9764 19963 9766
rect 19987 9764 20043 9766
rect 20067 9764 20123 9766
rect 20147 9764 20203 9766
rect 18602 8200 18658 8256
rect 19907 8730 19963 8732
rect 19987 8730 20043 8732
rect 20067 8730 20123 8732
rect 20147 8730 20203 8732
rect 19907 8678 19953 8730
rect 19953 8678 19963 8730
rect 19987 8678 20017 8730
rect 20017 8678 20029 8730
rect 20029 8678 20043 8730
rect 20067 8678 20081 8730
rect 20081 8678 20093 8730
rect 20093 8678 20123 8730
rect 20147 8678 20157 8730
rect 20157 8678 20203 8730
rect 19907 8676 19963 8678
rect 19987 8676 20043 8678
rect 20067 8676 20123 8678
rect 20147 8676 20203 8678
rect 19907 7642 19963 7644
rect 19987 7642 20043 7644
rect 20067 7642 20123 7644
rect 20147 7642 20203 7644
rect 19907 7590 19953 7642
rect 19953 7590 19963 7642
rect 19987 7590 20017 7642
rect 20017 7590 20029 7642
rect 20029 7590 20043 7642
rect 20067 7590 20081 7642
rect 20081 7590 20093 7642
rect 20093 7590 20123 7642
rect 20147 7590 20157 7642
rect 20157 7590 20203 7642
rect 19907 7588 19963 7590
rect 19987 7588 20043 7590
rect 20067 7588 20123 7590
rect 20147 7588 20203 7590
rect 19907 6554 19963 6556
rect 19987 6554 20043 6556
rect 20067 6554 20123 6556
rect 20147 6554 20203 6556
rect 19907 6502 19953 6554
rect 19953 6502 19963 6554
rect 19987 6502 20017 6554
rect 20017 6502 20029 6554
rect 20029 6502 20043 6554
rect 20067 6502 20081 6554
rect 20081 6502 20093 6554
rect 20093 6502 20123 6554
rect 20147 6502 20157 6554
rect 20157 6502 20203 6554
rect 19907 6500 19963 6502
rect 19987 6500 20043 6502
rect 20067 6500 20123 6502
rect 20147 6500 20203 6502
rect 21086 14864 21142 14920
rect 27342 32000 27398 32056
rect 26882 30640 26938 30696
rect 24645 25594 24701 25596
rect 24725 25594 24781 25596
rect 24805 25594 24861 25596
rect 24885 25594 24941 25596
rect 24645 25542 24691 25594
rect 24691 25542 24701 25594
rect 24725 25542 24755 25594
rect 24755 25542 24767 25594
rect 24767 25542 24781 25594
rect 24805 25542 24819 25594
rect 24819 25542 24831 25594
rect 24831 25542 24861 25594
rect 24885 25542 24895 25594
rect 24895 25542 24941 25594
rect 24645 25540 24701 25542
rect 24725 25540 24781 25542
rect 24805 25540 24861 25542
rect 24885 25540 24941 25542
rect 24645 24506 24701 24508
rect 24725 24506 24781 24508
rect 24805 24506 24861 24508
rect 24885 24506 24941 24508
rect 24645 24454 24691 24506
rect 24691 24454 24701 24506
rect 24725 24454 24755 24506
rect 24755 24454 24767 24506
rect 24767 24454 24781 24506
rect 24805 24454 24819 24506
rect 24819 24454 24831 24506
rect 24831 24454 24861 24506
rect 24885 24454 24895 24506
rect 24895 24454 24941 24506
rect 24645 24452 24701 24454
rect 24725 24452 24781 24454
rect 24805 24452 24861 24454
rect 24885 24452 24941 24454
rect 23754 20848 23810 20904
rect 23662 20304 23718 20360
rect 22098 15000 22154 15056
rect 22558 14864 22614 14920
rect 21914 13368 21970 13424
rect 19907 5466 19963 5468
rect 19987 5466 20043 5468
rect 20067 5466 20123 5468
rect 20147 5466 20203 5468
rect 19907 5414 19953 5466
rect 19953 5414 19963 5466
rect 19987 5414 20017 5466
rect 20017 5414 20029 5466
rect 20029 5414 20043 5466
rect 20067 5414 20081 5466
rect 20081 5414 20093 5466
rect 20093 5414 20123 5466
rect 20147 5414 20157 5466
rect 20157 5414 20203 5466
rect 19907 5412 19963 5414
rect 19987 5412 20043 5414
rect 20067 5412 20123 5414
rect 20147 5412 20203 5414
rect 18326 4140 18382 4176
rect 18326 4120 18328 4140
rect 18328 4120 18380 4140
rect 18380 4120 18382 4140
rect 18878 3732 18934 3768
rect 18878 3712 18880 3732
rect 18880 3712 18932 3732
rect 18932 3712 18934 3732
rect 18878 3304 18934 3360
rect 18970 3168 19026 3224
rect 19706 5072 19762 5128
rect 19614 3984 19670 4040
rect 19907 4378 19963 4380
rect 19987 4378 20043 4380
rect 20067 4378 20123 4380
rect 20147 4378 20203 4380
rect 19907 4326 19953 4378
rect 19953 4326 19963 4378
rect 19987 4326 20017 4378
rect 20017 4326 20029 4378
rect 20029 4326 20043 4378
rect 20067 4326 20081 4378
rect 20081 4326 20093 4378
rect 20093 4326 20123 4378
rect 20147 4326 20157 4378
rect 20157 4326 20203 4378
rect 19907 4324 19963 4326
rect 19987 4324 20043 4326
rect 20067 4324 20123 4326
rect 20147 4324 20203 4326
rect 19907 3290 19963 3292
rect 19987 3290 20043 3292
rect 20067 3290 20123 3292
rect 20147 3290 20203 3292
rect 19907 3238 19953 3290
rect 19953 3238 19963 3290
rect 19987 3238 20017 3290
rect 20017 3238 20029 3290
rect 20029 3238 20043 3290
rect 20067 3238 20081 3290
rect 20081 3238 20093 3290
rect 20093 3238 20123 3290
rect 20147 3238 20157 3290
rect 20157 3238 20203 3290
rect 19907 3236 19963 3238
rect 19987 3236 20043 3238
rect 20067 3236 20123 3238
rect 20147 3236 20203 3238
rect 19907 2202 19963 2204
rect 19987 2202 20043 2204
rect 20067 2202 20123 2204
rect 20147 2202 20203 2204
rect 19907 2150 19953 2202
rect 19953 2150 19963 2202
rect 19987 2150 20017 2202
rect 20017 2150 20029 2202
rect 20029 2150 20043 2202
rect 20067 2150 20081 2202
rect 20081 2150 20093 2202
rect 20093 2150 20123 2202
rect 20147 2150 20157 2202
rect 20157 2150 20203 2202
rect 19907 2148 19963 2150
rect 19987 2148 20043 2150
rect 20067 2148 20123 2150
rect 20147 2148 20203 2150
rect 23294 19760 23350 19816
rect 24645 23418 24701 23420
rect 24725 23418 24781 23420
rect 24805 23418 24861 23420
rect 24885 23418 24941 23420
rect 24645 23366 24691 23418
rect 24691 23366 24701 23418
rect 24725 23366 24755 23418
rect 24755 23366 24767 23418
rect 24767 23366 24781 23418
rect 24805 23366 24819 23418
rect 24819 23366 24831 23418
rect 24831 23366 24861 23418
rect 24885 23366 24895 23418
rect 24895 23366 24941 23418
rect 24645 23364 24701 23366
rect 24725 23364 24781 23366
rect 24805 23364 24861 23366
rect 24885 23364 24941 23366
rect 26698 24656 26754 24712
rect 24645 22330 24701 22332
rect 24725 22330 24781 22332
rect 24805 22330 24861 22332
rect 24885 22330 24941 22332
rect 24645 22278 24691 22330
rect 24691 22278 24701 22330
rect 24725 22278 24755 22330
rect 24755 22278 24767 22330
rect 24767 22278 24781 22330
rect 24805 22278 24819 22330
rect 24819 22278 24831 22330
rect 24831 22278 24861 22330
rect 24885 22278 24895 22330
rect 24895 22278 24941 22330
rect 24645 22276 24701 22278
rect 24725 22276 24781 22278
rect 24805 22276 24861 22278
rect 24885 22276 24941 22278
rect 27434 29144 27490 29200
rect 27526 27648 27582 27704
rect 27526 26152 27582 26208
rect 27434 23160 27490 23216
rect 24645 21242 24701 21244
rect 24725 21242 24781 21244
rect 24805 21242 24861 21244
rect 24885 21242 24941 21244
rect 24645 21190 24691 21242
rect 24691 21190 24701 21242
rect 24725 21190 24755 21242
rect 24755 21190 24767 21242
rect 24767 21190 24781 21242
rect 24805 21190 24819 21242
rect 24819 21190 24831 21242
rect 24831 21190 24861 21242
rect 24885 21190 24895 21242
rect 24895 21190 24941 21242
rect 24645 21188 24701 21190
rect 24725 21188 24781 21190
rect 24805 21188 24861 21190
rect 24885 21188 24941 21190
rect 24645 20154 24701 20156
rect 24725 20154 24781 20156
rect 24805 20154 24861 20156
rect 24885 20154 24941 20156
rect 24645 20102 24691 20154
rect 24691 20102 24701 20154
rect 24725 20102 24755 20154
rect 24755 20102 24767 20154
rect 24767 20102 24781 20154
rect 24805 20102 24819 20154
rect 24819 20102 24831 20154
rect 24831 20102 24861 20154
rect 24885 20102 24895 20154
rect 24895 20102 24941 20154
rect 24645 20100 24701 20102
rect 24725 20100 24781 20102
rect 24805 20100 24861 20102
rect 24885 20100 24941 20102
rect 25042 19796 25044 19816
rect 25044 19796 25096 19816
rect 25096 19796 25098 19816
rect 25042 19760 25098 19796
rect 24645 19066 24701 19068
rect 24725 19066 24781 19068
rect 24805 19066 24861 19068
rect 24885 19066 24941 19068
rect 24645 19014 24691 19066
rect 24691 19014 24701 19066
rect 24725 19014 24755 19066
rect 24755 19014 24767 19066
rect 24767 19014 24781 19066
rect 24805 19014 24819 19066
rect 24819 19014 24831 19066
rect 24831 19014 24861 19066
rect 24885 19014 24895 19066
rect 24895 19014 24941 19066
rect 24645 19012 24701 19014
rect 24725 19012 24781 19014
rect 24805 19012 24861 19014
rect 24885 19012 24941 19014
rect 24645 17978 24701 17980
rect 24725 17978 24781 17980
rect 24805 17978 24861 17980
rect 24885 17978 24941 17980
rect 24645 17926 24691 17978
rect 24691 17926 24701 17978
rect 24725 17926 24755 17978
rect 24755 17926 24767 17978
rect 24767 17926 24781 17978
rect 24805 17926 24819 17978
rect 24819 17926 24831 17978
rect 24831 17926 24861 17978
rect 24885 17926 24895 17978
rect 24895 17926 24941 17978
rect 24645 17924 24701 17926
rect 24725 17924 24781 17926
rect 24805 17924 24861 17926
rect 24885 17924 24941 17926
rect 24645 16890 24701 16892
rect 24725 16890 24781 16892
rect 24805 16890 24861 16892
rect 24885 16890 24941 16892
rect 24645 16838 24691 16890
rect 24691 16838 24701 16890
rect 24725 16838 24755 16890
rect 24755 16838 24767 16890
rect 24767 16838 24781 16890
rect 24805 16838 24819 16890
rect 24819 16838 24831 16890
rect 24831 16838 24861 16890
rect 24885 16838 24895 16890
rect 24895 16838 24941 16890
rect 24645 16836 24701 16838
rect 24725 16836 24781 16838
rect 24805 16836 24861 16838
rect 24885 16836 24941 16838
rect 24645 15802 24701 15804
rect 24725 15802 24781 15804
rect 24805 15802 24861 15804
rect 24885 15802 24941 15804
rect 24645 15750 24691 15802
rect 24691 15750 24701 15802
rect 24725 15750 24755 15802
rect 24755 15750 24767 15802
rect 24767 15750 24781 15802
rect 24805 15750 24819 15802
rect 24819 15750 24831 15802
rect 24831 15750 24861 15802
rect 24885 15750 24895 15802
rect 24895 15750 24941 15802
rect 24645 15748 24701 15750
rect 24725 15748 24781 15750
rect 24805 15748 24861 15750
rect 24885 15748 24941 15750
rect 24645 14714 24701 14716
rect 24725 14714 24781 14716
rect 24805 14714 24861 14716
rect 24885 14714 24941 14716
rect 24645 14662 24691 14714
rect 24691 14662 24701 14714
rect 24725 14662 24755 14714
rect 24755 14662 24767 14714
rect 24767 14662 24781 14714
rect 24805 14662 24819 14714
rect 24819 14662 24831 14714
rect 24831 14662 24861 14714
rect 24885 14662 24895 14714
rect 24895 14662 24941 14714
rect 24645 14660 24701 14662
rect 24725 14660 24781 14662
rect 24805 14660 24861 14662
rect 24885 14660 24941 14662
rect 24645 13626 24701 13628
rect 24725 13626 24781 13628
rect 24805 13626 24861 13628
rect 24885 13626 24941 13628
rect 24645 13574 24691 13626
rect 24691 13574 24701 13626
rect 24725 13574 24755 13626
rect 24755 13574 24767 13626
rect 24767 13574 24781 13626
rect 24805 13574 24819 13626
rect 24819 13574 24831 13626
rect 24831 13574 24861 13626
rect 24885 13574 24895 13626
rect 24895 13574 24941 13626
rect 24645 13572 24701 13574
rect 24725 13572 24781 13574
rect 24805 13572 24861 13574
rect 24885 13572 24941 13574
rect 24950 13368 25006 13424
rect 24645 12538 24701 12540
rect 24725 12538 24781 12540
rect 24805 12538 24861 12540
rect 24885 12538 24941 12540
rect 24645 12486 24691 12538
rect 24691 12486 24701 12538
rect 24725 12486 24755 12538
rect 24755 12486 24767 12538
rect 24767 12486 24781 12538
rect 24805 12486 24819 12538
rect 24819 12486 24831 12538
rect 24831 12486 24861 12538
rect 24885 12486 24895 12538
rect 24895 12486 24941 12538
rect 24645 12484 24701 12486
rect 24725 12484 24781 12486
rect 24805 12484 24861 12486
rect 24885 12484 24941 12486
rect 26422 20168 26478 20224
rect 24645 11450 24701 11452
rect 24725 11450 24781 11452
rect 24805 11450 24861 11452
rect 24885 11450 24941 11452
rect 24645 11398 24691 11450
rect 24691 11398 24701 11450
rect 24725 11398 24755 11450
rect 24755 11398 24767 11450
rect 24767 11398 24781 11450
rect 24805 11398 24819 11450
rect 24819 11398 24831 11450
rect 24831 11398 24861 11450
rect 24885 11398 24895 11450
rect 24895 11398 24941 11450
rect 24645 11396 24701 11398
rect 24725 11396 24781 11398
rect 24805 11396 24861 11398
rect 24885 11396 24941 11398
rect 24645 10362 24701 10364
rect 24725 10362 24781 10364
rect 24805 10362 24861 10364
rect 24885 10362 24941 10364
rect 24645 10310 24691 10362
rect 24691 10310 24701 10362
rect 24725 10310 24755 10362
rect 24755 10310 24767 10362
rect 24767 10310 24781 10362
rect 24805 10310 24819 10362
rect 24819 10310 24831 10362
rect 24831 10310 24861 10362
rect 24885 10310 24895 10362
rect 24895 10310 24941 10362
rect 24645 10308 24701 10310
rect 24725 10308 24781 10310
rect 24805 10308 24861 10310
rect 24885 10308 24941 10310
rect 24645 9274 24701 9276
rect 24725 9274 24781 9276
rect 24805 9274 24861 9276
rect 24885 9274 24941 9276
rect 24645 9222 24691 9274
rect 24691 9222 24701 9274
rect 24725 9222 24755 9274
rect 24755 9222 24767 9274
rect 24767 9222 24781 9274
rect 24805 9222 24819 9274
rect 24819 9222 24831 9274
rect 24831 9222 24861 9274
rect 24885 9222 24895 9274
rect 24895 9222 24941 9274
rect 24645 9220 24701 9222
rect 24725 9220 24781 9222
rect 24805 9220 24861 9222
rect 24885 9220 24941 9222
rect 24645 8186 24701 8188
rect 24725 8186 24781 8188
rect 24805 8186 24861 8188
rect 24885 8186 24941 8188
rect 24645 8134 24691 8186
rect 24691 8134 24701 8186
rect 24725 8134 24755 8186
rect 24755 8134 24767 8186
rect 24767 8134 24781 8186
rect 24805 8134 24819 8186
rect 24819 8134 24831 8186
rect 24831 8134 24861 8186
rect 24885 8134 24895 8186
rect 24895 8134 24941 8186
rect 24645 8132 24701 8134
rect 24725 8132 24781 8134
rect 24805 8132 24861 8134
rect 24885 8132 24941 8134
rect 24645 7098 24701 7100
rect 24725 7098 24781 7100
rect 24805 7098 24861 7100
rect 24885 7098 24941 7100
rect 24645 7046 24691 7098
rect 24691 7046 24701 7098
rect 24725 7046 24755 7098
rect 24755 7046 24767 7098
rect 24767 7046 24781 7098
rect 24805 7046 24819 7098
rect 24819 7046 24831 7098
rect 24831 7046 24861 7098
rect 24885 7046 24895 7098
rect 24895 7046 24941 7098
rect 24645 7044 24701 7046
rect 24725 7044 24781 7046
rect 24805 7044 24861 7046
rect 24885 7044 24941 7046
rect 26330 18672 26386 18728
rect 26330 17176 26386 17232
rect 28814 21684 28870 21720
rect 28814 21664 28816 21684
rect 28816 21664 28868 21684
rect 28868 21664 28870 21684
rect 24645 6010 24701 6012
rect 24725 6010 24781 6012
rect 24805 6010 24861 6012
rect 24885 6010 24941 6012
rect 24645 5958 24691 6010
rect 24691 5958 24701 6010
rect 24725 5958 24755 6010
rect 24755 5958 24767 6010
rect 24767 5958 24781 6010
rect 24805 5958 24819 6010
rect 24819 5958 24831 6010
rect 24831 5958 24861 6010
rect 24885 5958 24895 6010
rect 24895 5958 24941 6010
rect 24645 5956 24701 5958
rect 24725 5956 24781 5958
rect 24805 5956 24861 5958
rect 24885 5956 24941 5958
rect 24645 4922 24701 4924
rect 24725 4922 24781 4924
rect 24805 4922 24861 4924
rect 24885 4922 24941 4924
rect 24645 4870 24691 4922
rect 24691 4870 24701 4922
rect 24725 4870 24755 4922
rect 24755 4870 24767 4922
rect 24767 4870 24781 4922
rect 24805 4870 24819 4922
rect 24819 4870 24831 4922
rect 24831 4870 24861 4922
rect 24885 4870 24895 4922
rect 24895 4870 24941 4922
rect 24645 4868 24701 4870
rect 24725 4868 24781 4870
rect 24805 4868 24861 4870
rect 24885 4868 24941 4870
rect 24645 3834 24701 3836
rect 24725 3834 24781 3836
rect 24805 3834 24861 3836
rect 24885 3834 24941 3836
rect 24645 3782 24691 3834
rect 24691 3782 24701 3834
rect 24725 3782 24755 3834
rect 24755 3782 24767 3834
rect 24767 3782 24781 3834
rect 24805 3782 24819 3834
rect 24819 3782 24831 3834
rect 24831 3782 24861 3834
rect 24885 3782 24895 3834
rect 24895 3782 24941 3834
rect 24645 3780 24701 3782
rect 24725 3780 24781 3782
rect 24805 3780 24861 3782
rect 24885 3780 24941 3782
rect 26422 3440 26478 3496
rect 24645 2746 24701 2748
rect 24725 2746 24781 2748
rect 24805 2746 24861 2748
rect 24885 2746 24941 2748
rect 24645 2694 24691 2746
rect 24691 2694 24701 2746
rect 24725 2694 24755 2746
rect 24755 2694 24767 2746
rect 24767 2694 24781 2746
rect 24805 2694 24819 2746
rect 24819 2694 24831 2746
rect 24831 2694 24861 2746
rect 24885 2694 24895 2746
rect 24895 2694 24941 2746
rect 24645 2692 24701 2694
rect 24725 2692 24781 2694
rect 24805 2692 24861 2694
rect 24885 2692 24941 2694
rect 26606 5072 26662 5128
rect 27342 12688 27398 12744
rect 27526 11192 27582 11248
rect 27526 9696 27582 9752
rect 27434 6704 27490 6760
rect 29090 14184 29146 14240
rect 29090 8236 29092 8256
rect 29092 8236 29144 8256
rect 29144 8236 29146 8256
rect 29090 8200 29146 8236
rect 27526 5208 27582 5264
rect 27066 3712 27122 3768
rect 26514 2216 26570 2272
rect 27526 720 27582 776
<< metal3 >>
rect 0 32194 800 32224
rect 3877 32194 3943 32197
rect 29912 32194 30712 32224
rect 0 32192 3943 32194
rect 0 32136 3882 32192
rect 3938 32136 3943 32192
rect 0 32134 3943 32136
rect 0 32104 800 32134
rect 3877 32131 3943 32134
rect 27478 32134 30712 32194
rect 27337 32058 27403 32061
rect 27478 32058 27538 32134
rect 29912 32104 30712 32134
rect 27337 32056 27538 32058
rect 27337 32000 27342 32056
rect 27398 32000 27538 32056
rect 27337 31998 27538 32000
rect 27337 31995 27403 31998
rect 0 30834 800 30864
rect 4061 30834 4127 30837
rect 0 30832 4127 30834
rect 0 30776 4066 30832
rect 4122 30776 4127 30832
rect 0 30774 4127 30776
rect 0 30744 800 30774
rect 4061 30771 4127 30774
rect 26877 30698 26943 30701
rect 29912 30698 30712 30728
rect 26877 30696 30712 30698
rect 26877 30640 26882 30696
rect 26938 30640 30712 30696
rect 26877 30638 30712 30640
rect 26877 30635 26943 30638
rect 29912 30608 30712 30638
rect 10419 30496 10739 30497
rect 10419 30432 10427 30496
rect 10491 30432 10507 30496
rect 10571 30432 10587 30496
rect 10651 30432 10667 30496
rect 10731 30432 10739 30496
rect 10419 30431 10739 30432
rect 19895 30496 20215 30497
rect 19895 30432 19903 30496
rect 19967 30432 19983 30496
rect 20047 30432 20063 30496
rect 20127 30432 20143 30496
rect 20207 30432 20215 30496
rect 19895 30431 20215 30432
rect 5682 29952 6002 29953
rect 5682 29888 5690 29952
rect 5754 29888 5770 29952
rect 5834 29888 5850 29952
rect 5914 29888 5930 29952
rect 5994 29888 6002 29952
rect 5682 29887 6002 29888
rect 15157 29952 15477 29953
rect 15157 29888 15165 29952
rect 15229 29888 15245 29952
rect 15309 29888 15325 29952
rect 15389 29888 15405 29952
rect 15469 29888 15477 29952
rect 15157 29887 15477 29888
rect 24633 29952 24953 29953
rect 24633 29888 24641 29952
rect 24705 29888 24721 29952
rect 24785 29888 24801 29952
rect 24865 29888 24881 29952
rect 24945 29888 24953 29952
rect 24633 29887 24953 29888
rect 0 29474 800 29504
rect 4061 29474 4127 29477
rect 0 29472 4127 29474
rect 0 29416 4066 29472
rect 4122 29416 4127 29472
rect 0 29414 4127 29416
rect 0 29384 800 29414
rect 4061 29411 4127 29414
rect 14457 29474 14523 29477
rect 17585 29474 17651 29477
rect 14457 29472 17651 29474
rect 14457 29416 14462 29472
rect 14518 29416 17590 29472
rect 17646 29416 17651 29472
rect 14457 29414 17651 29416
rect 14457 29411 14523 29414
rect 17585 29411 17651 29414
rect 10419 29408 10739 29409
rect 10419 29344 10427 29408
rect 10491 29344 10507 29408
rect 10571 29344 10587 29408
rect 10651 29344 10667 29408
rect 10731 29344 10739 29408
rect 10419 29343 10739 29344
rect 19895 29408 20215 29409
rect 19895 29344 19903 29408
rect 19967 29344 19983 29408
rect 20047 29344 20063 29408
rect 20127 29344 20143 29408
rect 20207 29344 20215 29408
rect 19895 29343 20215 29344
rect 27429 29202 27495 29205
rect 29912 29202 30712 29232
rect 27429 29200 30712 29202
rect 27429 29144 27434 29200
rect 27490 29144 30712 29200
rect 27429 29142 30712 29144
rect 27429 29139 27495 29142
rect 29912 29112 30712 29142
rect 16573 29066 16639 29069
rect 17401 29066 17467 29069
rect 18781 29066 18847 29069
rect 16573 29064 18847 29066
rect 16573 29008 16578 29064
rect 16634 29008 17406 29064
rect 17462 29008 18786 29064
rect 18842 29008 18847 29064
rect 16573 29006 18847 29008
rect 16573 29003 16639 29006
rect 17401 29003 17467 29006
rect 18781 29003 18847 29006
rect 5682 28864 6002 28865
rect 5682 28800 5690 28864
rect 5754 28800 5770 28864
rect 5834 28800 5850 28864
rect 5914 28800 5930 28864
rect 5994 28800 6002 28864
rect 5682 28799 6002 28800
rect 15157 28864 15477 28865
rect 15157 28800 15165 28864
rect 15229 28800 15245 28864
rect 15309 28800 15325 28864
rect 15389 28800 15405 28864
rect 15469 28800 15477 28864
rect 15157 28799 15477 28800
rect 24633 28864 24953 28865
rect 24633 28800 24641 28864
rect 24705 28800 24721 28864
rect 24785 28800 24801 28864
rect 24865 28800 24881 28864
rect 24945 28800 24953 28864
rect 24633 28799 24953 28800
rect 9857 28522 9923 28525
rect 10593 28522 10659 28525
rect 9857 28520 10659 28522
rect 9857 28464 9862 28520
rect 9918 28464 10598 28520
rect 10654 28464 10659 28520
rect 9857 28462 10659 28464
rect 9857 28459 9923 28462
rect 10593 28459 10659 28462
rect 10777 28522 10843 28525
rect 12617 28522 12683 28525
rect 10777 28520 12683 28522
rect 10777 28464 10782 28520
rect 10838 28464 12622 28520
rect 12678 28464 12683 28520
rect 10777 28462 12683 28464
rect 10777 28459 10843 28462
rect 12617 28459 12683 28462
rect 10419 28320 10739 28321
rect 10419 28256 10427 28320
rect 10491 28256 10507 28320
rect 10571 28256 10587 28320
rect 10651 28256 10667 28320
rect 10731 28256 10739 28320
rect 10419 28255 10739 28256
rect 19895 28320 20215 28321
rect 19895 28256 19903 28320
rect 19967 28256 19983 28320
rect 20047 28256 20063 28320
rect 20127 28256 20143 28320
rect 20207 28256 20215 28320
rect 19895 28255 20215 28256
rect 0 28114 800 28144
rect 4061 28114 4127 28117
rect 0 28112 4127 28114
rect 0 28056 4066 28112
rect 4122 28056 4127 28112
rect 0 28054 4127 28056
rect 0 28024 800 28054
rect 4061 28051 4127 28054
rect 10317 27978 10383 27981
rect 16205 27978 16271 27981
rect 10317 27976 16271 27978
rect 10317 27920 10322 27976
rect 10378 27920 16210 27976
rect 16266 27920 16271 27976
rect 10317 27918 16271 27920
rect 10317 27915 10383 27918
rect 16205 27915 16271 27918
rect 5682 27776 6002 27777
rect 5682 27712 5690 27776
rect 5754 27712 5770 27776
rect 5834 27712 5850 27776
rect 5914 27712 5930 27776
rect 5994 27712 6002 27776
rect 5682 27711 6002 27712
rect 15157 27776 15477 27777
rect 15157 27712 15165 27776
rect 15229 27712 15245 27776
rect 15309 27712 15325 27776
rect 15389 27712 15405 27776
rect 15469 27712 15477 27776
rect 15157 27711 15477 27712
rect 24633 27776 24953 27777
rect 24633 27712 24641 27776
rect 24705 27712 24721 27776
rect 24785 27712 24801 27776
rect 24865 27712 24881 27776
rect 24945 27712 24953 27776
rect 24633 27711 24953 27712
rect 27521 27706 27587 27709
rect 29912 27706 30712 27736
rect 27521 27704 30712 27706
rect 27521 27648 27526 27704
rect 27582 27648 30712 27704
rect 27521 27646 30712 27648
rect 27521 27643 27587 27646
rect 29912 27616 30712 27646
rect 15377 27434 15443 27437
rect 16389 27434 16455 27437
rect 15377 27432 16455 27434
rect 15377 27376 15382 27432
rect 15438 27376 16394 27432
rect 16450 27376 16455 27432
rect 15377 27374 16455 27376
rect 15377 27371 15443 27374
rect 16389 27371 16455 27374
rect 13261 27300 13327 27301
rect 13261 27298 13308 27300
rect 13216 27296 13308 27298
rect 13216 27240 13266 27296
rect 13216 27238 13308 27240
rect 13261 27236 13308 27238
rect 13372 27236 13378 27300
rect 13261 27235 13327 27236
rect 10419 27232 10739 27233
rect 10419 27168 10427 27232
rect 10491 27168 10507 27232
rect 10571 27168 10587 27232
rect 10651 27168 10667 27232
rect 10731 27168 10739 27232
rect 10419 27167 10739 27168
rect 19895 27232 20215 27233
rect 19895 27168 19903 27232
rect 19967 27168 19983 27232
rect 20047 27168 20063 27232
rect 20127 27168 20143 27232
rect 20207 27168 20215 27232
rect 19895 27167 20215 27168
rect 11973 26890 12039 26893
rect 13353 26890 13419 26893
rect 11973 26888 13419 26890
rect 11973 26832 11978 26888
rect 12034 26832 13358 26888
rect 13414 26832 13419 26888
rect 11973 26830 13419 26832
rect 11973 26827 12039 26830
rect 13353 26827 13419 26830
rect 0 26754 800 26784
rect 4061 26754 4127 26757
rect 0 26752 4127 26754
rect 0 26696 4066 26752
rect 4122 26696 4127 26752
rect 0 26694 4127 26696
rect 0 26664 800 26694
rect 4061 26691 4127 26694
rect 5682 26688 6002 26689
rect 5682 26624 5690 26688
rect 5754 26624 5770 26688
rect 5834 26624 5850 26688
rect 5914 26624 5930 26688
rect 5994 26624 6002 26688
rect 5682 26623 6002 26624
rect 15157 26688 15477 26689
rect 15157 26624 15165 26688
rect 15229 26624 15245 26688
rect 15309 26624 15325 26688
rect 15389 26624 15405 26688
rect 15469 26624 15477 26688
rect 15157 26623 15477 26624
rect 24633 26688 24953 26689
rect 24633 26624 24641 26688
rect 24705 26624 24721 26688
rect 24785 26624 24801 26688
rect 24865 26624 24881 26688
rect 24945 26624 24953 26688
rect 24633 26623 24953 26624
rect 27521 26210 27587 26213
rect 29912 26210 30712 26240
rect 27521 26208 30712 26210
rect 27521 26152 27526 26208
rect 27582 26152 30712 26208
rect 27521 26150 30712 26152
rect 27521 26147 27587 26150
rect 10419 26144 10739 26145
rect 10419 26080 10427 26144
rect 10491 26080 10507 26144
rect 10571 26080 10587 26144
rect 10651 26080 10667 26144
rect 10731 26080 10739 26144
rect 10419 26079 10739 26080
rect 19895 26144 20215 26145
rect 19895 26080 19903 26144
rect 19967 26080 19983 26144
rect 20047 26080 20063 26144
rect 20127 26080 20143 26144
rect 20207 26080 20215 26144
rect 29912 26120 30712 26150
rect 19895 26079 20215 26080
rect 5682 25600 6002 25601
rect 5682 25536 5690 25600
rect 5754 25536 5770 25600
rect 5834 25536 5850 25600
rect 5914 25536 5930 25600
rect 5994 25536 6002 25600
rect 5682 25535 6002 25536
rect 15157 25600 15477 25601
rect 15157 25536 15165 25600
rect 15229 25536 15245 25600
rect 15309 25536 15325 25600
rect 15389 25536 15405 25600
rect 15469 25536 15477 25600
rect 15157 25535 15477 25536
rect 24633 25600 24953 25601
rect 24633 25536 24641 25600
rect 24705 25536 24721 25600
rect 24785 25536 24801 25600
rect 24865 25536 24881 25600
rect 24945 25536 24953 25600
rect 24633 25535 24953 25536
rect 0 25394 800 25424
rect 4061 25394 4127 25397
rect 0 25392 4127 25394
rect 0 25336 4066 25392
rect 4122 25336 4127 25392
rect 0 25334 4127 25336
rect 0 25304 800 25334
rect 4061 25331 4127 25334
rect 19609 25258 19675 25261
rect 20478 25258 20484 25260
rect 19609 25256 20484 25258
rect 19609 25200 19614 25256
rect 19670 25200 20484 25256
rect 19609 25198 20484 25200
rect 19609 25195 19675 25198
rect 20478 25196 20484 25198
rect 20548 25196 20554 25260
rect 10419 25056 10739 25057
rect 10419 24992 10427 25056
rect 10491 24992 10507 25056
rect 10571 24992 10587 25056
rect 10651 24992 10667 25056
rect 10731 24992 10739 25056
rect 10419 24991 10739 24992
rect 19895 25056 20215 25057
rect 19895 24992 19903 25056
rect 19967 24992 19983 25056
rect 20047 24992 20063 25056
rect 20127 24992 20143 25056
rect 20207 24992 20215 25056
rect 19895 24991 20215 24992
rect 26693 24714 26759 24717
rect 29912 24714 30712 24744
rect 26693 24712 30712 24714
rect 26693 24656 26698 24712
rect 26754 24656 30712 24712
rect 26693 24654 30712 24656
rect 26693 24651 26759 24654
rect 29912 24624 30712 24654
rect 5682 24512 6002 24513
rect 5682 24448 5690 24512
rect 5754 24448 5770 24512
rect 5834 24448 5850 24512
rect 5914 24448 5930 24512
rect 5994 24448 6002 24512
rect 5682 24447 6002 24448
rect 15157 24512 15477 24513
rect 15157 24448 15165 24512
rect 15229 24448 15245 24512
rect 15309 24448 15325 24512
rect 15389 24448 15405 24512
rect 15469 24448 15477 24512
rect 15157 24447 15477 24448
rect 24633 24512 24953 24513
rect 24633 24448 24641 24512
rect 24705 24448 24721 24512
rect 24785 24448 24801 24512
rect 24865 24448 24881 24512
rect 24945 24448 24953 24512
rect 24633 24447 24953 24448
rect 0 24034 800 24064
rect 4061 24034 4127 24037
rect 0 24032 4127 24034
rect 0 23976 4066 24032
rect 4122 23976 4127 24032
rect 0 23974 4127 23976
rect 0 23944 800 23974
rect 4061 23971 4127 23974
rect 10419 23968 10739 23969
rect 10419 23904 10427 23968
rect 10491 23904 10507 23968
rect 10571 23904 10587 23968
rect 10651 23904 10667 23968
rect 10731 23904 10739 23968
rect 10419 23903 10739 23904
rect 19895 23968 20215 23969
rect 19895 23904 19903 23968
rect 19967 23904 19983 23968
rect 20047 23904 20063 23968
rect 20127 23904 20143 23968
rect 20207 23904 20215 23968
rect 19895 23903 20215 23904
rect 18229 23762 18295 23765
rect 19333 23762 19399 23765
rect 18229 23760 19399 23762
rect 18229 23704 18234 23760
rect 18290 23704 19338 23760
rect 19394 23704 19399 23760
rect 18229 23702 19399 23704
rect 18229 23699 18295 23702
rect 19333 23699 19399 23702
rect 19742 23564 19748 23628
rect 19812 23626 19818 23628
rect 20161 23626 20227 23629
rect 19812 23624 20227 23626
rect 19812 23568 20166 23624
rect 20222 23568 20227 23624
rect 19812 23566 20227 23568
rect 19812 23564 19818 23566
rect 20161 23563 20227 23566
rect 12433 23490 12499 23493
rect 13670 23490 13676 23492
rect 12433 23488 13676 23490
rect 12433 23432 12438 23488
rect 12494 23432 13676 23488
rect 12433 23430 13676 23432
rect 12433 23427 12499 23430
rect 13670 23428 13676 23430
rect 13740 23428 13746 23492
rect 18689 23490 18755 23493
rect 19977 23490 20043 23493
rect 18689 23488 20043 23490
rect 18689 23432 18694 23488
rect 18750 23432 19982 23488
rect 20038 23432 20043 23488
rect 18689 23430 20043 23432
rect 18689 23427 18755 23430
rect 19977 23427 20043 23430
rect 5682 23424 6002 23425
rect 5682 23360 5690 23424
rect 5754 23360 5770 23424
rect 5834 23360 5850 23424
rect 5914 23360 5930 23424
rect 5994 23360 6002 23424
rect 5682 23359 6002 23360
rect 15157 23424 15477 23425
rect 15157 23360 15165 23424
rect 15229 23360 15245 23424
rect 15309 23360 15325 23424
rect 15389 23360 15405 23424
rect 15469 23360 15477 23424
rect 15157 23359 15477 23360
rect 24633 23424 24953 23425
rect 24633 23360 24641 23424
rect 24705 23360 24721 23424
rect 24785 23360 24801 23424
rect 24865 23360 24881 23424
rect 24945 23360 24953 23424
rect 24633 23359 24953 23360
rect 27429 23218 27495 23221
rect 29912 23218 30712 23248
rect 27429 23216 30712 23218
rect 27429 23160 27434 23216
rect 27490 23160 30712 23216
rect 27429 23158 30712 23160
rect 27429 23155 27495 23158
rect 29912 23128 30712 23158
rect 10419 22880 10739 22881
rect 10419 22816 10427 22880
rect 10491 22816 10507 22880
rect 10571 22816 10587 22880
rect 10651 22816 10667 22880
rect 10731 22816 10739 22880
rect 10419 22815 10739 22816
rect 19895 22880 20215 22881
rect 19895 22816 19903 22880
rect 19967 22816 19983 22880
rect 20047 22816 20063 22880
rect 20127 22816 20143 22880
rect 20207 22816 20215 22880
rect 19895 22815 20215 22816
rect 0 22674 800 22704
rect 3969 22674 4035 22677
rect 0 22672 4035 22674
rect 0 22616 3974 22672
rect 4030 22616 4035 22672
rect 0 22614 4035 22616
rect 0 22584 800 22614
rect 3969 22611 4035 22614
rect 5682 22336 6002 22337
rect 5682 22272 5690 22336
rect 5754 22272 5770 22336
rect 5834 22272 5850 22336
rect 5914 22272 5930 22336
rect 5994 22272 6002 22336
rect 5682 22271 6002 22272
rect 15157 22336 15477 22337
rect 15157 22272 15165 22336
rect 15229 22272 15245 22336
rect 15309 22272 15325 22336
rect 15389 22272 15405 22336
rect 15469 22272 15477 22336
rect 15157 22271 15477 22272
rect 24633 22336 24953 22337
rect 24633 22272 24641 22336
rect 24705 22272 24721 22336
rect 24785 22272 24801 22336
rect 24865 22272 24881 22336
rect 24945 22272 24953 22336
rect 24633 22271 24953 22272
rect 9765 21994 9831 21997
rect 10041 21994 10107 21997
rect 9765 21992 10107 21994
rect 9765 21936 9770 21992
rect 9826 21936 10046 21992
rect 10102 21936 10107 21992
rect 9765 21934 10107 21936
rect 9765 21931 9831 21934
rect 10041 21931 10107 21934
rect 10419 21792 10739 21793
rect 10419 21728 10427 21792
rect 10491 21728 10507 21792
rect 10571 21728 10587 21792
rect 10651 21728 10667 21792
rect 10731 21728 10739 21792
rect 10419 21727 10739 21728
rect 19895 21792 20215 21793
rect 19895 21728 19903 21792
rect 19967 21728 19983 21792
rect 20047 21728 20063 21792
rect 20127 21728 20143 21792
rect 20207 21728 20215 21792
rect 19895 21727 20215 21728
rect 15377 21722 15443 21725
rect 16297 21722 16363 21725
rect 15377 21720 16363 21722
rect 15377 21664 15382 21720
rect 15438 21664 16302 21720
rect 16358 21664 16363 21720
rect 15377 21662 16363 21664
rect 15377 21659 15443 21662
rect 16297 21659 16363 21662
rect 28809 21722 28875 21725
rect 29912 21722 30712 21752
rect 28809 21720 30712 21722
rect 28809 21664 28814 21720
rect 28870 21664 30712 21720
rect 28809 21662 30712 21664
rect 28809 21659 28875 21662
rect 29912 21632 30712 21662
rect 0 21314 800 21344
rect 4061 21314 4127 21317
rect 0 21312 4127 21314
rect 0 21256 4066 21312
rect 4122 21256 4127 21312
rect 0 21254 4127 21256
rect 0 21224 800 21254
rect 4061 21251 4127 21254
rect 5682 21248 6002 21249
rect 5682 21184 5690 21248
rect 5754 21184 5770 21248
rect 5834 21184 5850 21248
rect 5914 21184 5930 21248
rect 5994 21184 6002 21248
rect 5682 21183 6002 21184
rect 15157 21248 15477 21249
rect 15157 21184 15165 21248
rect 15229 21184 15245 21248
rect 15309 21184 15325 21248
rect 15389 21184 15405 21248
rect 15469 21184 15477 21248
rect 15157 21183 15477 21184
rect 24633 21248 24953 21249
rect 24633 21184 24641 21248
rect 24705 21184 24721 21248
rect 24785 21184 24801 21248
rect 24865 21184 24881 21248
rect 24945 21184 24953 21248
rect 24633 21183 24953 21184
rect 20161 20906 20227 20909
rect 21541 20906 21607 20909
rect 23749 20906 23815 20909
rect 20161 20904 23815 20906
rect 20161 20848 20166 20904
rect 20222 20848 21546 20904
rect 21602 20848 23754 20904
rect 23810 20848 23815 20904
rect 20161 20846 23815 20848
rect 20161 20843 20227 20846
rect 21541 20843 21607 20846
rect 23749 20843 23815 20846
rect 10419 20704 10739 20705
rect 10419 20640 10427 20704
rect 10491 20640 10507 20704
rect 10571 20640 10587 20704
rect 10651 20640 10667 20704
rect 10731 20640 10739 20704
rect 10419 20639 10739 20640
rect 19895 20704 20215 20705
rect 19895 20640 19903 20704
rect 19967 20640 19983 20704
rect 20047 20640 20063 20704
rect 20127 20640 20143 20704
rect 20207 20640 20215 20704
rect 19895 20639 20215 20640
rect 15009 20362 15075 20365
rect 23657 20362 23723 20365
rect 15009 20360 23723 20362
rect 15009 20304 15014 20360
rect 15070 20304 23662 20360
rect 23718 20304 23723 20360
rect 15009 20302 23723 20304
rect 15009 20299 15075 20302
rect 23657 20299 23723 20302
rect 26417 20226 26483 20229
rect 29912 20226 30712 20256
rect 26417 20224 30712 20226
rect 26417 20168 26422 20224
rect 26478 20168 30712 20224
rect 26417 20166 30712 20168
rect 26417 20163 26483 20166
rect 5682 20160 6002 20161
rect 5682 20096 5690 20160
rect 5754 20096 5770 20160
rect 5834 20096 5850 20160
rect 5914 20096 5930 20160
rect 5994 20096 6002 20160
rect 5682 20095 6002 20096
rect 15157 20160 15477 20161
rect 15157 20096 15165 20160
rect 15229 20096 15245 20160
rect 15309 20096 15325 20160
rect 15389 20096 15405 20160
rect 15469 20096 15477 20160
rect 15157 20095 15477 20096
rect 24633 20160 24953 20161
rect 24633 20096 24641 20160
rect 24705 20096 24721 20160
rect 24785 20096 24801 20160
rect 24865 20096 24881 20160
rect 24945 20096 24953 20160
rect 29912 20136 30712 20166
rect 24633 20095 24953 20096
rect 0 19954 800 19984
rect 9305 19954 9371 19957
rect 0 19952 9371 19954
rect 0 19896 9310 19952
rect 9366 19896 9371 19952
rect 0 19894 9371 19896
rect 0 19864 800 19894
rect 9305 19891 9371 19894
rect 14825 19954 14891 19957
rect 15469 19954 15535 19957
rect 14825 19952 15535 19954
rect 14825 19896 14830 19952
rect 14886 19896 15474 19952
rect 15530 19896 15535 19952
rect 14825 19894 15535 19896
rect 14825 19891 14891 19894
rect 15469 19891 15535 19894
rect 10225 19818 10291 19821
rect 18229 19818 18295 19821
rect 10225 19816 18295 19818
rect 10225 19760 10230 19816
rect 10286 19760 18234 19816
rect 18290 19760 18295 19816
rect 10225 19758 18295 19760
rect 10225 19755 10291 19758
rect 18229 19755 18295 19758
rect 23289 19818 23355 19821
rect 25037 19818 25103 19821
rect 23289 19816 25103 19818
rect 23289 19760 23294 19816
rect 23350 19760 25042 19816
rect 25098 19760 25103 19816
rect 23289 19758 25103 19760
rect 23289 19755 23355 19758
rect 25037 19755 25103 19758
rect 14549 19682 14615 19685
rect 19241 19682 19307 19685
rect 14549 19680 19307 19682
rect 14549 19624 14554 19680
rect 14610 19624 19246 19680
rect 19302 19624 19307 19680
rect 14549 19622 19307 19624
rect 14549 19619 14615 19622
rect 19241 19619 19307 19622
rect 10419 19616 10739 19617
rect 10419 19552 10427 19616
rect 10491 19552 10507 19616
rect 10571 19552 10587 19616
rect 10651 19552 10667 19616
rect 10731 19552 10739 19616
rect 10419 19551 10739 19552
rect 19895 19616 20215 19617
rect 19895 19552 19903 19616
rect 19967 19552 19983 19616
rect 20047 19552 20063 19616
rect 20127 19552 20143 19616
rect 20207 19552 20215 19616
rect 19895 19551 20215 19552
rect 16849 19546 16915 19549
rect 18689 19546 18755 19549
rect 16849 19544 18755 19546
rect 16849 19488 16854 19544
rect 16910 19488 18694 19544
rect 18750 19488 18755 19544
rect 16849 19486 18755 19488
rect 16849 19483 16915 19486
rect 18689 19483 18755 19486
rect 7925 19410 7991 19413
rect 19517 19410 19583 19413
rect 7925 19408 19583 19410
rect 7925 19352 7930 19408
rect 7986 19352 19522 19408
rect 19578 19352 19583 19408
rect 7925 19350 19583 19352
rect 7925 19347 7991 19350
rect 19517 19347 19583 19350
rect 5682 19072 6002 19073
rect 5682 19008 5690 19072
rect 5754 19008 5770 19072
rect 5834 19008 5850 19072
rect 5914 19008 5930 19072
rect 5994 19008 6002 19072
rect 5682 19007 6002 19008
rect 15157 19072 15477 19073
rect 15157 19008 15165 19072
rect 15229 19008 15245 19072
rect 15309 19008 15325 19072
rect 15389 19008 15405 19072
rect 15469 19008 15477 19072
rect 15157 19007 15477 19008
rect 24633 19072 24953 19073
rect 24633 19008 24641 19072
rect 24705 19008 24721 19072
rect 24785 19008 24801 19072
rect 24865 19008 24881 19072
rect 24945 19008 24953 19072
rect 24633 19007 24953 19008
rect 26325 18730 26391 18733
rect 29912 18730 30712 18760
rect 26325 18728 30712 18730
rect 26325 18672 26330 18728
rect 26386 18672 30712 18728
rect 26325 18670 30712 18672
rect 26325 18667 26391 18670
rect 29912 18640 30712 18670
rect 0 18594 800 18624
rect 3785 18594 3851 18597
rect 0 18592 3851 18594
rect 0 18536 3790 18592
rect 3846 18536 3851 18592
rect 0 18534 3851 18536
rect 0 18504 800 18534
rect 3785 18531 3851 18534
rect 10419 18528 10739 18529
rect 10419 18464 10427 18528
rect 10491 18464 10507 18528
rect 10571 18464 10587 18528
rect 10651 18464 10667 18528
rect 10731 18464 10739 18528
rect 10419 18463 10739 18464
rect 19895 18528 20215 18529
rect 19895 18464 19903 18528
rect 19967 18464 19983 18528
rect 20047 18464 20063 18528
rect 20127 18464 20143 18528
rect 20207 18464 20215 18528
rect 19895 18463 20215 18464
rect 5682 17984 6002 17985
rect 5682 17920 5690 17984
rect 5754 17920 5770 17984
rect 5834 17920 5850 17984
rect 5914 17920 5930 17984
rect 5994 17920 6002 17984
rect 5682 17919 6002 17920
rect 15157 17984 15477 17985
rect 15157 17920 15165 17984
rect 15229 17920 15245 17984
rect 15309 17920 15325 17984
rect 15389 17920 15405 17984
rect 15469 17920 15477 17984
rect 15157 17919 15477 17920
rect 24633 17984 24953 17985
rect 24633 17920 24641 17984
rect 24705 17920 24721 17984
rect 24785 17920 24801 17984
rect 24865 17920 24881 17984
rect 24945 17920 24953 17984
rect 24633 17919 24953 17920
rect 20478 17852 20484 17916
rect 20548 17914 20554 17916
rect 20621 17914 20687 17917
rect 20548 17912 20687 17914
rect 20548 17856 20626 17912
rect 20682 17856 20687 17912
rect 20548 17854 20687 17856
rect 20548 17852 20554 17854
rect 20621 17851 20687 17854
rect 12525 17506 12591 17509
rect 13721 17506 13787 17509
rect 12525 17504 13787 17506
rect 12525 17448 12530 17504
rect 12586 17448 13726 17504
rect 13782 17448 13787 17504
rect 12525 17446 13787 17448
rect 12525 17443 12591 17446
rect 13721 17443 13787 17446
rect 10419 17440 10739 17441
rect 10419 17376 10427 17440
rect 10491 17376 10507 17440
rect 10571 17376 10587 17440
rect 10651 17376 10667 17440
rect 10731 17376 10739 17440
rect 10419 17375 10739 17376
rect 19895 17440 20215 17441
rect 19895 17376 19903 17440
rect 19967 17376 19983 17440
rect 20047 17376 20063 17440
rect 20127 17376 20143 17440
rect 20207 17376 20215 17440
rect 19895 17375 20215 17376
rect 0 17234 800 17264
rect 4061 17234 4127 17237
rect 0 17232 4127 17234
rect 0 17176 4066 17232
rect 4122 17176 4127 17232
rect 0 17174 4127 17176
rect 0 17144 800 17174
rect 4061 17171 4127 17174
rect 26325 17234 26391 17237
rect 29912 17234 30712 17264
rect 26325 17232 30712 17234
rect 26325 17176 26330 17232
rect 26386 17176 30712 17232
rect 26325 17174 30712 17176
rect 26325 17171 26391 17174
rect 29912 17144 30712 17174
rect 19333 16962 19399 16965
rect 19742 16962 19748 16964
rect 19333 16960 19748 16962
rect 19333 16904 19338 16960
rect 19394 16904 19748 16960
rect 19333 16902 19748 16904
rect 19333 16899 19399 16902
rect 19742 16900 19748 16902
rect 19812 16900 19818 16964
rect 5682 16896 6002 16897
rect 5682 16832 5690 16896
rect 5754 16832 5770 16896
rect 5834 16832 5850 16896
rect 5914 16832 5930 16896
rect 5994 16832 6002 16896
rect 5682 16831 6002 16832
rect 15157 16896 15477 16897
rect 15157 16832 15165 16896
rect 15229 16832 15245 16896
rect 15309 16832 15325 16896
rect 15389 16832 15405 16896
rect 15469 16832 15477 16896
rect 15157 16831 15477 16832
rect 24633 16896 24953 16897
rect 24633 16832 24641 16896
rect 24705 16832 24721 16896
rect 24785 16832 24801 16896
rect 24865 16832 24881 16896
rect 24945 16832 24953 16896
rect 24633 16831 24953 16832
rect 10419 16352 10739 16353
rect 10419 16288 10427 16352
rect 10491 16288 10507 16352
rect 10571 16288 10587 16352
rect 10651 16288 10667 16352
rect 10731 16288 10739 16352
rect 10419 16287 10739 16288
rect 19895 16352 20215 16353
rect 19895 16288 19903 16352
rect 19967 16288 19983 16352
rect 20047 16288 20063 16352
rect 20127 16288 20143 16352
rect 20207 16288 20215 16352
rect 19895 16287 20215 16288
rect 3785 16146 3851 16149
rect 19517 16146 19583 16149
rect 3785 16144 19583 16146
rect 3785 16088 3790 16144
rect 3846 16088 19522 16144
rect 19578 16088 19583 16144
rect 3785 16086 19583 16088
rect 3785 16083 3851 16086
rect 19517 16083 19583 16086
rect 1301 16010 1367 16013
rect 15929 16010 15995 16013
rect 1301 16008 15995 16010
rect 1301 15952 1306 16008
rect 1362 15952 15934 16008
rect 15990 15952 15995 16008
rect 1301 15950 15995 15952
rect 1301 15947 1367 15950
rect 15929 15947 15995 15950
rect 5682 15808 6002 15809
rect 0 15738 800 15768
rect 5682 15744 5690 15808
rect 5754 15744 5770 15808
rect 5834 15744 5850 15808
rect 5914 15744 5930 15808
rect 5994 15744 6002 15808
rect 5682 15743 6002 15744
rect 15157 15808 15477 15809
rect 15157 15744 15165 15808
rect 15229 15744 15245 15808
rect 15309 15744 15325 15808
rect 15389 15744 15405 15808
rect 15469 15744 15477 15808
rect 15157 15743 15477 15744
rect 24633 15808 24953 15809
rect 24633 15744 24641 15808
rect 24705 15744 24721 15808
rect 24785 15744 24801 15808
rect 24865 15744 24881 15808
rect 24945 15744 24953 15808
rect 24633 15743 24953 15744
rect 4061 15738 4127 15741
rect 29912 15738 30712 15768
rect 0 15736 4127 15738
rect 0 15680 4066 15736
rect 4122 15680 4127 15736
rect 0 15678 4127 15680
rect 0 15648 800 15678
rect 4061 15675 4127 15678
rect 26006 15678 30712 15738
rect 9765 15602 9831 15605
rect 18505 15602 18571 15605
rect 18965 15602 19031 15605
rect 9765 15600 19031 15602
rect 9765 15544 9770 15600
rect 9826 15544 18510 15600
rect 18566 15544 18970 15600
rect 19026 15544 19031 15600
rect 9765 15542 19031 15544
rect 9765 15539 9831 15542
rect 18505 15539 18571 15542
rect 18965 15539 19031 15542
rect 13670 15404 13676 15468
rect 13740 15466 13746 15468
rect 26006 15466 26066 15678
rect 29912 15648 30712 15678
rect 13740 15406 26066 15466
rect 13740 15404 13746 15406
rect 10419 15264 10739 15265
rect 10419 15200 10427 15264
rect 10491 15200 10507 15264
rect 10571 15200 10587 15264
rect 10651 15200 10667 15264
rect 10731 15200 10739 15264
rect 10419 15199 10739 15200
rect 19895 15264 20215 15265
rect 19895 15200 19903 15264
rect 19967 15200 19983 15264
rect 20047 15200 20063 15264
rect 20127 15200 20143 15264
rect 20207 15200 20215 15264
rect 19895 15199 20215 15200
rect 4061 15058 4127 15061
rect 22093 15058 22159 15061
rect 4061 15056 22159 15058
rect 4061 15000 4066 15056
rect 4122 15000 22098 15056
rect 22154 15000 22159 15056
rect 4061 14998 22159 15000
rect 4061 14995 4127 14998
rect 22093 14995 22159 14998
rect 21081 14922 21147 14925
rect 22553 14922 22619 14925
rect 21081 14920 22619 14922
rect 21081 14864 21086 14920
rect 21142 14864 22558 14920
rect 22614 14864 22619 14920
rect 21081 14862 22619 14864
rect 21081 14859 21147 14862
rect 22553 14859 22619 14862
rect 5682 14720 6002 14721
rect 5682 14656 5690 14720
rect 5754 14656 5770 14720
rect 5834 14656 5850 14720
rect 5914 14656 5930 14720
rect 5994 14656 6002 14720
rect 5682 14655 6002 14656
rect 15157 14720 15477 14721
rect 15157 14656 15165 14720
rect 15229 14656 15245 14720
rect 15309 14656 15325 14720
rect 15389 14656 15405 14720
rect 15469 14656 15477 14720
rect 15157 14655 15477 14656
rect 24633 14720 24953 14721
rect 24633 14656 24641 14720
rect 24705 14656 24721 14720
rect 24785 14656 24801 14720
rect 24865 14656 24881 14720
rect 24945 14656 24953 14720
rect 24633 14655 24953 14656
rect 0 14378 800 14408
rect 4061 14378 4127 14381
rect 0 14376 4127 14378
rect 0 14320 4066 14376
rect 4122 14320 4127 14376
rect 0 14318 4127 14320
rect 0 14288 800 14318
rect 4061 14315 4127 14318
rect 29085 14242 29151 14245
rect 29912 14242 30712 14272
rect 29085 14240 30712 14242
rect 29085 14184 29090 14240
rect 29146 14184 30712 14240
rect 29085 14182 30712 14184
rect 29085 14179 29151 14182
rect 10419 14176 10739 14177
rect 10419 14112 10427 14176
rect 10491 14112 10507 14176
rect 10571 14112 10587 14176
rect 10651 14112 10667 14176
rect 10731 14112 10739 14176
rect 10419 14111 10739 14112
rect 19895 14176 20215 14177
rect 19895 14112 19903 14176
rect 19967 14112 19983 14176
rect 20047 14112 20063 14176
rect 20127 14112 20143 14176
rect 20207 14112 20215 14176
rect 29912 14152 30712 14182
rect 19895 14111 20215 14112
rect 12893 13970 12959 13973
rect 15653 13970 15719 13973
rect 12893 13968 15719 13970
rect 12893 13912 12898 13968
rect 12954 13912 15658 13968
rect 15714 13912 15719 13968
rect 12893 13910 15719 13912
rect 12893 13907 12959 13910
rect 15653 13907 15719 13910
rect 5682 13632 6002 13633
rect 5682 13568 5690 13632
rect 5754 13568 5770 13632
rect 5834 13568 5850 13632
rect 5914 13568 5930 13632
rect 5994 13568 6002 13632
rect 5682 13567 6002 13568
rect 15157 13632 15477 13633
rect 15157 13568 15165 13632
rect 15229 13568 15245 13632
rect 15309 13568 15325 13632
rect 15389 13568 15405 13632
rect 15469 13568 15477 13632
rect 15157 13567 15477 13568
rect 24633 13632 24953 13633
rect 24633 13568 24641 13632
rect 24705 13568 24721 13632
rect 24785 13568 24801 13632
rect 24865 13568 24881 13632
rect 24945 13568 24953 13632
rect 24633 13567 24953 13568
rect 21909 13426 21975 13429
rect 24945 13426 25011 13429
rect 21909 13424 25011 13426
rect 21909 13368 21914 13424
rect 21970 13368 24950 13424
rect 25006 13368 25011 13424
rect 21909 13366 25011 13368
rect 21909 13363 21975 13366
rect 24945 13363 25011 13366
rect 10419 13088 10739 13089
rect 0 13018 800 13048
rect 10419 13024 10427 13088
rect 10491 13024 10507 13088
rect 10571 13024 10587 13088
rect 10651 13024 10667 13088
rect 10731 13024 10739 13088
rect 10419 13023 10739 13024
rect 19895 13088 20215 13089
rect 19895 13024 19903 13088
rect 19967 13024 19983 13088
rect 20047 13024 20063 13088
rect 20127 13024 20143 13088
rect 20207 13024 20215 13088
rect 19895 13023 20215 13024
rect 3877 13018 3943 13021
rect 0 13016 3943 13018
rect 0 12960 3882 13016
rect 3938 12960 3943 13016
rect 0 12958 3943 12960
rect 0 12928 800 12958
rect 3877 12955 3943 12958
rect 4797 12882 4863 12885
rect 5441 12882 5507 12885
rect 4797 12880 5507 12882
rect 4797 12824 4802 12880
rect 4858 12824 5446 12880
rect 5502 12824 5507 12880
rect 4797 12822 5507 12824
rect 4797 12819 4863 12822
rect 5441 12819 5507 12822
rect 27337 12746 27403 12749
rect 29912 12746 30712 12776
rect 27337 12744 30712 12746
rect 27337 12688 27342 12744
rect 27398 12688 30712 12744
rect 27337 12686 30712 12688
rect 27337 12683 27403 12686
rect 29912 12656 30712 12686
rect 5257 12610 5323 12613
rect 5257 12608 5458 12610
rect 5257 12552 5262 12608
rect 5318 12552 5458 12608
rect 5257 12550 5458 12552
rect 5257 12547 5323 12550
rect 5398 12338 5458 12550
rect 5682 12544 6002 12545
rect 5682 12480 5690 12544
rect 5754 12480 5770 12544
rect 5834 12480 5850 12544
rect 5914 12480 5930 12544
rect 5994 12480 6002 12544
rect 5682 12479 6002 12480
rect 15157 12544 15477 12545
rect 15157 12480 15165 12544
rect 15229 12480 15245 12544
rect 15309 12480 15325 12544
rect 15389 12480 15405 12544
rect 15469 12480 15477 12544
rect 15157 12479 15477 12480
rect 24633 12544 24953 12545
rect 24633 12480 24641 12544
rect 24705 12480 24721 12544
rect 24785 12480 24801 12544
rect 24865 12480 24881 12544
rect 24945 12480 24953 12544
rect 24633 12479 24953 12480
rect 5901 12338 5967 12341
rect 5398 12336 5967 12338
rect 5398 12280 5906 12336
rect 5962 12280 5967 12336
rect 5398 12278 5967 12280
rect 5901 12275 5967 12278
rect 10419 12000 10739 12001
rect 10419 11936 10427 12000
rect 10491 11936 10507 12000
rect 10571 11936 10587 12000
rect 10651 11936 10667 12000
rect 10731 11936 10739 12000
rect 10419 11935 10739 11936
rect 19895 12000 20215 12001
rect 19895 11936 19903 12000
rect 19967 11936 19983 12000
rect 20047 11936 20063 12000
rect 20127 11936 20143 12000
rect 20207 11936 20215 12000
rect 19895 11935 20215 11936
rect 0 11658 800 11688
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11568 800 11598
rect 4061 11595 4127 11598
rect 5682 11456 6002 11457
rect 5682 11392 5690 11456
rect 5754 11392 5770 11456
rect 5834 11392 5850 11456
rect 5914 11392 5930 11456
rect 5994 11392 6002 11456
rect 5682 11391 6002 11392
rect 15157 11456 15477 11457
rect 15157 11392 15165 11456
rect 15229 11392 15245 11456
rect 15309 11392 15325 11456
rect 15389 11392 15405 11456
rect 15469 11392 15477 11456
rect 15157 11391 15477 11392
rect 24633 11456 24953 11457
rect 24633 11392 24641 11456
rect 24705 11392 24721 11456
rect 24785 11392 24801 11456
rect 24865 11392 24881 11456
rect 24945 11392 24953 11456
rect 24633 11391 24953 11392
rect 27521 11250 27587 11253
rect 29912 11250 30712 11280
rect 27521 11248 30712 11250
rect 27521 11192 27526 11248
rect 27582 11192 30712 11248
rect 27521 11190 30712 11192
rect 27521 11187 27587 11190
rect 29912 11160 30712 11190
rect 10685 11114 10751 11117
rect 10910 11114 10916 11116
rect 10685 11112 10916 11114
rect 10685 11056 10690 11112
rect 10746 11056 10916 11112
rect 10685 11054 10916 11056
rect 10685 11051 10751 11054
rect 10910 11052 10916 11054
rect 10980 11052 10986 11116
rect 10419 10912 10739 10913
rect 10419 10848 10427 10912
rect 10491 10848 10507 10912
rect 10571 10848 10587 10912
rect 10651 10848 10667 10912
rect 10731 10848 10739 10912
rect 10419 10847 10739 10848
rect 19895 10912 20215 10913
rect 19895 10848 19903 10912
rect 19967 10848 19983 10912
rect 20047 10848 20063 10912
rect 20127 10848 20143 10912
rect 20207 10848 20215 10912
rect 19895 10847 20215 10848
rect 10501 10706 10567 10709
rect 11145 10706 11211 10709
rect 10501 10704 11211 10706
rect 10501 10648 10506 10704
rect 10562 10648 11150 10704
rect 11206 10648 11211 10704
rect 10501 10646 11211 10648
rect 10501 10643 10567 10646
rect 11145 10643 11211 10646
rect 10685 10570 10751 10573
rect 10869 10572 10935 10573
rect 10869 10570 10916 10572
rect 10685 10568 10916 10570
rect 10980 10570 10986 10572
rect 10685 10512 10690 10568
rect 10746 10512 10874 10568
rect 10685 10510 10916 10512
rect 10685 10507 10751 10510
rect 10869 10508 10916 10510
rect 10980 10510 11026 10570
rect 10980 10508 10986 10510
rect 10869 10507 10935 10508
rect 5682 10368 6002 10369
rect 0 10298 800 10328
rect 5682 10304 5690 10368
rect 5754 10304 5770 10368
rect 5834 10304 5850 10368
rect 5914 10304 5930 10368
rect 5994 10304 6002 10368
rect 5682 10303 6002 10304
rect 15157 10368 15477 10369
rect 15157 10304 15165 10368
rect 15229 10304 15245 10368
rect 15309 10304 15325 10368
rect 15389 10304 15405 10368
rect 15469 10304 15477 10368
rect 15157 10303 15477 10304
rect 24633 10368 24953 10369
rect 24633 10304 24641 10368
rect 24705 10304 24721 10368
rect 24785 10304 24801 10368
rect 24865 10304 24881 10368
rect 24945 10304 24953 10368
rect 24633 10303 24953 10304
rect 3969 10298 4035 10301
rect 0 10296 4035 10298
rect 0 10240 3974 10296
rect 4030 10240 4035 10296
rect 0 10238 4035 10240
rect 0 10208 800 10238
rect 3969 10235 4035 10238
rect 10419 9824 10739 9825
rect 10419 9760 10427 9824
rect 10491 9760 10507 9824
rect 10571 9760 10587 9824
rect 10651 9760 10667 9824
rect 10731 9760 10739 9824
rect 10419 9759 10739 9760
rect 19895 9824 20215 9825
rect 19895 9760 19903 9824
rect 19967 9760 19983 9824
rect 20047 9760 20063 9824
rect 20127 9760 20143 9824
rect 20207 9760 20215 9824
rect 19895 9759 20215 9760
rect 27521 9754 27587 9757
rect 29912 9754 30712 9784
rect 27521 9752 30712 9754
rect 27521 9696 27526 9752
rect 27582 9696 30712 9752
rect 27521 9694 30712 9696
rect 27521 9691 27587 9694
rect 29912 9664 30712 9694
rect 5682 9280 6002 9281
rect 5682 9216 5690 9280
rect 5754 9216 5770 9280
rect 5834 9216 5850 9280
rect 5914 9216 5930 9280
rect 5994 9216 6002 9280
rect 5682 9215 6002 9216
rect 15157 9280 15477 9281
rect 15157 9216 15165 9280
rect 15229 9216 15245 9280
rect 15309 9216 15325 9280
rect 15389 9216 15405 9280
rect 15469 9216 15477 9280
rect 15157 9215 15477 9216
rect 24633 9280 24953 9281
rect 24633 9216 24641 9280
rect 24705 9216 24721 9280
rect 24785 9216 24801 9280
rect 24865 9216 24881 9280
rect 24945 9216 24953 9280
rect 24633 9215 24953 9216
rect 0 8938 800 8968
rect 3693 8938 3759 8941
rect 0 8936 3759 8938
rect 0 8880 3698 8936
rect 3754 8880 3759 8936
rect 0 8878 3759 8880
rect 0 8848 800 8878
rect 3693 8875 3759 8878
rect 17493 8938 17559 8941
rect 17493 8936 17602 8938
rect 17493 8880 17498 8936
rect 17554 8880 17602 8936
rect 17493 8875 17602 8880
rect 17542 8802 17602 8875
rect 17677 8802 17743 8805
rect 17542 8800 17743 8802
rect 17542 8744 17682 8800
rect 17738 8744 17743 8800
rect 17542 8742 17743 8744
rect 17677 8739 17743 8742
rect 10419 8736 10739 8737
rect 10419 8672 10427 8736
rect 10491 8672 10507 8736
rect 10571 8672 10587 8736
rect 10651 8672 10667 8736
rect 10731 8672 10739 8736
rect 10419 8671 10739 8672
rect 19895 8736 20215 8737
rect 19895 8672 19903 8736
rect 19967 8672 19983 8736
rect 20047 8672 20063 8736
rect 20127 8672 20143 8736
rect 20207 8672 20215 8736
rect 19895 8671 20215 8672
rect 15745 8394 15811 8397
rect 17769 8394 17835 8397
rect 15745 8392 17835 8394
rect 15745 8336 15750 8392
rect 15806 8336 17774 8392
rect 17830 8336 17835 8392
rect 15745 8334 17835 8336
rect 15745 8331 15811 8334
rect 17769 8331 17835 8334
rect 17125 8258 17191 8261
rect 18597 8258 18663 8261
rect 17125 8256 18663 8258
rect 17125 8200 17130 8256
rect 17186 8200 18602 8256
rect 18658 8200 18663 8256
rect 17125 8198 18663 8200
rect 17125 8195 17191 8198
rect 18597 8195 18663 8198
rect 29085 8258 29151 8261
rect 29912 8258 30712 8288
rect 29085 8256 30712 8258
rect 29085 8200 29090 8256
rect 29146 8200 30712 8256
rect 29085 8198 30712 8200
rect 29085 8195 29151 8198
rect 5682 8192 6002 8193
rect 5682 8128 5690 8192
rect 5754 8128 5770 8192
rect 5834 8128 5850 8192
rect 5914 8128 5930 8192
rect 5994 8128 6002 8192
rect 5682 8127 6002 8128
rect 15157 8192 15477 8193
rect 15157 8128 15165 8192
rect 15229 8128 15245 8192
rect 15309 8128 15325 8192
rect 15389 8128 15405 8192
rect 15469 8128 15477 8192
rect 15157 8127 15477 8128
rect 24633 8192 24953 8193
rect 24633 8128 24641 8192
rect 24705 8128 24721 8192
rect 24785 8128 24801 8192
rect 24865 8128 24881 8192
rect 24945 8128 24953 8192
rect 29912 8168 30712 8198
rect 24633 8127 24953 8128
rect 10419 7648 10739 7649
rect 0 7578 800 7608
rect 10419 7584 10427 7648
rect 10491 7584 10507 7648
rect 10571 7584 10587 7648
rect 10651 7584 10667 7648
rect 10731 7584 10739 7648
rect 10419 7583 10739 7584
rect 19895 7648 20215 7649
rect 19895 7584 19903 7648
rect 19967 7584 19983 7648
rect 20047 7584 20063 7648
rect 20127 7584 20143 7648
rect 20207 7584 20215 7648
rect 19895 7583 20215 7584
rect 4061 7578 4127 7581
rect 0 7576 4127 7578
rect 0 7520 4066 7576
rect 4122 7520 4127 7576
rect 0 7518 4127 7520
rect 0 7488 800 7518
rect 4061 7515 4127 7518
rect 5682 7104 6002 7105
rect 5682 7040 5690 7104
rect 5754 7040 5770 7104
rect 5834 7040 5850 7104
rect 5914 7040 5930 7104
rect 5994 7040 6002 7104
rect 5682 7039 6002 7040
rect 15157 7104 15477 7105
rect 15157 7040 15165 7104
rect 15229 7040 15245 7104
rect 15309 7040 15325 7104
rect 15389 7040 15405 7104
rect 15469 7040 15477 7104
rect 15157 7039 15477 7040
rect 24633 7104 24953 7105
rect 24633 7040 24641 7104
rect 24705 7040 24721 7104
rect 24785 7040 24801 7104
rect 24865 7040 24881 7104
rect 24945 7040 24953 7104
rect 24633 7039 24953 7040
rect 27429 6762 27495 6765
rect 29912 6762 30712 6792
rect 27429 6760 30712 6762
rect 27429 6704 27434 6760
rect 27490 6704 30712 6760
rect 27429 6702 30712 6704
rect 27429 6699 27495 6702
rect 29912 6672 30712 6702
rect 10419 6560 10739 6561
rect 10419 6496 10427 6560
rect 10491 6496 10507 6560
rect 10571 6496 10587 6560
rect 10651 6496 10667 6560
rect 10731 6496 10739 6560
rect 10419 6495 10739 6496
rect 19895 6560 20215 6561
rect 19895 6496 19903 6560
rect 19967 6496 19983 6560
rect 20047 6496 20063 6560
rect 20127 6496 20143 6560
rect 20207 6496 20215 6560
rect 19895 6495 20215 6496
rect 0 6218 800 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 800 6158
rect 4061 6155 4127 6158
rect 5682 6016 6002 6017
rect 5682 5952 5690 6016
rect 5754 5952 5770 6016
rect 5834 5952 5850 6016
rect 5914 5952 5930 6016
rect 5994 5952 6002 6016
rect 5682 5951 6002 5952
rect 15157 6016 15477 6017
rect 15157 5952 15165 6016
rect 15229 5952 15245 6016
rect 15309 5952 15325 6016
rect 15389 5952 15405 6016
rect 15469 5952 15477 6016
rect 15157 5951 15477 5952
rect 24633 6016 24953 6017
rect 24633 5952 24641 6016
rect 24705 5952 24721 6016
rect 24785 5952 24801 6016
rect 24865 5952 24881 6016
rect 24945 5952 24953 6016
rect 24633 5951 24953 5952
rect 10419 5472 10739 5473
rect 10419 5408 10427 5472
rect 10491 5408 10507 5472
rect 10571 5408 10587 5472
rect 10651 5408 10667 5472
rect 10731 5408 10739 5472
rect 10419 5407 10739 5408
rect 19895 5472 20215 5473
rect 19895 5408 19903 5472
rect 19967 5408 19983 5472
rect 20047 5408 20063 5472
rect 20127 5408 20143 5472
rect 20207 5408 20215 5472
rect 19895 5407 20215 5408
rect 27521 5266 27587 5269
rect 29912 5266 30712 5296
rect 27521 5264 30712 5266
rect 27521 5208 27526 5264
rect 27582 5208 30712 5264
rect 27521 5206 30712 5208
rect 27521 5203 27587 5206
rect 29912 5176 30712 5206
rect 19701 5130 19767 5133
rect 26601 5130 26667 5133
rect 19701 5128 26667 5130
rect 19701 5072 19706 5128
rect 19762 5072 26606 5128
rect 26662 5072 26667 5128
rect 19701 5070 26667 5072
rect 19701 5067 19767 5070
rect 26601 5067 26667 5070
rect 5682 4928 6002 4929
rect 0 4858 800 4888
rect 5682 4864 5690 4928
rect 5754 4864 5770 4928
rect 5834 4864 5850 4928
rect 5914 4864 5930 4928
rect 5994 4864 6002 4928
rect 5682 4863 6002 4864
rect 15157 4928 15477 4929
rect 15157 4864 15165 4928
rect 15229 4864 15245 4928
rect 15309 4864 15325 4928
rect 15389 4864 15405 4928
rect 15469 4864 15477 4928
rect 15157 4863 15477 4864
rect 24633 4928 24953 4929
rect 24633 4864 24641 4928
rect 24705 4864 24721 4928
rect 24785 4864 24801 4928
rect 24865 4864 24881 4928
rect 24945 4864 24953 4928
rect 24633 4863 24953 4864
rect 3877 4858 3943 4861
rect 0 4856 3943 4858
rect 0 4800 3882 4856
rect 3938 4800 3943 4856
rect 0 4798 3943 4800
rect 0 4768 800 4798
rect 3877 4795 3943 4798
rect 10419 4384 10739 4385
rect 10419 4320 10427 4384
rect 10491 4320 10507 4384
rect 10571 4320 10587 4384
rect 10651 4320 10667 4384
rect 10731 4320 10739 4384
rect 10419 4319 10739 4320
rect 19895 4384 20215 4385
rect 19895 4320 19903 4384
rect 19967 4320 19983 4384
rect 20047 4320 20063 4384
rect 20127 4320 20143 4384
rect 20207 4320 20215 4384
rect 19895 4319 20215 4320
rect 17769 4178 17835 4181
rect 18321 4178 18387 4181
rect 17769 4176 18387 4178
rect 17769 4120 17774 4176
rect 17830 4120 18326 4176
rect 18382 4120 18387 4176
rect 17769 4118 18387 4120
rect 17769 4115 17835 4118
rect 18321 4115 18387 4118
rect 13302 3980 13308 4044
rect 13372 4042 13378 4044
rect 19609 4042 19675 4045
rect 13372 4040 19675 4042
rect 13372 3984 19614 4040
rect 19670 3984 19675 4040
rect 13372 3982 19675 3984
rect 13372 3980 13378 3982
rect 19609 3979 19675 3982
rect 5682 3840 6002 3841
rect 5682 3776 5690 3840
rect 5754 3776 5770 3840
rect 5834 3776 5850 3840
rect 5914 3776 5930 3840
rect 5994 3776 6002 3840
rect 5682 3775 6002 3776
rect 15157 3840 15477 3841
rect 15157 3776 15165 3840
rect 15229 3776 15245 3840
rect 15309 3776 15325 3840
rect 15389 3776 15405 3840
rect 15469 3776 15477 3840
rect 15157 3775 15477 3776
rect 24633 3840 24953 3841
rect 24633 3776 24641 3840
rect 24705 3776 24721 3840
rect 24785 3776 24801 3840
rect 24865 3776 24881 3840
rect 24945 3776 24953 3840
rect 24633 3775 24953 3776
rect 17217 3770 17283 3773
rect 18873 3770 18939 3773
rect 17217 3768 18939 3770
rect 17217 3712 17222 3768
rect 17278 3712 18878 3768
rect 18934 3712 18939 3768
rect 17217 3710 18939 3712
rect 17217 3707 17283 3710
rect 18873 3707 18939 3710
rect 27061 3770 27127 3773
rect 29912 3770 30712 3800
rect 27061 3768 30712 3770
rect 27061 3712 27066 3768
rect 27122 3712 30712 3768
rect 27061 3710 30712 3712
rect 27061 3707 27127 3710
rect 29912 3680 30712 3710
rect 0 3498 800 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 800 3438
rect 1853 3435 1919 3438
rect 17585 3498 17651 3501
rect 26417 3498 26483 3501
rect 17585 3496 26483 3498
rect 17585 3440 17590 3496
rect 17646 3440 26422 3496
rect 26478 3440 26483 3496
rect 17585 3438 26483 3440
rect 17585 3435 17651 3438
rect 26417 3435 26483 3438
rect 16757 3362 16823 3365
rect 18873 3362 18939 3365
rect 16757 3360 18939 3362
rect 16757 3304 16762 3360
rect 16818 3304 18878 3360
rect 18934 3304 18939 3360
rect 16757 3302 18939 3304
rect 16757 3299 16823 3302
rect 18873 3299 18939 3302
rect 10419 3296 10739 3297
rect 10419 3232 10427 3296
rect 10491 3232 10507 3296
rect 10571 3232 10587 3296
rect 10651 3232 10667 3296
rect 10731 3232 10739 3296
rect 10419 3231 10739 3232
rect 19895 3296 20215 3297
rect 19895 3232 19903 3296
rect 19967 3232 19983 3296
rect 20047 3232 20063 3296
rect 20127 3232 20143 3296
rect 20207 3232 20215 3296
rect 19895 3231 20215 3232
rect 14457 3226 14523 3229
rect 18965 3226 19031 3229
rect 14457 3224 19031 3226
rect 14457 3168 14462 3224
rect 14518 3168 18970 3224
rect 19026 3168 19031 3224
rect 14457 3166 19031 3168
rect 14457 3163 14523 3166
rect 18965 3163 19031 3166
rect 5682 2752 6002 2753
rect 5682 2688 5690 2752
rect 5754 2688 5770 2752
rect 5834 2688 5850 2752
rect 5914 2688 5930 2752
rect 5994 2688 6002 2752
rect 5682 2687 6002 2688
rect 15157 2752 15477 2753
rect 15157 2688 15165 2752
rect 15229 2688 15245 2752
rect 15309 2688 15325 2752
rect 15389 2688 15405 2752
rect 15469 2688 15477 2752
rect 15157 2687 15477 2688
rect 24633 2752 24953 2753
rect 24633 2688 24641 2752
rect 24705 2688 24721 2752
rect 24785 2688 24801 2752
rect 24865 2688 24881 2752
rect 24945 2688 24953 2752
rect 24633 2687 24953 2688
rect 26509 2274 26575 2277
rect 29912 2274 30712 2304
rect 26509 2272 30712 2274
rect 26509 2216 26514 2272
rect 26570 2216 30712 2272
rect 26509 2214 30712 2216
rect 26509 2211 26575 2214
rect 10419 2208 10739 2209
rect 0 2138 800 2168
rect 10419 2144 10427 2208
rect 10491 2144 10507 2208
rect 10571 2144 10587 2208
rect 10651 2144 10667 2208
rect 10731 2144 10739 2208
rect 10419 2143 10739 2144
rect 19895 2208 20215 2209
rect 19895 2144 19903 2208
rect 19967 2144 19983 2208
rect 20047 2144 20063 2208
rect 20127 2144 20143 2208
rect 20207 2144 20215 2208
rect 29912 2184 30712 2214
rect 19895 2143 20215 2144
rect 3417 2138 3483 2141
rect 0 2136 3483 2138
rect 0 2080 3422 2136
rect 3478 2080 3483 2136
rect 0 2078 3483 2080
rect 0 2048 800 2078
rect 3417 2075 3483 2078
rect 0 778 800 808
rect 3141 778 3207 781
rect 0 776 3207 778
rect 0 720 3146 776
rect 3202 720 3207 776
rect 0 718 3207 720
rect 0 688 800 718
rect 3141 715 3207 718
rect 27521 778 27587 781
rect 29912 778 30712 808
rect 27521 776 30712 778
rect 27521 720 27526 776
rect 27582 720 30712 776
rect 27521 718 30712 720
rect 27521 715 27587 718
rect 29912 688 30712 718
<< via3 >>
rect 10427 30492 10491 30496
rect 10427 30436 10431 30492
rect 10431 30436 10487 30492
rect 10487 30436 10491 30492
rect 10427 30432 10491 30436
rect 10507 30492 10571 30496
rect 10507 30436 10511 30492
rect 10511 30436 10567 30492
rect 10567 30436 10571 30492
rect 10507 30432 10571 30436
rect 10587 30492 10651 30496
rect 10587 30436 10591 30492
rect 10591 30436 10647 30492
rect 10647 30436 10651 30492
rect 10587 30432 10651 30436
rect 10667 30492 10731 30496
rect 10667 30436 10671 30492
rect 10671 30436 10727 30492
rect 10727 30436 10731 30492
rect 10667 30432 10731 30436
rect 19903 30492 19967 30496
rect 19903 30436 19907 30492
rect 19907 30436 19963 30492
rect 19963 30436 19967 30492
rect 19903 30432 19967 30436
rect 19983 30492 20047 30496
rect 19983 30436 19987 30492
rect 19987 30436 20043 30492
rect 20043 30436 20047 30492
rect 19983 30432 20047 30436
rect 20063 30492 20127 30496
rect 20063 30436 20067 30492
rect 20067 30436 20123 30492
rect 20123 30436 20127 30492
rect 20063 30432 20127 30436
rect 20143 30492 20207 30496
rect 20143 30436 20147 30492
rect 20147 30436 20203 30492
rect 20203 30436 20207 30492
rect 20143 30432 20207 30436
rect 5690 29948 5754 29952
rect 5690 29892 5694 29948
rect 5694 29892 5750 29948
rect 5750 29892 5754 29948
rect 5690 29888 5754 29892
rect 5770 29948 5834 29952
rect 5770 29892 5774 29948
rect 5774 29892 5830 29948
rect 5830 29892 5834 29948
rect 5770 29888 5834 29892
rect 5850 29948 5914 29952
rect 5850 29892 5854 29948
rect 5854 29892 5910 29948
rect 5910 29892 5914 29948
rect 5850 29888 5914 29892
rect 5930 29948 5994 29952
rect 5930 29892 5934 29948
rect 5934 29892 5990 29948
rect 5990 29892 5994 29948
rect 5930 29888 5994 29892
rect 15165 29948 15229 29952
rect 15165 29892 15169 29948
rect 15169 29892 15225 29948
rect 15225 29892 15229 29948
rect 15165 29888 15229 29892
rect 15245 29948 15309 29952
rect 15245 29892 15249 29948
rect 15249 29892 15305 29948
rect 15305 29892 15309 29948
rect 15245 29888 15309 29892
rect 15325 29948 15389 29952
rect 15325 29892 15329 29948
rect 15329 29892 15385 29948
rect 15385 29892 15389 29948
rect 15325 29888 15389 29892
rect 15405 29948 15469 29952
rect 15405 29892 15409 29948
rect 15409 29892 15465 29948
rect 15465 29892 15469 29948
rect 15405 29888 15469 29892
rect 24641 29948 24705 29952
rect 24641 29892 24645 29948
rect 24645 29892 24701 29948
rect 24701 29892 24705 29948
rect 24641 29888 24705 29892
rect 24721 29948 24785 29952
rect 24721 29892 24725 29948
rect 24725 29892 24781 29948
rect 24781 29892 24785 29948
rect 24721 29888 24785 29892
rect 24801 29948 24865 29952
rect 24801 29892 24805 29948
rect 24805 29892 24861 29948
rect 24861 29892 24865 29948
rect 24801 29888 24865 29892
rect 24881 29948 24945 29952
rect 24881 29892 24885 29948
rect 24885 29892 24941 29948
rect 24941 29892 24945 29948
rect 24881 29888 24945 29892
rect 10427 29404 10491 29408
rect 10427 29348 10431 29404
rect 10431 29348 10487 29404
rect 10487 29348 10491 29404
rect 10427 29344 10491 29348
rect 10507 29404 10571 29408
rect 10507 29348 10511 29404
rect 10511 29348 10567 29404
rect 10567 29348 10571 29404
rect 10507 29344 10571 29348
rect 10587 29404 10651 29408
rect 10587 29348 10591 29404
rect 10591 29348 10647 29404
rect 10647 29348 10651 29404
rect 10587 29344 10651 29348
rect 10667 29404 10731 29408
rect 10667 29348 10671 29404
rect 10671 29348 10727 29404
rect 10727 29348 10731 29404
rect 10667 29344 10731 29348
rect 19903 29404 19967 29408
rect 19903 29348 19907 29404
rect 19907 29348 19963 29404
rect 19963 29348 19967 29404
rect 19903 29344 19967 29348
rect 19983 29404 20047 29408
rect 19983 29348 19987 29404
rect 19987 29348 20043 29404
rect 20043 29348 20047 29404
rect 19983 29344 20047 29348
rect 20063 29404 20127 29408
rect 20063 29348 20067 29404
rect 20067 29348 20123 29404
rect 20123 29348 20127 29404
rect 20063 29344 20127 29348
rect 20143 29404 20207 29408
rect 20143 29348 20147 29404
rect 20147 29348 20203 29404
rect 20203 29348 20207 29404
rect 20143 29344 20207 29348
rect 5690 28860 5754 28864
rect 5690 28804 5694 28860
rect 5694 28804 5750 28860
rect 5750 28804 5754 28860
rect 5690 28800 5754 28804
rect 5770 28860 5834 28864
rect 5770 28804 5774 28860
rect 5774 28804 5830 28860
rect 5830 28804 5834 28860
rect 5770 28800 5834 28804
rect 5850 28860 5914 28864
rect 5850 28804 5854 28860
rect 5854 28804 5910 28860
rect 5910 28804 5914 28860
rect 5850 28800 5914 28804
rect 5930 28860 5994 28864
rect 5930 28804 5934 28860
rect 5934 28804 5990 28860
rect 5990 28804 5994 28860
rect 5930 28800 5994 28804
rect 15165 28860 15229 28864
rect 15165 28804 15169 28860
rect 15169 28804 15225 28860
rect 15225 28804 15229 28860
rect 15165 28800 15229 28804
rect 15245 28860 15309 28864
rect 15245 28804 15249 28860
rect 15249 28804 15305 28860
rect 15305 28804 15309 28860
rect 15245 28800 15309 28804
rect 15325 28860 15389 28864
rect 15325 28804 15329 28860
rect 15329 28804 15385 28860
rect 15385 28804 15389 28860
rect 15325 28800 15389 28804
rect 15405 28860 15469 28864
rect 15405 28804 15409 28860
rect 15409 28804 15465 28860
rect 15465 28804 15469 28860
rect 15405 28800 15469 28804
rect 24641 28860 24705 28864
rect 24641 28804 24645 28860
rect 24645 28804 24701 28860
rect 24701 28804 24705 28860
rect 24641 28800 24705 28804
rect 24721 28860 24785 28864
rect 24721 28804 24725 28860
rect 24725 28804 24781 28860
rect 24781 28804 24785 28860
rect 24721 28800 24785 28804
rect 24801 28860 24865 28864
rect 24801 28804 24805 28860
rect 24805 28804 24861 28860
rect 24861 28804 24865 28860
rect 24801 28800 24865 28804
rect 24881 28860 24945 28864
rect 24881 28804 24885 28860
rect 24885 28804 24941 28860
rect 24941 28804 24945 28860
rect 24881 28800 24945 28804
rect 10427 28316 10491 28320
rect 10427 28260 10431 28316
rect 10431 28260 10487 28316
rect 10487 28260 10491 28316
rect 10427 28256 10491 28260
rect 10507 28316 10571 28320
rect 10507 28260 10511 28316
rect 10511 28260 10567 28316
rect 10567 28260 10571 28316
rect 10507 28256 10571 28260
rect 10587 28316 10651 28320
rect 10587 28260 10591 28316
rect 10591 28260 10647 28316
rect 10647 28260 10651 28316
rect 10587 28256 10651 28260
rect 10667 28316 10731 28320
rect 10667 28260 10671 28316
rect 10671 28260 10727 28316
rect 10727 28260 10731 28316
rect 10667 28256 10731 28260
rect 19903 28316 19967 28320
rect 19903 28260 19907 28316
rect 19907 28260 19963 28316
rect 19963 28260 19967 28316
rect 19903 28256 19967 28260
rect 19983 28316 20047 28320
rect 19983 28260 19987 28316
rect 19987 28260 20043 28316
rect 20043 28260 20047 28316
rect 19983 28256 20047 28260
rect 20063 28316 20127 28320
rect 20063 28260 20067 28316
rect 20067 28260 20123 28316
rect 20123 28260 20127 28316
rect 20063 28256 20127 28260
rect 20143 28316 20207 28320
rect 20143 28260 20147 28316
rect 20147 28260 20203 28316
rect 20203 28260 20207 28316
rect 20143 28256 20207 28260
rect 5690 27772 5754 27776
rect 5690 27716 5694 27772
rect 5694 27716 5750 27772
rect 5750 27716 5754 27772
rect 5690 27712 5754 27716
rect 5770 27772 5834 27776
rect 5770 27716 5774 27772
rect 5774 27716 5830 27772
rect 5830 27716 5834 27772
rect 5770 27712 5834 27716
rect 5850 27772 5914 27776
rect 5850 27716 5854 27772
rect 5854 27716 5910 27772
rect 5910 27716 5914 27772
rect 5850 27712 5914 27716
rect 5930 27772 5994 27776
rect 5930 27716 5934 27772
rect 5934 27716 5990 27772
rect 5990 27716 5994 27772
rect 5930 27712 5994 27716
rect 15165 27772 15229 27776
rect 15165 27716 15169 27772
rect 15169 27716 15225 27772
rect 15225 27716 15229 27772
rect 15165 27712 15229 27716
rect 15245 27772 15309 27776
rect 15245 27716 15249 27772
rect 15249 27716 15305 27772
rect 15305 27716 15309 27772
rect 15245 27712 15309 27716
rect 15325 27772 15389 27776
rect 15325 27716 15329 27772
rect 15329 27716 15385 27772
rect 15385 27716 15389 27772
rect 15325 27712 15389 27716
rect 15405 27772 15469 27776
rect 15405 27716 15409 27772
rect 15409 27716 15465 27772
rect 15465 27716 15469 27772
rect 15405 27712 15469 27716
rect 24641 27772 24705 27776
rect 24641 27716 24645 27772
rect 24645 27716 24701 27772
rect 24701 27716 24705 27772
rect 24641 27712 24705 27716
rect 24721 27772 24785 27776
rect 24721 27716 24725 27772
rect 24725 27716 24781 27772
rect 24781 27716 24785 27772
rect 24721 27712 24785 27716
rect 24801 27772 24865 27776
rect 24801 27716 24805 27772
rect 24805 27716 24861 27772
rect 24861 27716 24865 27772
rect 24801 27712 24865 27716
rect 24881 27772 24945 27776
rect 24881 27716 24885 27772
rect 24885 27716 24941 27772
rect 24941 27716 24945 27772
rect 24881 27712 24945 27716
rect 13308 27296 13372 27300
rect 13308 27240 13322 27296
rect 13322 27240 13372 27296
rect 13308 27236 13372 27240
rect 10427 27228 10491 27232
rect 10427 27172 10431 27228
rect 10431 27172 10487 27228
rect 10487 27172 10491 27228
rect 10427 27168 10491 27172
rect 10507 27228 10571 27232
rect 10507 27172 10511 27228
rect 10511 27172 10567 27228
rect 10567 27172 10571 27228
rect 10507 27168 10571 27172
rect 10587 27228 10651 27232
rect 10587 27172 10591 27228
rect 10591 27172 10647 27228
rect 10647 27172 10651 27228
rect 10587 27168 10651 27172
rect 10667 27228 10731 27232
rect 10667 27172 10671 27228
rect 10671 27172 10727 27228
rect 10727 27172 10731 27228
rect 10667 27168 10731 27172
rect 19903 27228 19967 27232
rect 19903 27172 19907 27228
rect 19907 27172 19963 27228
rect 19963 27172 19967 27228
rect 19903 27168 19967 27172
rect 19983 27228 20047 27232
rect 19983 27172 19987 27228
rect 19987 27172 20043 27228
rect 20043 27172 20047 27228
rect 19983 27168 20047 27172
rect 20063 27228 20127 27232
rect 20063 27172 20067 27228
rect 20067 27172 20123 27228
rect 20123 27172 20127 27228
rect 20063 27168 20127 27172
rect 20143 27228 20207 27232
rect 20143 27172 20147 27228
rect 20147 27172 20203 27228
rect 20203 27172 20207 27228
rect 20143 27168 20207 27172
rect 5690 26684 5754 26688
rect 5690 26628 5694 26684
rect 5694 26628 5750 26684
rect 5750 26628 5754 26684
rect 5690 26624 5754 26628
rect 5770 26684 5834 26688
rect 5770 26628 5774 26684
rect 5774 26628 5830 26684
rect 5830 26628 5834 26684
rect 5770 26624 5834 26628
rect 5850 26684 5914 26688
rect 5850 26628 5854 26684
rect 5854 26628 5910 26684
rect 5910 26628 5914 26684
rect 5850 26624 5914 26628
rect 5930 26684 5994 26688
rect 5930 26628 5934 26684
rect 5934 26628 5990 26684
rect 5990 26628 5994 26684
rect 5930 26624 5994 26628
rect 15165 26684 15229 26688
rect 15165 26628 15169 26684
rect 15169 26628 15225 26684
rect 15225 26628 15229 26684
rect 15165 26624 15229 26628
rect 15245 26684 15309 26688
rect 15245 26628 15249 26684
rect 15249 26628 15305 26684
rect 15305 26628 15309 26684
rect 15245 26624 15309 26628
rect 15325 26684 15389 26688
rect 15325 26628 15329 26684
rect 15329 26628 15385 26684
rect 15385 26628 15389 26684
rect 15325 26624 15389 26628
rect 15405 26684 15469 26688
rect 15405 26628 15409 26684
rect 15409 26628 15465 26684
rect 15465 26628 15469 26684
rect 15405 26624 15469 26628
rect 24641 26684 24705 26688
rect 24641 26628 24645 26684
rect 24645 26628 24701 26684
rect 24701 26628 24705 26684
rect 24641 26624 24705 26628
rect 24721 26684 24785 26688
rect 24721 26628 24725 26684
rect 24725 26628 24781 26684
rect 24781 26628 24785 26684
rect 24721 26624 24785 26628
rect 24801 26684 24865 26688
rect 24801 26628 24805 26684
rect 24805 26628 24861 26684
rect 24861 26628 24865 26684
rect 24801 26624 24865 26628
rect 24881 26684 24945 26688
rect 24881 26628 24885 26684
rect 24885 26628 24941 26684
rect 24941 26628 24945 26684
rect 24881 26624 24945 26628
rect 10427 26140 10491 26144
rect 10427 26084 10431 26140
rect 10431 26084 10487 26140
rect 10487 26084 10491 26140
rect 10427 26080 10491 26084
rect 10507 26140 10571 26144
rect 10507 26084 10511 26140
rect 10511 26084 10567 26140
rect 10567 26084 10571 26140
rect 10507 26080 10571 26084
rect 10587 26140 10651 26144
rect 10587 26084 10591 26140
rect 10591 26084 10647 26140
rect 10647 26084 10651 26140
rect 10587 26080 10651 26084
rect 10667 26140 10731 26144
rect 10667 26084 10671 26140
rect 10671 26084 10727 26140
rect 10727 26084 10731 26140
rect 10667 26080 10731 26084
rect 19903 26140 19967 26144
rect 19903 26084 19907 26140
rect 19907 26084 19963 26140
rect 19963 26084 19967 26140
rect 19903 26080 19967 26084
rect 19983 26140 20047 26144
rect 19983 26084 19987 26140
rect 19987 26084 20043 26140
rect 20043 26084 20047 26140
rect 19983 26080 20047 26084
rect 20063 26140 20127 26144
rect 20063 26084 20067 26140
rect 20067 26084 20123 26140
rect 20123 26084 20127 26140
rect 20063 26080 20127 26084
rect 20143 26140 20207 26144
rect 20143 26084 20147 26140
rect 20147 26084 20203 26140
rect 20203 26084 20207 26140
rect 20143 26080 20207 26084
rect 5690 25596 5754 25600
rect 5690 25540 5694 25596
rect 5694 25540 5750 25596
rect 5750 25540 5754 25596
rect 5690 25536 5754 25540
rect 5770 25596 5834 25600
rect 5770 25540 5774 25596
rect 5774 25540 5830 25596
rect 5830 25540 5834 25596
rect 5770 25536 5834 25540
rect 5850 25596 5914 25600
rect 5850 25540 5854 25596
rect 5854 25540 5910 25596
rect 5910 25540 5914 25596
rect 5850 25536 5914 25540
rect 5930 25596 5994 25600
rect 5930 25540 5934 25596
rect 5934 25540 5990 25596
rect 5990 25540 5994 25596
rect 5930 25536 5994 25540
rect 15165 25596 15229 25600
rect 15165 25540 15169 25596
rect 15169 25540 15225 25596
rect 15225 25540 15229 25596
rect 15165 25536 15229 25540
rect 15245 25596 15309 25600
rect 15245 25540 15249 25596
rect 15249 25540 15305 25596
rect 15305 25540 15309 25596
rect 15245 25536 15309 25540
rect 15325 25596 15389 25600
rect 15325 25540 15329 25596
rect 15329 25540 15385 25596
rect 15385 25540 15389 25596
rect 15325 25536 15389 25540
rect 15405 25596 15469 25600
rect 15405 25540 15409 25596
rect 15409 25540 15465 25596
rect 15465 25540 15469 25596
rect 15405 25536 15469 25540
rect 24641 25596 24705 25600
rect 24641 25540 24645 25596
rect 24645 25540 24701 25596
rect 24701 25540 24705 25596
rect 24641 25536 24705 25540
rect 24721 25596 24785 25600
rect 24721 25540 24725 25596
rect 24725 25540 24781 25596
rect 24781 25540 24785 25596
rect 24721 25536 24785 25540
rect 24801 25596 24865 25600
rect 24801 25540 24805 25596
rect 24805 25540 24861 25596
rect 24861 25540 24865 25596
rect 24801 25536 24865 25540
rect 24881 25596 24945 25600
rect 24881 25540 24885 25596
rect 24885 25540 24941 25596
rect 24941 25540 24945 25596
rect 24881 25536 24945 25540
rect 20484 25196 20548 25260
rect 10427 25052 10491 25056
rect 10427 24996 10431 25052
rect 10431 24996 10487 25052
rect 10487 24996 10491 25052
rect 10427 24992 10491 24996
rect 10507 25052 10571 25056
rect 10507 24996 10511 25052
rect 10511 24996 10567 25052
rect 10567 24996 10571 25052
rect 10507 24992 10571 24996
rect 10587 25052 10651 25056
rect 10587 24996 10591 25052
rect 10591 24996 10647 25052
rect 10647 24996 10651 25052
rect 10587 24992 10651 24996
rect 10667 25052 10731 25056
rect 10667 24996 10671 25052
rect 10671 24996 10727 25052
rect 10727 24996 10731 25052
rect 10667 24992 10731 24996
rect 19903 25052 19967 25056
rect 19903 24996 19907 25052
rect 19907 24996 19963 25052
rect 19963 24996 19967 25052
rect 19903 24992 19967 24996
rect 19983 25052 20047 25056
rect 19983 24996 19987 25052
rect 19987 24996 20043 25052
rect 20043 24996 20047 25052
rect 19983 24992 20047 24996
rect 20063 25052 20127 25056
rect 20063 24996 20067 25052
rect 20067 24996 20123 25052
rect 20123 24996 20127 25052
rect 20063 24992 20127 24996
rect 20143 25052 20207 25056
rect 20143 24996 20147 25052
rect 20147 24996 20203 25052
rect 20203 24996 20207 25052
rect 20143 24992 20207 24996
rect 5690 24508 5754 24512
rect 5690 24452 5694 24508
rect 5694 24452 5750 24508
rect 5750 24452 5754 24508
rect 5690 24448 5754 24452
rect 5770 24508 5834 24512
rect 5770 24452 5774 24508
rect 5774 24452 5830 24508
rect 5830 24452 5834 24508
rect 5770 24448 5834 24452
rect 5850 24508 5914 24512
rect 5850 24452 5854 24508
rect 5854 24452 5910 24508
rect 5910 24452 5914 24508
rect 5850 24448 5914 24452
rect 5930 24508 5994 24512
rect 5930 24452 5934 24508
rect 5934 24452 5990 24508
rect 5990 24452 5994 24508
rect 5930 24448 5994 24452
rect 15165 24508 15229 24512
rect 15165 24452 15169 24508
rect 15169 24452 15225 24508
rect 15225 24452 15229 24508
rect 15165 24448 15229 24452
rect 15245 24508 15309 24512
rect 15245 24452 15249 24508
rect 15249 24452 15305 24508
rect 15305 24452 15309 24508
rect 15245 24448 15309 24452
rect 15325 24508 15389 24512
rect 15325 24452 15329 24508
rect 15329 24452 15385 24508
rect 15385 24452 15389 24508
rect 15325 24448 15389 24452
rect 15405 24508 15469 24512
rect 15405 24452 15409 24508
rect 15409 24452 15465 24508
rect 15465 24452 15469 24508
rect 15405 24448 15469 24452
rect 24641 24508 24705 24512
rect 24641 24452 24645 24508
rect 24645 24452 24701 24508
rect 24701 24452 24705 24508
rect 24641 24448 24705 24452
rect 24721 24508 24785 24512
rect 24721 24452 24725 24508
rect 24725 24452 24781 24508
rect 24781 24452 24785 24508
rect 24721 24448 24785 24452
rect 24801 24508 24865 24512
rect 24801 24452 24805 24508
rect 24805 24452 24861 24508
rect 24861 24452 24865 24508
rect 24801 24448 24865 24452
rect 24881 24508 24945 24512
rect 24881 24452 24885 24508
rect 24885 24452 24941 24508
rect 24941 24452 24945 24508
rect 24881 24448 24945 24452
rect 10427 23964 10491 23968
rect 10427 23908 10431 23964
rect 10431 23908 10487 23964
rect 10487 23908 10491 23964
rect 10427 23904 10491 23908
rect 10507 23964 10571 23968
rect 10507 23908 10511 23964
rect 10511 23908 10567 23964
rect 10567 23908 10571 23964
rect 10507 23904 10571 23908
rect 10587 23964 10651 23968
rect 10587 23908 10591 23964
rect 10591 23908 10647 23964
rect 10647 23908 10651 23964
rect 10587 23904 10651 23908
rect 10667 23964 10731 23968
rect 10667 23908 10671 23964
rect 10671 23908 10727 23964
rect 10727 23908 10731 23964
rect 10667 23904 10731 23908
rect 19903 23964 19967 23968
rect 19903 23908 19907 23964
rect 19907 23908 19963 23964
rect 19963 23908 19967 23964
rect 19903 23904 19967 23908
rect 19983 23964 20047 23968
rect 19983 23908 19987 23964
rect 19987 23908 20043 23964
rect 20043 23908 20047 23964
rect 19983 23904 20047 23908
rect 20063 23964 20127 23968
rect 20063 23908 20067 23964
rect 20067 23908 20123 23964
rect 20123 23908 20127 23964
rect 20063 23904 20127 23908
rect 20143 23964 20207 23968
rect 20143 23908 20147 23964
rect 20147 23908 20203 23964
rect 20203 23908 20207 23964
rect 20143 23904 20207 23908
rect 19748 23564 19812 23628
rect 13676 23428 13740 23492
rect 5690 23420 5754 23424
rect 5690 23364 5694 23420
rect 5694 23364 5750 23420
rect 5750 23364 5754 23420
rect 5690 23360 5754 23364
rect 5770 23420 5834 23424
rect 5770 23364 5774 23420
rect 5774 23364 5830 23420
rect 5830 23364 5834 23420
rect 5770 23360 5834 23364
rect 5850 23420 5914 23424
rect 5850 23364 5854 23420
rect 5854 23364 5910 23420
rect 5910 23364 5914 23420
rect 5850 23360 5914 23364
rect 5930 23420 5994 23424
rect 5930 23364 5934 23420
rect 5934 23364 5990 23420
rect 5990 23364 5994 23420
rect 5930 23360 5994 23364
rect 15165 23420 15229 23424
rect 15165 23364 15169 23420
rect 15169 23364 15225 23420
rect 15225 23364 15229 23420
rect 15165 23360 15229 23364
rect 15245 23420 15309 23424
rect 15245 23364 15249 23420
rect 15249 23364 15305 23420
rect 15305 23364 15309 23420
rect 15245 23360 15309 23364
rect 15325 23420 15389 23424
rect 15325 23364 15329 23420
rect 15329 23364 15385 23420
rect 15385 23364 15389 23420
rect 15325 23360 15389 23364
rect 15405 23420 15469 23424
rect 15405 23364 15409 23420
rect 15409 23364 15465 23420
rect 15465 23364 15469 23420
rect 15405 23360 15469 23364
rect 24641 23420 24705 23424
rect 24641 23364 24645 23420
rect 24645 23364 24701 23420
rect 24701 23364 24705 23420
rect 24641 23360 24705 23364
rect 24721 23420 24785 23424
rect 24721 23364 24725 23420
rect 24725 23364 24781 23420
rect 24781 23364 24785 23420
rect 24721 23360 24785 23364
rect 24801 23420 24865 23424
rect 24801 23364 24805 23420
rect 24805 23364 24861 23420
rect 24861 23364 24865 23420
rect 24801 23360 24865 23364
rect 24881 23420 24945 23424
rect 24881 23364 24885 23420
rect 24885 23364 24941 23420
rect 24941 23364 24945 23420
rect 24881 23360 24945 23364
rect 10427 22876 10491 22880
rect 10427 22820 10431 22876
rect 10431 22820 10487 22876
rect 10487 22820 10491 22876
rect 10427 22816 10491 22820
rect 10507 22876 10571 22880
rect 10507 22820 10511 22876
rect 10511 22820 10567 22876
rect 10567 22820 10571 22876
rect 10507 22816 10571 22820
rect 10587 22876 10651 22880
rect 10587 22820 10591 22876
rect 10591 22820 10647 22876
rect 10647 22820 10651 22876
rect 10587 22816 10651 22820
rect 10667 22876 10731 22880
rect 10667 22820 10671 22876
rect 10671 22820 10727 22876
rect 10727 22820 10731 22876
rect 10667 22816 10731 22820
rect 19903 22876 19967 22880
rect 19903 22820 19907 22876
rect 19907 22820 19963 22876
rect 19963 22820 19967 22876
rect 19903 22816 19967 22820
rect 19983 22876 20047 22880
rect 19983 22820 19987 22876
rect 19987 22820 20043 22876
rect 20043 22820 20047 22876
rect 19983 22816 20047 22820
rect 20063 22876 20127 22880
rect 20063 22820 20067 22876
rect 20067 22820 20123 22876
rect 20123 22820 20127 22876
rect 20063 22816 20127 22820
rect 20143 22876 20207 22880
rect 20143 22820 20147 22876
rect 20147 22820 20203 22876
rect 20203 22820 20207 22876
rect 20143 22816 20207 22820
rect 5690 22332 5754 22336
rect 5690 22276 5694 22332
rect 5694 22276 5750 22332
rect 5750 22276 5754 22332
rect 5690 22272 5754 22276
rect 5770 22332 5834 22336
rect 5770 22276 5774 22332
rect 5774 22276 5830 22332
rect 5830 22276 5834 22332
rect 5770 22272 5834 22276
rect 5850 22332 5914 22336
rect 5850 22276 5854 22332
rect 5854 22276 5910 22332
rect 5910 22276 5914 22332
rect 5850 22272 5914 22276
rect 5930 22332 5994 22336
rect 5930 22276 5934 22332
rect 5934 22276 5990 22332
rect 5990 22276 5994 22332
rect 5930 22272 5994 22276
rect 15165 22332 15229 22336
rect 15165 22276 15169 22332
rect 15169 22276 15225 22332
rect 15225 22276 15229 22332
rect 15165 22272 15229 22276
rect 15245 22332 15309 22336
rect 15245 22276 15249 22332
rect 15249 22276 15305 22332
rect 15305 22276 15309 22332
rect 15245 22272 15309 22276
rect 15325 22332 15389 22336
rect 15325 22276 15329 22332
rect 15329 22276 15385 22332
rect 15385 22276 15389 22332
rect 15325 22272 15389 22276
rect 15405 22332 15469 22336
rect 15405 22276 15409 22332
rect 15409 22276 15465 22332
rect 15465 22276 15469 22332
rect 15405 22272 15469 22276
rect 24641 22332 24705 22336
rect 24641 22276 24645 22332
rect 24645 22276 24701 22332
rect 24701 22276 24705 22332
rect 24641 22272 24705 22276
rect 24721 22332 24785 22336
rect 24721 22276 24725 22332
rect 24725 22276 24781 22332
rect 24781 22276 24785 22332
rect 24721 22272 24785 22276
rect 24801 22332 24865 22336
rect 24801 22276 24805 22332
rect 24805 22276 24861 22332
rect 24861 22276 24865 22332
rect 24801 22272 24865 22276
rect 24881 22332 24945 22336
rect 24881 22276 24885 22332
rect 24885 22276 24941 22332
rect 24941 22276 24945 22332
rect 24881 22272 24945 22276
rect 10427 21788 10491 21792
rect 10427 21732 10431 21788
rect 10431 21732 10487 21788
rect 10487 21732 10491 21788
rect 10427 21728 10491 21732
rect 10507 21788 10571 21792
rect 10507 21732 10511 21788
rect 10511 21732 10567 21788
rect 10567 21732 10571 21788
rect 10507 21728 10571 21732
rect 10587 21788 10651 21792
rect 10587 21732 10591 21788
rect 10591 21732 10647 21788
rect 10647 21732 10651 21788
rect 10587 21728 10651 21732
rect 10667 21788 10731 21792
rect 10667 21732 10671 21788
rect 10671 21732 10727 21788
rect 10727 21732 10731 21788
rect 10667 21728 10731 21732
rect 19903 21788 19967 21792
rect 19903 21732 19907 21788
rect 19907 21732 19963 21788
rect 19963 21732 19967 21788
rect 19903 21728 19967 21732
rect 19983 21788 20047 21792
rect 19983 21732 19987 21788
rect 19987 21732 20043 21788
rect 20043 21732 20047 21788
rect 19983 21728 20047 21732
rect 20063 21788 20127 21792
rect 20063 21732 20067 21788
rect 20067 21732 20123 21788
rect 20123 21732 20127 21788
rect 20063 21728 20127 21732
rect 20143 21788 20207 21792
rect 20143 21732 20147 21788
rect 20147 21732 20203 21788
rect 20203 21732 20207 21788
rect 20143 21728 20207 21732
rect 5690 21244 5754 21248
rect 5690 21188 5694 21244
rect 5694 21188 5750 21244
rect 5750 21188 5754 21244
rect 5690 21184 5754 21188
rect 5770 21244 5834 21248
rect 5770 21188 5774 21244
rect 5774 21188 5830 21244
rect 5830 21188 5834 21244
rect 5770 21184 5834 21188
rect 5850 21244 5914 21248
rect 5850 21188 5854 21244
rect 5854 21188 5910 21244
rect 5910 21188 5914 21244
rect 5850 21184 5914 21188
rect 5930 21244 5994 21248
rect 5930 21188 5934 21244
rect 5934 21188 5990 21244
rect 5990 21188 5994 21244
rect 5930 21184 5994 21188
rect 15165 21244 15229 21248
rect 15165 21188 15169 21244
rect 15169 21188 15225 21244
rect 15225 21188 15229 21244
rect 15165 21184 15229 21188
rect 15245 21244 15309 21248
rect 15245 21188 15249 21244
rect 15249 21188 15305 21244
rect 15305 21188 15309 21244
rect 15245 21184 15309 21188
rect 15325 21244 15389 21248
rect 15325 21188 15329 21244
rect 15329 21188 15385 21244
rect 15385 21188 15389 21244
rect 15325 21184 15389 21188
rect 15405 21244 15469 21248
rect 15405 21188 15409 21244
rect 15409 21188 15465 21244
rect 15465 21188 15469 21244
rect 15405 21184 15469 21188
rect 24641 21244 24705 21248
rect 24641 21188 24645 21244
rect 24645 21188 24701 21244
rect 24701 21188 24705 21244
rect 24641 21184 24705 21188
rect 24721 21244 24785 21248
rect 24721 21188 24725 21244
rect 24725 21188 24781 21244
rect 24781 21188 24785 21244
rect 24721 21184 24785 21188
rect 24801 21244 24865 21248
rect 24801 21188 24805 21244
rect 24805 21188 24861 21244
rect 24861 21188 24865 21244
rect 24801 21184 24865 21188
rect 24881 21244 24945 21248
rect 24881 21188 24885 21244
rect 24885 21188 24941 21244
rect 24941 21188 24945 21244
rect 24881 21184 24945 21188
rect 10427 20700 10491 20704
rect 10427 20644 10431 20700
rect 10431 20644 10487 20700
rect 10487 20644 10491 20700
rect 10427 20640 10491 20644
rect 10507 20700 10571 20704
rect 10507 20644 10511 20700
rect 10511 20644 10567 20700
rect 10567 20644 10571 20700
rect 10507 20640 10571 20644
rect 10587 20700 10651 20704
rect 10587 20644 10591 20700
rect 10591 20644 10647 20700
rect 10647 20644 10651 20700
rect 10587 20640 10651 20644
rect 10667 20700 10731 20704
rect 10667 20644 10671 20700
rect 10671 20644 10727 20700
rect 10727 20644 10731 20700
rect 10667 20640 10731 20644
rect 19903 20700 19967 20704
rect 19903 20644 19907 20700
rect 19907 20644 19963 20700
rect 19963 20644 19967 20700
rect 19903 20640 19967 20644
rect 19983 20700 20047 20704
rect 19983 20644 19987 20700
rect 19987 20644 20043 20700
rect 20043 20644 20047 20700
rect 19983 20640 20047 20644
rect 20063 20700 20127 20704
rect 20063 20644 20067 20700
rect 20067 20644 20123 20700
rect 20123 20644 20127 20700
rect 20063 20640 20127 20644
rect 20143 20700 20207 20704
rect 20143 20644 20147 20700
rect 20147 20644 20203 20700
rect 20203 20644 20207 20700
rect 20143 20640 20207 20644
rect 5690 20156 5754 20160
rect 5690 20100 5694 20156
rect 5694 20100 5750 20156
rect 5750 20100 5754 20156
rect 5690 20096 5754 20100
rect 5770 20156 5834 20160
rect 5770 20100 5774 20156
rect 5774 20100 5830 20156
rect 5830 20100 5834 20156
rect 5770 20096 5834 20100
rect 5850 20156 5914 20160
rect 5850 20100 5854 20156
rect 5854 20100 5910 20156
rect 5910 20100 5914 20156
rect 5850 20096 5914 20100
rect 5930 20156 5994 20160
rect 5930 20100 5934 20156
rect 5934 20100 5990 20156
rect 5990 20100 5994 20156
rect 5930 20096 5994 20100
rect 15165 20156 15229 20160
rect 15165 20100 15169 20156
rect 15169 20100 15225 20156
rect 15225 20100 15229 20156
rect 15165 20096 15229 20100
rect 15245 20156 15309 20160
rect 15245 20100 15249 20156
rect 15249 20100 15305 20156
rect 15305 20100 15309 20156
rect 15245 20096 15309 20100
rect 15325 20156 15389 20160
rect 15325 20100 15329 20156
rect 15329 20100 15385 20156
rect 15385 20100 15389 20156
rect 15325 20096 15389 20100
rect 15405 20156 15469 20160
rect 15405 20100 15409 20156
rect 15409 20100 15465 20156
rect 15465 20100 15469 20156
rect 15405 20096 15469 20100
rect 24641 20156 24705 20160
rect 24641 20100 24645 20156
rect 24645 20100 24701 20156
rect 24701 20100 24705 20156
rect 24641 20096 24705 20100
rect 24721 20156 24785 20160
rect 24721 20100 24725 20156
rect 24725 20100 24781 20156
rect 24781 20100 24785 20156
rect 24721 20096 24785 20100
rect 24801 20156 24865 20160
rect 24801 20100 24805 20156
rect 24805 20100 24861 20156
rect 24861 20100 24865 20156
rect 24801 20096 24865 20100
rect 24881 20156 24945 20160
rect 24881 20100 24885 20156
rect 24885 20100 24941 20156
rect 24941 20100 24945 20156
rect 24881 20096 24945 20100
rect 10427 19612 10491 19616
rect 10427 19556 10431 19612
rect 10431 19556 10487 19612
rect 10487 19556 10491 19612
rect 10427 19552 10491 19556
rect 10507 19612 10571 19616
rect 10507 19556 10511 19612
rect 10511 19556 10567 19612
rect 10567 19556 10571 19612
rect 10507 19552 10571 19556
rect 10587 19612 10651 19616
rect 10587 19556 10591 19612
rect 10591 19556 10647 19612
rect 10647 19556 10651 19612
rect 10587 19552 10651 19556
rect 10667 19612 10731 19616
rect 10667 19556 10671 19612
rect 10671 19556 10727 19612
rect 10727 19556 10731 19612
rect 10667 19552 10731 19556
rect 19903 19612 19967 19616
rect 19903 19556 19907 19612
rect 19907 19556 19963 19612
rect 19963 19556 19967 19612
rect 19903 19552 19967 19556
rect 19983 19612 20047 19616
rect 19983 19556 19987 19612
rect 19987 19556 20043 19612
rect 20043 19556 20047 19612
rect 19983 19552 20047 19556
rect 20063 19612 20127 19616
rect 20063 19556 20067 19612
rect 20067 19556 20123 19612
rect 20123 19556 20127 19612
rect 20063 19552 20127 19556
rect 20143 19612 20207 19616
rect 20143 19556 20147 19612
rect 20147 19556 20203 19612
rect 20203 19556 20207 19612
rect 20143 19552 20207 19556
rect 5690 19068 5754 19072
rect 5690 19012 5694 19068
rect 5694 19012 5750 19068
rect 5750 19012 5754 19068
rect 5690 19008 5754 19012
rect 5770 19068 5834 19072
rect 5770 19012 5774 19068
rect 5774 19012 5830 19068
rect 5830 19012 5834 19068
rect 5770 19008 5834 19012
rect 5850 19068 5914 19072
rect 5850 19012 5854 19068
rect 5854 19012 5910 19068
rect 5910 19012 5914 19068
rect 5850 19008 5914 19012
rect 5930 19068 5994 19072
rect 5930 19012 5934 19068
rect 5934 19012 5990 19068
rect 5990 19012 5994 19068
rect 5930 19008 5994 19012
rect 15165 19068 15229 19072
rect 15165 19012 15169 19068
rect 15169 19012 15225 19068
rect 15225 19012 15229 19068
rect 15165 19008 15229 19012
rect 15245 19068 15309 19072
rect 15245 19012 15249 19068
rect 15249 19012 15305 19068
rect 15305 19012 15309 19068
rect 15245 19008 15309 19012
rect 15325 19068 15389 19072
rect 15325 19012 15329 19068
rect 15329 19012 15385 19068
rect 15385 19012 15389 19068
rect 15325 19008 15389 19012
rect 15405 19068 15469 19072
rect 15405 19012 15409 19068
rect 15409 19012 15465 19068
rect 15465 19012 15469 19068
rect 15405 19008 15469 19012
rect 24641 19068 24705 19072
rect 24641 19012 24645 19068
rect 24645 19012 24701 19068
rect 24701 19012 24705 19068
rect 24641 19008 24705 19012
rect 24721 19068 24785 19072
rect 24721 19012 24725 19068
rect 24725 19012 24781 19068
rect 24781 19012 24785 19068
rect 24721 19008 24785 19012
rect 24801 19068 24865 19072
rect 24801 19012 24805 19068
rect 24805 19012 24861 19068
rect 24861 19012 24865 19068
rect 24801 19008 24865 19012
rect 24881 19068 24945 19072
rect 24881 19012 24885 19068
rect 24885 19012 24941 19068
rect 24941 19012 24945 19068
rect 24881 19008 24945 19012
rect 10427 18524 10491 18528
rect 10427 18468 10431 18524
rect 10431 18468 10487 18524
rect 10487 18468 10491 18524
rect 10427 18464 10491 18468
rect 10507 18524 10571 18528
rect 10507 18468 10511 18524
rect 10511 18468 10567 18524
rect 10567 18468 10571 18524
rect 10507 18464 10571 18468
rect 10587 18524 10651 18528
rect 10587 18468 10591 18524
rect 10591 18468 10647 18524
rect 10647 18468 10651 18524
rect 10587 18464 10651 18468
rect 10667 18524 10731 18528
rect 10667 18468 10671 18524
rect 10671 18468 10727 18524
rect 10727 18468 10731 18524
rect 10667 18464 10731 18468
rect 19903 18524 19967 18528
rect 19903 18468 19907 18524
rect 19907 18468 19963 18524
rect 19963 18468 19967 18524
rect 19903 18464 19967 18468
rect 19983 18524 20047 18528
rect 19983 18468 19987 18524
rect 19987 18468 20043 18524
rect 20043 18468 20047 18524
rect 19983 18464 20047 18468
rect 20063 18524 20127 18528
rect 20063 18468 20067 18524
rect 20067 18468 20123 18524
rect 20123 18468 20127 18524
rect 20063 18464 20127 18468
rect 20143 18524 20207 18528
rect 20143 18468 20147 18524
rect 20147 18468 20203 18524
rect 20203 18468 20207 18524
rect 20143 18464 20207 18468
rect 5690 17980 5754 17984
rect 5690 17924 5694 17980
rect 5694 17924 5750 17980
rect 5750 17924 5754 17980
rect 5690 17920 5754 17924
rect 5770 17980 5834 17984
rect 5770 17924 5774 17980
rect 5774 17924 5830 17980
rect 5830 17924 5834 17980
rect 5770 17920 5834 17924
rect 5850 17980 5914 17984
rect 5850 17924 5854 17980
rect 5854 17924 5910 17980
rect 5910 17924 5914 17980
rect 5850 17920 5914 17924
rect 5930 17980 5994 17984
rect 5930 17924 5934 17980
rect 5934 17924 5990 17980
rect 5990 17924 5994 17980
rect 5930 17920 5994 17924
rect 15165 17980 15229 17984
rect 15165 17924 15169 17980
rect 15169 17924 15225 17980
rect 15225 17924 15229 17980
rect 15165 17920 15229 17924
rect 15245 17980 15309 17984
rect 15245 17924 15249 17980
rect 15249 17924 15305 17980
rect 15305 17924 15309 17980
rect 15245 17920 15309 17924
rect 15325 17980 15389 17984
rect 15325 17924 15329 17980
rect 15329 17924 15385 17980
rect 15385 17924 15389 17980
rect 15325 17920 15389 17924
rect 15405 17980 15469 17984
rect 15405 17924 15409 17980
rect 15409 17924 15465 17980
rect 15465 17924 15469 17980
rect 15405 17920 15469 17924
rect 24641 17980 24705 17984
rect 24641 17924 24645 17980
rect 24645 17924 24701 17980
rect 24701 17924 24705 17980
rect 24641 17920 24705 17924
rect 24721 17980 24785 17984
rect 24721 17924 24725 17980
rect 24725 17924 24781 17980
rect 24781 17924 24785 17980
rect 24721 17920 24785 17924
rect 24801 17980 24865 17984
rect 24801 17924 24805 17980
rect 24805 17924 24861 17980
rect 24861 17924 24865 17980
rect 24801 17920 24865 17924
rect 24881 17980 24945 17984
rect 24881 17924 24885 17980
rect 24885 17924 24941 17980
rect 24941 17924 24945 17980
rect 24881 17920 24945 17924
rect 20484 17852 20548 17916
rect 10427 17436 10491 17440
rect 10427 17380 10431 17436
rect 10431 17380 10487 17436
rect 10487 17380 10491 17436
rect 10427 17376 10491 17380
rect 10507 17436 10571 17440
rect 10507 17380 10511 17436
rect 10511 17380 10567 17436
rect 10567 17380 10571 17436
rect 10507 17376 10571 17380
rect 10587 17436 10651 17440
rect 10587 17380 10591 17436
rect 10591 17380 10647 17436
rect 10647 17380 10651 17436
rect 10587 17376 10651 17380
rect 10667 17436 10731 17440
rect 10667 17380 10671 17436
rect 10671 17380 10727 17436
rect 10727 17380 10731 17436
rect 10667 17376 10731 17380
rect 19903 17436 19967 17440
rect 19903 17380 19907 17436
rect 19907 17380 19963 17436
rect 19963 17380 19967 17436
rect 19903 17376 19967 17380
rect 19983 17436 20047 17440
rect 19983 17380 19987 17436
rect 19987 17380 20043 17436
rect 20043 17380 20047 17436
rect 19983 17376 20047 17380
rect 20063 17436 20127 17440
rect 20063 17380 20067 17436
rect 20067 17380 20123 17436
rect 20123 17380 20127 17436
rect 20063 17376 20127 17380
rect 20143 17436 20207 17440
rect 20143 17380 20147 17436
rect 20147 17380 20203 17436
rect 20203 17380 20207 17436
rect 20143 17376 20207 17380
rect 19748 16900 19812 16964
rect 5690 16892 5754 16896
rect 5690 16836 5694 16892
rect 5694 16836 5750 16892
rect 5750 16836 5754 16892
rect 5690 16832 5754 16836
rect 5770 16892 5834 16896
rect 5770 16836 5774 16892
rect 5774 16836 5830 16892
rect 5830 16836 5834 16892
rect 5770 16832 5834 16836
rect 5850 16892 5914 16896
rect 5850 16836 5854 16892
rect 5854 16836 5910 16892
rect 5910 16836 5914 16892
rect 5850 16832 5914 16836
rect 5930 16892 5994 16896
rect 5930 16836 5934 16892
rect 5934 16836 5990 16892
rect 5990 16836 5994 16892
rect 5930 16832 5994 16836
rect 15165 16892 15229 16896
rect 15165 16836 15169 16892
rect 15169 16836 15225 16892
rect 15225 16836 15229 16892
rect 15165 16832 15229 16836
rect 15245 16892 15309 16896
rect 15245 16836 15249 16892
rect 15249 16836 15305 16892
rect 15305 16836 15309 16892
rect 15245 16832 15309 16836
rect 15325 16892 15389 16896
rect 15325 16836 15329 16892
rect 15329 16836 15385 16892
rect 15385 16836 15389 16892
rect 15325 16832 15389 16836
rect 15405 16892 15469 16896
rect 15405 16836 15409 16892
rect 15409 16836 15465 16892
rect 15465 16836 15469 16892
rect 15405 16832 15469 16836
rect 24641 16892 24705 16896
rect 24641 16836 24645 16892
rect 24645 16836 24701 16892
rect 24701 16836 24705 16892
rect 24641 16832 24705 16836
rect 24721 16892 24785 16896
rect 24721 16836 24725 16892
rect 24725 16836 24781 16892
rect 24781 16836 24785 16892
rect 24721 16832 24785 16836
rect 24801 16892 24865 16896
rect 24801 16836 24805 16892
rect 24805 16836 24861 16892
rect 24861 16836 24865 16892
rect 24801 16832 24865 16836
rect 24881 16892 24945 16896
rect 24881 16836 24885 16892
rect 24885 16836 24941 16892
rect 24941 16836 24945 16892
rect 24881 16832 24945 16836
rect 10427 16348 10491 16352
rect 10427 16292 10431 16348
rect 10431 16292 10487 16348
rect 10487 16292 10491 16348
rect 10427 16288 10491 16292
rect 10507 16348 10571 16352
rect 10507 16292 10511 16348
rect 10511 16292 10567 16348
rect 10567 16292 10571 16348
rect 10507 16288 10571 16292
rect 10587 16348 10651 16352
rect 10587 16292 10591 16348
rect 10591 16292 10647 16348
rect 10647 16292 10651 16348
rect 10587 16288 10651 16292
rect 10667 16348 10731 16352
rect 10667 16292 10671 16348
rect 10671 16292 10727 16348
rect 10727 16292 10731 16348
rect 10667 16288 10731 16292
rect 19903 16348 19967 16352
rect 19903 16292 19907 16348
rect 19907 16292 19963 16348
rect 19963 16292 19967 16348
rect 19903 16288 19967 16292
rect 19983 16348 20047 16352
rect 19983 16292 19987 16348
rect 19987 16292 20043 16348
rect 20043 16292 20047 16348
rect 19983 16288 20047 16292
rect 20063 16348 20127 16352
rect 20063 16292 20067 16348
rect 20067 16292 20123 16348
rect 20123 16292 20127 16348
rect 20063 16288 20127 16292
rect 20143 16348 20207 16352
rect 20143 16292 20147 16348
rect 20147 16292 20203 16348
rect 20203 16292 20207 16348
rect 20143 16288 20207 16292
rect 5690 15804 5754 15808
rect 5690 15748 5694 15804
rect 5694 15748 5750 15804
rect 5750 15748 5754 15804
rect 5690 15744 5754 15748
rect 5770 15804 5834 15808
rect 5770 15748 5774 15804
rect 5774 15748 5830 15804
rect 5830 15748 5834 15804
rect 5770 15744 5834 15748
rect 5850 15804 5914 15808
rect 5850 15748 5854 15804
rect 5854 15748 5910 15804
rect 5910 15748 5914 15804
rect 5850 15744 5914 15748
rect 5930 15804 5994 15808
rect 5930 15748 5934 15804
rect 5934 15748 5990 15804
rect 5990 15748 5994 15804
rect 5930 15744 5994 15748
rect 15165 15804 15229 15808
rect 15165 15748 15169 15804
rect 15169 15748 15225 15804
rect 15225 15748 15229 15804
rect 15165 15744 15229 15748
rect 15245 15804 15309 15808
rect 15245 15748 15249 15804
rect 15249 15748 15305 15804
rect 15305 15748 15309 15804
rect 15245 15744 15309 15748
rect 15325 15804 15389 15808
rect 15325 15748 15329 15804
rect 15329 15748 15385 15804
rect 15385 15748 15389 15804
rect 15325 15744 15389 15748
rect 15405 15804 15469 15808
rect 15405 15748 15409 15804
rect 15409 15748 15465 15804
rect 15465 15748 15469 15804
rect 15405 15744 15469 15748
rect 24641 15804 24705 15808
rect 24641 15748 24645 15804
rect 24645 15748 24701 15804
rect 24701 15748 24705 15804
rect 24641 15744 24705 15748
rect 24721 15804 24785 15808
rect 24721 15748 24725 15804
rect 24725 15748 24781 15804
rect 24781 15748 24785 15804
rect 24721 15744 24785 15748
rect 24801 15804 24865 15808
rect 24801 15748 24805 15804
rect 24805 15748 24861 15804
rect 24861 15748 24865 15804
rect 24801 15744 24865 15748
rect 24881 15804 24945 15808
rect 24881 15748 24885 15804
rect 24885 15748 24941 15804
rect 24941 15748 24945 15804
rect 24881 15744 24945 15748
rect 13676 15404 13740 15468
rect 10427 15260 10491 15264
rect 10427 15204 10431 15260
rect 10431 15204 10487 15260
rect 10487 15204 10491 15260
rect 10427 15200 10491 15204
rect 10507 15260 10571 15264
rect 10507 15204 10511 15260
rect 10511 15204 10567 15260
rect 10567 15204 10571 15260
rect 10507 15200 10571 15204
rect 10587 15260 10651 15264
rect 10587 15204 10591 15260
rect 10591 15204 10647 15260
rect 10647 15204 10651 15260
rect 10587 15200 10651 15204
rect 10667 15260 10731 15264
rect 10667 15204 10671 15260
rect 10671 15204 10727 15260
rect 10727 15204 10731 15260
rect 10667 15200 10731 15204
rect 19903 15260 19967 15264
rect 19903 15204 19907 15260
rect 19907 15204 19963 15260
rect 19963 15204 19967 15260
rect 19903 15200 19967 15204
rect 19983 15260 20047 15264
rect 19983 15204 19987 15260
rect 19987 15204 20043 15260
rect 20043 15204 20047 15260
rect 19983 15200 20047 15204
rect 20063 15260 20127 15264
rect 20063 15204 20067 15260
rect 20067 15204 20123 15260
rect 20123 15204 20127 15260
rect 20063 15200 20127 15204
rect 20143 15260 20207 15264
rect 20143 15204 20147 15260
rect 20147 15204 20203 15260
rect 20203 15204 20207 15260
rect 20143 15200 20207 15204
rect 5690 14716 5754 14720
rect 5690 14660 5694 14716
rect 5694 14660 5750 14716
rect 5750 14660 5754 14716
rect 5690 14656 5754 14660
rect 5770 14716 5834 14720
rect 5770 14660 5774 14716
rect 5774 14660 5830 14716
rect 5830 14660 5834 14716
rect 5770 14656 5834 14660
rect 5850 14716 5914 14720
rect 5850 14660 5854 14716
rect 5854 14660 5910 14716
rect 5910 14660 5914 14716
rect 5850 14656 5914 14660
rect 5930 14716 5994 14720
rect 5930 14660 5934 14716
rect 5934 14660 5990 14716
rect 5990 14660 5994 14716
rect 5930 14656 5994 14660
rect 15165 14716 15229 14720
rect 15165 14660 15169 14716
rect 15169 14660 15225 14716
rect 15225 14660 15229 14716
rect 15165 14656 15229 14660
rect 15245 14716 15309 14720
rect 15245 14660 15249 14716
rect 15249 14660 15305 14716
rect 15305 14660 15309 14716
rect 15245 14656 15309 14660
rect 15325 14716 15389 14720
rect 15325 14660 15329 14716
rect 15329 14660 15385 14716
rect 15385 14660 15389 14716
rect 15325 14656 15389 14660
rect 15405 14716 15469 14720
rect 15405 14660 15409 14716
rect 15409 14660 15465 14716
rect 15465 14660 15469 14716
rect 15405 14656 15469 14660
rect 24641 14716 24705 14720
rect 24641 14660 24645 14716
rect 24645 14660 24701 14716
rect 24701 14660 24705 14716
rect 24641 14656 24705 14660
rect 24721 14716 24785 14720
rect 24721 14660 24725 14716
rect 24725 14660 24781 14716
rect 24781 14660 24785 14716
rect 24721 14656 24785 14660
rect 24801 14716 24865 14720
rect 24801 14660 24805 14716
rect 24805 14660 24861 14716
rect 24861 14660 24865 14716
rect 24801 14656 24865 14660
rect 24881 14716 24945 14720
rect 24881 14660 24885 14716
rect 24885 14660 24941 14716
rect 24941 14660 24945 14716
rect 24881 14656 24945 14660
rect 10427 14172 10491 14176
rect 10427 14116 10431 14172
rect 10431 14116 10487 14172
rect 10487 14116 10491 14172
rect 10427 14112 10491 14116
rect 10507 14172 10571 14176
rect 10507 14116 10511 14172
rect 10511 14116 10567 14172
rect 10567 14116 10571 14172
rect 10507 14112 10571 14116
rect 10587 14172 10651 14176
rect 10587 14116 10591 14172
rect 10591 14116 10647 14172
rect 10647 14116 10651 14172
rect 10587 14112 10651 14116
rect 10667 14172 10731 14176
rect 10667 14116 10671 14172
rect 10671 14116 10727 14172
rect 10727 14116 10731 14172
rect 10667 14112 10731 14116
rect 19903 14172 19967 14176
rect 19903 14116 19907 14172
rect 19907 14116 19963 14172
rect 19963 14116 19967 14172
rect 19903 14112 19967 14116
rect 19983 14172 20047 14176
rect 19983 14116 19987 14172
rect 19987 14116 20043 14172
rect 20043 14116 20047 14172
rect 19983 14112 20047 14116
rect 20063 14172 20127 14176
rect 20063 14116 20067 14172
rect 20067 14116 20123 14172
rect 20123 14116 20127 14172
rect 20063 14112 20127 14116
rect 20143 14172 20207 14176
rect 20143 14116 20147 14172
rect 20147 14116 20203 14172
rect 20203 14116 20207 14172
rect 20143 14112 20207 14116
rect 5690 13628 5754 13632
rect 5690 13572 5694 13628
rect 5694 13572 5750 13628
rect 5750 13572 5754 13628
rect 5690 13568 5754 13572
rect 5770 13628 5834 13632
rect 5770 13572 5774 13628
rect 5774 13572 5830 13628
rect 5830 13572 5834 13628
rect 5770 13568 5834 13572
rect 5850 13628 5914 13632
rect 5850 13572 5854 13628
rect 5854 13572 5910 13628
rect 5910 13572 5914 13628
rect 5850 13568 5914 13572
rect 5930 13628 5994 13632
rect 5930 13572 5934 13628
rect 5934 13572 5990 13628
rect 5990 13572 5994 13628
rect 5930 13568 5994 13572
rect 15165 13628 15229 13632
rect 15165 13572 15169 13628
rect 15169 13572 15225 13628
rect 15225 13572 15229 13628
rect 15165 13568 15229 13572
rect 15245 13628 15309 13632
rect 15245 13572 15249 13628
rect 15249 13572 15305 13628
rect 15305 13572 15309 13628
rect 15245 13568 15309 13572
rect 15325 13628 15389 13632
rect 15325 13572 15329 13628
rect 15329 13572 15385 13628
rect 15385 13572 15389 13628
rect 15325 13568 15389 13572
rect 15405 13628 15469 13632
rect 15405 13572 15409 13628
rect 15409 13572 15465 13628
rect 15465 13572 15469 13628
rect 15405 13568 15469 13572
rect 24641 13628 24705 13632
rect 24641 13572 24645 13628
rect 24645 13572 24701 13628
rect 24701 13572 24705 13628
rect 24641 13568 24705 13572
rect 24721 13628 24785 13632
rect 24721 13572 24725 13628
rect 24725 13572 24781 13628
rect 24781 13572 24785 13628
rect 24721 13568 24785 13572
rect 24801 13628 24865 13632
rect 24801 13572 24805 13628
rect 24805 13572 24861 13628
rect 24861 13572 24865 13628
rect 24801 13568 24865 13572
rect 24881 13628 24945 13632
rect 24881 13572 24885 13628
rect 24885 13572 24941 13628
rect 24941 13572 24945 13628
rect 24881 13568 24945 13572
rect 10427 13084 10491 13088
rect 10427 13028 10431 13084
rect 10431 13028 10487 13084
rect 10487 13028 10491 13084
rect 10427 13024 10491 13028
rect 10507 13084 10571 13088
rect 10507 13028 10511 13084
rect 10511 13028 10567 13084
rect 10567 13028 10571 13084
rect 10507 13024 10571 13028
rect 10587 13084 10651 13088
rect 10587 13028 10591 13084
rect 10591 13028 10647 13084
rect 10647 13028 10651 13084
rect 10587 13024 10651 13028
rect 10667 13084 10731 13088
rect 10667 13028 10671 13084
rect 10671 13028 10727 13084
rect 10727 13028 10731 13084
rect 10667 13024 10731 13028
rect 19903 13084 19967 13088
rect 19903 13028 19907 13084
rect 19907 13028 19963 13084
rect 19963 13028 19967 13084
rect 19903 13024 19967 13028
rect 19983 13084 20047 13088
rect 19983 13028 19987 13084
rect 19987 13028 20043 13084
rect 20043 13028 20047 13084
rect 19983 13024 20047 13028
rect 20063 13084 20127 13088
rect 20063 13028 20067 13084
rect 20067 13028 20123 13084
rect 20123 13028 20127 13084
rect 20063 13024 20127 13028
rect 20143 13084 20207 13088
rect 20143 13028 20147 13084
rect 20147 13028 20203 13084
rect 20203 13028 20207 13084
rect 20143 13024 20207 13028
rect 5690 12540 5754 12544
rect 5690 12484 5694 12540
rect 5694 12484 5750 12540
rect 5750 12484 5754 12540
rect 5690 12480 5754 12484
rect 5770 12540 5834 12544
rect 5770 12484 5774 12540
rect 5774 12484 5830 12540
rect 5830 12484 5834 12540
rect 5770 12480 5834 12484
rect 5850 12540 5914 12544
rect 5850 12484 5854 12540
rect 5854 12484 5910 12540
rect 5910 12484 5914 12540
rect 5850 12480 5914 12484
rect 5930 12540 5994 12544
rect 5930 12484 5934 12540
rect 5934 12484 5990 12540
rect 5990 12484 5994 12540
rect 5930 12480 5994 12484
rect 15165 12540 15229 12544
rect 15165 12484 15169 12540
rect 15169 12484 15225 12540
rect 15225 12484 15229 12540
rect 15165 12480 15229 12484
rect 15245 12540 15309 12544
rect 15245 12484 15249 12540
rect 15249 12484 15305 12540
rect 15305 12484 15309 12540
rect 15245 12480 15309 12484
rect 15325 12540 15389 12544
rect 15325 12484 15329 12540
rect 15329 12484 15385 12540
rect 15385 12484 15389 12540
rect 15325 12480 15389 12484
rect 15405 12540 15469 12544
rect 15405 12484 15409 12540
rect 15409 12484 15465 12540
rect 15465 12484 15469 12540
rect 15405 12480 15469 12484
rect 24641 12540 24705 12544
rect 24641 12484 24645 12540
rect 24645 12484 24701 12540
rect 24701 12484 24705 12540
rect 24641 12480 24705 12484
rect 24721 12540 24785 12544
rect 24721 12484 24725 12540
rect 24725 12484 24781 12540
rect 24781 12484 24785 12540
rect 24721 12480 24785 12484
rect 24801 12540 24865 12544
rect 24801 12484 24805 12540
rect 24805 12484 24861 12540
rect 24861 12484 24865 12540
rect 24801 12480 24865 12484
rect 24881 12540 24945 12544
rect 24881 12484 24885 12540
rect 24885 12484 24941 12540
rect 24941 12484 24945 12540
rect 24881 12480 24945 12484
rect 10427 11996 10491 12000
rect 10427 11940 10431 11996
rect 10431 11940 10487 11996
rect 10487 11940 10491 11996
rect 10427 11936 10491 11940
rect 10507 11996 10571 12000
rect 10507 11940 10511 11996
rect 10511 11940 10567 11996
rect 10567 11940 10571 11996
rect 10507 11936 10571 11940
rect 10587 11996 10651 12000
rect 10587 11940 10591 11996
rect 10591 11940 10647 11996
rect 10647 11940 10651 11996
rect 10587 11936 10651 11940
rect 10667 11996 10731 12000
rect 10667 11940 10671 11996
rect 10671 11940 10727 11996
rect 10727 11940 10731 11996
rect 10667 11936 10731 11940
rect 19903 11996 19967 12000
rect 19903 11940 19907 11996
rect 19907 11940 19963 11996
rect 19963 11940 19967 11996
rect 19903 11936 19967 11940
rect 19983 11996 20047 12000
rect 19983 11940 19987 11996
rect 19987 11940 20043 11996
rect 20043 11940 20047 11996
rect 19983 11936 20047 11940
rect 20063 11996 20127 12000
rect 20063 11940 20067 11996
rect 20067 11940 20123 11996
rect 20123 11940 20127 11996
rect 20063 11936 20127 11940
rect 20143 11996 20207 12000
rect 20143 11940 20147 11996
rect 20147 11940 20203 11996
rect 20203 11940 20207 11996
rect 20143 11936 20207 11940
rect 5690 11452 5754 11456
rect 5690 11396 5694 11452
rect 5694 11396 5750 11452
rect 5750 11396 5754 11452
rect 5690 11392 5754 11396
rect 5770 11452 5834 11456
rect 5770 11396 5774 11452
rect 5774 11396 5830 11452
rect 5830 11396 5834 11452
rect 5770 11392 5834 11396
rect 5850 11452 5914 11456
rect 5850 11396 5854 11452
rect 5854 11396 5910 11452
rect 5910 11396 5914 11452
rect 5850 11392 5914 11396
rect 5930 11452 5994 11456
rect 5930 11396 5934 11452
rect 5934 11396 5990 11452
rect 5990 11396 5994 11452
rect 5930 11392 5994 11396
rect 15165 11452 15229 11456
rect 15165 11396 15169 11452
rect 15169 11396 15225 11452
rect 15225 11396 15229 11452
rect 15165 11392 15229 11396
rect 15245 11452 15309 11456
rect 15245 11396 15249 11452
rect 15249 11396 15305 11452
rect 15305 11396 15309 11452
rect 15245 11392 15309 11396
rect 15325 11452 15389 11456
rect 15325 11396 15329 11452
rect 15329 11396 15385 11452
rect 15385 11396 15389 11452
rect 15325 11392 15389 11396
rect 15405 11452 15469 11456
rect 15405 11396 15409 11452
rect 15409 11396 15465 11452
rect 15465 11396 15469 11452
rect 15405 11392 15469 11396
rect 24641 11452 24705 11456
rect 24641 11396 24645 11452
rect 24645 11396 24701 11452
rect 24701 11396 24705 11452
rect 24641 11392 24705 11396
rect 24721 11452 24785 11456
rect 24721 11396 24725 11452
rect 24725 11396 24781 11452
rect 24781 11396 24785 11452
rect 24721 11392 24785 11396
rect 24801 11452 24865 11456
rect 24801 11396 24805 11452
rect 24805 11396 24861 11452
rect 24861 11396 24865 11452
rect 24801 11392 24865 11396
rect 24881 11452 24945 11456
rect 24881 11396 24885 11452
rect 24885 11396 24941 11452
rect 24941 11396 24945 11452
rect 24881 11392 24945 11396
rect 10916 11052 10980 11116
rect 10427 10908 10491 10912
rect 10427 10852 10431 10908
rect 10431 10852 10487 10908
rect 10487 10852 10491 10908
rect 10427 10848 10491 10852
rect 10507 10908 10571 10912
rect 10507 10852 10511 10908
rect 10511 10852 10567 10908
rect 10567 10852 10571 10908
rect 10507 10848 10571 10852
rect 10587 10908 10651 10912
rect 10587 10852 10591 10908
rect 10591 10852 10647 10908
rect 10647 10852 10651 10908
rect 10587 10848 10651 10852
rect 10667 10908 10731 10912
rect 10667 10852 10671 10908
rect 10671 10852 10727 10908
rect 10727 10852 10731 10908
rect 10667 10848 10731 10852
rect 19903 10908 19967 10912
rect 19903 10852 19907 10908
rect 19907 10852 19963 10908
rect 19963 10852 19967 10908
rect 19903 10848 19967 10852
rect 19983 10908 20047 10912
rect 19983 10852 19987 10908
rect 19987 10852 20043 10908
rect 20043 10852 20047 10908
rect 19983 10848 20047 10852
rect 20063 10908 20127 10912
rect 20063 10852 20067 10908
rect 20067 10852 20123 10908
rect 20123 10852 20127 10908
rect 20063 10848 20127 10852
rect 20143 10908 20207 10912
rect 20143 10852 20147 10908
rect 20147 10852 20203 10908
rect 20203 10852 20207 10908
rect 20143 10848 20207 10852
rect 10916 10568 10980 10572
rect 10916 10512 10930 10568
rect 10930 10512 10980 10568
rect 10916 10508 10980 10512
rect 5690 10364 5754 10368
rect 5690 10308 5694 10364
rect 5694 10308 5750 10364
rect 5750 10308 5754 10364
rect 5690 10304 5754 10308
rect 5770 10364 5834 10368
rect 5770 10308 5774 10364
rect 5774 10308 5830 10364
rect 5830 10308 5834 10364
rect 5770 10304 5834 10308
rect 5850 10364 5914 10368
rect 5850 10308 5854 10364
rect 5854 10308 5910 10364
rect 5910 10308 5914 10364
rect 5850 10304 5914 10308
rect 5930 10364 5994 10368
rect 5930 10308 5934 10364
rect 5934 10308 5990 10364
rect 5990 10308 5994 10364
rect 5930 10304 5994 10308
rect 15165 10364 15229 10368
rect 15165 10308 15169 10364
rect 15169 10308 15225 10364
rect 15225 10308 15229 10364
rect 15165 10304 15229 10308
rect 15245 10364 15309 10368
rect 15245 10308 15249 10364
rect 15249 10308 15305 10364
rect 15305 10308 15309 10364
rect 15245 10304 15309 10308
rect 15325 10364 15389 10368
rect 15325 10308 15329 10364
rect 15329 10308 15385 10364
rect 15385 10308 15389 10364
rect 15325 10304 15389 10308
rect 15405 10364 15469 10368
rect 15405 10308 15409 10364
rect 15409 10308 15465 10364
rect 15465 10308 15469 10364
rect 15405 10304 15469 10308
rect 24641 10364 24705 10368
rect 24641 10308 24645 10364
rect 24645 10308 24701 10364
rect 24701 10308 24705 10364
rect 24641 10304 24705 10308
rect 24721 10364 24785 10368
rect 24721 10308 24725 10364
rect 24725 10308 24781 10364
rect 24781 10308 24785 10364
rect 24721 10304 24785 10308
rect 24801 10364 24865 10368
rect 24801 10308 24805 10364
rect 24805 10308 24861 10364
rect 24861 10308 24865 10364
rect 24801 10304 24865 10308
rect 24881 10364 24945 10368
rect 24881 10308 24885 10364
rect 24885 10308 24941 10364
rect 24941 10308 24945 10364
rect 24881 10304 24945 10308
rect 10427 9820 10491 9824
rect 10427 9764 10431 9820
rect 10431 9764 10487 9820
rect 10487 9764 10491 9820
rect 10427 9760 10491 9764
rect 10507 9820 10571 9824
rect 10507 9764 10511 9820
rect 10511 9764 10567 9820
rect 10567 9764 10571 9820
rect 10507 9760 10571 9764
rect 10587 9820 10651 9824
rect 10587 9764 10591 9820
rect 10591 9764 10647 9820
rect 10647 9764 10651 9820
rect 10587 9760 10651 9764
rect 10667 9820 10731 9824
rect 10667 9764 10671 9820
rect 10671 9764 10727 9820
rect 10727 9764 10731 9820
rect 10667 9760 10731 9764
rect 19903 9820 19967 9824
rect 19903 9764 19907 9820
rect 19907 9764 19963 9820
rect 19963 9764 19967 9820
rect 19903 9760 19967 9764
rect 19983 9820 20047 9824
rect 19983 9764 19987 9820
rect 19987 9764 20043 9820
rect 20043 9764 20047 9820
rect 19983 9760 20047 9764
rect 20063 9820 20127 9824
rect 20063 9764 20067 9820
rect 20067 9764 20123 9820
rect 20123 9764 20127 9820
rect 20063 9760 20127 9764
rect 20143 9820 20207 9824
rect 20143 9764 20147 9820
rect 20147 9764 20203 9820
rect 20203 9764 20207 9820
rect 20143 9760 20207 9764
rect 5690 9276 5754 9280
rect 5690 9220 5694 9276
rect 5694 9220 5750 9276
rect 5750 9220 5754 9276
rect 5690 9216 5754 9220
rect 5770 9276 5834 9280
rect 5770 9220 5774 9276
rect 5774 9220 5830 9276
rect 5830 9220 5834 9276
rect 5770 9216 5834 9220
rect 5850 9276 5914 9280
rect 5850 9220 5854 9276
rect 5854 9220 5910 9276
rect 5910 9220 5914 9276
rect 5850 9216 5914 9220
rect 5930 9276 5994 9280
rect 5930 9220 5934 9276
rect 5934 9220 5990 9276
rect 5990 9220 5994 9276
rect 5930 9216 5994 9220
rect 15165 9276 15229 9280
rect 15165 9220 15169 9276
rect 15169 9220 15225 9276
rect 15225 9220 15229 9276
rect 15165 9216 15229 9220
rect 15245 9276 15309 9280
rect 15245 9220 15249 9276
rect 15249 9220 15305 9276
rect 15305 9220 15309 9276
rect 15245 9216 15309 9220
rect 15325 9276 15389 9280
rect 15325 9220 15329 9276
rect 15329 9220 15385 9276
rect 15385 9220 15389 9276
rect 15325 9216 15389 9220
rect 15405 9276 15469 9280
rect 15405 9220 15409 9276
rect 15409 9220 15465 9276
rect 15465 9220 15469 9276
rect 15405 9216 15469 9220
rect 24641 9276 24705 9280
rect 24641 9220 24645 9276
rect 24645 9220 24701 9276
rect 24701 9220 24705 9276
rect 24641 9216 24705 9220
rect 24721 9276 24785 9280
rect 24721 9220 24725 9276
rect 24725 9220 24781 9276
rect 24781 9220 24785 9276
rect 24721 9216 24785 9220
rect 24801 9276 24865 9280
rect 24801 9220 24805 9276
rect 24805 9220 24861 9276
rect 24861 9220 24865 9276
rect 24801 9216 24865 9220
rect 24881 9276 24945 9280
rect 24881 9220 24885 9276
rect 24885 9220 24941 9276
rect 24941 9220 24945 9276
rect 24881 9216 24945 9220
rect 10427 8732 10491 8736
rect 10427 8676 10431 8732
rect 10431 8676 10487 8732
rect 10487 8676 10491 8732
rect 10427 8672 10491 8676
rect 10507 8732 10571 8736
rect 10507 8676 10511 8732
rect 10511 8676 10567 8732
rect 10567 8676 10571 8732
rect 10507 8672 10571 8676
rect 10587 8732 10651 8736
rect 10587 8676 10591 8732
rect 10591 8676 10647 8732
rect 10647 8676 10651 8732
rect 10587 8672 10651 8676
rect 10667 8732 10731 8736
rect 10667 8676 10671 8732
rect 10671 8676 10727 8732
rect 10727 8676 10731 8732
rect 10667 8672 10731 8676
rect 19903 8732 19967 8736
rect 19903 8676 19907 8732
rect 19907 8676 19963 8732
rect 19963 8676 19967 8732
rect 19903 8672 19967 8676
rect 19983 8732 20047 8736
rect 19983 8676 19987 8732
rect 19987 8676 20043 8732
rect 20043 8676 20047 8732
rect 19983 8672 20047 8676
rect 20063 8732 20127 8736
rect 20063 8676 20067 8732
rect 20067 8676 20123 8732
rect 20123 8676 20127 8732
rect 20063 8672 20127 8676
rect 20143 8732 20207 8736
rect 20143 8676 20147 8732
rect 20147 8676 20203 8732
rect 20203 8676 20207 8732
rect 20143 8672 20207 8676
rect 5690 8188 5754 8192
rect 5690 8132 5694 8188
rect 5694 8132 5750 8188
rect 5750 8132 5754 8188
rect 5690 8128 5754 8132
rect 5770 8188 5834 8192
rect 5770 8132 5774 8188
rect 5774 8132 5830 8188
rect 5830 8132 5834 8188
rect 5770 8128 5834 8132
rect 5850 8188 5914 8192
rect 5850 8132 5854 8188
rect 5854 8132 5910 8188
rect 5910 8132 5914 8188
rect 5850 8128 5914 8132
rect 5930 8188 5994 8192
rect 5930 8132 5934 8188
rect 5934 8132 5990 8188
rect 5990 8132 5994 8188
rect 5930 8128 5994 8132
rect 15165 8188 15229 8192
rect 15165 8132 15169 8188
rect 15169 8132 15225 8188
rect 15225 8132 15229 8188
rect 15165 8128 15229 8132
rect 15245 8188 15309 8192
rect 15245 8132 15249 8188
rect 15249 8132 15305 8188
rect 15305 8132 15309 8188
rect 15245 8128 15309 8132
rect 15325 8188 15389 8192
rect 15325 8132 15329 8188
rect 15329 8132 15385 8188
rect 15385 8132 15389 8188
rect 15325 8128 15389 8132
rect 15405 8188 15469 8192
rect 15405 8132 15409 8188
rect 15409 8132 15465 8188
rect 15465 8132 15469 8188
rect 15405 8128 15469 8132
rect 24641 8188 24705 8192
rect 24641 8132 24645 8188
rect 24645 8132 24701 8188
rect 24701 8132 24705 8188
rect 24641 8128 24705 8132
rect 24721 8188 24785 8192
rect 24721 8132 24725 8188
rect 24725 8132 24781 8188
rect 24781 8132 24785 8188
rect 24721 8128 24785 8132
rect 24801 8188 24865 8192
rect 24801 8132 24805 8188
rect 24805 8132 24861 8188
rect 24861 8132 24865 8188
rect 24801 8128 24865 8132
rect 24881 8188 24945 8192
rect 24881 8132 24885 8188
rect 24885 8132 24941 8188
rect 24941 8132 24945 8188
rect 24881 8128 24945 8132
rect 10427 7644 10491 7648
rect 10427 7588 10431 7644
rect 10431 7588 10487 7644
rect 10487 7588 10491 7644
rect 10427 7584 10491 7588
rect 10507 7644 10571 7648
rect 10507 7588 10511 7644
rect 10511 7588 10567 7644
rect 10567 7588 10571 7644
rect 10507 7584 10571 7588
rect 10587 7644 10651 7648
rect 10587 7588 10591 7644
rect 10591 7588 10647 7644
rect 10647 7588 10651 7644
rect 10587 7584 10651 7588
rect 10667 7644 10731 7648
rect 10667 7588 10671 7644
rect 10671 7588 10727 7644
rect 10727 7588 10731 7644
rect 10667 7584 10731 7588
rect 19903 7644 19967 7648
rect 19903 7588 19907 7644
rect 19907 7588 19963 7644
rect 19963 7588 19967 7644
rect 19903 7584 19967 7588
rect 19983 7644 20047 7648
rect 19983 7588 19987 7644
rect 19987 7588 20043 7644
rect 20043 7588 20047 7644
rect 19983 7584 20047 7588
rect 20063 7644 20127 7648
rect 20063 7588 20067 7644
rect 20067 7588 20123 7644
rect 20123 7588 20127 7644
rect 20063 7584 20127 7588
rect 20143 7644 20207 7648
rect 20143 7588 20147 7644
rect 20147 7588 20203 7644
rect 20203 7588 20207 7644
rect 20143 7584 20207 7588
rect 5690 7100 5754 7104
rect 5690 7044 5694 7100
rect 5694 7044 5750 7100
rect 5750 7044 5754 7100
rect 5690 7040 5754 7044
rect 5770 7100 5834 7104
rect 5770 7044 5774 7100
rect 5774 7044 5830 7100
rect 5830 7044 5834 7100
rect 5770 7040 5834 7044
rect 5850 7100 5914 7104
rect 5850 7044 5854 7100
rect 5854 7044 5910 7100
rect 5910 7044 5914 7100
rect 5850 7040 5914 7044
rect 5930 7100 5994 7104
rect 5930 7044 5934 7100
rect 5934 7044 5990 7100
rect 5990 7044 5994 7100
rect 5930 7040 5994 7044
rect 15165 7100 15229 7104
rect 15165 7044 15169 7100
rect 15169 7044 15225 7100
rect 15225 7044 15229 7100
rect 15165 7040 15229 7044
rect 15245 7100 15309 7104
rect 15245 7044 15249 7100
rect 15249 7044 15305 7100
rect 15305 7044 15309 7100
rect 15245 7040 15309 7044
rect 15325 7100 15389 7104
rect 15325 7044 15329 7100
rect 15329 7044 15385 7100
rect 15385 7044 15389 7100
rect 15325 7040 15389 7044
rect 15405 7100 15469 7104
rect 15405 7044 15409 7100
rect 15409 7044 15465 7100
rect 15465 7044 15469 7100
rect 15405 7040 15469 7044
rect 24641 7100 24705 7104
rect 24641 7044 24645 7100
rect 24645 7044 24701 7100
rect 24701 7044 24705 7100
rect 24641 7040 24705 7044
rect 24721 7100 24785 7104
rect 24721 7044 24725 7100
rect 24725 7044 24781 7100
rect 24781 7044 24785 7100
rect 24721 7040 24785 7044
rect 24801 7100 24865 7104
rect 24801 7044 24805 7100
rect 24805 7044 24861 7100
rect 24861 7044 24865 7100
rect 24801 7040 24865 7044
rect 24881 7100 24945 7104
rect 24881 7044 24885 7100
rect 24885 7044 24941 7100
rect 24941 7044 24945 7100
rect 24881 7040 24945 7044
rect 10427 6556 10491 6560
rect 10427 6500 10431 6556
rect 10431 6500 10487 6556
rect 10487 6500 10491 6556
rect 10427 6496 10491 6500
rect 10507 6556 10571 6560
rect 10507 6500 10511 6556
rect 10511 6500 10567 6556
rect 10567 6500 10571 6556
rect 10507 6496 10571 6500
rect 10587 6556 10651 6560
rect 10587 6500 10591 6556
rect 10591 6500 10647 6556
rect 10647 6500 10651 6556
rect 10587 6496 10651 6500
rect 10667 6556 10731 6560
rect 10667 6500 10671 6556
rect 10671 6500 10727 6556
rect 10727 6500 10731 6556
rect 10667 6496 10731 6500
rect 19903 6556 19967 6560
rect 19903 6500 19907 6556
rect 19907 6500 19963 6556
rect 19963 6500 19967 6556
rect 19903 6496 19967 6500
rect 19983 6556 20047 6560
rect 19983 6500 19987 6556
rect 19987 6500 20043 6556
rect 20043 6500 20047 6556
rect 19983 6496 20047 6500
rect 20063 6556 20127 6560
rect 20063 6500 20067 6556
rect 20067 6500 20123 6556
rect 20123 6500 20127 6556
rect 20063 6496 20127 6500
rect 20143 6556 20207 6560
rect 20143 6500 20147 6556
rect 20147 6500 20203 6556
rect 20203 6500 20207 6556
rect 20143 6496 20207 6500
rect 5690 6012 5754 6016
rect 5690 5956 5694 6012
rect 5694 5956 5750 6012
rect 5750 5956 5754 6012
rect 5690 5952 5754 5956
rect 5770 6012 5834 6016
rect 5770 5956 5774 6012
rect 5774 5956 5830 6012
rect 5830 5956 5834 6012
rect 5770 5952 5834 5956
rect 5850 6012 5914 6016
rect 5850 5956 5854 6012
rect 5854 5956 5910 6012
rect 5910 5956 5914 6012
rect 5850 5952 5914 5956
rect 5930 6012 5994 6016
rect 5930 5956 5934 6012
rect 5934 5956 5990 6012
rect 5990 5956 5994 6012
rect 5930 5952 5994 5956
rect 15165 6012 15229 6016
rect 15165 5956 15169 6012
rect 15169 5956 15225 6012
rect 15225 5956 15229 6012
rect 15165 5952 15229 5956
rect 15245 6012 15309 6016
rect 15245 5956 15249 6012
rect 15249 5956 15305 6012
rect 15305 5956 15309 6012
rect 15245 5952 15309 5956
rect 15325 6012 15389 6016
rect 15325 5956 15329 6012
rect 15329 5956 15385 6012
rect 15385 5956 15389 6012
rect 15325 5952 15389 5956
rect 15405 6012 15469 6016
rect 15405 5956 15409 6012
rect 15409 5956 15465 6012
rect 15465 5956 15469 6012
rect 15405 5952 15469 5956
rect 24641 6012 24705 6016
rect 24641 5956 24645 6012
rect 24645 5956 24701 6012
rect 24701 5956 24705 6012
rect 24641 5952 24705 5956
rect 24721 6012 24785 6016
rect 24721 5956 24725 6012
rect 24725 5956 24781 6012
rect 24781 5956 24785 6012
rect 24721 5952 24785 5956
rect 24801 6012 24865 6016
rect 24801 5956 24805 6012
rect 24805 5956 24861 6012
rect 24861 5956 24865 6012
rect 24801 5952 24865 5956
rect 24881 6012 24945 6016
rect 24881 5956 24885 6012
rect 24885 5956 24941 6012
rect 24941 5956 24945 6012
rect 24881 5952 24945 5956
rect 10427 5468 10491 5472
rect 10427 5412 10431 5468
rect 10431 5412 10487 5468
rect 10487 5412 10491 5468
rect 10427 5408 10491 5412
rect 10507 5468 10571 5472
rect 10507 5412 10511 5468
rect 10511 5412 10567 5468
rect 10567 5412 10571 5468
rect 10507 5408 10571 5412
rect 10587 5468 10651 5472
rect 10587 5412 10591 5468
rect 10591 5412 10647 5468
rect 10647 5412 10651 5468
rect 10587 5408 10651 5412
rect 10667 5468 10731 5472
rect 10667 5412 10671 5468
rect 10671 5412 10727 5468
rect 10727 5412 10731 5468
rect 10667 5408 10731 5412
rect 19903 5468 19967 5472
rect 19903 5412 19907 5468
rect 19907 5412 19963 5468
rect 19963 5412 19967 5468
rect 19903 5408 19967 5412
rect 19983 5468 20047 5472
rect 19983 5412 19987 5468
rect 19987 5412 20043 5468
rect 20043 5412 20047 5468
rect 19983 5408 20047 5412
rect 20063 5468 20127 5472
rect 20063 5412 20067 5468
rect 20067 5412 20123 5468
rect 20123 5412 20127 5468
rect 20063 5408 20127 5412
rect 20143 5468 20207 5472
rect 20143 5412 20147 5468
rect 20147 5412 20203 5468
rect 20203 5412 20207 5468
rect 20143 5408 20207 5412
rect 5690 4924 5754 4928
rect 5690 4868 5694 4924
rect 5694 4868 5750 4924
rect 5750 4868 5754 4924
rect 5690 4864 5754 4868
rect 5770 4924 5834 4928
rect 5770 4868 5774 4924
rect 5774 4868 5830 4924
rect 5830 4868 5834 4924
rect 5770 4864 5834 4868
rect 5850 4924 5914 4928
rect 5850 4868 5854 4924
rect 5854 4868 5910 4924
rect 5910 4868 5914 4924
rect 5850 4864 5914 4868
rect 5930 4924 5994 4928
rect 5930 4868 5934 4924
rect 5934 4868 5990 4924
rect 5990 4868 5994 4924
rect 5930 4864 5994 4868
rect 15165 4924 15229 4928
rect 15165 4868 15169 4924
rect 15169 4868 15225 4924
rect 15225 4868 15229 4924
rect 15165 4864 15229 4868
rect 15245 4924 15309 4928
rect 15245 4868 15249 4924
rect 15249 4868 15305 4924
rect 15305 4868 15309 4924
rect 15245 4864 15309 4868
rect 15325 4924 15389 4928
rect 15325 4868 15329 4924
rect 15329 4868 15385 4924
rect 15385 4868 15389 4924
rect 15325 4864 15389 4868
rect 15405 4924 15469 4928
rect 15405 4868 15409 4924
rect 15409 4868 15465 4924
rect 15465 4868 15469 4924
rect 15405 4864 15469 4868
rect 24641 4924 24705 4928
rect 24641 4868 24645 4924
rect 24645 4868 24701 4924
rect 24701 4868 24705 4924
rect 24641 4864 24705 4868
rect 24721 4924 24785 4928
rect 24721 4868 24725 4924
rect 24725 4868 24781 4924
rect 24781 4868 24785 4924
rect 24721 4864 24785 4868
rect 24801 4924 24865 4928
rect 24801 4868 24805 4924
rect 24805 4868 24861 4924
rect 24861 4868 24865 4924
rect 24801 4864 24865 4868
rect 24881 4924 24945 4928
rect 24881 4868 24885 4924
rect 24885 4868 24941 4924
rect 24941 4868 24945 4924
rect 24881 4864 24945 4868
rect 10427 4380 10491 4384
rect 10427 4324 10431 4380
rect 10431 4324 10487 4380
rect 10487 4324 10491 4380
rect 10427 4320 10491 4324
rect 10507 4380 10571 4384
rect 10507 4324 10511 4380
rect 10511 4324 10567 4380
rect 10567 4324 10571 4380
rect 10507 4320 10571 4324
rect 10587 4380 10651 4384
rect 10587 4324 10591 4380
rect 10591 4324 10647 4380
rect 10647 4324 10651 4380
rect 10587 4320 10651 4324
rect 10667 4380 10731 4384
rect 10667 4324 10671 4380
rect 10671 4324 10727 4380
rect 10727 4324 10731 4380
rect 10667 4320 10731 4324
rect 19903 4380 19967 4384
rect 19903 4324 19907 4380
rect 19907 4324 19963 4380
rect 19963 4324 19967 4380
rect 19903 4320 19967 4324
rect 19983 4380 20047 4384
rect 19983 4324 19987 4380
rect 19987 4324 20043 4380
rect 20043 4324 20047 4380
rect 19983 4320 20047 4324
rect 20063 4380 20127 4384
rect 20063 4324 20067 4380
rect 20067 4324 20123 4380
rect 20123 4324 20127 4380
rect 20063 4320 20127 4324
rect 20143 4380 20207 4384
rect 20143 4324 20147 4380
rect 20147 4324 20203 4380
rect 20203 4324 20207 4380
rect 20143 4320 20207 4324
rect 13308 3980 13372 4044
rect 5690 3836 5754 3840
rect 5690 3780 5694 3836
rect 5694 3780 5750 3836
rect 5750 3780 5754 3836
rect 5690 3776 5754 3780
rect 5770 3836 5834 3840
rect 5770 3780 5774 3836
rect 5774 3780 5830 3836
rect 5830 3780 5834 3836
rect 5770 3776 5834 3780
rect 5850 3836 5914 3840
rect 5850 3780 5854 3836
rect 5854 3780 5910 3836
rect 5910 3780 5914 3836
rect 5850 3776 5914 3780
rect 5930 3836 5994 3840
rect 5930 3780 5934 3836
rect 5934 3780 5990 3836
rect 5990 3780 5994 3836
rect 5930 3776 5994 3780
rect 15165 3836 15229 3840
rect 15165 3780 15169 3836
rect 15169 3780 15225 3836
rect 15225 3780 15229 3836
rect 15165 3776 15229 3780
rect 15245 3836 15309 3840
rect 15245 3780 15249 3836
rect 15249 3780 15305 3836
rect 15305 3780 15309 3836
rect 15245 3776 15309 3780
rect 15325 3836 15389 3840
rect 15325 3780 15329 3836
rect 15329 3780 15385 3836
rect 15385 3780 15389 3836
rect 15325 3776 15389 3780
rect 15405 3836 15469 3840
rect 15405 3780 15409 3836
rect 15409 3780 15465 3836
rect 15465 3780 15469 3836
rect 15405 3776 15469 3780
rect 24641 3836 24705 3840
rect 24641 3780 24645 3836
rect 24645 3780 24701 3836
rect 24701 3780 24705 3836
rect 24641 3776 24705 3780
rect 24721 3836 24785 3840
rect 24721 3780 24725 3836
rect 24725 3780 24781 3836
rect 24781 3780 24785 3836
rect 24721 3776 24785 3780
rect 24801 3836 24865 3840
rect 24801 3780 24805 3836
rect 24805 3780 24861 3836
rect 24861 3780 24865 3836
rect 24801 3776 24865 3780
rect 24881 3836 24945 3840
rect 24881 3780 24885 3836
rect 24885 3780 24941 3836
rect 24941 3780 24945 3836
rect 24881 3776 24945 3780
rect 10427 3292 10491 3296
rect 10427 3236 10431 3292
rect 10431 3236 10487 3292
rect 10487 3236 10491 3292
rect 10427 3232 10491 3236
rect 10507 3292 10571 3296
rect 10507 3236 10511 3292
rect 10511 3236 10567 3292
rect 10567 3236 10571 3292
rect 10507 3232 10571 3236
rect 10587 3292 10651 3296
rect 10587 3236 10591 3292
rect 10591 3236 10647 3292
rect 10647 3236 10651 3292
rect 10587 3232 10651 3236
rect 10667 3292 10731 3296
rect 10667 3236 10671 3292
rect 10671 3236 10727 3292
rect 10727 3236 10731 3292
rect 10667 3232 10731 3236
rect 19903 3292 19967 3296
rect 19903 3236 19907 3292
rect 19907 3236 19963 3292
rect 19963 3236 19967 3292
rect 19903 3232 19967 3236
rect 19983 3292 20047 3296
rect 19983 3236 19987 3292
rect 19987 3236 20043 3292
rect 20043 3236 20047 3292
rect 19983 3232 20047 3236
rect 20063 3292 20127 3296
rect 20063 3236 20067 3292
rect 20067 3236 20123 3292
rect 20123 3236 20127 3292
rect 20063 3232 20127 3236
rect 20143 3292 20207 3296
rect 20143 3236 20147 3292
rect 20147 3236 20203 3292
rect 20203 3236 20207 3292
rect 20143 3232 20207 3236
rect 5690 2748 5754 2752
rect 5690 2692 5694 2748
rect 5694 2692 5750 2748
rect 5750 2692 5754 2748
rect 5690 2688 5754 2692
rect 5770 2748 5834 2752
rect 5770 2692 5774 2748
rect 5774 2692 5830 2748
rect 5830 2692 5834 2748
rect 5770 2688 5834 2692
rect 5850 2748 5914 2752
rect 5850 2692 5854 2748
rect 5854 2692 5910 2748
rect 5910 2692 5914 2748
rect 5850 2688 5914 2692
rect 5930 2748 5994 2752
rect 5930 2692 5934 2748
rect 5934 2692 5990 2748
rect 5990 2692 5994 2748
rect 5930 2688 5994 2692
rect 15165 2748 15229 2752
rect 15165 2692 15169 2748
rect 15169 2692 15225 2748
rect 15225 2692 15229 2748
rect 15165 2688 15229 2692
rect 15245 2748 15309 2752
rect 15245 2692 15249 2748
rect 15249 2692 15305 2748
rect 15305 2692 15309 2748
rect 15245 2688 15309 2692
rect 15325 2748 15389 2752
rect 15325 2692 15329 2748
rect 15329 2692 15385 2748
rect 15385 2692 15389 2748
rect 15325 2688 15389 2692
rect 15405 2748 15469 2752
rect 15405 2692 15409 2748
rect 15409 2692 15465 2748
rect 15465 2692 15469 2748
rect 15405 2688 15469 2692
rect 24641 2748 24705 2752
rect 24641 2692 24645 2748
rect 24645 2692 24701 2748
rect 24701 2692 24705 2748
rect 24641 2688 24705 2692
rect 24721 2748 24785 2752
rect 24721 2692 24725 2748
rect 24725 2692 24781 2748
rect 24781 2692 24785 2748
rect 24721 2688 24785 2692
rect 24801 2748 24865 2752
rect 24801 2692 24805 2748
rect 24805 2692 24861 2748
rect 24861 2692 24865 2748
rect 24801 2688 24865 2692
rect 24881 2748 24945 2752
rect 24881 2692 24885 2748
rect 24885 2692 24941 2748
rect 24941 2692 24945 2748
rect 24881 2688 24945 2692
rect 10427 2204 10491 2208
rect 10427 2148 10431 2204
rect 10431 2148 10487 2204
rect 10487 2148 10491 2204
rect 10427 2144 10491 2148
rect 10507 2204 10571 2208
rect 10507 2148 10511 2204
rect 10511 2148 10567 2204
rect 10567 2148 10571 2204
rect 10507 2144 10571 2148
rect 10587 2204 10651 2208
rect 10587 2148 10591 2204
rect 10591 2148 10647 2204
rect 10647 2148 10651 2204
rect 10587 2144 10651 2148
rect 10667 2204 10731 2208
rect 10667 2148 10671 2204
rect 10671 2148 10727 2204
rect 10727 2148 10731 2204
rect 10667 2144 10731 2148
rect 19903 2204 19967 2208
rect 19903 2148 19907 2204
rect 19907 2148 19963 2204
rect 19963 2148 19967 2204
rect 19903 2144 19967 2148
rect 19983 2204 20047 2208
rect 19983 2148 19987 2204
rect 19987 2148 20043 2204
rect 20043 2148 20047 2204
rect 19983 2144 20047 2148
rect 20063 2204 20127 2208
rect 20063 2148 20067 2204
rect 20067 2148 20123 2204
rect 20123 2148 20127 2204
rect 20063 2144 20127 2148
rect 20143 2204 20207 2208
rect 20143 2148 20147 2204
rect 20147 2148 20203 2204
rect 20203 2148 20207 2204
rect 20143 2144 20207 2148
<< metal4 >>
rect 5681 29952 6002 30512
rect 5681 29888 5690 29952
rect 5754 29888 5770 29952
rect 5834 29888 5850 29952
rect 5914 29888 5930 29952
rect 5994 29888 6002 29952
rect 5681 28864 6002 29888
rect 5681 28800 5690 28864
rect 5754 28800 5770 28864
rect 5834 28800 5850 28864
rect 5914 28800 5930 28864
rect 5994 28800 6002 28864
rect 5681 27776 6002 28800
rect 5681 27712 5690 27776
rect 5754 27712 5770 27776
rect 5834 27712 5850 27776
rect 5914 27712 5930 27776
rect 5994 27712 6002 27776
rect 5681 26688 6002 27712
rect 5681 26624 5690 26688
rect 5754 26624 5770 26688
rect 5834 26624 5850 26688
rect 5914 26624 5930 26688
rect 5994 26624 6002 26688
rect 5681 25600 6002 26624
rect 5681 25536 5690 25600
rect 5754 25536 5770 25600
rect 5834 25536 5850 25600
rect 5914 25536 5930 25600
rect 5994 25536 6002 25600
rect 5681 24512 6002 25536
rect 5681 24448 5690 24512
rect 5754 24448 5770 24512
rect 5834 24448 5850 24512
rect 5914 24448 5930 24512
rect 5994 24448 6002 24512
rect 5681 23424 6002 24448
rect 5681 23360 5690 23424
rect 5754 23360 5770 23424
rect 5834 23360 5850 23424
rect 5914 23360 5930 23424
rect 5994 23360 6002 23424
rect 5681 22336 6002 23360
rect 5681 22272 5690 22336
rect 5754 22272 5770 22336
rect 5834 22272 5850 22336
rect 5914 22272 5930 22336
rect 5994 22272 6002 22336
rect 5681 21248 6002 22272
rect 5681 21184 5690 21248
rect 5754 21184 5770 21248
rect 5834 21184 5850 21248
rect 5914 21184 5930 21248
rect 5994 21184 6002 21248
rect 5681 20160 6002 21184
rect 5681 20096 5690 20160
rect 5754 20096 5770 20160
rect 5834 20096 5850 20160
rect 5914 20096 5930 20160
rect 5994 20096 6002 20160
rect 5681 19072 6002 20096
rect 5681 19008 5690 19072
rect 5754 19008 5770 19072
rect 5834 19008 5850 19072
rect 5914 19008 5930 19072
rect 5994 19008 6002 19072
rect 5681 17984 6002 19008
rect 5681 17920 5690 17984
rect 5754 17920 5770 17984
rect 5834 17920 5850 17984
rect 5914 17920 5930 17984
rect 5994 17920 6002 17984
rect 5681 16896 6002 17920
rect 5681 16832 5690 16896
rect 5754 16832 5770 16896
rect 5834 16832 5850 16896
rect 5914 16832 5930 16896
rect 5994 16832 6002 16896
rect 5681 15808 6002 16832
rect 5681 15744 5690 15808
rect 5754 15744 5770 15808
rect 5834 15744 5850 15808
rect 5914 15744 5930 15808
rect 5994 15744 6002 15808
rect 5681 14720 6002 15744
rect 5681 14656 5690 14720
rect 5754 14656 5770 14720
rect 5834 14656 5850 14720
rect 5914 14656 5930 14720
rect 5994 14656 6002 14720
rect 5681 13632 6002 14656
rect 5681 13568 5690 13632
rect 5754 13568 5770 13632
rect 5834 13568 5850 13632
rect 5914 13568 5930 13632
rect 5994 13568 6002 13632
rect 5681 12544 6002 13568
rect 5681 12480 5690 12544
rect 5754 12480 5770 12544
rect 5834 12480 5850 12544
rect 5914 12480 5930 12544
rect 5994 12480 6002 12544
rect 5681 11456 6002 12480
rect 5681 11392 5690 11456
rect 5754 11392 5770 11456
rect 5834 11392 5850 11456
rect 5914 11392 5930 11456
rect 5994 11392 6002 11456
rect 5681 10368 6002 11392
rect 5681 10304 5690 10368
rect 5754 10304 5770 10368
rect 5834 10304 5850 10368
rect 5914 10304 5930 10368
rect 5994 10304 6002 10368
rect 5681 9280 6002 10304
rect 5681 9216 5690 9280
rect 5754 9216 5770 9280
rect 5834 9216 5850 9280
rect 5914 9216 5930 9280
rect 5994 9216 6002 9280
rect 5681 8192 6002 9216
rect 5681 8128 5690 8192
rect 5754 8128 5770 8192
rect 5834 8128 5850 8192
rect 5914 8128 5930 8192
rect 5994 8128 6002 8192
rect 5681 7104 6002 8128
rect 5681 7040 5690 7104
rect 5754 7040 5770 7104
rect 5834 7040 5850 7104
rect 5914 7040 5930 7104
rect 5994 7040 6002 7104
rect 5681 6016 6002 7040
rect 5681 5952 5690 6016
rect 5754 5952 5770 6016
rect 5834 5952 5850 6016
rect 5914 5952 5930 6016
rect 5994 5952 6002 6016
rect 5681 4928 6002 5952
rect 5681 4864 5690 4928
rect 5754 4864 5770 4928
rect 5834 4864 5850 4928
rect 5914 4864 5930 4928
rect 5994 4864 6002 4928
rect 5681 3840 6002 4864
rect 5681 3776 5690 3840
rect 5754 3776 5770 3840
rect 5834 3776 5850 3840
rect 5914 3776 5930 3840
rect 5994 3776 6002 3840
rect 5681 2752 6002 3776
rect 5681 2688 5690 2752
rect 5754 2688 5770 2752
rect 5834 2688 5850 2752
rect 5914 2688 5930 2752
rect 5994 2688 6002 2752
rect 5681 2128 6002 2688
rect 10419 30496 10739 30512
rect 10419 30432 10427 30496
rect 10491 30432 10507 30496
rect 10571 30432 10587 30496
rect 10651 30432 10667 30496
rect 10731 30432 10739 30496
rect 10419 29408 10739 30432
rect 10419 29344 10427 29408
rect 10491 29344 10507 29408
rect 10571 29344 10587 29408
rect 10651 29344 10667 29408
rect 10731 29344 10739 29408
rect 10419 28320 10739 29344
rect 10419 28256 10427 28320
rect 10491 28256 10507 28320
rect 10571 28256 10587 28320
rect 10651 28256 10667 28320
rect 10731 28256 10739 28320
rect 10419 27232 10739 28256
rect 15157 29952 15477 30512
rect 15157 29888 15165 29952
rect 15229 29888 15245 29952
rect 15309 29888 15325 29952
rect 15389 29888 15405 29952
rect 15469 29888 15477 29952
rect 15157 28864 15477 29888
rect 15157 28800 15165 28864
rect 15229 28800 15245 28864
rect 15309 28800 15325 28864
rect 15389 28800 15405 28864
rect 15469 28800 15477 28864
rect 15157 27776 15477 28800
rect 15157 27712 15165 27776
rect 15229 27712 15245 27776
rect 15309 27712 15325 27776
rect 15389 27712 15405 27776
rect 15469 27712 15477 27776
rect 13307 27300 13373 27301
rect 13307 27236 13308 27300
rect 13372 27236 13373 27300
rect 13307 27235 13373 27236
rect 10419 27168 10427 27232
rect 10491 27168 10507 27232
rect 10571 27168 10587 27232
rect 10651 27168 10667 27232
rect 10731 27168 10739 27232
rect 10419 26144 10739 27168
rect 10419 26080 10427 26144
rect 10491 26080 10507 26144
rect 10571 26080 10587 26144
rect 10651 26080 10667 26144
rect 10731 26080 10739 26144
rect 10419 25056 10739 26080
rect 10419 24992 10427 25056
rect 10491 24992 10507 25056
rect 10571 24992 10587 25056
rect 10651 24992 10667 25056
rect 10731 24992 10739 25056
rect 10419 23968 10739 24992
rect 10419 23904 10427 23968
rect 10491 23904 10507 23968
rect 10571 23904 10587 23968
rect 10651 23904 10667 23968
rect 10731 23904 10739 23968
rect 10419 22880 10739 23904
rect 10419 22816 10427 22880
rect 10491 22816 10507 22880
rect 10571 22816 10587 22880
rect 10651 22816 10667 22880
rect 10731 22816 10739 22880
rect 10419 21792 10739 22816
rect 10419 21728 10427 21792
rect 10491 21728 10507 21792
rect 10571 21728 10587 21792
rect 10651 21728 10667 21792
rect 10731 21728 10739 21792
rect 10419 20704 10739 21728
rect 10419 20640 10427 20704
rect 10491 20640 10507 20704
rect 10571 20640 10587 20704
rect 10651 20640 10667 20704
rect 10731 20640 10739 20704
rect 10419 19616 10739 20640
rect 10419 19552 10427 19616
rect 10491 19552 10507 19616
rect 10571 19552 10587 19616
rect 10651 19552 10667 19616
rect 10731 19552 10739 19616
rect 10419 18528 10739 19552
rect 10419 18464 10427 18528
rect 10491 18464 10507 18528
rect 10571 18464 10587 18528
rect 10651 18464 10667 18528
rect 10731 18464 10739 18528
rect 10419 17440 10739 18464
rect 10419 17376 10427 17440
rect 10491 17376 10507 17440
rect 10571 17376 10587 17440
rect 10651 17376 10667 17440
rect 10731 17376 10739 17440
rect 10419 16352 10739 17376
rect 10419 16288 10427 16352
rect 10491 16288 10507 16352
rect 10571 16288 10587 16352
rect 10651 16288 10667 16352
rect 10731 16288 10739 16352
rect 10419 15264 10739 16288
rect 10419 15200 10427 15264
rect 10491 15200 10507 15264
rect 10571 15200 10587 15264
rect 10651 15200 10667 15264
rect 10731 15200 10739 15264
rect 10419 14176 10739 15200
rect 10419 14112 10427 14176
rect 10491 14112 10507 14176
rect 10571 14112 10587 14176
rect 10651 14112 10667 14176
rect 10731 14112 10739 14176
rect 10419 13088 10739 14112
rect 10419 13024 10427 13088
rect 10491 13024 10507 13088
rect 10571 13024 10587 13088
rect 10651 13024 10667 13088
rect 10731 13024 10739 13088
rect 10419 12000 10739 13024
rect 10419 11936 10427 12000
rect 10491 11936 10507 12000
rect 10571 11936 10587 12000
rect 10651 11936 10667 12000
rect 10731 11936 10739 12000
rect 10419 10912 10739 11936
rect 10915 11116 10981 11117
rect 10915 11052 10916 11116
rect 10980 11052 10981 11116
rect 10915 11051 10981 11052
rect 10419 10848 10427 10912
rect 10491 10848 10507 10912
rect 10571 10848 10587 10912
rect 10651 10848 10667 10912
rect 10731 10848 10739 10912
rect 10419 9824 10739 10848
rect 10918 10573 10978 11051
rect 10915 10572 10981 10573
rect 10915 10508 10916 10572
rect 10980 10508 10981 10572
rect 10915 10507 10981 10508
rect 10419 9760 10427 9824
rect 10491 9760 10507 9824
rect 10571 9760 10587 9824
rect 10651 9760 10667 9824
rect 10731 9760 10739 9824
rect 10419 8736 10739 9760
rect 10419 8672 10427 8736
rect 10491 8672 10507 8736
rect 10571 8672 10587 8736
rect 10651 8672 10667 8736
rect 10731 8672 10739 8736
rect 10419 7648 10739 8672
rect 10419 7584 10427 7648
rect 10491 7584 10507 7648
rect 10571 7584 10587 7648
rect 10651 7584 10667 7648
rect 10731 7584 10739 7648
rect 10419 6560 10739 7584
rect 10419 6496 10427 6560
rect 10491 6496 10507 6560
rect 10571 6496 10587 6560
rect 10651 6496 10667 6560
rect 10731 6496 10739 6560
rect 10419 5472 10739 6496
rect 10419 5408 10427 5472
rect 10491 5408 10507 5472
rect 10571 5408 10587 5472
rect 10651 5408 10667 5472
rect 10731 5408 10739 5472
rect 10419 4384 10739 5408
rect 10419 4320 10427 4384
rect 10491 4320 10507 4384
rect 10571 4320 10587 4384
rect 10651 4320 10667 4384
rect 10731 4320 10739 4384
rect 10419 3296 10739 4320
rect 13310 4045 13370 27235
rect 15157 26688 15477 27712
rect 15157 26624 15165 26688
rect 15229 26624 15245 26688
rect 15309 26624 15325 26688
rect 15389 26624 15405 26688
rect 15469 26624 15477 26688
rect 15157 25600 15477 26624
rect 15157 25536 15165 25600
rect 15229 25536 15245 25600
rect 15309 25536 15325 25600
rect 15389 25536 15405 25600
rect 15469 25536 15477 25600
rect 15157 24512 15477 25536
rect 15157 24448 15165 24512
rect 15229 24448 15245 24512
rect 15309 24448 15325 24512
rect 15389 24448 15405 24512
rect 15469 24448 15477 24512
rect 13675 23492 13741 23493
rect 13675 23428 13676 23492
rect 13740 23428 13741 23492
rect 13675 23427 13741 23428
rect 13678 15469 13738 23427
rect 15157 23424 15477 24448
rect 19895 30496 20215 30512
rect 19895 30432 19903 30496
rect 19967 30432 19983 30496
rect 20047 30432 20063 30496
rect 20127 30432 20143 30496
rect 20207 30432 20215 30496
rect 19895 29408 20215 30432
rect 19895 29344 19903 29408
rect 19967 29344 19983 29408
rect 20047 29344 20063 29408
rect 20127 29344 20143 29408
rect 20207 29344 20215 29408
rect 19895 28320 20215 29344
rect 19895 28256 19903 28320
rect 19967 28256 19983 28320
rect 20047 28256 20063 28320
rect 20127 28256 20143 28320
rect 20207 28256 20215 28320
rect 19895 27232 20215 28256
rect 19895 27168 19903 27232
rect 19967 27168 19983 27232
rect 20047 27168 20063 27232
rect 20127 27168 20143 27232
rect 20207 27168 20215 27232
rect 19895 26144 20215 27168
rect 19895 26080 19903 26144
rect 19967 26080 19983 26144
rect 20047 26080 20063 26144
rect 20127 26080 20143 26144
rect 20207 26080 20215 26144
rect 19895 25056 20215 26080
rect 24633 29952 24953 30512
rect 24633 29888 24641 29952
rect 24705 29888 24721 29952
rect 24785 29888 24801 29952
rect 24865 29888 24881 29952
rect 24945 29888 24953 29952
rect 24633 28864 24953 29888
rect 24633 28800 24641 28864
rect 24705 28800 24721 28864
rect 24785 28800 24801 28864
rect 24865 28800 24881 28864
rect 24945 28800 24953 28864
rect 24633 27776 24953 28800
rect 24633 27712 24641 27776
rect 24705 27712 24721 27776
rect 24785 27712 24801 27776
rect 24865 27712 24881 27776
rect 24945 27712 24953 27776
rect 24633 26688 24953 27712
rect 24633 26624 24641 26688
rect 24705 26624 24721 26688
rect 24785 26624 24801 26688
rect 24865 26624 24881 26688
rect 24945 26624 24953 26688
rect 24633 25600 24953 26624
rect 24633 25536 24641 25600
rect 24705 25536 24721 25600
rect 24785 25536 24801 25600
rect 24865 25536 24881 25600
rect 24945 25536 24953 25600
rect 20483 25260 20549 25261
rect 20483 25196 20484 25260
rect 20548 25196 20549 25260
rect 20483 25195 20549 25196
rect 19895 24992 19903 25056
rect 19967 24992 19983 25056
rect 20047 24992 20063 25056
rect 20127 24992 20143 25056
rect 20207 24992 20215 25056
rect 19895 23968 20215 24992
rect 19895 23904 19903 23968
rect 19967 23904 19983 23968
rect 20047 23904 20063 23968
rect 20127 23904 20143 23968
rect 20207 23904 20215 23968
rect 19747 23628 19813 23629
rect 19747 23564 19748 23628
rect 19812 23564 19813 23628
rect 19747 23563 19813 23564
rect 15157 23360 15165 23424
rect 15229 23360 15245 23424
rect 15309 23360 15325 23424
rect 15389 23360 15405 23424
rect 15469 23360 15477 23424
rect 15157 22336 15477 23360
rect 15157 22272 15165 22336
rect 15229 22272 15245 22336
rect 15309 22272 15325 22336
rect 15389 22272 15405 22336
rect 15469 22272 15477 22336
rect 15157 21248 15477 22272
rect 15157 21184 15165 21248
rect 15229 21184 15245 21248
rect 15309 21184 15325 21248
rect 15389 21184 15405 21248
rect 15469 21184 15477 21248
rect 15157 20160 15477 21184
rect 15157 20096 15165 20160
rect 15229 20096 15245 20160
rect 15309 20096 15325 20160
rect 15389 20096 15405 20160
rect 15469 20096 15477 20160
rect 15157 19072 15477 20096
rect 15157 19008 15165 19072
rect 15229 19008 15245 19072
rect 15309 19008 15325 19072
rect 15389 19008 15405 19072
rect 15469 19008 15477 19072
rect 15157 17984 15477 19008
rect 15157 17920 15165 17984
rect 15229 17920 15245 17984
rect 15309 17920 15325 17984
rect 15389 17920 15405 17984
rect 15469 17920 15477 17984
rect 15157 16896 15477 17920
rect 19750 16965 19810 23563
rect 19895 22880 20215 23904
rect 19895 22816 19903 22880
rect 19967 22816 19983 22880
rect 20047 22816 20063 22880
rect 20127 22816 20143 22880
rect 20207 22816 20215 22880
rect 19895 21792 20215 22816
rect 19895 21728 19903 21792
rect 19967 21728 19983 21792
rect 20047 21728 20063 21792
rect 20127 21728 20143 21792
rect 20207 21728 20215 21792
rect 19895 20704 20215 21728
rect 19895 20640 19903 20704
rect 19967 20640 19983 20704
rect 20047 20640 20063 20704
rect 20127 20640 20143 20704
rect 20207 20640 20215 20704
rect 19895 19616 20215 20640
rect 19895 19552 19903 19616
rect 19967 19552 19983 19616
rect 20047 19552 20063 19616
rect 20127 19552 20143 19616
rect 20207 19552 20215 19616
rect 19895 18528 20215 19552
rect 19895 18464 19903 18528
rect 19967 18464 19983 18528
rect 20047 18464 20063 18528
rect 20127 18464 20143 18528
rect 20207 18464 20215 18528
rect 19895 17440 20215 18464
rect 20486 17917 20546 25195
rect 24633 24512 24953 25536
rect 24633 24448 24641 24512
rect 24705 24448 24721 24512
rect 24785 24448 24801 24512
rect 24865 24448 24881 24512
rect 24945 24448 24953 24512
rect 24633 23424 24953 24448
rect 24633 23360 24641 23424
rect 24705 23360 24721 23424
rect 24785 23360 24801 23424
rect 24865 23360 24881 23424
rect 24945 23360 24953 23424
rect 24633 22336 24953 23360
rect 24633 22272 24641 22336
rect 24705 22272 24721 22336
rect 24785 22272 24801 22336
rect 24865 22272 24881 22336
rect 24945 22272 24953 22336
rect 24633 21248 24953 22272
rect 24633 21184 24641 21248
rect 24705 21184 24721 21248
rect 24785 21184 24801 21248
rect 24865 21184 24881 21248
rect 24945 21184 24953 21248
rect 24633 20160 24953 21184
rect 24633 20096 24641 20160
rect 24705 20096 24721 20160
rect 24785 20096 24801 20160
rect 24865 20096 24881 20160
rect 24945 20096 24953 20160
rect 24633 19072 24953 20096
rect 24633 19008 24641 19072
rect 24705 19008 24721 19072
rect 24785 19008 24801 19072
rect 24865 19008 24881 19072
rect 24945 19008 24953 19072
rect 24633 17984 24953 19008
rect 24633 17920 24641 17984
rect 24705 17920 24721 17984
rect 24785 17920 24801 17984
rect 24865 17920 24881 17984
rect 24945 17920 24953 17984
rect 20483 17916 20549 17917
rect 20483 17852 20484 17916
rect 20548 17852 20549 17916
rect 20483 17851 20549 17852
rect 19895 17376 19903 17440
rect 19967 17376 19983 17440
rect 20047 17376 20063 17440
rect 20127 17376 20143 17440
rect 20207 17376 20215 17440
rect 19747 16964 19813 16965
rect 19747 16900 19748 16964
rect 19812 16900 19813 16964
rect 19747 16899 19813 16900
rect 15157 16832 15165 16896
rect 15229 16832 15245 16896
rect 15309 16832 15325 16896
rect 15389 16832 15405 16896
rect 15469 16832 15477 16896
rect 15157 15808 15477 16832
rect 15157 15744 15165 15808
rect 15229 15744 15245 15808
rect 15309 15744 15325 15808
rect 15389 15744 15405 15808
rect 15469 15744 15477 15808
rect 13675 15468 13741 15469
rect 13675 15404 13676 15468
rect 13740 15404 13741 15468
rect 13675 15403 13741 15404
rect 15157 14720 15477 15744
rect 15157 14656 15165 14720
rect 15229 14656 15245 14720
rect 15309 14656 15325 14720
rect 15389 14656 15405 14720
rect 15469 14656 15477 14720
rect 15157 13632 15477 14656
rect 15157 13568 15165 13632
rect 15229 13568 15245 13632
rect 15309 13568 15325 13632
rect 15389 13568 15405 13632
rect 15469 13568 15477 13632
rect 15157 12544 15477 13568
rect 15157 12480 15165 12544
rect 15229 12480 15245 12544
rect 15309 12480 15325 12544
rect 15389 12480 15405 12544
rect 15469 12480 15477 12544
rect 15157 11456 15477 12480
rect 15157 11392 15165 11456
rect 15229 11392 15245 11456
rect 15309 11392 15325 11456
rect 15389 11392 15405 11456
rect 15469 11392 15477 11456
rect 15157 10368 15477 11392
rect 15157 10304 15165 10368
rect 15229 10304 15245 10368
rect 15309 10304 15325 10368
rect 15389 10304 15405 10368
rect 15469 10304 15477 10368
rect 15157 9280 15477 10304
rect 15157 9216 15165 9280
rect 15229 9216 15245 9280
rect 15309 9216 15325 9280
rect 15389 9216 15405 9280
rect 15469 9216 15477 9280
rect 15157 8192 15477 9216
rect 15157 8128 15165 8192
rect 15229 8128 15245 8192
rect 15309 8128 15325 8192
rect 15389 8128 15405 8192
rect 15469 8128 15477 8192
rect 15157 7104 15477 8128
rect 15157 7040 15165 7104
rect 15229 7040 15245 7104
rect 15309 7040 15325 7104
rect 15389 7040 15405 7104
rect 15469 7040 15477 7104
rect 15157 6016 15477 7040
rect 15157 5952 15165 6016
rect 15229 5952 15245 6016
rect 15309 5952 15325 6016
rect 15389 5952 15405 6016
rect 15469 5952 15477 6016
rect 15157 4928 15477 5952
rect 15157 4864 15165 4928
rect 15229 4864 15245 4928
rect 15309 4864 15325 4928
rect 15389 4864 15405 4928
rect 15469 4864 15477 4928
rect 13307 4044 13373 4045
rect 13307 3980 13308 4044
rect 13372 3980 13373 4044
rect 13307 3979 13373 3980
rect 10419 3232 10427 3296
rect 10491 3232 10507 3296
rect 10571 3232 10587 3296
rect 10651 3232 10667 3296
rect 10731 3232 10739 3296
rect 10419 2208 10739 3232
rect 10419 2144 10427 2208
rect 10491 2144 10507 2208
rect 10571 2144 10587 2208
rect 10651 2144 10667 2208
rect 10731 2144 10739 2208
rect 10419 2128 10739 2144
rect 15157 3840 15477 4864
rect 15157 3776 15165 3840
rect 15229 3776 15245 3840
rect 15309 3776 15325 3840
rect 15389 3776 15405 3840
rect 15469 3776 15477 3840
rect 15157 2752 15477 3776
rect 15157 2688 15165 2752
rect 15229 2688 15245 2752
rect 15309 2688 15325 2752
rect 15389 2688 15405 2752
rect 15469 2688 15477 2752
rect 15157 2128 15477 2688
rect 19895 16352 20215 17376
rect 19895 16288 19903 16352
rect 19967 16288 19983 16352
rect 20047 16288 20063 16352
rect 20127 16288 20143 16352
rect 20207 16288 20215 16352
rect 19895 15264 20215 16288
rect 19895 15200 19903 15264
rect 19967 15200 19983 15264
rect 20047 15200 20063 15264
rect 20127 15200 20143 15264
rect 20207 15200 20215 15264
rect 19895 14176 20215 15200
rect 19895 14112 19903 14176
rect 19967 14112 19983 14176
rect 20047 14112 20063 14176
rect 20127 14112 20143 14176
rect 20207 14112 20215 14176
rect 19895 13088 20215 14112
rect 19895 13024 19903 13088
rect 19967 13024 19983 13088
rect 20047 13024 20063 13088
rect 20127 13024 20143 13088
rect 20207 13024 20215 13088
rect 19895 12000 20215 13024
rect 19895 11936 19903 12000
rect 19967 11936 19983 12000
rect 20047 11936 20063 12000
rect 20127 11936 20143 12000
rect 20207 11936 20215 12000
rect 19895 10912 20215 11936
rect 19895 10848 19903 10912
rect 19967 10848 19983 10912
rect 20047 10848 20063 10912
rect 20127 10848 20143 10912
rect 20207 10848 20215 10912
rect 19895 9824 20215 10848
rect 19895 9760 19903 9824
rect 19967 9760 19983 9824
rect 20047 9760 20063 9824
rect 20127 9760 20143 9824
rect 20207 9760 20215 9824
rect 19895 8736 20215 9760
rect 19895 8672 19903 8736
rect 19967 8672 19983 8736
rect 20047 8672 20063 8736
rect 20127 8672 20143 8736
rect 20207 8672 20215 8736
rect 19895 7648 20215 8672
rect 19895 7584 19903 7648
rect 19967 7584 19983 7648
rect 20047 7584 20063 7648
rect 20127 7584 20143 7648
rect 20207 7584 20215 7648
rect 19895 6560 20215 7584
rect 19895 6496 19903 6560
rect 19967 6496 19983 6560
rect 20047 6496 20063 6560
rect 20127 6496 20143 6560
rect 20207 6496 20215 6560
rect 19895 5472 20215 6496
rect 19895 5408 19903 5472
rect 19967 5408 19983 5472
rect 20047 5408 20063 5472
rect 20127 5408 20143 5472
rect 20207 5408 20215 5472
rect 19895 4384 20215 5408
rect 19895 4320 19903 4384
rect 19967 4320 19983 4384
rect 20047 4320 20063 4384
rect 20127 4320 20143 4384
rect 20207 4320 20215 4384
rect 19895 3296 20215 4320
rect 19895 3232 19903 3296
rect 19967 3232 19983 3296
rect 20047 3232 20063 3296
rect 20127 3232 20143 3296
rect 20207 3232 20215 3296
rect 19895 2208 20215 3232
rect 19895 2144 19903 2208
rect 19967 2144 19983 2208
rect 20047 2144 20063 2208
rect 20127 2144 20143 2208
rect 20207 2144 20215 2208
rect 19895 2128 20215 2144
rect 24633 16896 24953 17920
rect 24633 16832 24641 16896
rect 24705 16832 24721 16896
rect 24785 16832 24801 16896
rect 24865 16832 24881 16896
rect 24945 16832 24953 16896
rect 24633 15808 24953 16832
rect 24633 15744 24641 15808
rect 24705 15744 24721 15808
rect 24785 15744 24801 15808
rect 24865 15744 24881 15808
rect 24945 15744 24953 15808
rect 24633 14720 24953 15744
rect 24633 14656 24641 14720
rect 24705 14656 24721 14720
rect 24785 14656 24801 14720
rect 24865 14656 24881 14720
rect 24945 14656 24953 14720
rect 24633 13632 24953 14656
rect 24633 13568 24641 13632
rect 24705 13568 24721 13632
rect 24785 13568 24801 13632
rect 24865 13568 24881 13632
rect 24945 13568 24953 13632
rect 24633 12544 24953 13568
rect 24633 12480 24641 12544
rect 24705 12480 24721 12544
rect 24785 12480 24801 12544
rect 24865 12480 24881 12544
rect 24945 12480 24953 12544
rect 24633 11456 24953 12480
rect 24633 11392 24641 11456
rect 24705 11392 24721 11456
rect 24785 11392 24801 11456
rect 24865 11392 24881 11456
rect 24945 11392 24953 11456
rect 24633 10368 24953 11392
rect 24633 10304 24641 10368
rect 24705 10304 24721 10368
rect 24785 10304 24801 10368
rect 24865 10304 24881 10368
rect 24945 10304 24953 10368
rect 24633 9280 24953 10304
rect 24633 9216 24641 9280
rect 24705 9216 24721 9280
rect 24785 9216 24801 9280
rect 24865 9216 24881 9280
rect 24945 9216 24953 9280
rect 24633 8192 24953 9216
rect 24633 8128 24641 8192
rect 24705 8128 24721 8192
rect 24785 8128 24801 8192
rect 24865 8128 24881 8192
rect 24945 8128 24953 8192
rect 24633 7104 24953 8128
rect 24633 7040 24641 7104
rect 24705 7040 24721 7104
rect 24785 7040 24801 7104
rect 24865 7040 24881 7104
rect 24945 7040 24953 7104
rect 24633 6016 24953 7040
rect 24633 5952 24641 6016
rect 24705 5952 24721 6016
rect 24785 5952 24801 6016
rect 24865 5952 24881 6016
rect 24945 5952 24953 6016
rect 24633 4928 24953 5952
rect 24633 4864 24641 4928
rect 24705 4864 24721 4928
rect 24785 4864 24801 4928
rect 24865 4864 24881 4928
rect 24945 4864 24953 4928
rect 24633 3840 24953 4864
rect 24633 3776 24641 3840
rect 24705 3776 24721 3840
rect 24785 3776 24801 3840
rect 24865 3776 24881 3840
rect 24945 3776 24953 3840
rect 24633 2752 24953 3776
rect 24633 2688 24641 2752
rect 24705 2688 24721 2752
rect 24785 2688 24801 2752
rect 24865 2688 24881 2752
rect 24945 2688 24953 2752
rect 24633 2128 24953 2688
use sky130_fd_sc_hd__decap_12  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1640608721
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1640608721
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1640608721
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1640608721
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp 1640608721
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1788_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 4324 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1824_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 4140 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1640608721
transform 1 0 5152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1640608721
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1640608721
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1640608721
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1603_
timestamp 1640608721
transform -1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1610_
timestamp 1640608721
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1787_
timestamp 1640608721
transform 1 0 6440 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1825_
timestamp 1640608721
transform 1 0 6348 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_0_67
timestamp 1640608721
transform 1 0 7268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1640608721
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1640608721
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1640608721
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1625_
timestamp 1640608721
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1784_
timestamp 1640608721
transform 1 0 8924 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1828_
timestamp 1640608721
transform 1 0 8556 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106
timestamp 1640608721
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1640608721
transform 1 0 9752 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_102
timestamp 1640608721
transform 1 0 10488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_98
timestamp 1640608721
transform 1 0 10120 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1613_
timestamp 1640608721
transform 1 0 10580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_122
timestamp 1640608721
transform 1 0 12328 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_130
timestamp 1640608721
transform 1 0 13064 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1640608721
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1640608721
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1786_
timestamp 1640608721
transform 1 0 11500 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1826_
timestamp 1640608721
transform -1 0 13064 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1640608721
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1640608721
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_142 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 14168 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_150
timestamp 1640608721
transform 1 0 14904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1640608721
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1816_
timestamp 1640608721
transform 1 0 14996 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1640608721
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1640608721
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1640608721
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_174
timestamp 1640608721
transform 1 0 17112 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1640608721
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1640608721
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 16652 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_0_175
timestamp 1640608721
transform 1 0 17204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1640608721
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1640608721
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1640608721
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1813_
timestamp 1640608721
transform 1 0 18768 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1817_
timestamp 1640608721
transform 1 0 17204 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1640608721
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1640608721
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1504_
timestamp 1640608721
transform 1 0 20976 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _1506_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 20332 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1640608721
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1640608721
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1640608721
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1640608721
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_233
timestamp 1640608721
transform 1 0 22540 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1640608721
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1640608721
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1507_
timestamp 1640608721
transform 1 0 22264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1508_
timestamp 1640608721
transform -1 0 22264 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1640608721
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1640608721
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1640608721
transform 1 0 23644 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1640608721
transform 1 0 24748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1640608721
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1640608721
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1640608721
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1640608721
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1640608721
transform 1 0 25852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1640608721
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1640608721
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1640608721
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1640608721
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1640608721
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_305
timestamp 1640608721
transform 1 0 29164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1640608721
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_305
timestamp 1640608721
transform 1 0 29164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1640608721
transform -1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1640608721
transform -1 0 29532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1640608721
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1640608721
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1640608721
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1640608721
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1640608721
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_41
timestamp 1640608721
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1640608721
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1604_
timestamp 1640608721
transform -1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_55
timestamp 1640608721
transform 1 0 6164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 5428 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1608_
timestamp 1640608721
transform -1 0 7268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1609_
timestamp 1640608721
transform -1 0 6992 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 7268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1640608721
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1640608721
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1606_
timestamp 1640608721
transform 1 0 8188 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1607_
timestamp 1640608721
transform 1 0 7452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1624_
timestamp 1640608721
transform -1 0 9476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_101
timestamp 1640608721
transform 1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 10396 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1612_
timestamp 1640608721
transform 1 0 10672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1623_
timestamp 1640608721
transform -1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_120
timestamp 1640608721
transform 1 0 12144 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1611_
timestamp 1640608721
transform 1 0 11408 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1616_
timestamp 1640608721
transform 1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1640608721
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1640608721
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1640608721
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_153
timestamp 1640608721
transform 1 0 15180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_159
timestamp 1640608721
transform 1 0 15732 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1513_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 16652 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1757_
timestamp 1640608721
transform -1 0 16652 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1640608721
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1640608721
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1512_
timestamp 1640608721
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 19044 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _1518_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 17572 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_200
timestamp 1640608721
transform 1 0 19504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_210
timestamp 1640608721
transform 1 0 20424 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1517_
timestamp 1640608721
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1755_
timestamp 1640608721
transform 1 0 19596 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1814_
timestamp 1640608721
transform 1 0 20516 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_2_238
timestamp 1640608721
transform 1 0 23000 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1505_
timestamp 1640608721
transform 1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1509_
timestamp 1640608721
transform 1 0 22080 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_2_242
timestamp 1640608721
transform 1 0 23368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1640608721
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1640608721
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1801_
timestamp 1640608721
transform 1 0 23460 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1640608721
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1640608721
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1640608721
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_301
timestamp 1640608721
transform 1 0 28796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_305
timestamp 1640608721
transform 1 0 29164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1640608721
transform -1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_21
timestamp 1640608721
transform 1 0 3036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1640608721
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_9
timestamp 1640608721
transform 1 0 1932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1640608721
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1700_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_29
timestamp 1640608721
transform 1 0 3772 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_41
timestamp 1640608721
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 1640608721
transform 1 0 4048 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1640608721
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_63
timestamp 1640608721
transform 1 0 6900 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1640608721
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1640608721
transform 1 0 8004 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_82
timestamp 1640608721
transform 1 0 8648 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1223_
timestamp 1640608721
transform 1 0 8188 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_3_100
timestamp 1640608721
transform 1 0 10304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1640608721
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1640608721
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_2  _1618_
timestamp 1640608721
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1622_
timestamp 1640608721
transform 1 0 9200 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1640608721
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1640608721
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1640608721
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_137
timestamp 1640608721
transform 1 0 13708 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1815_
timestamp 1640608721
transform 1 0 14260 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_3_160
timestamp 1640608721
transform 1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1640608721
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 1640608721
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1640608721
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1511_
timestamp 1640608721
transform -1 0 16468 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1756_
timestamp 1640608721
transform 1 0 16744 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_179
timestamp 1640608721
transform 1 0 17572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_191
timestamp 1640608721
transform 1 0 18676 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1754_
timestamp 1640608721
transform -1 0 18676 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1640608721
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1812_
timestamp 1640608721
transform 1 0 19412 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_3_234
timestamp 1640608721
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1640608721
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_2  _1305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 21804 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1549_
timestamp 1640608721
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1833_
timestamp 1640608721
transform 1 0 23184 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_3_257
timestamp 1640608721
transform 1 0 24748 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_265
timestamp 1640608721
transform 1 0 25484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1640608721
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1640608721
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1640608721
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1640608721
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 25760 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1640608721
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_305
timestamp 1640608721
transform 1 0 29164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1640608721
transform -1 0 29532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1640608721
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1640608721
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1640608721
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1640608721
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1640608721
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1601_
timestamp 1640608721
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1823_
timestamp 1640608721
transform 1 0 4048 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_4_57
timestamp 1640608721
transform 1 0 6348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_65
timestamp 1640608721
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1228_
timestamp 1640608721
transform 1 0 6440 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1597_
timestamp 1640608721
transform 1 0 5612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_73
timestamp 1640608721
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1640608721
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1640608721
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1640608721
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1626_
timestamp 1640608721
transform 1 0 8924 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1628_
timestamp 1640608721
transform 1 0 8096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_104
timestamp 1640608721
transform 1 0 10672 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp 1640608721
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_90
timestamp 1640608721
transform 1 0 9384 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1617_
timestamp 1640608721
transform -1 0 10672 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1619_
timestamp 1640608721
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_129
timestamp 1640608721
transform 1 0 12972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1827_
timestamp 1640608721
transform -1 0 12972 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1640608721
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1640608721
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1640608721
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_153
timestamp 1640608721
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_164
timestamp 1640608721
transform 1 0 16192 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1510_
timestamp 1640608721
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_176
timestamp 1640608721
transform 1 0 17296 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_182
timestamp 1640608721
transform 1 0 17848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_186
timestamp 1640608721
transform 1 0 18216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1640608721
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1640608721
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1640608721
transform -1 0 18216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1640608721
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_209
timestamp 1640608721
transform 1 0 20332 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_217
timestamp 1640608721
transform 1 0 21068 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1306_
timestamp 1640608721
transform -1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_221
timestamp 1640608721
transform 1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_234
timestamp 1640608721
transform 1 0 22632 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1758_
timestamp 1640608721
transform 1 0 21804 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1640608721
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1640608721
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1545_
timestamp 1640608721
transform 1 0 24380 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1546_
timestamp 1640608721
transform -1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1548_
timestamp 1640608721
transform -1 0 24196 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1792_
timestamp 1640608721
transform -1 0 25944 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1842_
timestamp 1640608721
transform 1 0 25944 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_4_296
timestamp 1640608721
transform 1 0 28336 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_304
timestamp 1640608721
transform 1 0 29072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_2  _1299_
timestamp 1640608721
transform -1 0 28336 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1640608721
transform -1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1640608721
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1640608721
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1809_
timestamp 1640608721
transform 1 0 1932 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_5_26
timestamp 1640608721
transform 1 0 3496 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_38
timestamp 1640608721
transform 1 0 4600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_43
timestamp 1640608721
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1598_
timestamp 1640608721
transform -1 0 5060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1600_
timestamp 1640608721
transform -1 0 4600 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1640608721
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1640608721
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1596_
timestamp 1640608721
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1829_
timestamp 1640608721
transform -1 0 8372 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1783_
timestamp 1640608721
transform 1 0 8372 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_101
timestamp 1640608721
transform 1 0 10396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_105
timestamp 1640608721
transform 1 0 10764 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1224_
timestamp 1640608721
transform 1 0 9844 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1620_
timestamp 1640608721
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1627_
timestamp 1640608721
transform -1 0 9844 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1640608721
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1640608721
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1621_
timestamp 1640608721
transform -1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1785_
timestamp 1640608721
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1640608721
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_149
timestamp 1640608721
transform 1 0 14812 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1640608721
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1640608721
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1292_
timestamp 1640608721
transform 1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1728_
timestamp 1640608721
transform 1 0 15364 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1739_
timestamp 1640608721
transform 1 0 16652 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_178
timestamp 1640608721
transform 1 0 17480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1293_
timestamp 1640608721
transform 1 0 18400 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1725_
timestamp 1640608721
transform 1 0 18952 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1729_
timestamp 1640608721
transform 1 0 17572 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1640608721
transform 1 0 20884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1307_
timestamp 1640608721
transform -1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1724_
timestamp 1640608721
transform 1 0 19780 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_234
timestamp 1640608721
transform 1 0 22632 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1640608721
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1655_
timestamp 1640608721
transform 1 0 21252 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 1640608721
transform 1 0 21804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1802_
timestamp 1640608721
transform 1 0 23000 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_247
timestamp 1640608721
transform 1 0 23828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_259
timestamp 1640608721
transform 1 0 24932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_263
timestamp 1640608721
transform 1 0 25300 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_272
timestamp 1640608721
transform 1 0 26128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1640608721
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1640608721
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1640608721
transform -1 0 26128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1587_
timestamp 1640608721
transform 1 0 25392 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1640608721
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_305
timestamp 1640608721
transform 1 0 29164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1640608721
transform -1 0 29532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_20
timestamp 1640608721
transform 1 0 2944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1640608721
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1640608721
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1640608721
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1640608721
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1528_
timestamp 1640608721
transform 1 0 2852 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1808_
timestamp 1640608721
transform 1 0 1380 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1714_
timestamp 1640608721
transform 1 0 3496 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _1530_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1529_
timestamp 1640608721
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1640608721
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_24
timestamp 1640608721
transform 1 0 3312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1527_
timestamp 1640608721
transform -1 0 4600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1526_
timestamp 1640608721
transform 1 0 4508 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_7_38
timestamp 1640608721
transform 1 0 4600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1640608721
transform 1 0 4968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1821_
timestamp 1640608721
transform 1 0 4692 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_6_55
timestamp 1640608721
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_60
timestamp 1640608721
transform 1 0 6624 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1640608721
transform 1 0 6808 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1640608721
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1220_
timestamp 1640608721
transform -1 0 6808 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1227_
timestamp 1640608721
transform -1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1229_
timestamp 1640608721
transform -1 0 7544 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1791_
timestamp 1640608721
transform 1 0 5336 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_72
timestamp 1640608721
transform 1 0 7728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1640608721
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1640608721
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_70
timestamp 1640608721
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_74
timestamp 1640608721
transform 1 0 7912 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1640608721
transform 1 0 8464 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1640608721
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1629_
timestamp 1640608721
transform 1 0 7820 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1634_
timestamp 1640608721
transform 1 0 8004 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_7_92
timestamp 1640608721
transform 1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1630_
timestamp 1640608721
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 9292 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1632_
timestamp 1640608721
transform 1 0 11040 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1782_
timestamp 1640608721
transform -1 0 11040 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1830_
timestamp 1640608721
transform -1 0 11408 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_6_114
timestamp 1640608721
transform 1 0 11592 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_126
timestamp 1640608721
transform 1 0 12696 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1640608721
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1640608721
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1640608721
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1640608721
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_141
timestamp 1640608721
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_149
timestamp 1640608721
transform 1 0 14812 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1640608721
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_149
timestamp 1640608721
transform 1 0 14812 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1640608721
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1727_
timestamp 1640608721
transform 1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1640608721
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1640608721
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp 1640608721
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1640608721
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1289_
timestamp 1640608721
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1673_
timestamp 1640608721
transform 1 0 16652 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1674_
timestamp 1640608721
transform -1 0 17388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1675_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 15732 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_7_177
timestamp 1640608721
transform 1 0 17388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_187
timestamp 1640608721
transform 1 0 18308 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1640608721
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1660_
timestamp 1640608721
transform -1 0 19320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1676_
timestamp 1640608721
transform 1 0 17572 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1677_
timestamp 1640608721
transform 1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1678_
timestamp 1640608721
transform 1 0 17388 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1716_
timestamp 1640608721
transform 1 0 18308 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_198
timestamp 1640608721
transform 1 0 19320 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_210
timestamp 1640608721
transform 1 0 20424 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_2  _1308_
timestamp 1640608721
transform 1 0 19228 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1309_
timestamp 1640608721
transform -1 0 20148 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1659_
timestamp 1640608721
transform 1 0 20148 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1726_
timestamp 1640608721
transform 1 0 21068 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1640608721
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_228
timestamp 1640608721
transform 1 0 22080 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1640608721
transform 1 0 23184 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1640608721
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1290_
timestamp 1640608721
transform 1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1547_
timestamp 1640608721
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1656_
timestamp 1640608721
transform 1 0 22172 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1832_
timestamp 1640608721
transform 1 0 22448 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1640608721
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_247
timestamp 1640608721
transform 1 0 23828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_253
timestamp 1640608721
transform 1 0 24380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_259
timestamp 1640608721
transform 1 0 24932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1640608721
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1295_
timestamp 1640608721
transform 1 0 24472 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1301_
timestamp 1640608721
transform 1 0 25116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1540_
timestamp 1640608721
transform -1 0 23828 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _1544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_267
timestamp 1640608721
transform 1 0 25668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_282
timestamp 1640608721
transform 1 0 27048 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1640608721
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1543_
timestamp 1640608721
transform 1 0 25392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1585_
timestamp 1640608721
transform -1 0 27048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1586_
timestamp 1640608721
transform 1 0 26956 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1793_
timestamp 1640608721
transform 1 0 25944 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1841_
timestamp 1640608721
transform 1 0 25300 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_6_294
timestamp 1640608721
transform 1 0 28152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_286
timestamp 1640608721
transform 1 0 27416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_298
timestamp 1640608721
transform 1 0 28520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1640608721
transform -1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1640608721
transform -1 0 29532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_17
timestamp 1640608721
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1640608721
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1640608721
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1691_
timestamp 1640608721
transform -1 0 2668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1737_
timestamp 1640608721
transform 1 0 1564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1640608721
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_38
timestamp 1640608721
transform 1 0 4600 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1640608721
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1713_
timestamp 1640608721
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_55
timestamp 1640608721
transform 1 0 6164 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_65
timestamp 1640608721
transform 1 0 7084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1589_
timestamp 1640608721
transform -1 0 6164 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _1591_
timestamp 1640608721
transform 1 0 6348 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_71
timestamp 1640608721
transform 1 0 7636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1640608721
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1640608721
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_2  _1225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 9016 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1226_
timestamp 1640608721
transform -1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1230_
timestamp 1640608721
transform -1 0 7636 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1781_
timestamp 1640608721
transform -1 0 8832 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp 1640608721
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1640608721
transform 1 0 10764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_95
timestamp 1640608721
transform 1 0 9844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1633_
timestamp 1640608721
transform -1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1640608721
transform 1 0 11868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp 1640608721
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1640608721
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1640608721
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1640608721
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_153
timestamp 1640608721
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_173
timestamp 1640608721
transform 1 0 17020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1669_
timestamp 1640608721
transform 1 0 16560 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1712_
timestamp 1640608721
transform 1 0 15732 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1640608721
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1662_
timestamp 1640608721
transform 1 0 18676 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1664_
timestamp 1640608721
transform 1 0 18124 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1665__A1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp 1640608721
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_203
timestamp 1640608721
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_206
timestamp 1640608721
transform 1 0 20056 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_210
timestamp 1640608721
transform 1 0 20424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1658_
timestamp 1640608721
transform -1 0 21068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1661_
timestamp 1640608721
transform -1 0 21344 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_234
timestamp 1640608721
transform 1 0 22632 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1666_
timestamp 1640608721
transform -1 0 22632 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1761_
timestamp 1640608721
transform 1 0 21344 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1800_
timestamp 1640608721
transform 1 0 22908 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1640608721
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1640608721
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1640608721
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1302_
timestamp 1640608721
transform 1 0 24748 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_8_264
timestamp 1640608721
transform 1 0 25392 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_270
timestamp 1640608721
transform 1 0 25944 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1303_
timestamp 1640608721
transform -1 0 26680 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1584_
timestamp 1640608721
transform 1 0 26680 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_8_285
timestamp 1640608721
transform 1 0 27324 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1840_
timestamp 1640608721
transform 1 0 27692 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1640608721
transform -1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_12
timestamp 1640608721
transform 1 0 2208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1640608721
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1640608721
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1690_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 1564 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1738_
timestamp 1640608721
transform 1 0 2300 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_25
timestamp 1640608721
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_37
timestamp 1640608721
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1693_
timestamp 1640608721
transform -1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1640608721
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1640608721
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1640608721
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1640608721
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1590_
timestamp 1640608721
transform -1 0 7268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1592_
timestamp 1640608721
transform 1 0 6532 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_9_67
timestamp 1640608721
transform 1 0 7268 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_75
timestamp 1640608721
transform 1 0 8004 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1831_
timestamp 1640608721
transform 1 0 8188 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1640608721
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1640608721
transform 1 0 9752 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1640608721
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1640608721
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1640608721
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_137
timestamp 1640608721
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_145
timestamp 1640608721
transform 1 0 14444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1671_
timestamp 1640608721
transform 1 0 14720 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1640608721
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp 1640608721
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1640608721
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1310_
timestamp 1640608721
transform 1 0 16744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1670_
timestamp 1640608721
transform -1 0 16468 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1672_
timestamp 1640608721
transform 1 0 15272 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1747_
timestamp 1640608721
transform -1 0 17848 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1640608721
transform 1 0 17848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_2  _1665_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 18768 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1749_
timestamp 1640608721
transform -1 0 18768 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _1667_
timestamp 1640608721
transform 1 0 19872 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_2  _1668_
timestamp 1640608721
transform 1 0 20516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1640608721
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1640608721
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1640608721
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1552_
timestamp 1640608721
transform 1 0 22356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1834_
timestamp 1640608721
transform 1 0 22908 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_2  _1296_
timestamp 1640608721
transform 1 0 25208 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1550_
timestamp 1640608721
transform 1 0 24472 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_272
timestamp 1640608721
transform 1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1640608721
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1297_
timestamp 1640608721
transform 1 0 25668 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _1298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 27876 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_9_299
timestamp 1640608721
transform 1 0 28612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_305
timestamp 1640608721
transform 1 0 29164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1580_
timestamp 1640608721
transform -1 0 28612 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1640608721
transform -1 0 29532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1640608721
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1640608721
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1640608721
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1640608721
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1692_
timestamp 1640608721
transform 1 0 2208 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1640608721
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp 1640608721
transform 1 0 4784 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1640608721
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1218_
timestamp 1640608721
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _1523_
timestamp 1640608721
transform 1 0 4968 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1524_
timestamp 1640608721
transform -1 0 4784 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_10_50
timestamp 1640608721
transform 1 0 5704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_58
timestamp 1640608721
transform 1 0 6440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1790_
timestamp 1640608721
transform 1 0 6716 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1640608721
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1640608721
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1640608721
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1593_
timestamp 1640608721
transform -1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1595_
timestamp 1640608721
transform -1 0 8096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_92
timestamp 1640608721
transform 1 0 9568 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1640608721
transform -1 0 9568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1905_
timestamp 1640608721
transform -1 0 11684 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_10_115
timestamp 1640608721
transform 1 0 11684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_127
timestamp 1640608721
transform 1 0 12788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1640608721
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1640608721
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1640608721
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1640608721
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1640608721
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1640608721
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1640608721
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1640608721
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1541_
timestamp 1640608721
transform 1 0 17572 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1663_
timestamp 1640608721
transform -1 0 19136 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1640608721
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_209
timestamp 1640608721
transform 1 0 20332 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1657_
timestamp 1640608721
transform -1 0 21344 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__A
timestamp 1640608721
transform 1 0 22908 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_220
timestamp 1640608721
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_226
timestamp 1640608721
transform 1 0 21896 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_234
timestamp 1640608721
transform 1 0 22632 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1539_
timestamp 1640608721
transform 1 0 21620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1553_
timestamp 1640608721
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_242
timestamp 1640608721
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1640608721
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_253
timestamp 1640608721
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_262
timestamp 1640608721
transform 1 0 25208 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1640608721
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1551_
timestamp 1640608721
transform -1 0 23920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1555_
timestamp 1640608721
transform 1 0 24472 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1556_
timestamp 1640608721
transform -1 0 24196 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_270
timestamp 1640608721
transform 1 0 25944 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_274
timestamp 1640608721
transform 1 0 26312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_278
timestamp 1640608721
transform 1 0 26680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1554_
timestamp 1640608721
transform -1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1575_
timestamp 1640608721
transform 1 0 26772 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_10_284
timestamp 1640608721
transform 1 0 27232 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_290
timestamp 1640608721
transform 1 0 27784 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_304
timestamp 1640608721
transform 1 0 29072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1579_
timestamp 1640608721
transform -1 0 27784 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1581_
timestamp 1640608721
transform -1 0 29072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1794_
timestamp 1640608721
transform 1 0 27968 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1640608721
transform -1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_17
timestamp 1640608721
transform 1 0 2668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1640608721
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1640608721
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1640608721
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1733_
timestamp 1640608721
transform 1 0 1840 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp 1640608721
transform 1 0 4876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1521_
timestamp 1640608721
transform -1 0 4140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1525_
timestamp 1640608721
transform 1 0 4140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1718_
timestamp 1640608721
transform 1 0 4968 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1640608721
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1522_
timestamp 1640608721
transform 1 0 5796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1822_
timestamp 1640608721
transform 1 0 6348 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1640608721
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1906_
timestamp 1640608721
transform -1 0 9660 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__o221a_2  _1201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 10488 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _1206_
timestamp 1640608721
transform 1 0 10488 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A1
timestamp 1640608721
transform -1 0 11960 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1640608721
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_129
timestamp 1640608721
transform 1 0 12972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1640608721
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1202_
timestamp 1640608721
transform -1 0 12972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1205_
timestamp 1640608721
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1269_
timestamp 1640608721
transform 1 0 11960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_141
timestamp 1640608721
transform 1 0 14076 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_153
timestamp 1640608721
transform 1 0 15180 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1640608721
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 1640608721
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1640608721
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1647_
timestamp 1640608721
transform -1 0 17296 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1730_
timestamp 1640608721
transform -1 0 16284 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1640608721
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1640608721
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1286_
timestamp 1640608721
transform 1 0 17296 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1760_
timestamp 1640608721
transform 1 0 19044 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1760__A1
timestamp 1640608721
transform 1 0 19872 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_206
timestamp 1640608721
transform 1 0 20056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_218
timestamp 1640608721
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1648_
timestamp 1640608721
transform 1 0 20424 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1650_
timestamp 1640608721
transform 1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__A
timestamp 1640608721
transform 1 0 22908 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1753__A1
timestamp 1640608721
transform 1 0 23092 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_225
timestamp 1640608721
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1640608721
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1470_
timestamp 1640608721
transform 1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1538_
timestamp 1640608721
transform -1 0 21712 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1542_
timestamp 1640608721
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_258
timestamp 1640608721
transform 1 0 24840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_262
timestamp 1640608721
transform 1 0 25208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1835_
timestamp 1640608721
transform 1 0 23276 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_11_272
timestamp 1640608721
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1640608721
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1640608721
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1796_
timestamp 1640608721
transform 1 0 25300 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_289
timestamp 1640608721
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_300
timestamp 1640608721
transform 1 0 28704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_304
timestamp 1640608721
transform 1 0 29072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__and2_2  _1582_
timestamp 1640608721
transform 1 0 27876 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1583_
timestamp 1640608721
transform -1 0 28704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 29072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1640608721
transform -1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1640608721
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1684_
timestamp 1640608721
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1804_
timestamp 1640608721
transform 1 0 1656 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_12_38
timestamp 1640608721
transform 1 0 4600 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1640608721
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_2  _1231_
timestamp 1640608721
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _1520_
timestamp 1640608721
transform 1 0 3220 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_12_50
timestamp 1640608721
transform 1 0 5704 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_62
timestamp 1640608721
transform 1 0 6808 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1594_
timestamp 1640608721
transform 1 0 6992 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_12_69
timestamp 1640608721
transform 1 0 7452 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_73
timestamp 1640608721
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1640608721
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1640608721
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1640608721
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1588_
timestamp 1640608721
transform 1 0 7544 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1640608721
transform 1 0 10028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_2  _1204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 11040 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1803_
timestamp 1640608721
transform 1 0 10212 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_116
timestamp 1640608721
transform 1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1897_
timestamp 1640608721
transform 1 0 11960 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1640608721
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1640608721
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1640608721
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1819_
timestamp 1640608721
transform -1 0 15640 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 1640608721
transform 1 0 16744 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_2  _1654_
timestamp 1640608721
transform 1 0 15640 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1721_
timestamp 1640608721
transform 1 0 17020 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1640608721
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1640608721
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_2  _1651_
timestamp 1640608721
transform -1 0 19136 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A
timestamp 1640608721
transform 1 0 20056 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_208
timestamp 1640608721
transform 1 0 20240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_212
timestamp 1640608721
transform 1 0 20608 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1705_
timestamp 1640608721
transform 1 0 20700 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1759_
timestamp 1640608721
transform 1 0 19228 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_234
timestamp 1640608721
transform 1 0 22632 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1469_
timestamp 1640608721
transform 1 0 22356 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1557_
timestamp 1640608721
transform 1 0 22724 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1753_
timestamp 1640608721
transform 1 0 21528 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1640608721
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1640608721
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_257
timestamp 1640608721
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1640608721
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1799_
timestamp 1640608721
transform 1 0 23276 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1838_
timestamp 1640608721
transform 1 0 24840 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_12_282
timestamp 1640608721
transform 1 0 27048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1571_
timestamp 1640608721
transform 1 0 26404 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1576_
timestamp 1640608721
transform 1 0 27140 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_12_290
timestamp 1640608721
transform 1 0 27784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_300
timestamp 1640608721
transform 1 0 28704 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1795_
timestamp 1640608721
transform 1 0 27876 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1640608721
transform -1 0 29532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1734_
timestamp 1640608721
transform 1 0 1840 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _1683_
timestamp 1640608721
transform -1 0 2300 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1640608721
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1640608721
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1640608721
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1640608721
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1640608721
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1232_
timestamp 1640608721
transform -1 0 3680 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_14_17
timestamp 1640608721
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_13
timestamp 1640608721
transform 1 0 2300 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_25
timestamp 1640608721
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_31
timestamp 1640608721
transform 1 0 3956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1640608721
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1219_
timestamp 1640608721
transform 1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1711_
timestamp 1640608721
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1717_
timestamp 1640608721
transform 1 0 4600 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1806_
timestamp 1640608721
transform 1 0 4692 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1640608721
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_63
timestamp 1640608721
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_56
timestamp 1640608721
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1640608721
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1599_
timestamp 1640608721
transform -1 0 7268 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1735_
timestamp 1640608721
transform 1 0 5428 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1859_
timestamp 1640608721
transform 1 0 6440 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 6900 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_67
timestamp 1640608721
transform 1 0 7268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_75
timestamp 1640608721
transform 1 0 8004 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_80
timestamp 1640608721
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1640608721
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1640608721
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1456_
timestamp 1640608721
transform -1 0 8464 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1614_
timestamp 1640608721
transform 1 0 8188 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1940_
timestamp 1640608721
transform 1 0 8924 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_13_103
timestamp 1640608721
transform 1 0 10580 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_108
timestamp 1640608721
transform 1 0 11040 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_92
timestamp 1640608721
transform 1 0 9568 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1640608721
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1120_
timestamp 1640608721
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1128_
timestamp 1640608721
transform 1 0 10304 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1129_
timestamp 1640608721
transform 1 0 10488 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_clk_i
timestamp 1640608721
transform -1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1203_
timestamp 1640608721
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1640608721
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_113
timestamp 1640608721
transform 1 0 11500 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A
timestamp 1640608721
transform 1 0 11316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _1270_
timestamp 1640608721
transform -1 0 12512 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1640608721
transform -1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1118_
timestamp 1640608721
transform 1 0 12512 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_14_121
timestamp 1640608721
transform 1 0 12236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_131
timestamp 1640608721
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_127
timestamp 1640608721
transform 1 0 12788 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1282_
timestamp 1640608721
transform 1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1640608721
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1640608721
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_135
timestamp 1640608721
transform 1 0 13524 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A
timestamp 1640608721
transform 1 0 13800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1281_
timestamp 1640608721
transform -1 0 14720 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1640608721
transform -1 0 15088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_152
timestamp 1640608721
transform 1 0 15088 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_148
timestamp 1640608721
transform 1 0 14720 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1820_
timestamp 1640608721
transform -1 0 15640 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1640608721
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1640608721
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_158
timestamp 1640608721
transform 1 0 15640 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_173
timestamp 1640608721
transform 1 0 17020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1640608721
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1280_
timestamp 1640608721
transform 1 0 16744 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1652_
timestamp 1640608721
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1653_
timestamp 1640608721
transform -1 0 15916 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1722_
timestamp 1640608721
transform 1 0 15916 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _1642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 17204 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1287_
timestamp 1640608721
transform 1 0 17756 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1643_
timestamp 1640608721
transform -1 0 18492 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1283_
timestamp 1640608721
transform 1 0 18216 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_185
timestamp 1640608721
transform 1 0 18124 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1317_
timestamp 1640608721
transform 1 0 18860 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1316_
timestamp 1640608721
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_192
timestamp 1640608721
transform 1 0 18768 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_189
timestamp 1640608721
transform 1 0 18492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1640608721
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_198
timestamp 1640608721
transform 1 0 19320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1640608721
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_208
timestamp 1640608721
transform 1 0 20240 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1284_
timestamp 1640608721
transform 1 0 19320 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1288_
timestamp 1640608721
transform 1 0 19412 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1311_
timestamp 1640608721
transform 1 0 19596 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1646_
timestamp 1640608721
transform 1 0 19872 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_2  _1649_
timestamp 1640608721
transform 1 0 20148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1704_
timestamp 1640608721
transform 1 0 21804 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1645_
timestamp 1640608721
transform 1 0 21344 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1315_
timestamp 1640608721
transform 1 0 21988 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1640608721
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_223
timestamp 1640608721
transform 1 0 21620 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1640608721
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1640608721
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1562_
timestamp 1640608721
transform 1 0 22724 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_240
timestamp 1640608721
transform 1 0 23184 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_234
timestamp 1640608721
transform 1 0 22632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1557__A
timestamp 1640608721
transform -1 0 23184 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_237
timestamp 1640608721
transform 1 0 22908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_246
timestamp 1640608721
transform 1 0 23736 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_258
timestamp 1640608721
transform 1 0 24840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1640608721
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_259
timestamp 1640608721
transform 1 0 24932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1640608721
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1558_
timestamp 1640608721
transform 1 0 23460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1568_
timestamp 1640608721
transform -1 0 24932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_274
timestamp 1640608721
transform 1 0 26312 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_281
timestamp 1640608721
transform 1 0 26956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1640608721
transform 1 0 26036 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_282
timestamp 1640608721
transform 1 0 27048 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1640608721
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1294_
timestamp 1640608721
transform -1 0 27048 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1570_
timestamp 1640608721
transform 1 0 26404 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1572_
timestamp 1640608721
transform -1 0 26312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1573_
timestamp 1640608721
transform -1 0 26036 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_13_287
timestamp 1640608721
transform 1 0 27508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_288
timestamp 1640608721
transform 1 0 27600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_298
timestamp 1640608721
transform 1 0 28520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1574_
timestamp 1640608721
transform -1 0 27508 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1577_
timestamp 1640608721
transform 1 0 27692 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1578_
timestamp 1640608721
transform 1 0 28244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1839_
timestamp 1640608721
transform 1 0 27692 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1640608721
transform -1 0 29532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1640608721
transform -1 0 29532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1640608721
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1640608721
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1686_
timestamp 1640608721
transform 1 0 1472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1805_
timestamp 1640608721
transform 1 0 1748 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_15_24
timestamp 1640608721
transform 1 0 3312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_30
timestamp 1640608721
transform 1 0 3864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_34
timestamp 1640608721
transform 1 0 4232 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_42
timestamp 1640608721
transform 1 0 4968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1233_
timestamp 1640608721
transform 1 0 3956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1640608721
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_60
timestamp 1640608721
transform 1 0 6624 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1640608721
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1245_
timestamp 1640608721
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1687_
timestamp 1640608721
transform 1 0 5244 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__B1
timestamp 1640608721
transform -1 0 9108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_68
timestamp 1640608721
transform 1 0 7360 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_78
timestamp 1640608721
transform 1 0 8280 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_84
timestamp 1640608721
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o311a_2  _1130_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 9108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1246_
timestamp 1640608721
transform -1 0 8280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1248_
timestamp 1640608721
transform -1 0 8004 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _1117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 11408 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _1121_
timestamp 1640608721
transform 1 0 9936 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_123
timestamp 1640608721
transform 1 0 12420 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_129
timestamp 1640608721
transform 1 0 12972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1640608721
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1115_
timestamp 1640608721
transform -1 0 11960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1126_
timestamp 1640608721
transform -1 0 13340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1133_
timestamp 1640608721
transform 1 0 11960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_15_133
timestamp 1640608721
transform 1 0 13340 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1640608721
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1640608721
transform -1 0 14904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1029_
timestamp 1640608721
transform 1 0 14904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1640608721
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1640608721
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1640608721
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1640608721
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1278_
timestamp 1640608721
transform 1 0 15180 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1279_
timestamp 1640608721
transform 1 0 15640 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_184
timestamp 1640608721
transform 1 0 18032 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_191
timestamp 1640608721
transform 1 0 18676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1277_
timestamp 1640608721
transform 1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1503_
timestamp 1640608721
transform -1 0 18676 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1720_
timestamp 1640608721
transform -1 0 18032 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_197
timestamp 1640608721
transform 1 0 19228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_202
timestamp 1640608721
transform 1 0 19688 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_214
timestamp 1640608721
transform 1 0 20792 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__o31a_2  _1314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 21712 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_clk_i
timestamp 1640608721
transform -1 0 19688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 1640608721
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_229
timestamp 1640608721
transform 1 0 22172 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1640608721
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1896_
timestamp 1640608721
transform 1 0 22264 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_15_247
timestamp 1640608721
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_251
timestamp 1640608721
transform 1 0 24196 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1567_
timestamp 1640608721
transform -1 0 25392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1797_
timestamp 1640608721
transform 1 0 24288 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1640608721
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1640608721
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1640608721
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1559_
timestamp 1640608721
transform -1 0 26772 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1560_
timestamp 1640608721
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1566_
timestamp 1640608721
transform 1 0 25576 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_292
timestamp 1640608721
transform 1 0 27968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_304
timestamp 1640608721
transform 1 0 29072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1564_
timestamp 1640608721
transform -1 0 27968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1640608721
transform -1 0 29532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_13
timestamp 1640608721
transform 1 0 2300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1640608721
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1640608721
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1685_
timestamp 1640608721
transform -1 0 2300 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1640608721
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1640608721
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_41
timestamp 1640608721
transform 1 0 4876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1640608721
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1723_
timestamp 1640608721
transform -1 0 5796 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_59
timestamp 1640608721
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_65
timestamp 1640608721
transform 1 0 7084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1433_
timestamp 1640608721
transform -1 0 7084 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1688_
timestamp 1640608721
transform 1 0 5796 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B
timestamp 1640608721
transform 1 0 8556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__C
timestamp 1640608721
transform -1 0 8556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1640608721
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1640608721
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1640608721
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1047_
timestamp 1640608721
transform -1 0 9476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 8372 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1519_
timestamp 1640608721
transform -1 0 7452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A
timestamp 1640608721
transform -1 0 9936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A2
timestamp 1640608721
transform -1 0 10304 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__B2
timestamp 1640608721
transform -1 0 10120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_103
timestamp 1640608721
transform 1 0 10580 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1111_
timestamp 1640608721
transform 1 0 10304 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1640608721
transform 1 0 9476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1116_
timestamp 1640608721
transform -1 0 11316 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_2  _1134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 12144 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1939_
timestamp 1640608721
transform -1 0 13708 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A
timestamp 1640608721
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_143
timestamp 1640608721
transform 1 0 14260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1640608721
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0903_
timestamp 1640608721
transform 1 0 14628 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1046_
timestamp 1640608721
transform 1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1125_
timestamp 1640608721
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_164
timestamp 1640608721
transform 1 0 16192 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_168
timestamp 1640608721
transform 1 0 16560 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__and3_2  _1030_
timestamp 1640608721
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1275_
timestamp 1640608721
transform 1 0 15732 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1276_
timestamp 1640608721
transform 1 0 16284 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1818_
timestamp 1640608721
transform -1 0 18216 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_16_186
timestamp 1640608721
transform 1 0 18216 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1640608721
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1640608721
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_205
timestamp 1640608721
transform 1 0 19964 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_209
timestamp 1640608721
transform 1 0 20332 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1322_
timestamp 1640608721
transform -1 0 20332 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1326_
timestamp 1640608721
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1644_
timestamp 1640608721
transform 1 0 20884 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_222
timestamp 1640608721
transform 1 0 21528 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_233
timestamp 1640608721
transform 1 0 22540 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_239
timestamp 1640608721
transform 1 0 23092 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1271_
timestamp 1640608721
transform -1 0 23092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1274_
timestamp 1640608721
transform 1 0 22264 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1640608721
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1569_
timestamp 1640608721
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1837_
timestamp 1640608721
transform 1 0 24380 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_clk_i
timestamp 1640608721
transform -1 0 24012 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_270
timestamp 1640608721
transform 1 0 25944 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_276
timestamp 1640608721
transform 1 0 26496 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_280
timestamp 1640608721
transform 1 0 26864 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1561_
timestamp 1640608721
transform 1 0 26956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1565_
timestamp 1640608721
transform -1 0 26496 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_16_299
timestamp 1640608721
transform 1 0 28612 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_305
timestamp 1640608721
transform 1 0 29164 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1563_
timestamp 1640608721
transform 1 0 28060 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1798_
timestamp 1640608721
transform 1 0 27232 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1640608721
transform -1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp 1640608721
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1640608721
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1640608721
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1682_
timestamp 1640608721
transform 1 0 4876 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _1689_
timestamp 1640608721
transform 1 0 3220 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1719_
timestamp 1640608721
transform 1 0 4048 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1640608721
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1680_
timestamp 1640608721
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1870_
timestamp 1640608721
transform 1 0 6348 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_17_84
timestamp 1640608721
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1048_
timestamp 1640608721
transform 1 0 8924 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1234_
timestamp 1640608721
transform -1 0 8832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1247_
timestamp 1640608721
transform 1 0 8280 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clk_i
timestamp 1640608721
transform -1 0 8280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1640608721
transform 1 0 9568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_i_A
timestamp 1640608721
transform -1 0 9936 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_i_A
timestamp 1640608721
transform -1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1122_
timestamp 1640608721
transform 1 0 9936 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1123_
timestamp 1640608721
transform 1 0 10764 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clk_i
timestamp 1640608721
transform 1 0 10396 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1640608721
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1640608721
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_126
timestamp 1640608721
transform 1 0 12696 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1640608721
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1113_
timestamp 1640608721
transform -1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1640608721
transform 1 0 12420 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1135_
timestamp 1640608721
transform 1 0 11960 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_17_132
timestamp 1640608721
transform 1 0 13248 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_138
timestamp 1640608721
transform 1 0 13800 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_150
timestamp 1640608721
transform 1 0 14904 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1432_
timestamp 1640608721
transform -1 0 13800 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1640608721
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1640608721
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1640608721
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_174
timestamp 1640608721
transform 1 0 17112 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1640608721
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1022_
timestamp 1640608721
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1031_
timestamp 1640608721
transform -1 0 15732 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1640608721
transform -1 0 15456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_186
timestamp 1640608721
transform 1 0 18216 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1893_
timestamp 1640608721
transform 1 0 18400 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_17_205
timestamp 1640608721
transform 1 0 19964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1273_
timestamp 1640608721
transform 1 0 20884 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1323_
timestamp 1640608721
transform -1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1640608721
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1640608721
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_240
timestamp 1640608721
transform 1 0 23184 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1640608721
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1312_
timestamp 1640608721
transform -1 0 21620 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1313_
timestamp 1640608721
transform 1 0 22632 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _1319_
timestamp 1640608721
transform 1 0 21896 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_252
timestamp 1640608721
transform 1 0 24288 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_264
timestamp 1640608721
transform 1 0 25392 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1640608721
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1640608721
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1836_
timestamp 1640608721
transform 1 0 26956 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_17_298
timestamp 1640608721
transform 1 0 28520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1640608721
transform -1 0 29532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1640608721
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1640608721
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1807_
timestamp 1640608721
transform 1 0 1564 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1640608721
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_38
timestamp 1640608721
transform 1 0 4600 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1640608721
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1736_
timestamp 1640608721
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_44
timestamp 1640608721
transform 1 0 5152 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_54
timestamp 1640608721
transform 1 0 6072 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1710_
timestamp 1640608721
transform -1 0 6072 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_66
timestamp 1640608721
transform 1 0 7176 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1640608721
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1903_
timestamp 1640608721
transform 1 0 7268 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 9660 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_2  _1127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 9660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1136_
timestamp 1640608721
transform -1 0 11224 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_18_110
timestamp 1640608721
transform 1 0 11224 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_125
timestamp 1640608721
transform 1 0 12604 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1640608721
transform 1 0 12328 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1640608721
transform 1 0 12052 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1131_
timestamp 1640608721
transform 1 0 11776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_133
timestamp 1640608721
transform 1 0 13340 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1640608721
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_151
timestamp 1640608721
transform 1 0 14996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1640608721
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1038_
timestamp 1640608721
transform -1 0 13984 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_2  _1051_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 14168 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1439_
timestamp 1640608721
transform 1 0 13432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_160
timestamp 1640608721
transform 1 0 15824 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_166
timestamp 1640608721
transform 1 0 16376 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_170
timestamp 1640608721
transform 1 0 16744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1640608721
transform -1 0 16744 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1443_
timestamp 1640608721
transform 1 0 15548 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1950_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 16836 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_18_192
timestamp 1640608721
transform 1 0 18768 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1640608721
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1325_
timestamp 1640608721
transform -1 0 19136 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_i_A
timestamp 1640608721
transform 1 0 19504 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1318_
timestamp 1640608721
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1321_
timestamp 1640608721
transform -1 0 21252 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1324_
timestamp 1640608721
transform 1 0 20056 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clk_i
timestamp 1640608721
transform -1 0 20056 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1640608721
transform 1 0 21252 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o22ai_2  _1320_
timestamp 1640608721
transform 1 0 21344 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_2  _1895_
timestamp 1640608721
transform -1 0 23828 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1640608721
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1640608721
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1640608721
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_257
timestamp 1640608721
transform 1 0 24748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1640608721
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1015_
timestamp 1640608721
transform 1 0 24840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1016_
timestamp 1640608721
transform 1 0 25116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_264
timestamp 1640608721
transform 1 0 25392 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1640608721
transform 1 0 26496 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_288
timestamp 1640608721
transform 1 0 27600 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_300
timestamp 1640608721
transform 1 0 28704 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1640608721
transform -1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_11
timestamp 1640608721
transform 1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1640608721
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1640608721
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1640608721
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1466_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 3404 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _1467_
timestamp 1640608721
transform 1 0 2392 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1851_
timestamp 1640608721
transform -1 0 2944 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_1  _1243_
timestamp 1640608721
transform -1 0 3772 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _1236_
timestamp 1640608721
transform 1 0 3864 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1209_
timestamp 1640608721
transform -1 0 3680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1640608721
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1640608721
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_29
timestamp 1640608721
transform 1 0 3772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_23
timestamp 1640608721
transform 1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _1681_
timestamp 1640608721
transform -1 0 5612 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1235_
timestamp 1640608721
transform -1 0 4784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1217_
timestamp 1640608721
transform -1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1740_
timestamp 1640608721
transform 1 0 4968 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1640608721
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1640608721
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_61
timestamp 1640608721
transform 1 0 6716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1640608721
transform 1 0 5612 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1640608721
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1731_
timestamp 1640608721
transform -1 0 6624 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1810_
timestamp 1640608721
transform 1 0 6624 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_clk_i
timestamp 1640608721
transform -1 0 6716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_73
timestamp 1640608721
transform 1 0 7820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_85
timestamp 1640608721
transform 1 0 8924 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_77
timestamp 1640608721
transform 1 0 8188 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1640608721
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1640608721
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1640608721
transform -1 0 9200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1207_
timestamp 1640608721
transform 1 0 8280 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1640608721
transform -1 0 9384 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1640608721
transform 1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_102
timestamp 1640608721
transform 1 0 10488 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_90
timestamp 1640608721
transform 1 0 9384 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1941_
timestamp 1640608721
transform 1 0 9844 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1640608721
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_123
timestamp 1640608721
transform 1 0 12420 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_114
timestamp 1640608721
transform 1 0 11592 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1640608721
transform 1 0 12420 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1640608721
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1340_
timestamp 1640608721
transform 1 0 11592 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1483_
timestamp 1640608721
transform 1 0 11868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _1867_
timestamp 1640608721
transform 1 0 12512 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_clk_i
timestamp 1640608721
transform 1 0 12052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1640608721
transform 1 0 14444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_135
timestamp 1640608721
transform 1 0 13524 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1640608721
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1640608721
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1640608721
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1440_
timestamp 1640608721
transform 1 0 13616 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _1865_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 14628 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1640608721
transform 1 0 16928 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_153
timestamp 1640608721
transform 1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_158
timestamp 1640608721
transform 1 0 15640 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1640608721
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_2  _1040_
timestamp 1640608721
transform -1 0 17572 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1444_
timestamp 1640608721
transform -1 0 16928 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1496_
timestamp 1640608721
transform -1 0 15640 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_184
timestamp 1640608721
transform 1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_190
timestamp 1640608721
transform 1 0 18584 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_187
timestamp 1640608721
transform 1 0 18308 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1640608721
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1640608721
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1019_
timestamp 1640608721
transform -1 0 18584 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1039_
timestamp 1640608721
transform -1 0 18032 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1437_
timestamp 1640608721
transform 1 0 18032 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1438_
timestamp 1640608721
transform 1 0 18492 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_198
timestamp 1640608721
transform 1 0 19320 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1640608721
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1640608721
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_209
timestamp 1640608721
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1887_
timestamp 1640608721
transform 1 0 20516 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_2  _1894_
timestamp 1640608721
transform 1 0 19596 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_i_A
timestamp 1640608721
transform 1 0 22724 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 1640608721
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_234
timestamp 1640608721
transform 1 0 22632 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_232
timestamp 1640608721
transform 1 0 22448 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1640608721
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1018_
timestamp 1640608721
transform -1 0 23276 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1272_
timestamp 1640608721
transform 1 0 22356 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clk_i
timestamp 1640608721
transform 1 0 22908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_241
timestamp 1640608721
transform 1 0 23276 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_249
timestamp 1640608721
transform 1 0 24012 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1640608721
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1640608721
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1008_
timestamp 1640608721
transform -1 0 23552 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1011_
timestamp 1640608721
transform 1 0 24748 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1017_
timestamp 1640608721
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1951_
timestamp 1640608721
transform 1 0 24104 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1640608721
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1640608721
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1640608721
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1009_
timestamp 1640608721
transform 1 0 26036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1010_
timestamp 1640608721
transform 1 0 26312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1953_
timestamp 1640608721
transform 1 0 25484 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1640608721
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_305
timestamp 1640608721
transform 1 0 29164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_286
timestamp 1640608721
transform 1 0 27416 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_298
timestamp 1640608721
transform 1 0 28520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1640608721
transform -1 0 29532 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1640608721
transform -1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_15
timestamp 1640608721
transform 1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_21
timestamp 1640608721
transform 1 0 3036 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1640608721
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1640608721
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_25
timestamp 1640608721
transform 1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1210_
timestamp 1640608721
transform 1 0 3680 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1213_
timestamp 1640608721
transform 1 0 4876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _1237_
timestamp 1640608721
transform 1 0 4140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1244_
timestamp 1640608721
transform 1 0 3128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_44
timestamp 1640608721
transform 1 0 5152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1640608721
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1640608721
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1732_
timestamp 1640608721
transform -1 0 6256 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1811_
timestamp 1640608721
transform 1 0 6624 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_21_77
timestamp 1640608721
transform 1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0913_
timestamp 1640608721
transform 1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1020_
timestamp 1640608721
transform 1 0 8372 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _1892_
timestamp 1640608721
transform 1 0 9108 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1640608721
transform 1 0 11040 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1640608721
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1640608721
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_126
timestamp 1640608721
transform 1 0 12696 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1640608721
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_2  _1334_
timestamp 1640608721
transform -1 0 12696 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _1484_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 12788 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_21_134
timestamp 1640608721
transform 1 0 13432 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_140
timestamp 1640608721
transform 1 0 13984 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_144
timestamp 1640608721
transform 1 0 14352 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1062_
timestamp 1640608721
transform 1 0 15088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1333_
timestamp 1640608721
transform -1 0 15088 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1482_
timestamp 1640608721
transform 1 0 14076 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B
timestamp 1640608721
transform 1 0 15732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_158
timestamp 1640608721
transform 1 0 15640 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1640608721
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_172
timestamp 1640608721
transform 1 0 16928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1640608721
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1052_
timestamp 1640608721
transform -1 0 16928 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1066_
timestamp 1640608721
transform 1 0 15916 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1332_
timestamp 1640608721
transform -1 0 15640 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1534_
timestamp 1640608721
transform 1 0 17020 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1868_
timestamp 1640608721
transform 1 0 17756 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1640608721
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1348_
timestamp 1640608721
transform 1 0 20056 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1349_
timestamp 1640608721
transform 1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1360_
timestamp 1640608721
transform -1 0 21068 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__A1
timestamp 1640608721
transform 1 0 21344 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1640608721
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1640608721
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_229
timestamp 1640608721
transform 1 0 22172 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1640608721
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1952_
timestamp 1640608721
transform -1 0 24196 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_21_254
timestamp 1640608721
transform 1 0 24472 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1013_
timestamp 1640608721
transform -1 0 24472 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_266
timestamp 1640608721
transform 1 0 25576 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_274
timestamp 1640608721
transform 1 0 26312 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1640608721
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1640608721
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1640608721
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1003_
timestamp 1640608721
transform 1 0 26404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1957_
timestamp 1640608721
transform 1 0 27324 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1640608721
transform -1 0 29532 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_11
timestamp 1640608721
transform 1 0 2116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_19
timestamp 1640608721
transform 1 0 2852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1640608721
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1640608721
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1640608721
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1260_
timestamp 1640608721
transform -1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1640608721
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1640608721
transform 1 0 4048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1640608721
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1211_
timestamp 1640608721
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1255_
timestamp 1640608721
transform 1 0 3128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_44
timestamp 1640608721
transform 1 0 5152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_48
timestamp 1640608721
transform 1 0 5520 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1640608721
transform 1 0 6072 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1679_
timestamp 1640608721
transform 1 0 5612 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_22_66
timestamp 1640608721
transform 1 0 7176 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_74
timestamp 1640608721
transform 1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1640608721
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1640608721
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1640608721
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _1208_
timestamp 1640608721
transform -1 0 8648 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1640608721
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1640608721
transform 1 0 10212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1328_
timestamp 1640608721
transform 1 0 9936 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1335_
timestamp 1640608721
transform -1 0 13340 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _1336_
timestamp 1640608721
transform 1 0 12236 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_2  _1337_
timestamp 1640608721
transform 1 0 11316 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1640608721
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_147
timestamp 1640608721
transform 1 0 14628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_151
timestamp 1640608721
transform 1 0 14996 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1640608721
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1053_
timestamp 1640608721
transform -1 0 14628 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1640608721
transform -1 0 13616 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1495_
timestamp 1640608721
transform -1 0 15548 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_22_174
timestamp 1640608721
transform 1 0 17112 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _1068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 16376 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _1069_
timestamp 1640608721
transform 1 0 15548 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_183
timestamp 1640608721
transform 1 0 17940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1640608721
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1640608721
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1640608721
transform -1 0 17940 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1533_
timestamp 1640608721
transform -1 0 17664 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_22_204
timestamp 1640608721
transform 1 0 19872 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_210
timestamp 1640608721
transform 1 0 20424 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1640608721
transform 1 0 21160 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__or3b_2  _1346_
timestamp 1640608721
transform -1 0 19872 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1347_
timestamp 1640608721
transform 1 0 20148 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A1
timestamp 1640608721
transform -1 0 23184 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_223
timestamp 1640608721
transform 1 0 21620 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_235
timestamp 1640608721
transform 1 0 22724 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1012_
timestamp 1640608721
transform 1 0 23184 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1359_
timestamp 1640608721
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_243
timestamp 1640608721
transform 1 0 23460 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1640608721
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1007_
timestamp 1640608721
transform 1 0 24748 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1014_
timestamp 1640608721
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_clk_i
timestamp 1640608721
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1954_
timestamp 1640608721
transform 1 0 25484 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_22_286
timestamp 1640608721
transform 1 0 27416 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_295
timestamp 1640608721
transform 1 0 28244 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_299
timestamp 1640608721
transform 1 0 28612 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_305
timestamp 1640608721
transform 1 0 29164 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0994_
timestamp 1640608721
transform 1 0 27968 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0995_
timestamp 1640608721
transform 1 0 28336 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1640608721
transform -1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1640608721
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1257_
timestamp 1640608721
transform 1 0 2944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1901_
timestamp 1640608721
transform 1 0 1380 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_23_28
timestamp 1640608721
transform 1 0 3680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_36
timestamp 1640608721
transform 1 0 4416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_42
timestamp 1640608721
transform 1 0 4968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1216_
timestamp 1640608721
transform -1 0 4968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1253_
timestamp 1640608721
transform 1 0 3864 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1640608721
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1640608721
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1640608721
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1251_
timestamp 1640608721
transform 1 0 5704 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1465_
timestamp 1640608721
transform -1 0 5704 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _1891_
timestamp 1640608721
transform 1 0 7452 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1640608721
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_90
timestamp 1640608721
transform 1 0 9384 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_96
timestamp 1640608721
transform 1 0 9936 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1327_
timestamp 1640608721
transform 1 0 9660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1436_
timestamp 1640608721
transform 1 0 10488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1442_
timestamp 1640608721
transform 1 0 10764 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1640608721
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1640608721
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1063_
timestamp 1640608721
transform -1 0 13432 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1330_
timestamp 1640608721
transform -1 0 13156 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_2  _1341_
timestamp 1640608721
transform 1 0 12052 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_2  _1064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 14536 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o2111ai_2  _1071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 13432 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1640608721
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1640608721
transform 1 0 16928 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1640608721
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1640608721
transform -1 0 16928 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_2  _1070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 16376 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A
timestamp 1640608721
transform -1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1640608721
transform 1 0 18032 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1344_
timestamp 1640608721
transform 1 0 18952 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__A1
timestamp 1640608721
transform -1 0 19412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_202
timestamp 1640608721
transform 1 0 19688 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_207
timestamp 1640608721
transform 1 0 20148 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_216
timestamp 1640608721
transform 1 0 20976 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1345_
timestamp 1640608721
transform 1 0 19412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1350_
timestamp 1640608721
transform 1 0 20240 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1358_
timestamp 1640608721
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_clk_i
timestamp 1640608721
transform 1 0 19780 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A1
timestamp 1640608721
transform -1 0 21712 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_220
timestamp 1640608721
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_236
timestamp 1640608721
transform 1 0 22816 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1640608721
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1352_
timestamp 1640608721
transform 1 0 22540 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1354_
timestamp 1640608721
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_248
timestamp 1640608721
transform 1 0 23920 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_261
timestamp 1640608721
transform 1 0 25116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1640608721
transform 1 0 24288 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1005_
timestamp 1640608721
transform 1 0 24564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1006_
timestamp 1640608721
transform -1 0 25116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_269
timestamp 1640608721
transform 1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_275
timestamp 1640608721
transform 1 0 26404 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1640608721
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1640608721
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1640608721
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0993_
timestamp 1640608721
transform 1 0 26128 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1004_
timestamp 1640608721
transform 1 0 26496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1640608721
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_305
timestamp 1640608721
transform 1 0 29164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1640608721
transform -1 0 29532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_15
timestamp 1640608721
transform 1 0 2484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1640608721
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1640608721
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_2  _1259_
timestamp 1640608721
transform 1 0 2576 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1640608721
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1640608721
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_43
timestamp 1640608721
transform 1 0 5060 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1640608721
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1215_
timestamp 1640608721
transform 1 0 4508 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _1252_
timestamp 1640608721
transform 1 0 3864 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1464_
timestamp 1640608721
transform 1 0 5152 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1852_
timestamp 1640608721
transform -1 0 7452 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1640608721
transform 1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_73
timestamp 1640608721
transform 1 0 7820 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1640608721
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1640608721
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1640608721
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1640608721
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1338_
timestamp 1640608721
transform 1 0 9016 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1343_
timestamp 1640608721
transform -1 0 8188 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_92
timestamp 1640608721
transform 1 0 9568 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1339_
timestamp 1640608721
transform -1 0 9568 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1866_
timestamp 1640608721
transform 1 0 9660 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_24_114
timestamp 1640608721
transform 1 0 11592 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_126
timestamp 1640608721
transform 1 0 12696 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1640608721
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_146
timestamp 1640608721
transform 1 0 14536 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1640608721
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1054_
timestamp 1640608721
transform 1 0 14076 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_24_168
timestamp 1640608721
transform 1 0 16560 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1032_
timestamp 1640608721
transform 1 0 15640 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1067_
timestamp 1640608721
transform -1 0 16560 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _1268_
timestamp 1640608721
transform 1 0 17112 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_183
timestamp 1640608721
transform 1 0 17940 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1640608721
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1640608721
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1265_
timestamp 1640608721
transform -1 0 18768 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1266_
timestamp 1640608721
transform -1 0 19044 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1267_
timestamp 1640608721
transform 1 0 18216 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_218
timestamp 1640608721
transform 1 0 21160 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1890_
timestamp 1640608721
transform -1 0 21160 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _1353_
timestamp 1640608721
transform -1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1889_
timestamp 1640608721
transform -1 0 23184 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_24_243
timestamp 1640608721
transform 1 0 23460 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1640608721
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1640608721
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_253
timestamp 1640608721
transform 1 0 24380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_257
timestamp 1640608721
transform 1 0 24748 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1640608721
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0991_
timestamp 1640608721
transform 1 0 24472 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0999_
timestamp 1640608721
transform -1 0 25760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1355_
timestamp 1640608721
transform 1 0 23552 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B1
timestamp 1640608721
transform 1 0 26956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A1
timestamp 1640608721
transform 1 0 25760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_270
timestamp 1640608721
transform 1 0 25944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_280
timestamp 1640608721
transform 1 0 26864 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0996_
timestamp 1640608721
transform 1 0 27140 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0997_
timestamp 1640608721
transform 1 0 26312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0998_
timestamp 1640608721
transform -1 0 26864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_291
timestamp 1640608721
transform 1 0 27876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_296
timestamp 1640608721
transform 1 0 28336 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_300
timestamp 1640608721
transform 1 0 28704 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1000_
timestamp 1640608721
transform 1 0 28060 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1001_
timestamp 1640608721
transform 1 0 28428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1640608721
transform -1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1640608721
transform 1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1640608721
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1640608721
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_2  _1262_
timestamp 1640608721
transform 1 0 2300 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_32
timestamp 1640608721
transform 1 0 4048 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1238_
timestamp 1640608721
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1239_
timestamp 1640608721
transform 1 0 4600 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1256_
timestamp 1640608721
transform -1 0 4048 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1258_
timestamp 1640608721
transform 1 0 4876 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1261_
timestamp 1640608721
transform 1 0 3128 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1640608721
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1640608721
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1640608721
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_72
timestamp 1640608721
transform 1 0 7728 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_2  _1109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 7912 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1110_
timestamp 1640608721
transform -1 0 7728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1342_
timestamp 1640608721
transform 1 0 8740 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1640608721
transform 1 0 10304 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 1640608721
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_92
timestamp 1640608721
transform 1 0 9568 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1441_
timestamp 1640608721
transform 1 0 10488 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1491_
timestamp 1640608721
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1640608721
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1640608721
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1640608721
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1060_
timestamp 1640608721
transform 1 0 12604 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_2  _1493_
timestamp 1640608721
transform 1 0 11776 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_134
timestamp 1640608721
transform 1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__o221ai_2  _1494_
timestamp 1640608721
transform -1 0 15824 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1635_
timestamp 1640608721
transform 1 0 14444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1715_
timestamp 1640608721
transform 1 0 13616 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__B
timestamp 1640608721
transform 1 0 15824 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1640608721
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1034_
timestamp 1640608721
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _1035_
timestamp 1640608721
transform -1 0 17296 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_2  _1898_
timestamp 1640608721
transform 1 0 17296 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__A
timestamp 1640608721
transform 1 0 20240 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_197
timestamp 1640608721
transform 1 0 19228 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_205
timestamp 1640608721
transform 1 0 19964 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_213
timestamp 1640608721
transform 1 0 20700 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1351_
timestamp 1640608721
transform 1 0 20424 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1640608721
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_225
timestamp 1640608721
transform 1 0 21804 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1640608721
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1357_
timestamp 1640608721
transform 1 0 21896 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1888_
timestamp 1640608721
transform 1 0 22632 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_25_258
timestamp 1640608721
transform 1 0 24840 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0989_
timestamp 1640608721
transform 1 0 24564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1956_
timestamp 1640608721
transform 1 0 24932 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_25_281
timestamp 1640608721
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1640608721
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1955_
timestamp 1640608721
transform 1 0 27324 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1640608721
transform -1 0 29532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_15
timestamp 1640608721
transform 1 0 2484 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_21
timestamp 1640608721
transform 1 0 3036 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1640608721
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1640608721
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1640608721
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1214_
timestamp 1640608721
transform 1 0 2944 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1900_
timestamp 1640608721
transform 1 0 1380 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1640608721
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 1640608721
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_43
timestamp 1640608721
transform 1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1640608721
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1250_
timestamp 1640608721
transform 1 0 4784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1254_
timestamp 1640608721
transform 1 0 4048 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1853_
timestamp 1640608721
transform 1 0 4692 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1902_
timestamp 1640608721
transform -1 0 4692 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_26_62
timestamp 1640608721
transform 1 0 6808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1640608721
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1640608721
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1463_
timestamp 1640608721
transform 1 0 5244 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1780_
timestamp 1640608721
transform 1 0 5980 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1942_
timestamp 1640608721
transform 1 0 6900 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1640608721
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_72
timestamp 1640608721
transform 1 0 7728 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_76
timestamp 1640608721
transform 1 0 8096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1640608721
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1640608721
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1107_
timestamp 1640608721
transform 1 0 7452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1108_
timestamp 1640608721
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1861_
timestamp 1640608721
transform 1 0 9016 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1640608721
transform 1 0 9660 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_97
timestamp 1640608721
transform 1 0 10028 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1640608721
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1453_
timestamp 1640608721
transform 1 0 9752 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1502_
timestamp 1640608721
transform -1 0 11500 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o2111a_2  _1501_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 11592 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or3_2  _1492_
timestamp 1640608721
transform 1 0 11500 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1059_
timestamp 1640608721
transform 1 0 12052 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1640608721
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1640608721
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1640608721
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_2  _1487_
timestamp 1640608721
transform 1 0 12788 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1640608721
transform 1 0 12604 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_124
timestamp 1640608721
transform 1 0 12512 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_128
timestamp 1640608721
transform 1 0 12880 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1640608721
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1640608721
transform 1 0 14812 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_139
timestamp 1640608721
transform 1 0 13892 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1640608721
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1640608721
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1074_
timestamp 1640608721
transform -1 0 13892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1331_
timestamp 1640608721
transform -1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1531_
timestamp 1640608721
transform 1 0 14812 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 16836 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_i_A
timestamp 1640608721
transform -1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1640608721
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1640608721
transform 1 0 16928 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1640608721
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _0988_
timestamp 1640608721
transform 1 0 15732 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1640608721
transform 1 0 16192 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1640608721
transform -1 0 17296 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1050_
timestamp 1640608721
transform -1 0 16928 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1640608721
transform 1 0 18584 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_176
timestamp 1640608721
transform 1 0 17296 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1640608721
transform 1 0 18400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1640608721
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1640608721
transform 1 0 18032 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1640608721
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0924_
timestamp 1640608721
transform 1 0 18768 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1971_
timestamp 1640608721
transform -1 0 20056 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_26_200
timestamp 1640608721
transform 1 0 19504 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_204
timestamp 1640608721
transform 1 0 19872 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_209
timestamp 1640608721
transform 1 0 20332 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0920_
timestamp 1640608721
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0921_
timestamp 1640608721
transform 1 0 20424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0923_
timestamp 1640608721
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0925_
timestamp 1640608721
transform -1 0 19504 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1972_
timestamp 1640608721
transform -1 0 21896 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_26_226
timestamp 1640608721
transform 1 0 21896 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_238
timestamp 1640608721
transform 1 0 23000 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1640608721
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1640608721
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1640608721
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1959_
timestamp 1640608721
transform -1 0 23920 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _1356_
timestamp 1640608721
transform 1 0 23644 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0982_
timestamp 1640608721
transform -1 0 24196 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_251
timestamp 1640608721
transform 1 0 24196 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1640608721
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_244
timestamp 1640608721
transform 1 0 23552 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0992_
timestamp 1640608721
transform 1 0 24472 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1640608721
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_253
timestamp 1640608721
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A1
timestamp 1640608721
transform 1 0 25208 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1958_
timestamp 1640608721
transform -1 0 26312 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_26_264
timestamp 1640608721
transform 1 0 25392 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_276
timestamp 1640608721
transform 1 0 26496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_281
timestamp 1640608721
transform 1 0 26956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1640608721
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1640608721
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1002_
timestamp 1640608721
transform 1 0 27140 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1361_
timestamp 1640608721
transform 1 0 26680 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1886_
timestamp 1640608721
transform 1 0 26956 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_26_294
timestamp 1640608721
transform 1 0 28152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_302
timestamp 1640608721
transform 1 0 28888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1362_
timestamp 1640608721
transform 1 0 27876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1640608721
transform -1 0 29532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1640608721
transform -1 0 29532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1640608721
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1264_
timestamp 1640608721
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1899_
timestamp 1640608721
transform 1 0 1380 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_28_37
timestamp 1640608721
transform 1 0 4508 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1640608721
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1241_
timestamp 1640608721
transform -1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1263_
timestamp 1640608721
transform 1 0 3772 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_28_49
timestamp 1640608721
transform 1 0 5612 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_62
timestamp 1640608721
transform 1 0 6808 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1779_
timestamp 1640608721
transform 1 0 5980 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1640608721
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1640608721
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1640608721
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1103_
timestamp 1640608721
transform -1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1105_
timestamp 1640608721
transform 1 0 7728 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1106_
timestamp 1640608721
transform -1 0 7452 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1640608721
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1640608721
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1448_
timestamp 1640608721
transform 1 0 9476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1452_
timestamp 1640608721
transform -1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1485_
timestamp 1640608721
transform 1 0 13064 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1488_
timestamp 1640608721
transform -1 0 13064 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_133
timestamp 1640608721
transform 1 0 13340 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_150
timestamp 1640608721
transform 1 0 14904 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1640608721
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1061_
timestamp 1640608721
transform 1 0 13524 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _1641_
timestamp 1640608721
transform 1 0 14076 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_162
timestamp 1640608721
transform 1 0 16008 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1869_
timestamp 1640608721
transform 1 0 16192 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1640608721
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1640608721
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1435_
timestamp 1640608721
transform -1 0 18400 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1640608721
transform -1 0 20884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A1
timestamp 1640608721
transform -1 0 21068 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A1
timestamp 1640608721
transform -1 0 19964 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1640608721
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_217
timestamp 1640608721
transform 1 0 21068 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0927_
timestamp 1640608721
transform -1 0 20700 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A1
timestamp 1640608721
transform -1 0 22172 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_225
timestamp 1640608721
transform 1 0 21804 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_237
timestamp 1640608721
transform 1 0 22908 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0981_
timestamp 1640608721
transform 1 0 23092 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0983_
timestamp 1640608721
transform 1 0 22172 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A1
timestamp 1640608721
transform 1 0 24932 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1640608721
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1640608721
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_253
timestamp 1640608721
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1640608721
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0974_
timestamp 1640608721
transform 1 0 23368 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0984_
timestamp 1640608721
transform 1 0 24656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0985_
timestamp 1640608721
transform -1 0 25392 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_264
timestamp 1640608721
transform 1 0 25392 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_276
timestamp 1640608721
transform 1 0 26496 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1368_
timestamp 1640608721
transform 1 0 26772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__A1
timestamp 1640608721
transform -1 0 27692 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1640608721
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_301
timestamp 1640608721
transform 1 0 28796 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_305
timestamp 1640608721
transform 1 0 29164 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1640608721
transform -1 0 29532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_11
timestamp 1640608721
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1640608721
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1640608721
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1240_
timestamp 1640608721
transform 1 0 2392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1904_
timestamp 1640608721
transform 1 0 2668 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_29_34
timestamp 1640608721
transform 1 0 4232 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_40
timestamp 1640608721
transform 1 0 4784 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1458_
timestamp 1640608721
transform -1 0 4784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1640608721
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1640608721
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1640608721
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1462_
timestamp 1640608721
transform 1 0 5152 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1943_
timestamp 1640608721
transform 1 0 6624 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_29_81
timestamp 1640608721
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _1863_
timestamp 1640608721
transform 1 0 8924 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_29_106
timestamp 1640608721
transform 1 0 10856 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1500_
timestamp 1640608721
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1640608721
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1640608721
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 1640608721
transform 1 0 12420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_127
timestamp 1640608721
transform 1 0 12788 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1640608721
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1056_
timestamp 1640608721
transform -1 0 13340 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1058_
timestamp 1640608721
transform -1 0 12420 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_133
timestamp 1640608721
transform 1 0 13340 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_139
timestamp 1640608721
transform 1 0 13892 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_145
timestamp 1640608721
transform 1 0 14444 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_151
timestamp 1640608721
transform 1 0 14996 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0904_
timestamp 1640608721
transform 1 0 13984 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1640608721
transform 1 0 14720 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1640608721
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1640608721
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1640608721
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1707_
timestamp 1640608721
transform 1 0 15364 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_183
timestamp 1640608721
transform 1 0 17940 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1426_
timestamp 1640608721
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1434_
timestamp 1640608721
transform 1 0 17664 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1873_
timestamp 1640608721
transform 1 0 18124 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1640608721
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_210
timestamp 1640608721
transform 1 0 20424 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_218
timestamp 1640608721
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _1026_
timestamp 1640608721
transform -1 0 21160 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1640608721
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 1640608721
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1640608721
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0975_
timestamp 1640608721
transform 1 0 23092 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_245
timestamp 1640608721
transform 1 0 23644 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_249
timestamp 1640608721
transform 1 0 24012 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_258
timestamp 1640608721
transform 1 0 24840 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0973_
timestamp 1640608721
transform 1 0 24104 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0976_
timestamp 1640608721
transform -1 0 23644 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1962_
timestamp 1640608721
transform 1 0 24932 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1640608721
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1640608721
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1379_
timestamp 1640608721
transform 1 0 27140 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__A1
timestamp 1640608721
transform 1 0 27876 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1640608721
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_305
timestamp 1640608721
transform 1 0 29164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1640608721
transform -1 0 29532 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_15
timestamp 1640608721
transform 1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_21
timestamp 1640608721
transform 1 0 3036 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1640608721
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1640608721
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_37
timestamp 1640608721
transform 1 0 4508 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1640608721
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1212_
timestamp 1640608721
transform -1 0 3680 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _1242_
timestamp 1640608721
transform -1 0 4508 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1854_
timestamp 1640608721
transform 1 0 4876 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_30_58
timestamp 1640608721
transform 1 0 6440 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_66
timestamp 1640608721
transform 1 0 7176 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_72
timestamp 1640608721
transform 1 0 7728 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1640608721
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1640608721
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1104_
timestamp 1640608721
transform 1 0 7452 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_104
timestamp 1640608721
transform 1 0 10672 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_96
timestamp 1640608721
transform 1 0 9936 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1449_
timestamp 1640608721
transform 1 0 9660 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1537_
timestamp 1640608721
transform 1 0 10764 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_30_122
timestamp 1640608721
transform 1 0 12328 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1329_
timestamp 1640608721
transform 1 0 13064 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1486_
timestamp 1640608721
transform 1 0 11684 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1497_
timestamp 1640608721
transform -1 0 13064 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1640608721
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1640608721
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_150
timestamp 1640608721
transform 1 0 14904 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1640608721
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__and4b_2  _0987_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 14076 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_163
timestamp 1640608721
transform 1 0 16100 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1706_
timestamp 1640608721
transform 1 0 15272 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1872_
timestamp 1640608721
transform -1 0 18400 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_30_191
timestamp 1640608721
transform 1 0 18676 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1640608721
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1640608721
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1423_
timestamp 1640608721
transform 1 0 18400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1424_
timestamp 1640608721
transform 1 0 18768 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 1640608721
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1844_
timestamp 1640608721
transform 1 0 19964 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_30_225
timestamp 1640608721
transform 1 0 21804 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1393_
timestamp 1640608721
transform -1 0 21804 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1961_
timestamp 1640608721
transform 1 0 22080 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1640608721
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_253
timestamp 1640608721
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1640608721
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0972_
timestamp 1640608721
transform -1 0 24748 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0978_
timestamp 1640608721
transform 1 0 24748 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0979_
timestamp 1640608721
transform 1 0 25024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_263
timestamp 1640608721
transform 1 0 25300 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_271
timestamp 1640608721
transform 1 0 26036 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_276
timestamp 1640608721
transform 1 0 26496 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1640608721
transform -1 0 26496 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_284
timestamp 1640608721
transform 1 0 27232 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1883_
timestamp 1640608721
transform 1 0 27324 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1640608721
transform -1 0 29532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1640608721
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1457_
timestamp 1640608721
transform 1 0 2944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1858_
timestamp 1640608721
transform 1 0 1380 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_31_37
timestamp 1640608721
transform 1 0 4508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _1461_
timestamp 1640608721
transform 1 0 4876 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1774_
timestamp 1640608721
transform 1 0 3680 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1640608721
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1640608721
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1640608721
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1778_
timestamp 1640608721
transform 1 0 6348 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A
timestamp 1640608721
transform 1 0 7820 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_66
timestamp 1640608721
transform 1 0 7176 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_75
timestamp 1640608721
transform 1 0 8004 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_87
timestamp 1640608721
transform 1 0 9108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1093_
timestamp 1640608721
transform 1 0 7268 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1094_
timestamp 1640608721
transform 1 0 7544 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_101
timestamp 1640608721
transform 1 0 10396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1640608721
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1445_
timestamp 1640608721
transform 1 0 9568 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1446_
timestamp 1640608721
transform 1 0 9844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1450_
timestamp 1640608721
transform 1 0 9292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1451_
timestamp 1640608721
transform -1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1640608721
transform 1 0 12420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1640608721
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__o22ai_2  _1489_
timestamp 1640608721
transform 1 0 11500 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or3_2  _1498_
timestamp 1640608721
transform -1 0 13340 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_136
timestamp 1640608721
transform 1 0 13616 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_151
timestamp 1640608721
transform 1 0 14996 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0905_
timestamp 1640608721
transform -1 0 14996 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0952_
timestamp 1640608721
transform 1 0 14168 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1402_
timestamp 1640608721
transform 1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_159
timestamp 1640608721
transform 1 0 15732 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1640608721
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1640608721
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1428_
timestamp 1640608721
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1532_
timestamp 1640608721
transform -1 0 16468 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__A1
timestamp 1640608721
transform 1 0 18860 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_177
timestamp 1640608721
transform 1 0 17388 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1640608721
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_195
timestamp 1640608721
transform 1 0 19044 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _1425_
timestamp 1640608721
transform -1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1427_
timestamp 1640608721
transform -1 0 17756 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_207
timestamp 1640608721
transform 1 0 20148 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_215
timestamp 1640608721
transform 1 0 20884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1640608721
transform -1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _1027_
timestamp 1640608721
transform 1 0 20240 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A1
timestamp 1640608721
transform 1 0 22908 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_228
timestamp 1640608721
transform 1 0 22080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_239
timestamp 1640608721
transform 1 0 23092 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1640608721
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0942_
timestamp 1640608721
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0946_
timestamp 1640608721
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0977_
timestamp 1640608721
transform -1 0 22908 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0971_
timestamp 1640608721
transform 1 0 23276 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0980_
timestamp 1640608721
transform 1 0 23552 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1960_
timestamp 1640608721
transform 1 0 24288 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_31_273
timestamp 1640608721
transform 1 0 26220 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1640608721
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1640608721
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1640608721
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0963_
timestamp 1640608721
transform 1 0 27140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1640608721
transform -1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_289
timestamp 1640608721
transform 1 0 27692 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_298
timestamp 1640608721
transform 1 0 28520 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0964_
timestamp 1640608721
transform 1 0 27416 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1378_
timestamp 1640608721
transform 1 0 28244 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1640608721
transform -1 0 29532 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1640608721
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1640608721
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1640608721
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1640608721
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1640608721
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_37
timestamp 1640608721
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1640608721
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1855_
timestamp 1640608721
transform 1 0 4600 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_32_55
timestamp 1640608721
transform 1 0 6164 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_59
timestamp 1640608721
transform 1 0 6532 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1944_
timestamp 1640608721
transform -1 0 8556 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1640608721
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1100_
timestamp 1640608721
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1862_
timestamp 1640608721
transform -1 0 10856 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1640608721
transform 1 0 10856 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_118
timestamp 1640608721
transform 1 0 11960 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_131
timestamp 1640608721
transform 1 0 13156 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_2  _1536_
timestamp 1640608721
transform -1 0 13156 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1640608721
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_144
timestamp 1640608721
transform 1 0 14352 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1640608721
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0951_
timestamp 1640608721
transform 1 0 13432 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1363_
timestamp 1640608721
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1420_
timestamp 1640608721
transform 1 0 14904 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__A1
timestamp 1640608721
transform -1 0 16652 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_164
timestamp 1640608721
transform 1 0 16192 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_169
timestamp 1640608721
transform 1 0 16652 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1419_
timestamp 1640608721
transform 1 0 15916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1638_
timestamp 1640608721
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__A1
timestamp 1640608721
transform 1 0 17572 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_177
timestamp 1640608721
transform 1 0 17388 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1640608721
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1640608721
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1640608721
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1421_
timestamp 1640608721
transform 1 0 17756 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1640608721
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 1640608721
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_212
timestamp 1640608721
transform 1 0 20608 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_218
timestamp 1640608721
transform 1 0 21160 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1480_
timestamp 1640608721
transform 1 0 19872 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_222
timestamp 1640608721
transform 1 0 21528 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_230
timestamp 1640608721
transform 1 0 22264 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_236
timestamp 1640608721
transform 1 0 22816 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0958_
timestamp 1640608721
transform 1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1397_
timestamp 1640608721
transform -1 0 21528 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1640608721
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1640608721
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_257
timestamp 1640608721
transform 1 0 24748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1640608721
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1640608721
transform -1 0 25116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0955_
timestamp 1640608721
transform 1 0 25116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_267
timestamp 1640608721
transform 1 0 25668 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_271
timestamp 1640608721
transform 1 0 26036 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_275
timestamp 1640608721
transform 1 0 26404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0953_
timestamp 1640608721
transform 1 0 25392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0959_
timestamp 1640608721
transform 1 0 26128 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1964_
timestamp 1640608721
transform 1 0 26588 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_32_301
timestamp 1640608721
transform 1 0 28796 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_305
timestamp 1640608721
transform 1 0 29164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1377_
timestamp 1640608721
transform -1 0 28796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1640608721
transform -1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_15
timestamp 1640608721
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1640608721
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1640608721
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1640608721
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1459_
timestamp 1640608721
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 1640608721
transform -1 0 3496 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1857_
timestamp 1640608721
transform 1 0 1380 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_33_34
timestamp 1640608721
transform 1 0 4232 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_42
timestamp 1640608721
transform 1 0 4968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1640608721
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1460_
timestamp 1640608721
transform -1 0 4232 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1856_
timestamp 1640608721
transform 1 0 3772 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_clk_i
timestamp 1640608721
transform -1 0 5520 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1777_
timestamp 1640608721
transform 1 0 5428 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_46
timestamp 1640608721
transform 1 0 5336 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1640608721
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clk_i
timestamp 1640608721
transform -1 0 6900 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1640608721
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_56
timestamp 1640608721
transform 1 0 6256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_65
timestamp 1640608721
transform 1 0 7084 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1640608721
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_i_A
timestamp 1640608721
transform 1 0 6900 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2ai_2  _1098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 6440 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_73
timestamp 1640608721
transform 1 0 7820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_70
timestamp 1640608721
transform 1 0 7544 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1640608721
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1640608721
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0914_
timestamp 1640608721
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1640608721
transform 1 0 8924 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1095_
timestamp 1640608721
transform -1 0 7820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1099_
timestamp 1640608721
transform 1 0 7268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_clk_i
timestamp 1640608721
transform 1 0 10120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1160_
timestamp 1640608721
transform -1 0 9844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0918_
timestamp 1640608721
transform 1 0 9200 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_97
timestamp 1640608721
transform 1 0 10028 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1640608721
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_88
timestamp 1640608721
transform 1 0 9200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_i_A
timestamp 1640608721
transform 1 0 9844 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__A
timestamp 1640608721
transform 1 0 9292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1145_
timestamp 1640608721
transform 1 0 10948 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0919_
timestamp 1640608721
transform -1 0 10764 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_105
timestamp 1640608721
transform 1 0 10764 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1864_
timestamp 1640608721
transform -1 0 11408 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _1447_
timestamp 1640608721
transform -1 0 11500 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1640608721
transform 1 0 11868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1640608721
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_113
timestamp 1640608721
transform 1 0 11500 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_120
timestamp 1640608721
transform 1 0 12144 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1640608721
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1535_
timestamp 1640608721
transform 1 0 12236 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1499_
timestamp 1640608721
transform -1 0 13064 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_130
timestamp 1640608721
transform 1 0 13064 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_2  _1860_
timestamp 1640608721
transform 1 0 12052 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_33_138
timestamp 1640608721
transform 1 0 13800 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_141
timestamp 1640608721
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_149
timestamp 1640608721
transform 1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1640608721
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0906_
timestamp 1640608721
transform 1 0 14076 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1364_
timestamp 1640608721
transform 1 0 14628 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1403_
timestamp 1640608721
transform -1 0 15364 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1637_
timestamp 1640608721
transform 1 0 15088 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__A1
timestamp 1640608721
transform -1 0 16560 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_155
timestamp 1640608721
transform 1 0 15364 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1640608721
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1640608721
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1429_
timestamp 1640608721
transform -1 0 17296 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1431_
timestamp 1640608721
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1871_
timestamp 1640608721
transform 1 0 15824 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_33_176
timestamp 1640608721
transform 1 0 17296 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_181
timestamp 1640608721
transform 1 0 17756 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_185
timestamp 1640608721
transform 1 0 18124 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1640608721
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1640608721
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1418_
timestamp 1640608721
transform -1 0 19044 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1422_
timestamp 1640608721
transform -1 0 18124 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1874_
timestamp 1640608721
transform -1 0 19504 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_clk_i
timestamp 1640608721
transform -1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _1481_
timestamp 1640608721
transform 1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1477_
timestamp 1640608721
transform 1 0 19596 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1471_
timestamp 1640608721
transform -1 0 19504 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1041_
timestamp 1640608721
transform -1 0 19872 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_204
timestamp 1640608721
transform 1 0 19872 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_200
timestamp 1640608721
transform 1 0 19504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_204
timestamp 1640608721
transform 1 0 19872 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_200
timestamp 1640608721
transform 1 0 19504 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1476_
timestamp 1640608721
transform -1 0 20976 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_216
timestamp 1640608721
transform 1 0 20976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1843_
timestamp 1640608721
transform 1 0 20148 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__A1
timestamp 1640608721
transform -1 0 22448 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1640608721
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_235
timestamp 1640608721
transform 1 0 22724 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1640608721
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1369_
timestamp 1640608721
transform -1 0 22264 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1395_
timestamp 1640608721
transform 1 0 22448 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1398_
timestamp 1640608721
transform 1 0 22816 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1879_
timestamp 1640608721
transform -1 0 23644 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_2  _1394_
timestamp 1640608721
transform 1 0 23552 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1382_
timestamp 1640608721
transform 1 0 23644 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1370_
timestamp 1640608721
transform 1 0 23920 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1640608721
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1392_
timestamp 1640608721
transform 1 0 24840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1640608721
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_261
timestamp 1640608721
transform 1 0 25116 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_254
timestamp 1640608721
transform 1 0 24472 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__A1
timestamp 1640608721
transform 1 0 24288 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1880_
timestamp 1640608721
transform -1 0 26312 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _1384_
timestamp 1640608721
transform -1 0 26036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_267
timestamp 1640608721
transform 1 0 25668 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1367_
timestamp 1640608721
transform 1 0 26588 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1366_
timestamp 1640608721
transform -1 0 26588 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1365_
timestamp 1640608721
transform 1 0 26496 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1640608721
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_275
timestamp 1640608721
transform 1 0 26404 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_271
timestamp 1640608721
transform 1 0 26036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0965_
timestamp 1640608721
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1640608721
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_280
timestamp 1640608721
transform 1 0 26864 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A1
timestamp 1640608721
transform 1 0 27692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_291
timestamp 1640608721
transform 1 0 27876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_303
timestamp 1640608721
transform 1 0 28980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_284
timestamp 1640608721
transform 1 0 27232 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_288
timestamp 1640608721
transform 1 0 27600 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_293
timestamp 1640608721
transform 1 0 28060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_305
timestamp 1640608721
transform 1 0 29164 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0966_
timestamp 1640608721
transform 1 0 27324 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0967_
timestamp 1640608721
transform 1 0 27784 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1640608721
transform -1 0 29532 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1640608721
transform -1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_15
timestamp 1640608721
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1640608721
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1640608721
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1776_
timestamp 1640608721
transform -1 0 3864 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_35_30
timestamp 1640608721
transform 1 0 3864 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_39
timestamp 1640608721
transform 1 0 4692 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_2  _1082_
timestamp 1640608721
transform 1 0 4876 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1083_
timestamp 1640608721
transform -1 0 4692 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A
timestamp 1640608721
transform 1 0 5980 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1640608721
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1640608721
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1640608721
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1042_
timestamp 1640608721
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1945_
timestamp 1640608721
transform -1 0 8648 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_35_85
timestamp 1640608721
transform 1 0 8924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1072_
timestamp 1640608721
transform -1 0 8924 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1198_
timestamp 1640608721
transform -1 0 9292 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B1
timestamp 1640608721
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_104
timestamp 1640608721
transform 1 0 10672 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _1175_
timestamp 1640608721
transform 1 0 9844 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clk_i
timestamp 1640608721
transform 1 0 9292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_113
timestamp 1640608721
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_121
timestamp 1640608721
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_129
timestamp 1640608721
transform 1 0 12972 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1640608721
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1454_
timestamp 1640608721
transform 1 0 12420 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1455_
timestamp 1640608721
transform 1 0 12696 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_135
timestamp 1640608721
transform 1 0 13524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_144
timestamp 1640608721
transform 1 0 14352 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_150
timestamp 1640608721
transform 1 0 14904 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1490_
timestamp 1640608721
transform 1 0 13248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1636_
timestamp 1640608721
transform 1 0 14076 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1708_
timestamp 1640608721
transform 1 0 14996 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1640608721
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_169
timestamp 1640608721
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1640608721
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1430_
timestamp 1640608721
transform -1 0 17204 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_175
timestamp 1640608721
transform 1 0 17204 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1640608721
transform 1 0 18308 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1405_
timestamp 1640608721
transform -1 0 18032 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1417_
timestamp 1640608721
transform 1 0 18032 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_202
timestamp 1640608721
transform 1 0 19688 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1640608721
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1468_
timestamp 1640608721
transform -1 0 19688 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1479_
timestamp 1640608721
transform 1 0 20424 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_225
timestamp 1640608721
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_233
timestamp 1640608721
transform 1 0 22540 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_237
timestamp 1640608721
transform 1 0 22908 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1640608721
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1396_
timestamp 1640608721
transform -1 0 22908 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_245
timestamp 1640608721
transform 1 0 23644 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_258
timestamp 1640608721
transform 1 0 24840 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1386_
timestamp 1640608721
transform 1 0 24288 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1391_
timestamp 1640608721
transform 1 0 24564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_clk_i
timestamp 1640608721
transform 1 0 23920 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_266
timestamp 1640608721
transform 1 0 25576 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_281
timestamp 1640608721
transform 1 0 26956 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1640608721
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0960_
timestamp 1640608721
transform 1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0968_
timestamp 1640608721
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1963_
timestamp 1640608721
transform 1 0 27048 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_35_303
timestamp 1640608721
transform 1 0 28980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1640608721
transform -1 0 29532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_14
timestamp 1640608721
transform 1 0 2392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_18
timestamp 1640608721
transform 1 0 2760 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1640608721
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1640608721
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1640608721
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1084_
timestamp 1640608721
transform -1 0 2392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1086_
timestamp 1640608721
transform 1 0 2852 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1087_
timestamp 1640608721
transform -1 0 2116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 1640608721
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1640608721
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1948_
timestamp 1640608721
transform 1 0 3864 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_36_51
timestamp 1640608721
transform 1 0 5796 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1096_
timestamp 1640608721
transform 1 0 6164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_2  _1102_
timestamp 1640608721
transform 1 0 6440 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_70
timestamp 1640608721
transform 1 0 7544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1640608721
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1640608721
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1920_
timestamp 1640608721
transform -1 0 10488 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1921_
timestamp 1640608721
transform 1 0 10488 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_36_128
timestamp 1640608721
transform 1 0 12880 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__a22oi_2  _1101_
timestamp 1640608721
transform 1 0 13064 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1762_
timestamp 1640608721
transform 1 0 12052 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_36_150
timestamp 1640608721
transform 1 0 14904 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1640608721
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1401_
timestamp 1640608721
transform -1 0 15364 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1709_
timestamp 1640608721
transform 1 0 14076 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_36_155
timestamp 1640608721
transform 1 0 15364 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _1876_
timestamp 1640608721
transform 1 0 15456 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1640608721
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1640608721
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1640608721
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1640608721
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_197
timestamp 1640608721
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_203
timestamp 1640608721
transform 1 0 19780 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_215
timestamp 1640608721
transform 1 0 20884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1640608721
transform 1 0 19872 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1478_
timestamp 1640608721
transform 1 0 20148 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1845_
timestamp 1640608721
transform 1 0 21160 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_i_A
timestamp 1640608721
transform -1 0 23276 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clk_i
timestamp 1640608721
transform 1 0 22724 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_241
timestamp 1640608721
transform 1 0 23276 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1640608721
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_256
timestamp 1640608721
transform 1 0 24656 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_262
timestamp 1640608721
transform 1 0 25208 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1640608721
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1387_
timestamp 1640608721
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1390_
timestamp 1640608721
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1965_
timestamp 1640608721
transform -1 0 27232 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_36_284
timestamp 1640608721
transform 1 0 27232 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_296
timestamp 1640608721
transform 1 0 28336 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_304
timestamp 1640608721
transform 1 0 29072 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1640608721
transform -1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1640608721
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1947_
timestamp 1640608721
transform 1 0 1380 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_37_24
timestamp 1640608721
transform 1 0 3312 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_36
timestamp 1640608721
transform 1 0 4416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1080_
timestamp 1640608721
transform 1 0 4692 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1081_
timestamp 1640608721
transform 1 0 4968 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__B1
timestamp 1640608721
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1640608721
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_53
timestamp 1640608721
transform 1 0 5980 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1640608721
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1199_
timestamp 1640608721
transform -1 0 7176 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_37_66
timestamp 1640608721
transform 1 0 7176 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1912_
timestamp 1640608721
transform 1 0 7912 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_37_100
timestamp 1640608721
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _1176_
timestamp 1640608721
transform 1 0 9476 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_130
timestamp 1640608721
transform 1 0 13064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1640608721
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1913_
timestamp 1640608721
transform 1 0 11500 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_37_134
timestamp 1640608721
transform 1 0 13432 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_141
timestamp 1640608721
transform 1 0 14076 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_149
timestamp 1640608721
transform 1 0 14812 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1075_
timestamp 1640608721
transform 1 0 13524 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1077_
timestamp 1640608721
transform -1 0 14076 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1413_
timestamp 1640608721
transform 1 0 14996 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1640608721
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1640608721
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1410_
timestamp 1640608721
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1411_
timestamp 1640608721
transform -1 0 17204 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1639_
timestamp 1640608721
transform 1 0 15732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1640608721
transform 1 0 17204 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_2  _1475_
timestamp 1640608721
transform 1 0 17388 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1847_
timestamp 1640608721
transform 1 0 18124 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_37_212
timestamp 1640608721
transform 1 0 20608 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_2  _1024_
timestamp 1640608721
transform 1 0 19688 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1090_
timestamp 1640608721
transform -1 0 20608 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1640608721
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_235
timestamp 1640608721
transform 1 0 22724 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1640608721
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0937_
timestamp 1640608721
transform 1 0 22448 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1383_
timestamp 1640608721
transform 1 0 22172 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1385_
timestamp 1640608721
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1389_
timestamp 1640608721
transform -1 0 22172 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1881_
timestamp 1640608721
transform 1 0 23644 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1640608721
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1640608721
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1640608721
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0961_
timestamp 1640608721
transform -1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0962_
timestamp 1640608721
transform 1 0 25576 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_296
timestamp 1640608721
transform 1 0 28336 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_300
timestamp 1640608721
transform 1 0 28704 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1374_
timestamp 1640608721
transform 1 0 28060 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1375_
timestamp 1640608721
transform 1 0 28428 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1640608721
transform -1 0 29532 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_11
timestamp 1640608721
transform 1 0 2116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1640608721
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1640608721
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1640608721
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1085_
timestamp 1640608721
transform 1 0 2208 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1088_
timestamp 1640608721
transform 1 0 2484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1089_
timestamp 1640608721
transform -1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__B1
timestamp 1640608721
transform -1 0 4784 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1640608721
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_32
timestamp 1640608721
transform 1 0 4048 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1640608721
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1073_
timestamp 1640608721
transform -1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1185_
timestamp 1640608721
transform -1 0 5612 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_38_49
timestamp 1640608721
transform 1 0 5612 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_54
timestamp 1640608721
transform 1 0 6072 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1907_
timestamp 1640608721
transform 1 0 6164 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_clk_i
timestamp 1640608721
transform -1 0 6072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B1
timestamp 1640608721
transform -1 0 8004 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_72
timestamp 1640608721
transform 1 0 7728 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1640608721
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1640608721
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1190_
timestamp 1640608721
transform 1 0 8004 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__B1
timestamp 1640608721
transform -1 0 9476 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_100
timestamp 1640608721
transform 1 0 10304 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_108
timestamp 1640608721
transform 1 0 11040 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1741_
timestamp 1640608721
transform -1 0 10304 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__B1
timestamp 1640608721
transform -1 0 12236 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1640608721
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _1189_
timestamp 1640608721
transform 1 0 11224 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1640608721
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1640608721
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1640608721
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_2  _1097_
timestamp 1640608721
transform 1 0 14076 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _1416_
timestamp 1640608721
transform 1 0 14996 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__A1
timestamp 1640608721
transform -1 0 15916 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_161
timestamp 1640608721
transform 1 0 15916 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_173
timestamp 1640608721
transform 1 0 17020 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_177
timestamp 1640608721
transform 1 0 17388 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1640608721
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1640608721
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1848_
timestamp 1640608721
transform 1 0 17480 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1640608721
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0922_
timestamp 1640608721
transform 1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1025_
timestamp 1640608721
transform 1 0 20148 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _1065_
timestamp 1640608721
transform 1 0 19504 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1846_
timestamp 1640608721
transform 1 0 20976 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_38_236
timestamp 1640608721
transform 1 0 22816 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0931_
timestamp 1640608721
transform 1 0 22540 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__B1
timestamp 1640608721
transform 1 0 25208 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1640608721
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1640608721
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_258
timestamp 1640608721
transform 1 0 24840 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1640608721
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1388_
timestamp 1640608721
transform 1 0 24564 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A1
timestamp 1640608721
transform -1 0 25576 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_266
timestamp 1640608721
transform 1 0 25576 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_274
timestamp 1640608721
transform 1 0 26312 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1376_
timestamp 1640608721
transform 1 0 26588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1884_
timestamp 1640608721
transform 1 0 27324 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1640608721
transform -1 0 29532 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1640608721
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_11
timestamp 1640608721
transform 1 0 2116 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_18
timestamp 1640608721
transform 1 0 2760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_3
timestamp 1640608721
transform 1 0 1380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1640608721
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1640608721
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1043_
timestamp 1640608721
transform 1 0 2208 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1044_
timestamp 1640608721
transform 1 0 2484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1946_
timestamp 1640608721
transform 1 0 1564 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1640608721
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1640608721
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_41
timestamp 1640608721
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1640608721
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2ai_2  _1092_
timestamp 1640608721
transform 1 0 3496 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1915_
timestamp 1640608721
transform 1 0 4600 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1640608721
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_57
timestamp 1640608721
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_49
timestamp 1640608721
transform 1 0 5612 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_54
timestamp 1640608721
transform 1 0 6072 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1640608721
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1180_
timestamp 1640608721
transform -1 0 6072 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1194_
timestamp 1640608721
transform 1 0 6164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1196_
timestamp 1640608721
transform -1 0 7268 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1701_
timestamp 1640608721
transform -1 0 7728 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_40_69
timestamp 1640608721
transform 1 0 7452 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__B1
timestamp 1640608721
transform -1 0 7452 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _1192_
timestamp 1640608721
transform 1 0 8924 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1187_
timestamp 1640608721
transform 1 0 8464 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1640608721
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1640608721
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_77
timestamp 1640608721
transform 1 0 8188 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_84
timestamp 1640608721
transform 1 0 8832 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__B1
timestamp 1640608721
transform -1 0 8464 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_72
timestamp 1640608721
transform 1 0 7728 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B1
timestamp 1640608721
transform 1 0 10856 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1640608721
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_88
timestamp 1640608721
transform 1 0 9200 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1640608721
transform 1 0 9844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1172_
timestamp 1640608721
transform -1 0 10028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1173_
timestamp 1640608721
transform 1 0 9568 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1174_
timestamp 1640608721
transform 1 0 10028 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1184_
timestamp 1640608721
transform -1 0 9568 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1922_
timestamp 1640608721
transform 1 0 10028 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__B1
timestamp 1640608721
transform 1 0 12328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_124
timestamp 1640608721
transform 1 0 12512 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_131
timestamp 1640608721
transform 1 0 13156 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1640608721
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1188_
timestamp 1640608721
transform 1 0 11500 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1914_
timestamp 1640608721
transform 1 0 11592 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_39_132
timestamp 1640608721
transform 1 0 13248 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_143
timestamp 1640608721
transform 1 0 14260 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_151
timestamp 1640608721
transform 1 0 14996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1640608721
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_2  _1078_
timestamp 1640608721
transform 1 0 14076 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a22oi_2  _1091_
timestamp 1640608721
transform 1 0 13340 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _1640_
timestamp 1640608721
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1875_
timestamp 1640608721
transform -1 0 16560 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_40_163
timestamp 1640608721
transform 1 0 16100 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_170
timestamp 1640608721
transform 1 0 16744 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1640608721
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1406_
timestamp 1640608721
transform 1 0 16468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1414_
timestamp 1640608721
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1415_
timestamp 1640608721
transform -1 0 17204 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1474_
timestamp 1640608721
transform -1 0 18308 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1473_
timestamp 1640608721
transform 1 0 17756 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_178
timestamp 1640608721
transform 1 0 17480 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_175
timestamp 1640608721
transform 1 0 17204 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_clk_i
timestamp 1640608721
transform -1 0 18860 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1412_
timestamp 1640608721
transform -1 0 18584 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_190
timestamp 1640608721
transform 1 0 18584 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1408_
timestamp 1640608721
transform -1 0 19136 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1640608721
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_196
timestamp 1640608721
transform 1 0 19136 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__B1
timestamp 1640608721
transform 1 0 20332 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_i_A
timestamp 1640608721
transform 1 0 20516 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_213
timestamp 1640608721
transform 1 0 20700 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1640608721
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0908_
timestamp 1640608721
transform 1 0 21068 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1640608721
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1472_
timestamp 1640608721
transform 1 0 19228 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1850_
timestamp 1640608721
transform 1 0 19688 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clk_i
timestamp 1640608721
transform -1 0 20332 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1399_
timestamp 1640608721
transform -1 0 22448 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0943_
timestamp 1640608721
transform 1 0 21620 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0907_
timestamp 1640608721
transform -1 0 21528 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1640608721
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_222
timestamp 1640608721
transform 1 0 21528 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1640608721
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1640608721
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_clk_i
timestamp 1640608721
transform -1 0 23368 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_232
timestamp 1640608721
transform 1 0 22448 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _1968_
timestamp 1640608721
transform 1 0 22356 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_39_242
timestamp 1640608721
transform 1 0 23368 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_257
timestamp 1640608721
transform 1 0 24748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1640608721
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1380_
timestamp 1640608721
transform 1 0 24472 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1882_
timestamp 1640608721
transform 1 0 24380 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1966_
timestamp 1640608721
transform 1 0 24932 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__B1
timestamp 1640608721
transform 1 0 27048 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_281
timestamp 1640608721
transform 1 0 26956 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1640608721
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0956_
timestamp 1640608721
transform -1 0 27048 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1373_
timestamp 1640608721
transform 1 0 27048 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_290
timestamp 1640608721
transform 1 0 27784 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_299
timestamp 1640608721
transform 1 0 28612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_305
timestamp 1640608721
transform 1 0 29164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_284
timestamp 1640608721
transform 1 0 27232 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1371_
timestamp 1640608721
transform 1 0 28060 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1372_
timestamp 1640608721
transform 1 0 28336 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1885_
timestamp 1640608721
transform 1 0 27324 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1640608721
transform -1 0 29532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1640608721
transform -1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1640608721
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1640608721
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1949_
timestamp 1640608721
transform 1 0 1748 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_41_40
timestamp 1640608721
transform 1 0 4784 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2ai_2  _1079_
timestamp 1640608721
transform 1 0 3680 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1640608721
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1640608721
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1909_
timestamp 1640608721
transform 1 0 6348 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_41_74
timestamp 1640608721
transform 1 0 7912 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1911_
timestamp 1640608721
transform 1 0 8648 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_41_103
timestamp 1640608721
transform 1 0 10580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_clk_i
timestamp 1640608721
transform 1 0 10212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1640608721
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_113
timestamp 1640608721
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_117
timestamp 1640608721
transform 1 0 11868 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_127
timestamp 1640608721
transform 1 0 12788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1640608721
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1750_
timestamp 1640608721
transform -1 0 12788 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_139
timestamp 1640608721
transform 1 0 13892 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_143
timestamp 1640608721
transform 1 0 14260 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1404_
timestamp 1640608721
transform 1 0 15088 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1409_
timestamp 1640608721
transform 1 0 14352 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp 1640608721
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_172
timestamp 1640608721
transform 1 0 16928 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1640608721
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1407_
timestamp 1640608721
transform -1 0 16928 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_180
timestamp 1640608721
transform 1 0 17664 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1849_
timestamp 1640608721
transform 1 0 17940 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_41_200
timestamp 1640608721
transform 1 0 19504 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_207
timestamp 1640608721
transform 1 0 20148 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1640608721
transform 1 0 20884 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0910_
timestamp 1640608721
transform -1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0916_
timestamp 1640608721
transform 1 0 19872 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1076_
timestamp 1640608721
transform -1 0 19872 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A1
timestamp 1640608721
transform -1 0 22540 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_233
timestamp 1640608721
transform 1 0 22540 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_239
timestamp 1640608721
transform 1 0 23092 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1640608721
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0930_
timestamp 1640608721
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0932_
timestamp 1640608721
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0939_
timestamp 1640608721
transform 1 0 23184 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1400_
timestamp 1640608721
transform -1 0 22356 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_246
timestamp 1640608721
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0940_
timestamp 1640608721
transform 1 0 23460 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0948_
timestamp 1640608721
transform 1 0 24840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1381_
timestamp 1640608721
transform 1 0 25116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_264
timestamp 1640608721
transform 1 0 25392 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_270
timestamp 1640608721
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1640608721
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1640608721
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1640608721
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0949_
timestamp 1640608721
transform 1 0 25668 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1640608721
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_305
timestamp 1640608721
transform 1 0 29164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1640608721
transform -1 0 29532 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1640608721
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1640608721
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1640608721
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1640608721
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_29
timestamp 1640608721
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1640608721
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1917_
timestamp 1640608721
transform 1 0 4140 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_42_50
timestamp 1640608721
transform 1 0 5704 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_55
timestamp 1640608721
transform 1 0 6164 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_59
timestamp 1640608721
transform 1 0 6532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_65
timestamp 1640608721
transform 1 0 7084 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1179_
timestamp 1640608721
transform -1 0 6164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1193_
timestamp 1640608721
transform -1 0 6532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1640608721
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1640608721
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1640608721
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1186_
timestamp 1640608721
transform -1 0 9200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1744_
timestamp 1640608721
transform -1 0 8004 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__B1
timestamp 1640608721
transform 1 0 10764 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_107
timestamp 1640608721
transform 1 0 10948 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_88
timestamp 1640608721
transform 1 0 9200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_92
timestamp 1640608721
transform 1 0 9568 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1171_
timestamp 1640608721
transform 1 0 9660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1178_
timestamp 1640608721
transform 1 0 9936 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_42_119
timestamp 1640608721
transform 1 0 12052 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_125
timestamp 1640608721
transform 1 0 12604 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1751_
timestamp 1640608721
transform -1 0 13524 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1768_
timestamp 1640608721
transform -1 0 12052 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 1640608721
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1640608721
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_150
timestamp 1640608721
transform 1 0 14904 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1640608721
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1752_
timestamp 1640608721
transform -1 0 14904 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _1877_
timestamp 1640608721
transform 1 0 15180 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1878_
timestamp 1640608721
transform 1 0 17112 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1640608721
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1640608721
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1640608721
transform -1 0 19688 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_197
timestamp 1640608721
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_208
timestamp 1640608721
transform 1 0 20240 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0928_
timestamp 1640608721
transform 1 0 19688 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0929_
timestamp 1640608721
transform -1 0 20240 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0933_
timestamp 1640608721
transform -1 0 21528 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1640608721
transform 1 0 21804 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A1
timestamp 1640608721
transform -1 0 23276 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_222
timestamp 1640608721
transform 1 0 21528 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_230
timestamp 1640608721
transform 1 0 22264 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0934_
timestamp 1640608721
transform 1 0 21988 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0935_
timestamp 1640608721
transform 1 0 22540 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0936_
timestamp 1640608721
transform 1 0 22816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_241
timestamp 1640608721
transform 1 0 23276 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1640608721
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_256
timestamp 1640608721
transform 1 0 24656 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1640608721
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0944_
timestamp 1640608721
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_268
timestamp 1640608721
transform 1 0 25760 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_280
timestamp 1640608721
transform 1 0 26864 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_292
timestamp 1640608721
transform 1 0 27968 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_304
timestamp 1640608721
transform 1 0 29072 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1640608721
transform -1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1640608721
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1640608721
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1640608721
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__B1
timestamp 1640608721
transform 1 0 4416 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_27
timestamp 1640608721
transform 1 0 3588 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_35
timestamp 1640608721
transform 1 0 4324 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1182_
timestamp 1640608721
transform -1 0 5428 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__B1
timestamp 1640608721
transform -1 0 5888 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_47
timestamp 1640608721
transform 1 0 5428 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1640608721
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1640608721
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1640608721
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1195_
timestamp 1640608721
transform 1 0 6716 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__B1
timestamp 1640608721
transform 1 0 7544 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_72
timestamp 1640608721
transform 1 0 7728 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_78
timestamp 1640608721
transform 1 0 8280 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1745_
timestamp 1640608721
transform -1 0 9200 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A
timestamp 1640608721
transform 1 0 9476 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_93
timestamp 1640608721
transform 1 0 9660 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1191_
timestamp 1640608721
transform -1 0 9476 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1919_
timestamp 1640608721
transform 1 0 9844 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1640608721
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_126
timestamp 1640608721
transform 1 0 12696 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1640608721
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1763_
timestamp 1640608721
transform -1 0 12696 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_43_134
timestamp 1640608721
transform 1 0 13432 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 1640608721
transform 1 0 13708 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1764_
timestamp 1640608721
transform 1 0 14536 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_43_155
timestamp 1640608721
transform 1 0 15364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1640608721
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1640608721
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1640608721
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__B1
timestamp 1640608721
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_179
timestamp 1640608721
transform 1 0 17572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_191
timestamp 1640608721
transform 1 0 18676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_218
timestamp 1640608721
transform 1 0 21160 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _1970_
timestamp 1640608721
transform -1 0 21160 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_43_233
timestamp 1640608721
transform 1 0 22540 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1640608721
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0938_
timestamp 1640608721
transform -1 0 22540 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0947_
timestamp 1640608721
transform 1 0 22632 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _1967_
timestamp 1640608721
transform 1 0 23368 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_43_263
timestamp 1640608721
transform 1 0 25300 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1640608721
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1640608721
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1640608721
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1640608721
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1640608721
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_305
timestamp 1640608721
transform 1 0 29164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1640608721
transform -1 0 29532 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1640608721
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1640608721
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1640608721
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1640608721
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_29
timestamp 1640608721
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_37
timestamp 1640608721
transform 1 0 4508 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1640608721
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1183_
timestamp 1640608721
transform -1 0 5612 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__B1
timestamp 1640608721
transform -1 0 5796 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_51
timestamp 1640608721
transform 1 0 5796 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_61
timestamp 1640608721
transform 1 0 6716 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1197_
timestamp 1640608721
transform -1 0 6716 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1910_
timestamp 1640608721
transform 1 0 6992 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1640608721
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1640608721
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1640608721
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_102
timestamp 1640608721
transform 1 0 10488 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1640608721
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1170_
timestamp 1640608721
transform -1 0 10488 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1702_
timestamp 1640608721
transform -1 0 10212 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_44_114
timestamp 1640608721
transform 1 0 11592 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1742_
timestamp 1640608721
transform -1 0 13524 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1640608721
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1640608721
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1640608721
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1640608721
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_153
timestamp 1640608721
transform 1 0 15180 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_164
timestamp 1640608721
transform 1 0 16192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _1151_
timestamp 1640608721
transform 1 0 16560 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1743_
timestamp 1640608721
transform -1 0 16192 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1640608721
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1640608721
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1933_
timestamp 1640608721
transform -1 0 18952 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1640608721
transform -1 0 19688 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_202
timestamp 1640608721
transform 1 0 19688 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_214
timestamp 1640608721
transform 1 0 20792 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0915_
timestamp 1640608721
transform -1 0 19504 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_222
timestamp 1640608721
transform 1 0 21528 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _1969_
timestamp 1640608721
transform 1 0 21712 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1640608721
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1640608721
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_256
timestamp 1640608721
transform 1 0 24656 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1640608721
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0945_
timestamp 1640608721
transform -1 0 24656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_268
timestamp 1640608721
transform 1 0 25760 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_280
timestamp 1640608721
transform 1 0 26864 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_292
timestamp 1640608721
transform 1 0 27968 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_304
timestamp 1640608721
transform 1 0 29072 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1640608721
transform -1 0 29532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_15
timestamp 1640608721
transform 1 0 2484 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_21
timestamp 1640608721
transform 1 0 3036 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1640608721
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1640608721
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1908_
timestamp 1640608721
transform 1 0 4692 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1916_
timestamp 1640608721
transform 1 0 3128 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1640608721
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1765_
timestamp 1640608721
transform -1 0 7176 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_45_66
timestamp 1640608721
transform 1 0 7176 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_78
timestamp 1640608721
transform 1 0 8280 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1772_
timestamp 1640608721
transform -1 0 9292 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__B1
timestamp 1640608721
transform -1 0 10212 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_89
timestamp 1640608721
transform 1 0 9292 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_99
timestamp 1640608721
transform 1 0 10212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 1640608721
transform 1 0 9752 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1177_
timestamp 1640608721
transform 1 0 9476 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1640608721
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1640608721
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_126
timestamp 1640608721
transform 1 0 12696 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1640608721
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1769_
timestamp 1640608721
transform -1 0 12696 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_45_138
timestamp 1640608721
transform 1 0 13800 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_149
timestamp 1640608721
transform 1 0 14812 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1770_
timestamp 1640608721
transform 1 0 13984 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1640608721
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1640608721
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_174
timestamp 1640608721
transform 1 0 17112 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1640608721
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1146_
timestamp 1640608721
transform -1 0 17112 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1703_
timestamp 1640608721
transform 1 0 15364 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__B1
timestamp 1640608721
transform -1 0 17572 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_179
timestamp 1640608721
transform 1 0 17572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_191
timestamp 1640608721
transform 1 0 18676 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__B1
timestamp 1640608721
transform 1 0 20792 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_203
timestamp 1640608721
transform 1 0 19780 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0911_
timestamp 1640608721
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0917_
timestamp 1640608721
transform -1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1640608721
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1640608721
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1640608721
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1640608721
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1640608721
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1640608721
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1640608721
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1640608721
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1640608721
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1640608721
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_305
timestamp 1640608721
transform 1 0 29164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1640608721
transform -1 0 29532 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1640608721
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1640608721
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1640608721
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1640608721
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1640608721
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1640608721
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1640608721
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1640608721
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1640608721
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1640608721
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_39
timestamp 1640608721
transform 1 0 4692 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1640608721
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__B1
timestamp 1640608721
transform -1 0 6440 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp 1640608721
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_58
timestamp 1640608721
transform 1 0 6440 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1640608721
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1181_
timestamp 1640608721
transform 1 0 5428 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1918_
timestamp 1640608721
transform 1 0 6348 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_46_66
timestamp 1640608721
transform 1 0 7176 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1640608721
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1640608721
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1640608721
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1165_
timestamp 1640608721
transform -1 0 9752 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1771_
timestamp 1640608721
transform -1 0 8188 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1926_
timestamp 1640608721
transform 1 0 7912 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_1  _1168_
timestamp 1640608721
transform 1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1161_
timestamp 1640608721
transform -1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1138_
timestamp 1640608721
transform 1 0 9844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_91
timestamp 1640608721
transform 1 0 9476 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_94
timestamp 1640608721
transform 1 0 9752 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1766_
timestamp 1640608721
transform -1 0 11040 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _1162_
timestamp 1640608721
transform 1 0 10580 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_99
timestamp 1640608721
transform 1 0 10212 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_98
timestamp 1640608721
transform 1 0 10120 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__B1
timestamp 1640608721
transform -1 0 10580 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1140_
timestamp 1640608721
transform 1 0 11040 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_111
timestamp 1640608721
transform 1 0 11316 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_118
timestamp 1640608721
transform 1 0 11960 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_122
timestamp 1640608721
transform 1 0 12328 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1640608721
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1156_
timestamp 1640608721
transform -1 0 11960 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1159_
timestamp 1640608721
transform 1 0 12420 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1927_
timestamp 1640608721
transform 1 0 11500 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1928_
timestamp 1640608721
transform -1 0 14628 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1773_
timestamp 1640608721
transform -1 0 14904 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1153_
timestamp 1640608721
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1640608721
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_134
timestamp 1640608721
transform 1 0 13432 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__B1
timestamp 1640608721
transform -1 0 13432 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _1154_
timestamp 1640608721
transform 1 0 15088 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1148_
timestamp 1640608721
transform 1 0 14720 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_147
timestamp 1640608721
transform 1 0 14628 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_150
timestamp 1640608721
transform 1 0 14904 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1931_
timestamp 1640608721
transform -1 0 16560 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__B1
timestamp 1640608721
transform 1 0 15916 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_163
timestamp 1640608721
transform 1 0 16100 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_167
timestamp 1640608721
transform 1 0 16468 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1640608721
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1640608721
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1150_
timestamp 1640608721
transform 1 0 16928 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _1152_
timestamp 1640608721
transform 1 0 16560 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1640608721
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1640608721
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1932_
timestamp 1640608721
transform -1 0 18952 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1934_
timestamp 1640608721
transform -1 0 19320 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_47_198
timestamp 1640608721
transform 1 0 19320 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_210
timestamp 1640608721
transform 1 0 20424 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_217
timestamp 1640608721
transform 1 0 21068 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1694_
timestamp 1640608721
transform 1 0 20792 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1973_
timestamp 1640608721
transform -1 0 21160 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1974_
timestamp 1640608721
transform 1 0 21160 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_46_239
timestamp 1640608721
transform 1 0 23092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1640608721
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1640608721
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1640608721
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1695_
timestamp 1640608721
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1640608721
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1640608721
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1640608721
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1640608721
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1640608721
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1640608721
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1640608721
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1640608721
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1640608721
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1640608721
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1640608721
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1640608721
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_301
timestamp 1640608721
transform 1 0 28796 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_305
timestamp 1640608721
transform 1 0 29164 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1640608721
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_305
timestamp 1640608721
transform 1 0 29164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1640608721
transform -1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1640608721
transform -1 0 29532 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1640608721
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1640608721
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1640608721
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1640608721
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1640608721
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1640608721
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1640608721
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1640608721
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1640608721
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1640608721
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1640608721
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1640608721
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1640608721
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__B1
timestamp 1640608721
transform 1 0 11132 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_93
timestamp 1640608721
transform 1 0 9660 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1163_
timestamp 1640608721
transform -1 0 10856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1164_
timestamp 1640608721
transform -1 0 11132 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1167_
timestamp 1640608721
transform -1 0 10580 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_48_111
timestamp 1640608721
transform 1 0 11316 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_126
timestamp 1640608721
transform 1 0 12696 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1155_
timestamp 1640608721
transform -1 0 12696 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1640608721
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1640608721
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1640608721
transform 1 0 14444 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1640608721
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1139_
timestamp 1640608721
transform -1 0 14812 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1141_
timestamp 1640608721
transform -1 0 15088 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1149_
timestamp 1640608721
transform 1 0 15088 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_155
timestamp 1640608721
transform 1 0 15364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_166
timestamp 1640608721
transform 1 0 16376 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1767_
timestamp 1640608721
transform 1 0 15548 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__B1
timestamp 1640608721
transform 1 0 17756 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_178
timestamp 1640608721
transform 1 0 17480 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_183
timestamp 1640608721
transform 1 0 17940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1640608721
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1640608721
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1640608721
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1640608721
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1640608721
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1640608721
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1640608721
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1640608721
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1640608721
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1640608721
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1640608721
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1640608721
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1640608721
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_301
timestamp 1640608721
transform 1 0 28796 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_305
timestamp 1640608721
transform 1 0 29164 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1640608721
transform -1 0 29532 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1640608721
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1640608721
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1640608721
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1640608721
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1640608721
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1640608721
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1640608721
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1640608721
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1640608721
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__B1
timestamp 1640608721
transform 1 0 7728 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_69
timestamp 1640608721
transform 1 0 7452 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_83
timestamp 1640608721
transform 1 0 8740 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _1166_
timestamp 1640608721
transform -1 0 8740 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_49_91
timestamp 1640608721
transform 1 0 9476 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1924_
timestamp 1640608721
transform 1 0 9660 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1640608721
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1640608721
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1640608721
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1930_
timestamp 1640608721
transform 1 0 12236 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__B1
timestamp 1640608721
transform -1 0 14076 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_138
timestamp 1640608721
transform 1 0 13800 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1142_
timestamp 1640608721
transform -1 0 14904 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1937_
timestamp 1640608721
transform -1 0 16468 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1640608721
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1640608721
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1144_
timestamp 1640608721
transform -1 0 17480 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__B1
timestamp 1640608721
transform -1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_180
timestamp 1640608721
transform 1 0 17664 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_192
timestamp 1640608721
transform 1 0 18768 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_204
timestamp 1640608721
transform 1 0 19872 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_216
timestamp 1640608721
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1640608721
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1640608721
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1640608721
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1640608721
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1640608721
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1640608721
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1640608721
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1640608721
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1640608721
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1640608721
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_305
timestamp 1640608721
transform 1 0 29164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1640608721
transform -1 0 29532 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_15
timestamp 1640608721
transform 1 0 2484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_19
timestamp 1640608721
transform 1 0 2852 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1640608721
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1640608721
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1696_
timestamp 1640608721
transform 1 0 2944 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1640608721
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1640608721
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_29
timestamp 1640608721
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_33
timestamp 1640608721
transform 1 0 4140 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_37
timestamp 1640608721
transform 1 0 4508 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1640608721
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1697_
timestamp 1640608721
transform 1 0 4232 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_49
timestamp 1640608721
transform 1 0 5612 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_57
timestamp 1640608721
transform 1 0 6348 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_63
timestamp 1640608721
transform 1 0 6900 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _1698_
timestamp 1640608721
transform 1 0 6624 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1925_
timestamp 1640608721
transform 1 0 7084 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1640608721
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1640608721
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1923_
timestamp 1640608721
transform -1 0 10488 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_50_102
timestamp 1640608721
transform 1 0 10488 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_106
timestamp 1640608721
transform 1 0 10856 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1929_
timestamp 1640608721
transform 1 0 10948 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__o221a_2  _1157_
timestamp 1640608721
transform -1 0 13340 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__B1
timestamp 1640608721
transform 1 0 13340 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_135
timestamp 1640608721
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1640608721
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1640608721
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1938_
timestamp 1640608721
transform -1 0 15640 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_50_158
timestamp 1640608721
transform 1 0 15640 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1936_
timestamp 1640608721
transform -1 0 17480 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1640608721
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1640608721
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1935_
timestamp 1640608721
transform -1 0 19044 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1640608721
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1640608721
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1640608721
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1640608721
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1640608721
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1640608721
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1640608721
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1640608721
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1640608721
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1640608721
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1640608721
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_301
timestamp 1640608721
transform 1 0 28796 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_305
timestamp 1640608721
transform 1 0 29164 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1640608721
transform -1 0 29532 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1640608721
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1640608721
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1640608721
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_27
timestamp 1640608721
transform 1 0 3588 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_29
timestamp 1640608721
transform 1 0 3772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_41
timestamp 1640608721
transform 1 0 4876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1640608721
transform 1 0 3680 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1640608721
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1640608721
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1640608721
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1640608721
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_81
timestamp 1640608721
transform 1 0 8556 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_85
timestamp 1640608721
transform 1 0 8924 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1640608721
transform 1 0 8832 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__B1
timestamp 1640608721
transform -1 0 10396 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_101
timestamp 1640608721
transform 1 0 10396 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_109
timestamp 1640608721
transform 1 0 11132 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_89
timestamp 1640608721
transform 1 0 9292 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1169_
timestamp 1640608721
transform -1 0 10212 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__B1
timestamp 1640608721
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_122
timestamp 1640608721
transform 1 0 12328 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1640608721
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1158_
timestamp 1640608721
transform -1 0 12328 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__B1
timestamp 1640608721
transform -1 0 14444 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_134
timestamp 1640608721
transform 1 0 13432 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_141
timestamp 1640608721
transform 1 0 14076 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1640608721
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1143_
timestamp 1640608721
transform 1 0 14444 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_51_154
timestamp 1640608721
transform 1 0 15272 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1640608721
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1640608721
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1640608721
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1147_
timestamp 1640608721
transform 1 0 16928 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B1
timestamp 1640608721
transform -1 0 17940 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_183
timestamp 1640608721
transform 1 0 17940 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_195
timestamp 1640608721
transform 1 0 19044 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1640608721
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_197
timestamp 1640608721
transform 1 0 19228 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_209
timestamp 1640608721
transform 1 0 20332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1640608721
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1640608721
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1640608721
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1640608721
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_249
timestamp 1640608721
transform 1 0 24012 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_253
timestamp 1640608721
transform 1 0 24380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1640608721
transform 1 0 24288 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_265
timestamp 1640608721
transform 1 0 25484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1640608721
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1640608721
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1640608721
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1640608721
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_305
timestamp 1640608721
transform 1 0 29164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1640608721
transform -1 0 29532 0 -1 30464
box -38 -48 314 592
<< labels >>
rlabel metal3 s 29912 688 30712 808 6 clk_i
port 0 nsew signal input
rlabel metal2 s 1766 32056 1822 32856 6 data_addr_o[0]
port 1 nsew signal tristate
rlabel metal3 s 0 15648 800 15768 6 data_addr_o[10]
port 2 nsew signal tristate
rlabel metal3 s 0 18504 800 18624 6 data_addr_o[11]
port 3 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 data_addr_o[1]
port 4 nsew signal tristate
rlabel metal3 s 29912 5176 30712 5296 6 data_addr_o[2]
port 5 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 data_addr_o[3]
port 6 nsew signal tristate
rlabel metal2 s 7930 32056 7986 32856 6 data_addr_o[4]
port 7 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 data_addr_o[5]
port 8 nsew signal tristate
rlabel metal2 s 9126 32056 9182 32856 6 data_addr_o[6]
port 9 nsew signal tristate
rlabel metal2 s 10322 32056 10378 32856 6 data_addr_o[7]
port 10 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 data_addr_o[8]
port 11 nsew signal tristate
rlabel metal3 s 29912 17144 30712 17264 6 data_addr_o[9]
port 12 nsew signal tristate
rlabel metal2 s 2962 32056 3018 32856 6 data_be_o[0]
port 13 nsew signal tristate
rlabel metal2 s 4250 32056 4306 32856 6 data_be_o[1]
port 14 nsew signal tristate
rlabel metal2 s 6642 32056 6698 32856 6 data_be_o[2]
port 15 nsew signal tristate
rlabel metal3 s 29912 8168 30712 8288 6 data_be_o[3]
port 16 nsew signal tristate
rlabel metal2 s 846 0 902 800 6 data_gnt_i
port 17 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 data_rdata_i[0]
port 18 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 data_rdata_i[10]
port 19 nsew signal input
rlabel metal2 s 14002 32056 14058 32856 6 data_rdata_i[11]
port 20 nsew signal input
rlabel metal2 s 15290 32056 15346 32856 6 data_rdata_i[12]
port 21 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 data_rdata_i[13]
port 22 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 data_rdata_i[14]
port 23 nsew signal input
rlabel metal3 s 29912 23128 30712 23248 6 data_rdata_i[15]
port 24 nsew signal input
rlabel metal2 s 16486 32056 16542 32856 6 data_rdata_i[16]
port 25 nsew signal input
rlabel metal2 s 17774 32056 17830 32856 6 data_rdata_i[17]
port 26 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 data_rdata_i[18]
port 27 nsew signal input
rlabel metal3 s 29912 27616 30712 27736 6 data_rdata_i[19]
port 28 nsew signal input
rlabel metal2 s 5446 32056 5502 32856 6 data_rdata_i[1]
port 29 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 data_rdata_i[20]
port 30 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 data_rdata_i[21]
port 31 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 data_rdata_i[22]
port 32 nsew signal input
rlabel metal2 s 21454 32056 21510 32856 6 data_rdata_i[23]
port 33 nsew signal input
rlabel metal3 s 29912 29112 30712 29232 6 data_rdata_i[24]
port 34 nsew signal input
rlabel metal2 s 23846 32056 23902 32856 6 data_rdata_i[25]
port 35 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 data_rdata_i[26]
port 36 nsew signal input
rlabel metal2 s 26330 32056 26386 32856 6 data_rdata_i[27]
port 37 nsew signal input
rlabel metal2 s 27526 32056 27582 32856 6 data_rdata_i[28]
port 38 nsew signal input
rlabel metal2 s 28814 32056 28870 32856 6 data_rdata_i[29]
port 39 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 data_rdata_i[2]
port 40 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 data_rdata_i[30]
port 41 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 data_rdata_i[31]
port 42 nsew signal input
rlabel metal3 s 29912 9664 30712 9784 6 data_rdata_i[3]
port 43 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 data_rdata_i[4]
port 44 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 data_rdata_i[5]
port 45 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 data_rdata_i[6]
port 46 nsew signal input
rlabel metal3 s 29912 15648 30712 15768 6 data_rdata_i[7]
port 47 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 data_rdata_i[8]
port 48 nsew signal input
rlabel metal3 s 29912 18640 30712 18760 6 data_rdata_i[9]
port 49 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 data_req_o
port 50 nsew signal tristate
rlabel metal3 s 0 688 800 808 6 data_rvalid_i
port 51 nsew signal input
rlabel metal3 s 29912 3680 30712 3800 6 data_wdata_o[0]
port 52 nsew signal tristate
rlabel metal2 s 12806 32056 12862 32856 6 data_wdata_o[10]
port 53 nsew signal tristate
rlabel metal2 s 14462 0 14518 800 6 data_wdata_o[11]
port 54 nsew signal tristate
rlabel metal3 s 29912 21632 30712 21752 6 data_wdata_o[12]
port 55 nsew signal tristate
rlabel metal2 s 16210 0 16266 800 6 data_wdata_o[13]
port 56 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 data_wdata_o[14]
port 57 nsew signal tristate
rlabel metal3 s 29912 24624 30712 24744 6 data_wdata_o[15]
port 58 nsew signal tristate
rlabel metal3 s 29912 26120 30712 26240 6 data_wdata_o[16]
port 59 nsew signal tristate
rlabel metal3 s 0 23944 800 24064 6 data_wdata_o[17]
port 60 nsew signal tristate
rlabel metal3 s 0 26664 800 26784 6 data_wdata_o[18]
port 61 nsew signal tristate
rlabel metal2 s 18970 32056 19026 32856 6 data_wdata_o[19]
port 62 nsew signal tristate
rlabel metal2 s 7654 0 7710 800 6 data_wdata_o[1]
port 63 nsew signal tristate
rlabel metal2 s 17866 0 17922 800 6 data_wdata_o[20]
port 64 nsew signal tristate
rlabel metal2 s 21270 0 21326 800 6 data_wdata_o[21]
port 65 nsew signal tristate
rlabel metal2 s 20166 32056 20222 32856 6 data_wdata_o[22]
port 66 nsew signal tristate
rlabel metal2 s 22650 32056 22706 32856 6 data_wdata_o[23]
port 67 nsew signal tristate
rlabel metal2 s 23018 0 23074 800 6 data_wdata_o[24]
port 68 nsew signal tristate
rlabel metal2 s 24674 0 24730 800 6 data_wdata_o[25]
port 69 nsew signal tristate
rlabel metal2 s 25134 32056 25190 32856 6 data_wdata_o[26]
port 70 nsew signal tristate
rlabel metal3 s 29912 30608 30712 30728 6 data_wdata_o[27]
port 71 nsew signal tristate
rlabel metal2 s 28078 0 28134 800 6 data_wdata_o[28]
port 72 nsew signal tristate
rlabel metal2 s 30010 32056 30066 32856 6 data_wdata_o[29]
port 73 nsew signal tristate
rlabel metal3 s 29912 6672 30712 6792 6 data_wdata_o[2]
port 74 nsew signal tristate
rlabel metal3 s 29912 32104 30712 32224 6 data_wdata_o[30]
port 75 nsew signal tristate
rlabel metal2 s 29826 0 29882 800 6 data_wdata_o[31]
port 76 nsew signal tristate
rlabel metal3 s 29912 11160 30712 11280 6 data_wdata_o[3]
port 77 nsew signal tristate
rlabel metal3 s 29912 12656 30712 12776 6 data_wdata_o[4]
port 78 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 data_wdata_o[5]
port 79 nsew signal tristate
rlabel metal3 s 29912 14152 30712 14272 6 data_wdata_o[6]
port 80 nsew signal tristate
rlabel metal2 s 11610 32056 11666 32856 6 data_wdata_o[7]
port 81 nsew signal tristate
rlabel metal3 s 0 14288 800 14408 6 data_wdata_o[8]
port 82 nsew signal tristate
rlabel metal3 s 29912 20136 30712 20256 6 data_wdata_o[9]
port 83 nsew signal tristate
rlabel metal2 s 4250 0 4306 800 6 data_we_o
port 84 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 rst_i
port 85 nsew signal input
rlabel metal3 s 29912 2184 30712 2304 6 rx_i
port 86 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 tx_o
port 87 nsew signal tristate
rlabel metal2 s 570 32056 626 32856 6 uart_error
port 88 nsew signal tristate
rlabel metal4 s 5681 2128 6001 30512 6 vccd1
port 89 nsew power input
rlabel metal4 s 15157 2128 15477 30512 6 vccd1
port 89 nsew power input
rlabel metal4 s 24633 2128 24953 30512 6 vccd1
port 89 nsew power input
rlabel metal4 s 10419 2128 10739 30512 6 vssd1
port 90 nsew ground input
rlabel metal4 s 19895 2128 20215 30512 6 vssd1
port 90 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 30712 32856
<< end >>
