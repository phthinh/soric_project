magic
tech sky130A
magscale 1 2
timestamp 1640346924
<< obsli1 >>
rect 1104 2159 238987 237745
<< obsm1 >>
rect 14 1368 239554 237856
<< metal2 >>
rect 478 239200 534 240000
rect 1490 239200 1546 240000
rect 2502 239200 2558 240000
rect 3514 239200 3570 240000
rect 4526 239200 4582 240000
rect 5538 239200 5594 240000
rect 6550 239200 6606 240000
rect 7654 239200 7710 240000
rect 8666 239200 8722 240000
rect 9678 239200 9734 240000
rect 10690 239200 10746 240000
rect 11702 239200 11758 240000
rect 12714 239200 12770 240000
rect 13726 239200 13782 240000
rect 14830 239200 14886 240000
rect 15842 239200 15898 240000
rect 16854 239200 16910 240000
rect 17866 239200 17922 240000
rect 18878 239200 18934 240000
rect 19890 239200 19946 240000
rect 20902 239200 20958 240000
rect 22006 239200 22062 240000
rect 23018 239200 23074 240000
rect 24030 239200 24086 240000
rect 25042 239200 25098 240000
rect 26054 239200 26110 240000
rect 27066 239200 27122 240000
rect 28170 239200 28226 240000
rect 29182 239200 29238 240000
rect 30194 239200 30250 240000
rect 31206 239200 31262 240000
rect 32218 239200 32274 240000
rect 33230 239200 33286 240000
rect 34242 239200 34298 240000
rect 35346 239200 35402 240000
rect 36358 239200 36414 240000
rect 37370 239200 37426 240000
rect 38382 239200 38438 240000
rect 39394 239200 39450 240000
rect 40406 239200 40462 240000
rect 41418 239200 41474 240000
rect 42522 239200 42578 240000
rect 43534 239200 43590 240000
rect 44546 239200 44602 240000
rect 45558 239200 45614 240000
rect 46570 239200 46626 240000
rect 47582 239200 47638 240000
rect 48686 239200 48742 240000
rect 49698 239200 49754 240000
rect 50710 239200 50766 240000
rect 51722 239200 51778 240000
rect 52734 239200 52790 240000
rect 53746 239200 53802 240000
rect 54758 239200 54814 240000
rect 55862 239200 55918 240000
rect 56874 239200 56930 240000
rect 57886 239200 57942 240000
rect 58898 239200 58954 240000
rect 59910 239200 59966 240000
rect 60922 239200 60978 240000
rect 61934 239200 61990 240000
rect 63038 239200 63094 240000
rect 64050 239200 64106 240000
rect 65062 239200 65118 240000
rect 66074 239200 66130 240000
rect 67086 239200 67142 240000
rect 68098 239200 68154 240000
rect 69202 239200 69258 240000
rect 70214 239200 70270 240000
rect 71226 239200 71282 240000
rect 72238 239200 72294 240000
rect 73250 239200 73306 240000
rect 74262 239200 74318 240000
rect 75274 239200 75330 240000
rect 76378 239200 76434 240000
rect 77390 239200 77446 240000
rect 78402 239200 78458 240000
rect 79414 239200 79470 240000
rect 80426 239200 80482 240000
rect 81438 239200 81494 240000
rect 82450 239200 82506 240000
rect 83554 239200 83610 240000
rect 84566 239200 84622 240000
rect 85578 239200 85634 240000
rect 86590 239200 86646 240000
rect 87602 239200 87658 240000
rect 88614 239200 88670 240000
rect 89718 239200 89774 240000
rect 90730 239200 90786 240000
rect 91742 239200 91798 240000
rect 92754 239200 92810 240000
rect 93766 239200 93822 240000
rect 94778 239200 94834 240000
rect 95790 239200 95846 240000
rect 96894 239200 96950 240000
rect 97906 239200 97962 240000
rect 98918 239200 98974 240000
rect 99930 239200 99986 240000
rect 100942 239200 100998 240000
rect 101954 239200 102010 240000
rect 102966 239200 103022 240000
rect 104070 239200 104126 240000
rect 105082 239200 105138 240000
rect 106094 239200 106150 240000
rect 107106 239200 107162 240000
rect 108118 239200 108174 240000
rect 109130 239200 109186 240000
rect 110234 239200 110290 240000
rect 111246 239200 111302 240000
rect 112258 239200 112314 240000
rect 113270 239200 113326 240000
rect 114282 239200 114338 240000
rect 115294 239200 115350 240000
rect 116306 239200 116362 240000
rect 117410 239200 117466 240000
rect 118422 239200 118478 240000
rect 119434 239200 119490 240000
rect 120446 239200 120502 240000
rect 121458 239200 121514 240000
rect 122470 239200 122526 240000
rect 123482 239200 123538 240000
rect 124586 239200 124642 240000
rect 125598 239200 125654 240000
rect 126610 239200 126666 240000
rect 127622 239200 127678 240000
rect 128634 239200 128690 240000
rect 129646 239200 129702 240000
rect 130658 239200 130714 240000
rect 131762 239200 131818 240000
rect 132774 239200 132830 240000
rect 133786 239200 133842 240000
rect 134798 239200 134854 240000
rect 135810 239200 135866 240000
rect 136822 239200 136878 240000
rect 137926 239200 137982 240000
rect 138938 239200 138994 240000
rect 139950 239200 140006 240000
rect 140962 239200 141018 240000
rect 141974 239200 142030 240000
rect 142986 239200 143042 240000
rect 143998 239200 144054 240000
rect 145102 239200 145158 240000
rect 146114 239200 146170 240000
rect 147126 239200 147182 240000
rect 148138 239200 148194 240000
rect 149150 239200 149206 240000
rect 150162 239200 150218 240000
rect 151174 239200 151230 240000
rect 152278 239200 152334 240000
rect 153290 239200 153346 240000
rect 154302 239200 154358 240000
rect 155314 239200 155370 240000
rect 156326 239200 156382 240000
rect 157338 239200 157394 240000
rect 158442 239200 158498 240000
rect 159454 239200 159510 240000
rect 160466 239200 160522 240000
rect 161478 239200 161534 240000
rect 162490 239200 162546 240000
rect 163502 239200 163558 240000
rect 164514 239200 164570 240000
rect 165618 239200 165674 240000
rect 166630 239200 166686 240000
rect 167642 239200 167698 240000
rect 168654 239200 168710 240000
rect 169666 239200 169722 240000
rect 170678 239200 170734 240000
rect 171690 239200 171746 240000
rect 172794 239200 172850 240000
rect 173806 239200 173862 240000
rect 174818 239200 174874 240000
rect 175830 239200 175886 240000
rect 176842 239200 176898 240000
rect 177854 239200 177910 240000
rect 178958 239200 179014 240000
rect 179970 239200 180026 240000
rect 180982 239200 181038 240000
rect 181994 239200 182050 240000
rect 183006 239200 183062 240000
rect 184018 239200 184074 240000
rect 185030 239200 185086 240000
rect 186134 239200 186190 240000
rect 187146 239200 187202 240000
rect 188158 239200 188214 240000
rect 189170 239200 189226 240000
rect 190182 239200 190238 240000
rect 191194 239200 191250 240000
rect 192206 239200 192262 240000
rect 193310 239200 193366 240000
rect 194322 239200 194378 240000
rect 195334 239200 195390 240000
rect 196346 239200 196402 240000
rect 197358 239200 197414 240000
rect 198370 239200 198426 240000
rect 199474 239200 199530 240000
rect 200486 239200 200542 240000
rect 201498 239200 201554 240000
rect 202510 239200 202566 240000
rect 203522 239200 203578 240000
rect 204534 239200 204590 240000
rect 205546 239200 205602 240000
rect 206650 239200 206706 240000
rect 207662 239200 207718 240000
rect 208674 239200 208730 240000
rect 209686 239200 209742 240000
rect 210698 239200 210754 240000
rect 211710 239200 211766 240000
rect 212722 239200 212778 240000
rect 213826 239200 213882 240000
rect 214838 239200 214894 240000
rect 215850 239200 215906 240000
rect 216862 239200 216918 240000
rect 217874 239200 217930 240000
rect 218886 239200 218942 240000
rect 219990 239200 220046 240000
rect 221002 239200 221058 240000
rect 222014 239200 222070 240000
rect 223026 239200 223082 240000
rect 224038 239200 224094 240000
rect 225050 239200 225106 240000
rect 226062 239200 226118 240000
rect 227166 239200 227222 240000
rect 228178 239200 228234 240000
rect 229190 239200 229246 240000
rect 230202 239200 230258 240000
rect 231214 239200 231270 240000
rect 232226 239200 232282 240000
rect 233238 239200 233294 240000
rect 234342 239200 234398 240000
rect 235354 239200 235410 240000
rect 236366 239200 236422 240000
rect 237378 239200 237434 240000
rect 238390 239200 238446 240000
rect 239402 239200 239458 240000
rect 386 0 442 800
rect 1214 0 1270 800
rect 2134 0 2190 800
rect 3054 0 3110 800
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 6734 0 6790 800
rect 7654 0 7710 800
rect 8574 0 8630 800
rect 9494 0 9550 800
rect 10414 0 10470 800
rect 11334 0 11390 800
rect 12254 0 12310 800
rect 13174 0 13230 800
rect 14094 0 14150 800
rect 15014 0 15070 800
rect 15934 0 15990 800
rect 16854 0 16910 800
rect 17774 0 17830 800
rect 18694 0 18750 800
rect 19614 0 19670 800
rect 20534 0 20590 800
rect 21454 0 21510 800
rect 22282 0 22338 800
rect 23202 0 23258 800
rect 24122 0 24178 800
rect 25042 0 25098 800
rect 25962 0 26018 800
rect 26882 0 26938 800
rect 27802 0 27858 800
rect 28722 0 28778 800
rect 29642 0 29698 800
rect 30562 0 30618 800
rect 31482 0 31538 800
rect 32402 0 32458 800
rect 33322 0 33378 800
rect 34242 0 34298 800
rect 35162 0 35218 800
rect 36082 0 36138 800
rect 37002 0 37058 800
rect 37922 0 37978 800
rect 38842 0 38898 800
rect 39762 0 39818 800
rect 40682 0 40738 800
rect 41602 0 41658 800
rect 42522 0 42578 800
rect 43442 0 43498 800
rect 44270 0 44326 800
rect 45190 0 45246 800
rect 46110 0 46166 800
rect 47030 0 47086 800
rect 47950 0 48006 800
rect 48870 0 48926 800
rect 49790 0 49846 800
rect 50710 0 50766 800
rect 51630 0 51686 800
rect 52550 0 52606 800
rect 53470 0 53526 800
rect 54390 0 54446 800
rect 55310 0 55366 800
rect 56230 0 56286 800
rect 57150 0 57206 800
rect 58070 0 58126 800
rect 58990 0 59046 800
rect 59910 0 59966 800
rect 60830 0 60886 800
rect 61750 0 61806 800
rect 62670 0 62726 800
rect 63590 0 63646 800
rect 64510 0 64566 800
rect 65430 0 65486 800
rect 66258 0 66314 800
rect 67178 0 67234 800
rect 68098 0 68154 800
rect 69018 0 69074 800
rect 69938 0 69994 800
rect 70858 0 70914 800
rect 71778 0 71834 800
rect 72698 0 72754 800
rect 73618 0 73674 800
rect 74538 0 74594 800
rect 75458 0 75514 800
rect 76378 0 76434 800
rect 77298 0 77354 800
rect 78218 0 78274 800
rect 79138 0 79194 800
rect 80058 0 80114 800
rect 80978 0 81034 800
rect 81898 0 81954 800
rect 82818 0 82874 800
rect 83738 0 83794 800
rect 84658 0 84714 800
rect 85578 0 85634 800
rect 86498 0 86554 800
rect 87418 0 87474 800
rect 88246 0 88302 800
rect 89166 0 89222 800
rect 90086 0 90142 800
rect 91006 0 91062 800
rect 91926 0 91982 800
rect 92846 0 92902 800
rect 93766 0 93822 800
rect 94686 0 94742 800
rect 95606 0 95662 800
rect 96526 0 96582 800
rect 97446 0 97502 800
rect 98366 0 98422 800
rect 99286 0 99342 800
rect 100206 0 100262 800
rect 101126 0 101182 800
rect 102046 0 102102 800
rect 102966 0 103022 800
rect 103886 0 103942 800
rect 104806 0 104862 800
rect 105726 0 105782 800
rect 106646 0 106702 800
rect 107566 0 107622 800
rect 108486 0 108542 800
rect 109406 0 109462 800
rect 110234 0 110290 800
rect 111154 0 111210 800
rect 112074 0 112130 800
rect 112994 0 113050 800
rect 113914 0 113970 800
rect 114834 0 114890 800
rect 115754 0 115810 800
rect 116674 0 116730 800
rect 117594 0 117650 800
rect 118514 0 118570 800
rect 119434 0 119490 800
rect 120354 0 120410 800
rect 121274 0 121330 800
rect 122194 0 122250 800
rect 123114 0 123170 800
rect 124034 0 124090 800
rect 124954 0 125010 800
rect 125874 0 125930 800
rect 126794 0 126850 800
rect 127714 0 127770 800
rect 128634 0 128690 800
rect 129554 0 129610 800
rect 130474 0 130530 800
rect 131302 0 131358 800
rect 132222 0 132278 800
rect 133142 0 133198 800
rect 134062 0 134118 800
rect 134982 0 135038 800
rect 135902 0 135958 800
rect 136822 0 136878 800
rect 137742 0 137798 800
rect 138662 0 138718 800
rect 139582 0 139638 800
rect 140502 0 140558 800
rect 141422 0 141478 800
rect 142342 0 142398 800
rect 143262 0 143318 800
rect 144182 0 144238 800
rect 145102 0 145158 800
rect 146022 0 146078 800
rect 146942 0 146998 800
rect 147862 0 147918 800
rect 148782 0 148838 800
rect 149702 0 149758 800
rect 150622 0 150678 800
rect 151542 0 151598 800
rect 152462 0 152518 800
rect 153290 0 153346 800
rect 154210 0 154266 800
rect 155130 0 155186 800
rect 156050 0 156106 800
rect 156970 0 157026 800
rect 157890 0 157946 800
rect 158810 0 158866 800
rect 159730 0 159786 800
rect 160650 0 160706 800
rect 161570 0 161626 800
rect 162490 0 162546 800
rect 163410 0 163466 800
rect 164330 0 164386 800
rect 165250 0 165306 800
rect 166170 0 166226 800
rect 167090 0 167146 800
rect 168010 0 168066 800
rect 168930 0 168986 800
rect 169850 0 169906 800
rect 170770 0 170826 800
rect 171690 0 171746 800
rect 172610 0 172666 800
rect 173530 0 173586 800
rect 174450 0 174506 800
rect 175278 0 175334 800
rect 176198 0 176254 800
rect 177118 0 177174 800
rect 178038 0 178094 800
rect 178958 0 179014 800
rect 179878 0 179934 800
rect 180798 0 180854 800
rect 181718 0 181774 800
rect 182638 0 182694 800
rect 183558 0 183614 800
rect 184478 0 184534 800
rect 185398 0 185454 800
rect 186318 0 186374 800
rect 187238 0 187294 800
rect 188158 0 188214 800
rect 189078 0 189134 800
rect 189998 0 190054 800
rect 190918 0 190974 800
rect 191838 0 191894 800
rect 192758 0 192814 800
rect 193678 0 193734 800
rect 194598 0 194654 800
rect 195518 0 195574 800
rect 196438 0 196494 800
rect 197266 0 197322 800
rect 198186 0 198242 800
rect 199106 0 199162 800
rect 200026 0 200082 800
rect 200946 0 201002 800
rect 201866 0 201922 800
rect 202786 0 202842 800
rect 203706 0 203762 800
rect 204626 0 204682 800
rect 205546 0 205602 800
rect 206466 0 206522 800
rect 207386 0 207442 800
rect 208306 0 208362 800
rect 209226 0 209282 800
rect 210146 0 210202 800
rect 211066 0 211122 800
rect 211986 0 212042 800
rect 212906 0 212962 800
rect 213826 0 213882 800
rect 214746 0 214802 800
rect 215666 0 215722 800
rect 216586 0 216642 800
rect 217506 0 217562 800
rect 218426 0 218482 800
rect 219254 0 219310 800
rect 220174 0 220230 800
rect 221094 0 221150 800
rect 222014 0 222070 800
rect 222934 0 222990 800
rect 223854 0 223910 800
rect 224774 0 224830 800
rect 225694 0 225750 800
rect 226614 0 226670 800
rect 227534 0 227590 800
rect 228454 0 228510 800
rect 229374 0 229430 800
rect 230294 0 230350 800
rect 231214 0 231270 800
rect 232134 0 232190 800
rect 233054 0 233110 800
rect 233974 0 234030 800
rect 234894 0 234950 800
rect 235814 0 235870 800
rect 236734 0 236790 800
rect 237654 0 237710 800
rect 238574 0 238630 800
rect 239494 0 239550 800
<< obsm2 >>
rect 20 239144 422 239306
rect 590 239144 1434 239306
rect 1602 239144 2446 239306
rect 2614 239144 3458 239306
rect 3626 239144 4470 239306
rect 4638 239144 5482 239306
rect 5650 239144 6494 239306
rect 6662 239144 7598 239306
rect 7766 239144 8610 239306
rect 8778 239144 9622 239306
rect 9790 239144 10634 239306
rect 10802 239144 11646 239306
rect 11814 239144 12658 239306
rect 12826 239144 13670 239306
rect 13838 239144 14774 239306
rect 14942 239144 15786 239306
rect 15954 239144 16798 239306
rect 16966 239144 17810 239306
rect 17978 239144 18822 239306
rect 18990 239144 19834 239306
rect 20002 239144 20846 239306
rect 21014 239144 21950 239306
rect 22118 239144 22962 239306
rect 23130 239144 23974 239306
rect 24142 239144 24986 239306
rect 25154 239144 25998 239306
rect 26166 239144 27010 239306
rect 27178 239144 28114 239306
rect 28282 239144 29126 239306
rect 29294 239144 30138 239306
rect 30306 239144 31150 239306
rect 31318 239144 32162 239306
rect 32330 239144 33174 239306
rect 33342 239144 34186 239306
rect 34354 239144 35290 239306
rect 35458 239144 36302 239306
rect 36470 239144 37314 239306
rect 37482 239144 38326 239306
rect 38494 239144 39338 239306
rect 39506 239144 40350 239306
rect 40518 239144 41362 239306
rect 41530 239144 42466 239306
rect 42634 239144 43478 239306
rect 43646 239144 44490 239306
rect 44658 239144 45502 239306
rect 45670 239144 46514 239306
rect 46682 239144 47526 239306
rect 47694 239144 48630 239306
rect 48798 239144 49642 239306
rect 49810 239144 50654 239306
rect 50822 239144 51666 239306
rect 51834 239144 52678 239306
rect 52846 239144 53690 239306
rect 53858 239144 54702 239306
rect 54870 239144 55806 239306
rect 55974 239144 56818 239306
rect 56986 239144 57830 239306
rect 57998 239144 58842 239306
rect 59010 239144 59854 239306
rect 60022 239144 60866 239306
rect 61034 239144 61878 239306
rect 62046 239144 62982 239306
rect 63150 239144 63994 239306
rect 64162 239144 65006 239306
rect 65174 239144 66018 239306
rect 66186 239144 67030 239306
rect 67198 239144 68042 239306
rect 68210 239144 69146 239306
rect 69314 239144 70158 239306
rect 70326 239144 71170 239306
rect 71338 239144 72182 239306
rect 72350 239144 73194 239306
rect 73362 239144 74206 239306
rect 74374 239144 75218 239306
rect 75386 239144 76322 239306
rect 76490 239144 77334 239306
rect 77502 239144 78346 239306
rect 78514 239144 79358 239306
rect 79526 239144 80370 239306
rect 80538 239144 81382 239306
rect 81550 239144 82394 239306
rect 82562 239144 83498 239306
rect 83666 239144 84510 239306
rect 84678 239144 85522 239306
rect 85690 239144 86534 239306
rect 86702 239144 87546 239306
rect 87714 239144 88558 239306
rect 88726 239144 89662 239306
rect 89830 239144 90674 239306
rect 90842 239144 91686 239306
rect 91854 239144 92698 239306
rect 92866 239144 93710 239306
rect 93878 239144 94722 239306
rect 94890 239144 95734 239306
rect 95902 239144 96838 239306
rect 97006 239144 97850 239306
rect 98018 239144 98862 239306
rect 99030 239144 99874 239306
rect 100042 239144 100886 239306
rect 101054 239144 101898 239306
rect 102066 239144 102910 239306
rect 103078 239144 104014 239306
rect 104182 239144 105026 239306
rect 105194 239144 106038 239306
rect 106206 239144 107050 239306
rect 107218 239144 108062 239306
rect 108230 239144 109074 239306
rect 109242 239144 110178 239306
rect 110346 239144 111190 239306
rect 111358 239144 112202 239306
rect 112370 239144 113214 239306
rect 113382 239144 114226 239306
rect 114394 239144 115238 239306
rect 115406 239144 116250 239306
rect 116418 239144 117354 239306
rect 117522 239144 118366 239306
rect 118534 239144 119378 239306
rect 119546 239144 120390 239306
rect 120558 239144 121402 239306
rect 121570 239144 122414 239306
rect 122582 239144 123426 239306
rect 123594 239144 124530 239306
rect 124698 239144 125542 239306
rect 125710 239144 126554 239306
rect 126722 239144 127566 239306
rect 127734 239144 128578 239306
rect 128746 239144 129590 239306
rect 129758 239144 130602 239306
rect 130770 239144 131706 239306
rect 131874 239144 132718 239306
rect 132886 239144 133730 239306
rect 133898 239144 134742 239306
rect 134910 239144 135754 239306
rect 135922 239144 136766 239306
rect 136934 239144 137870 239306
rect 138038 239144 138882 239306
rect 139050 239144 139894 239306
rect 140062 239144 140906 239306
rect 141074 239144 141918 239306
rect 142086 239144 142930 239306
rect 143098 239144 143942 239306
rect 144110 239144 145046 239306
rect 145214 239144 146058 239306
rect 146226 239144 147070 239306
rect 147238 239144 148082 239306
rect 148250 239144 149094 239306
rect 149262 239144 150106 239306
rect 150274 239144 151118 239306
rect 151286 239144 152222 239306
rect 152390 239144 153234 239306
rect 153402 239144 154246 239306
rect 154414 239144 155258 239306
rect 155426 239144 156270 239306
rect 156438 239144 157282 239306
rect 157450 239144 158386 239306
rect 158554 239144 159398 239306
rect 159566 239144 160410 239306
rect 160578 239144 161422 239306
rect 161590 239144 162434 239306
rect 162602 239144 163446 239306
rect 163614 239144 164458 239306
rect 164626 239144 165562 239306
rect 165730 239144 166574 239306
rect 166742 239144 167586 239306
rect 167754 239144 168598 239306
rect 168766 239144 169610 239306
rect 169778 239144 170622 239306
rect 170790 239144 171634 239306
rect 171802 239144 172738 239306
rect 172906 239144 173750 239306
rect 173918 239144 174762 239306
rect 174930 239144 175774 239306
rect 175942 239144 176786 239306
rect 176954 239144 177798 239306
rect 177966 239144 178902 239306
rect 179070 239144 179914 239306
rect 180082 239144 180926 239306
rect 181094 239144 181938 239306
rect 182106 239144 182950 239306
rect 183118 239144 183962 239306
rect 184130 239144 184974 239306
rect 185142 239144 186078 239306
rect 186246 239144 187090 239306
rect 187258 239144 188102 239306
rect 188270 239144 189114 239306
rect 189282 239144 190126 239306
rect 190294 239144 191138 239306
rect 191306 239144 192150 239306
rect 192318 239144 193254 239306
rect 193422 239144 194266 239306
rect 194434 239144 195278 239306
rect 195446 239144 196290 239306
rect 196458 239144 197302 239306
rect 197470 239144 198314 239306
rect 198482 239144 199418 239306
rect 199586 239144 200430 239306
rect 200598 239144 201442 239306
rect 201610 239144 202454 239306
rect 202622 239144 203466 239306
rect 203634 239144 204478 239306
rect 204646 239144 205490 239306
rect 205658 239144 206594 239306
rect 206762 239144 207606 239306
rect 207774 239144 208618 239306
rect 208786 239144 209630 239306
rect 209798 239144 210642 239306
rect 210810 239144 211654 239306
rect 211822 239144 212666 239306
rect 212834 239144 213770 239306
rect 213938 239144 214782 239306
rect 214950 239144 215794 239306
rect 215962 239144 216806 239306
rect 216974 239144 217818 239306
rect 217986 239144 218830 239306
rect 218998 239144 219934 239306
rect 220102 239144 220946 239306
rect 221114 239144 221958 239306
rect 222126 239144 222970 239306
rect 223138 239144 223982 239306
rect 224150 239144 224994 239306
rect 225162 239144 226006 239306
rect 226174 239144 227110 239306
rect 227278 239144 228122 239306
rect 228290 239144 229134 239306
rect 229302 239144 230146 239306
rect 230314 239144 231158 239306
rect 231326 239144 232170 239306
rect 232338 239144 233182 239306
rect 233350 239144 234286 239306
rect 234454 239144 235298 239306
rect 235466 239144 236310 239306
rect 236478 239144 237322 239306
rect 237490 239144 238334 239306
rect 238502 239144 239346 239306
rect 239514 239144 239548 239306
rect 20 856 239548 239144
rect 20 439 330 856
rect 498 439 1158 856
rect 1326 439 2078 856
rect 2246 439 2998 856
rect 3166 439 3918 856
rect 4086 439 4838 856
rect 5006 439 5758 856
rect 5926 439 6678 856
rect 6846 439 7598 856
rect 7766 439 8518 856
rect 8686 439 9438 856
rect 9606 439 10358 856
rect 10526 439 11278 856
rect 11446 439 12198 856
rect 12366 439 13118 856
rect 13286 439 14038 856
rect 14206 439 14958 856
rect 15126 439 15878 856
rect 16046 439 16798 856
rect 16966 439 17718 856
rect 17886 439 18638 856
rect 18806 439 19558 856
rect 19726 439 20478 856
rect 20646 439 21398 856
rect 21566 439 22226 856
rect 22394 439 23146 856
rect 23314 439 24066 856
rect 24234 439 24986 856
rect 25154 439 25906 856
rect 26074 439 26826 856
rect 26994 439 27746 856
rect 27914 439 28666 856
rect 28834 439 29586 856
rect 29754 439 30506 856
rect 30674 439 31426 856
rect 31594 439 32346 856
rect 32514 439 33266 856
rect 33434 439 34186 856
rect 34354 439 35106 856
rect 35274 439 36026 856
rect 36194 439 36946 856
rect 37114 439 37866 856
rect 38034 439 38786 856
rect 38954 439 39706 856
rect 39874 439 40626 856
rect 40794 439 41546 856
rect 41714 439 42466 856
rect 42634 439 43386 856
rect 43554 439 44214 856
rect 44382 439 45134 856
rect 45302 439 46054 856
rect 46222 439 46974 856
rect 47142 439 47894 856
rect 48062 439 48814 856
rect 48982 439 49734 856
rect 49902 439 50654 856
rect 50822 439 51574 856
rect 51742 439 52494 856
rect 52662 439 53414 856
rect 53582 439 54334 856
rect 54502 439 55254 856
rect 55422 439 56174 856
rect 56342 439 57094 856
rect 57262 439 58014 856
rect 58182 439 58934 856
rect 59102 439 59854 856
rect 60022 439 60774 856
rect 60942 439 61694 856
rect 61862 439 62614 856
rect 62782 439 63534 856
rect 63702 439 64454 856
rect 64622 439 65374 856
rect 65542 439 66202 856
rect 66370 439 67122 856
rect 67290 439 68042 856
rect 68210 439 68962 856
rect 69130 439 69882 856
rect 70050 439 70802 856
rect 70970 439 71722 856
rect 71890 439 72642 856
rect 72810 439 73562 856
rect 73730 439 74482 856
rect 74650 439 75402 856
rect 75570 439 76322 856
rect 76490 439 77242 856
rect 77410 439 78162 856
rect 78330 439 79082 856
rect 79250 439 80002 856
rect 80170 439 80922 856
rect 81090 439 81842 856
rect 82010 439 82762 856
rect 82930 439 83682 856
rect 83850 439 84602 856
rect 84770 439 85522 856
rect 85690 439 86442 856
rect 86610 439 87362 856
rect 87530 439 88190 856
rect 88358 439 89110 856
rect 89278 439 90030 856
rect 90198 439 90950 856
rect 91118 439 91870 856
rect 92038 439 92790 856
rect 92958 439 93710 856
rect 93878 439 94630 856
rect 94798 439 95550 856
rect 95718 439 96470 856
rect 96638 439 97390 856
rect 97558 439 98310 856
rect 98478 439 99230 856
rect 99398 439 100150 856
rect 100318 439 101070 856
rect 101238 439 101990 856
rect 102158 439 102910 856
rect 103078 439 103830 856
rect 103998 439 104750 856
rect 104918 439 105670 856
rect 105838 439 106590 856
rect 106758 439 107510 856
rect 107678 439 108430 856
rect 108598 439 109350 856
rect 109518 439 110178 856
rect 110346 439 111098 856
rect 111266 439 112018 856
rect 112186 439 112938 856
rect 113106 439 113858 856
rect 114026 439 114778 856
rect 114946 439 115698 856
rect 115866 439 116618 856
rect 116786 439 117538 856
rect 117706 439 118458 856
rect 118626 439 119378 856
rect 119546 439 120298 856
rect 120466 439 121218 856
rect 121386 439 122138 856
rect 122306 439 123058 856
rect 123226 439 123978 856
rect 124146 439 124898 856
rect 125066 439 125818 856
rect 125986 439 126738 856
rect 126906 439 127658 856
rect 127826 439 128578 856
rect 128746 439 129498 856
rect 129666 439 130418 856
rect 130586 439 131246 856
rect 131414 439 132166 856
rect 132334 439 133086 856
rect 133254 439 134006 856
rect 134174 439 134926 856
rect 135094 439 135846 856
rect 136014 439 136766 856
rect 136934 439 137686 856
rect 137854 439 138606 856
rect 138774 439 139526 856
rect 139694 439 140446 856
rect 140614 439 141366 856
rect 141534 439 142286 856
rect 142454 439 143206 856
rect 143374 439 144126 856
rect 144294 439 145046 856
rect 145214 439 145966 856
rect 146134 439 146886 856
rect 147054 439 147806 856
rect 147974 439 148726 856
rect 148894 439 149646 856
rect 149814 439 150566 856
rect 150734 439 151486 856
rect 151654 439 152406 856
rect 152574 439 153234 856
rect 153402 439 154154 856
rect 154322 439 155074 856
rect 155242 439 155994 856
rect 156162 439 156914 856
rect 157082 439 157834 856
rect 158002 439 158754 856
rect 158922 439 159674 856
rect 159842 439 160594 856
rect 160762 439 161514 856
rect 161682 439 162434 856
rect 162602 439 163354 856
rect 163522 439 164274 856
rect 164442 439 165194 856
rect 165362 439 166114 856
rect 166282 439 167034 856
rect 167202 439 167954 856
rect 168122 439 168874 856
rect 169042 439 169794 856
rect 169962 439 170714 856
rect 170882 439 171634 856
rect 171802 439 172554 856
rect 172722 439 173474 856
rect 173642 439 174394 856
rect 174562 439 175222 856
rect 175390 439 176142 856
rect 176310 439 177062 856
rect 177230 439 177982 856
rect 178150 439 178902 856
rect 179070 439 179822 856
rect 179990 439 180742 856
rect 180910 439 181662 856
rect 181830 439 182582 856
rect 182750 439 183502 856
rect 183670 439 184422 856
rect 184590 439 185342 856
rect 185510 439 186262 856
rect 186430 439 187182 856
rect 187350 439 188102 856
rect 188270 439 189022 856
rect 189190 439 189942 856
rect 190110 439 190862 856
rect 191030 439 191782 856
rect 191950 439 192702 856
rect 192870 439 193622 856
rect 193790 439 194542 856
rect 194710 439 195462 856
rect 195630 439 196382 856
rect 196550 439 197210 856
rect 197378 439 198130 856
rect 198298 439 199050 856
rect 199218 439 199970 856
rect 200138 439 200890 856
rect 201058 439 201810 856
rect 201978 439 202730 856
rect 202898 439 203650 856
rect 203818 439 204570 856
rect 204738 439 205490 856
rect 205658 439 206410 856
rect 206578 439 207330 856
rect 207498 439 208250 856
rect 208418 439 209170 856
rect 209338 439 210090 856
rect 210258 439 211010 856
rect 211178 439 211930 856
rect 212098 439 212850 856
rect 213018 439 213770 856
rect 213938 439 214690 856
rect 214858 439 215610 856
rect 215778 439 216530 856
rect 216698 439 217450 856
rect 217618 439 218370 856
rect 218538 439 219198 856
rect 219366 439 220118 856
rect 220286 439 221038 856
rect 221206 439 221958 856
rect 222126 439 222878 856
rect 223046 439 223798 856
rect 223966 439 224718 856
rect 224886 439 225638 856
rect 225806 439 226558 856
rect 226726 439 227478 856
rect 227646 439 228398 856
rect 228566 439 229318 856
rect 229486 439 230238 856
rect 230406 439 231158 856
rect 231326 439 232078 856
rect 232246 439 232998 856
rect 233166 439 233918 856
rect 234086 439 234838 856
rect 235006 439 235758 856
rect 235926 439 236678 856
rect 236846 439 237598 856
rect 237766 439 238518 856
rect 238686 439 239438 856
<< metal3 >>
rect 0 239368 800 239488
rect 239200 239368 240000 239488
rect 0 238280 800 238400
rect 239200 238280 240000 238400
rect 0 237192 800 237312
rect 239200 237192 240000 237312
rect 0 236240 800 236360
rect 239200 236240 240000 236360
rect 0 235152 800 235272
rect 239200 235152 240000 235272
rect 0 234064 800 234184
rect 239200 234064 240000 234184
rect 0 233112 800 233232
rect 239200 233112 240000 233232
rect 0 232024 800 232144
rect 239200 232024 240000 232144
rect 0 230936 800 231056
rect 239200 230936 240000 231056
rect 0 229848 800 229968
rect 239200 229848 240000 229968
rect 0 228896 800 229016
rect 239200 228896 240000 229016
rect 0 227808 800 227928
rect 239200 227808 240000 227928
rect 0 226720 800 226840
rect 239200 226720 240000 226840
rect 0 225768 800 225888
rect 239200 225768 240000 225888
rect 0 224680 800 224800
rect 239200 224680 240000 224800
rect 0 223592 800 223712
rect 239200 223592 240000 223712
rect 0 222504 800 222624
rect 239200 222504 240000 222624
rect 0 221552 800 221672
rect 239200 221552 240000 221672
rect 0 220464 800 220584
rect 239200 220464 240000 220584
rect 0 219376 800 219496
rect 239200 219376 240000 219496
rect 0 218424 800 218544
rect 239200 218424 240000 218544
rect 0 217336 800 217456
rect 239200 217336 240000 217456
rect 0 216248 800 216368
rect 239200 216248 240000 216368
rect 0 215296 800 215416
rect 239200 215296 240000 215416
rect 0 214208 800 214328
rect 239200 214208 240000 214328
rect 0 213120 800 213240
rect 239200 213120 240000 213240
rect 0 212032 800 212152
rect 239200 212032 240000 212152
rect 0 211080 800 211200
rect 239200 211080 240000 211200
rect 0 209992 800 210112
rect 239200 209992 240000 210112
rect 0 208904 800 209024
rect 239200 208904 240000 209024
rect 0 207952 800 208072
rect 239200 207952 240000 208072
rect 0 206864 800 206984
rect 239200 206864 240000 206984
rect 0 205776 800 205896
rect 239200 205776 240000 205896
rect 0 204688 800 204808
rect 239200 204688 240000 204808
rect 0 203736 800 203856
rect 239200 203736 240000 203856
rect 0 202648 800 202768
rect 239200 202648 240000 202768
rect 0 201560 800 201680
rect 239200 201560 240000 201680
rect 0 200608 800 200728
rect 239200 200608 240000 200728
rect 0 199520 800 199640
rect 239200 199520 240000 199640
rect 0 198432 800 198552
rect 239200 198432 240000 198552
rect 0 197344 800 197464
rect 239200 197344 240000 197464
rect 0 196392 800 196512
rect 239200 196392 240000 196512
rect 0 195304 800 195424
rect 239200 195304 240000 195424
rect 0 194216 800 194336
rect 239200 194216 240000 194336
rect 0 193264 800 193384
rect 239200 193264 240000 193384
rect 0 192176 800 192296
rect 239200 192176 240000 192296
rect 0 191088 800 191208
rect 239200 191088 240000 191208
rect 0 190136 800 190256
rect 239200 190136 240000 190256
rect 0 189048 800 189168
rect 239200 189048 240000 189168
rect 0 187960 800 188080
rect 239200 187960 240000 188080
rect 0 186872 800 186992
rect 239200 186872 240000 186992
rect 0 185920 800 186040
rect 239200 185920 240000 186040
rect 0 184832 800 184952
rect 239200 184832 240000 184952
rect 0 183744 800 183864
rect 239200 183744 240000 183864
rect 0 182792 800 182912
rect 239200 182792 240000 182912
rect 0 181704 800 181824
rect 239200 181704 240000 181824
rect 0 180616 800 180736
rect 239200 180616 240000 180736
rect 0 179528 800 179648
rect 239200 179528 240000 179648
rect 0 178576 800 178696
rect 239200 178576 240000 178696
rect 0 177488 800 177608
rect 239200 177488 240000 177608
rect 0 176400 800 176520
rect 239200 176400 240000 176520
rect 0 175448 800 175568
rect 239200 175448 240000 175568
rect 0 174360 800 174480
rect 239200 174360 240000 174480
rect 0 173272 800 173392
rect 239200 173272 240000 173392
rect 0 172320 800 172440
rect 239200 172320 240000 172440
rect 0 171232 800 171352
rect 239200 171232 240000 171352
rect 0 170144 800 170264
rect 239200 170144 240000 170264
rect 0 169056 800 169176
rect 239200 169056 240000 169176
rect 0 168104 800 168224
rect 239200 168104 240000 168224
rect 0 167016 800 167136
rect 239200 167016 240000 167136
rect 0 165928 800 166048
rect 239200 165928 240000 166048
rect 0 164976 800 165096
rect 239200 164976 240000 165096
rect 0 163888 800 164008
rect 239200 163888 240000 164008
rect 0 162800 800 162920
rect 239200 162800 240000 162920
rect 0 161712 800 161832
rect 239200 161712 240000 161832
rect 0 160760 800 160880
rect 239200 160760 240000 160880
rect 0 159672 800 159792
rect 239200 159672 240000 159792
rect 0 158584 800 158704
rect 239200 158584 240000 158704
rect 0 157632 800 157752
rect 239200 157632 240000 157752
rect 0 156544 800 156664
rect 239200 156544 240000 156664
rect 0 155456 800 155576
rect 239200 155456 240000 155576
rect 0 154368 800 154488
rect 239200 154368 240000 154488
rect 0 153416 800 153536
rect 239200 153416 240000 153536
rect 0 152328 800 152448
rect 239200 152328 240000 152448
rect 0 151240 800 151360
rect 239200 151240 240000 151360
rect 0 150288 800 150408
rect 239200 150288 240000 150408
rect 0 149200 800 149320
rect 239200 149200 240000 149320
rect 0 148112 800 148232
rect 239200 148112 240000 148232
rect 0 147160 800 147280
rect 239200 147160 240000 147280
rect 0 146072 800 146192
rect 239200 146072 240000 146192
rect 0 144984 800 145104
rect 239200 144984 240000 145104
rect 0 143896 800 144016
rect 239200 143896 240000 144016
rect 0 142944 800 143064
rect 239200 142944 240000 143064
rect 0 141856 800 141976
rect 239200 141856 240000 141976
rect 0 140768 800 140888
rect 239200 140768 240000 140888
rect 0 139816 800 139936
rect 239200 139816 240000 139936
rect 0 138728 800 138848
rect 239200 138728 240000 138848
rect 0 137640 800 137760
rect 239200 137640 240000 137760
rect 0 136552 800 136672
rect 239200 136552 240000 136672
rect 0 135600 800 135720
rect 239200 135600 240000 135720
rect 0 134512 800 134632
rect 239200 134512 240000 134632
rect 0 133424 800 133544
rect 239200 133424 240000 133544
rect 0 132472 800 132592
rect 239200 132472 240000 132592
rect 0 131384 800 131504
rect 239200 131384 240000 131504
rect 0 130296 800 130416
rect 239200 130296 240000 130416
rect 0 129344 800 129464
rect 239200 129344 240000 129464
rect 0 128256 800 128376
rect 239200 128256 240000 128376
rect 0 127168 800 127288
rect 239200 127168 240000 127288
rect 0 126080 800 126200
rect 239200 126080 240000 126200
rect 0 125128 800 125248
rect 239200 125128 240000 125248
rect 0 124040 800 124160
rect 239200 124040 240000 124160
rect 0 122952 800 123072
rect 239200 122952 240000 123072
rect 0 122000 800 122120
rect 239200 122000 240000 122120
rect 0 120912 800 121032
rect 239200 120912 240000 121032
rect 0 119824 800 119944
rect 239200 119824 240000 119944
rect 0 118736 800 118856
rect 239200 118736 240000 118856
rect 0 117784 800 117904
rect 239200 117784 240000 117904
rect 0 116696 800 116816
rect 239200 116696 240000 116816
rect 0 115608 800 115728
rect 239200 115608 240000 115728
rect 0 114656 800 114776
rect 239200 114656 240000 114776
rect 0 113568 800 113688
rect 239200 113568 240000 113688
rect 0 112480 800 112600
rect 239200 112480 240000 112600
rect 0 111392 800 111512
rect 239200 111392 240000 111512
rect 0 110440 800 110560
rect 239200 110440 240000 110560
rect 0 109352 800 109472
rect 239200 109352 240000 109472
rect 0 108264 800 108384
rect 239200 108264 240000 108384
rect 0 107312 800 107432
rect 239200 107312 240000 107432
rect 0 106224 800 106344
rect 239200 106224 240000 106344
rect 0 105136 800 105256
rect 239200 105136 240000 105256
rect 0 104184 800 104304
rect 239200 104184 240000 104304
rect 0 103096 800 103216
rect 239200 103096 240000 103216
rect 0 102008 800 102128
rect 239200 102008 240000 102128
rect 0 100920 800 101040
rect 239200 100920 240000 101040
rect 0 99968 800 100088
rect 239200 99968 240000 100088
rect 0 98880 800 99000
rect 239200 98880 240000 99000
rect 0 97792 800 97912
rect 239200 97792 240000 97912
rect 0 96840 800 96960
rect 239200 96840 240000 96960
rect 0 95752 800 95872
rect 239200 95752 240000 95872
rect 0 94664 800 94784
rect 239200 94664 240000 94784
rect 0 93576 800 93696
rect 239200 93576 240000 93696
rect 0 92624 800 92744
rect 239200 92624 240000 92744
rect 0 91536 800 91656
rect 239200 91536 240000 91656
rect 0 90448 800 90568
rect 239200 90448 240000 90568
rect 0 89496 800 89616
rect 239200 89496 240000 89616
rect 0 88408 800 88528
rect 239200 88408 240000 88528
rect 0 87320 800 87440
rect 239200 87320 240000 87440
rect 0 86368 800 86488
rect 239200 86368 240000 86488
rect 0 85280 800 85400
rect 239200 85280 240000 85400
rect 0 84192 800 84312
rect 239200 84192 240000 84312
rect 0 83104 800 83224
rect 239200 83104 240000 83224
rect 0 82152 800 82272
rect 239200 82152 240000 82272
rect 0 81064 800 81184
rect 239200 81064 240000 81184
rect 0 79976 800 80096
rect 239200 79976 240000 80096
rect 0 79024 800 79144
rect 239200 79024 240000 79144
rect 0 77936 800 78056
rect 239200 77936 240000 78056
rect 0 76848 800 76968
rect 239200 76848 240000 76968
rect 0 75760 800 75880
rect 239200 75760 240000 75880
rect 0 74808 800 74928
rect 239200 74808 240000 74928
rect 0 73720 800 73840
rect 239200 73720 240000 73840
rect 0 72632 800 72752
rect 239200 72632 240000 72752
rect 0 71680 800 71800
rect 239200 71680 240000 71800
rect 0 70592 800 70712
rect 239200 70592 240000 70712
rect 0 69504 800 69624
rect 239200 69504 240000 69624
rect 0 68416 800 68536
rect 239200 68416 240000 68536
rect 0 67464 800 67584
rect 239200 67464 240000 67584
rect 0 66376 800 66496
rect 239200 66376 240000 66496
rect 0 65288 800 65408
rect 239200 65288 240000 65408
rect 0 64336 800 64456
rect 239200 64336 240000 64456
rect 0 63248 800 63368
rect 239200 63248 240000 63368
rect 0 62160 800 62280
rect 239200 62160 240000 62280
rect 0 61208 800 61328
rect 239200 61208 240000 61328
rect 0 60120 800 60240
rect 239200 60120 240000 60240
rect 0 59032 800 59152
rect 239200 59032 240000 59152
rect 0 57944 800 58064
rect 239200 57944 240000 58064
rect 0 56992 800 57112
rect 239200 56992 240000 57112
rect 0 55904 800 56024
rect 239200 55904 240000 56024
rect 0 54816 800 54936
rect 239200 54816 240000 54936
rect 0 53864 800 53984
rect 239200 53864 240000 53984
rect 0 52776 800 52896
rect 239200 52776 240000 52896
rect 0 51688 800 51808
rect 239200 51688 240000 51808
rect 0 50600 800 50720
rect 239200 50600 240000 50720
rect 0 49648 800 49768
rect 239200 49648 240000 49768
rect 0 48560 800 48680
rect 239200 48560 240000 48680
rect 0 47472 800 47592
rect 239200 47472 240000 47592
rect 0 46520 800 46640
rect 239200 46520 240000 46640
rect 0 45432 800 45552
rect 239200 45432 240000 45552
rect 0 44344 800 44464
rect 239200 44344 240000 44464
rect 0 43392 800 43512
rect 239200 43392 240000 43512
rect 0 42304 800 42424
rect 239200 42304 240000 42424
rect 0 41216 800 41336
rect 239200 41216 240000 41336
rect 0 40128 800 40248
rect 239200 40128 240000 40248
rect 0 39176 800 39296
rect 239200 39176 240000 39296
rect 0 38088 800 38208
rect 239200 38088 240000 38208
rect 0 37000 800 37120
rect 239200 37000 240000 37120
rect 0 36048 800 36168
rect 239200 36048 240000 36168
rect 0 34960 800 35080
rect 239200 34960 240000 35080
rect 0 33872 800 33992
rect 239200 33872 240000 33992
rect 0 32784 800 32904
rect 239200 32784 240000 32904
rect 0 31832 800 31952
rect 239200 31832 240000 31952
rect 0 30744 800 30864
rect 239200 30744 240000 30864
rect 0 29656 800 29776
rect 239200 29656 240000 29776
rect 0 28704 800 28824
rect 239200 28704 240000 28824
rect 0 27616 800 27736
rect 239200 27616 240000 27736
rect 0 26528 800 26648
rect 239200 26528 240000 26648
rect 0 25440 800 25560
rect 239200 25440 240000 25560
rect 0 24488 800 24608
rect 239200 24488 240000 24608
rect 0 23400 800 23520
rect 239200 23400 240000 23520
rect 0 22312 800 22432
rect 239200 22312 240000 22432
rect 0 21360 800 21480
rect 239200 21360 240000 21480
rect 0 20272 800 20392
rect 239200 20272 240000 20392
rect 0 19184 800 19304
rect 239200 19184 240000 19304
rect 0 18232 800 18352
rect 239200 18232 240000 18352
rect 0 17144 800 17264
rect 239200 17144 240000 17264
rect 0 16056 800 16176
rect 239200 16056 240000 16176
rect 0 14968 800 15088
rect 239200 14968 240000 15088
rect 0 14016 800 14136
rect 239200 14016 240000 14136
rect 0 12928 800 13048
rect 239200 12928 240000 13048
rect 0 11840 800 11960
rect 239200 11840 240000 11960
rect 0 10888 800 11008
rect 239200 10888 240000 11008
rect 0 9800 800 9920
rect 239200 9800 240000 9920
rect 0 8712 800 8832
rect 239200 8712 240000 8832
rect 0 7624 800 7744
rect 239200 7624 240000 7744
rect 0 6672 800 6792
rect 239200 6672 240000 6792
rect 0 5584 800 5704
rect 239200 5584 240000 5704
rect 0 4496 800 4616
rect 239200 4496 240000 4616
rect 0 3544 800 3664
rect 239200 3544 240000 3664
rect 0 2456 800 2576
rect 239200 2456 240000 2576
rect 0 1368 800 1488
rect 239200 1368 240000 1488
rect 0 416 800 536
rect 239200 416 240000 536
<< obsm3 >>
rect 880 238200 239120 238373
rect 800 237392 239322 238200
rect 880 237112 239120 237392
rect 800 236440 239322 237112
rect 880 236160 239120 236440
rect 800 235352 239322 236160
rect 880 235072 239120 235352
rect 800 234264 239322 235072
rect 880 233984 239120 234264
rect 800 233312 239322 233984
rect 880 233032 239120 233312
rect 800 232224 239322 233032
rect 880 231944 239120 232224
rect 800 231136 239322 231944
rect 880 230856 239120 231136
rect 800 230048 239322 230856
rect 880 229768 239120 230048
rect 800 229096 239322 229768
rect 880 228816 239120 229096
rect 800 228008 239322 228816
rect 880 227728 239120 228008
rect 800 226920 239322 227728
rect 880 226640 239120 226920
rect 800 225968 239322 226640
rect 880 225688 239120 225968
rect 800 224880 239322 225688
rect 880 224600 239120 224880
rect 800 223792 239322 224600
rect 880 223512 239120 223792
rect 800 222704 239322 223512
rect 880 222424 239120 222704
rect 800 221752 239322 222424
rect 880 221472 239120 221752
rect 800 220664 239322 221472
rect 880 220384 239120 220664
rect 800 219576 239322 220384
rect 880 219296 239120 219576
rect 800 218624 239322 219296
rect 880 218344 239120 218624
rect 800 217536 239322 218344
rect 880 217256 239120 217536
rect 800 216448 239322 217256
rect 880 216168 239120 216448
rect 800 215496 239322 216168
rect 880 215216 239120 215496
rect 800 214408 239322 215216
rect 880 214128 239120 214408
rect 800 213320 239322 214128
rect 880 213040 239120 213320
rect 800 212232 239322 213040
rect 880 211952 239120 212232
rect 800 211280 239322 211952
rect 880 211000 239120 211280
rect 800 210192 239322 211000
rect 880 209912 239120 210192
rect 800 209104 239322 209912
rect 880 208824 239120 209104
rect 800 208152 239322 208824
rect 880 207872 239120 208152
rect 800 207064 239322 207872
rect 880 206784 239120 207064
rect 800 205976 239322 206784
rect 880 205696 239120 205976
rect 800 204888 239322 205696
rect 880 204608 239120 204888
rect 800 203936 239322 204608
rect 880 203656 239120 203936
rect 800 202848 239322 203656
rect 880 202568 239120 202848
rect 800 201760 239322 202568
rect 880 201480 239120 201760
rect 800 200808 239322 201480
rect 880 200528 239120 200808
rect 800 199720 239322 200528
rect 880 199440 239120 199720
rect 800 198632 239322 199440
rect 880 198352 239120 198632
rect 800 197544 239322 198352
rect 880 197264 239120 197544
rect 800 196592 239322 197264
rect 880 196312 239120 196592
rect 800 195504 239322 196312
rect 880 195224 239120 195504
rect 800 194416 239322 195224
rect 880 194136 239120 194416
rect 800 193464 239322 194136
rect 880 193184 239120 193464
rect 800 192376 239322 193184
rect 880 192096 239120 192376
rect 800 191288 239322 192096
rect 880 191008 239120 191288
rect 800 190336 239322 191008
rect 880 190056 239120 190336
rect 800 189248 239322 190056
rect 880 188968 239120 189248
rect 800 188160 239322 188968
rect 880 187880 239120 188160
rect 800 187072 239322 187880
rect 880 186792 239120 187072
rect 800 186120 239322 186792
rect 880 185840 239120 186120
rect 800 185032 239322 185840
rect 880 184752 239120 185032
rect 800 183944 239322 184752
rect 880 183664 239120 183944
rect 800 182992 239322 183664
rect 880 182712 239120 182992
rect 800 181904 239322 182712
rect 880 181624 239120 181904
rect 800 180816 239322 181624
rect 880 180536 239120 180816
rect 800 179728 239322 180536
rect 880 179448 239120 179728
rect 800 178776 239322 179448
rect 880 178496 239120 178776
rect 800 177688 239322 178496
rect 880 177408 239120 177688
rect 800 176600 239322 177408
rect 880 176320 239120 176600
rect 800 175648 239322 176320
rect 880 175368 239120 175648
rect 800 174560 239322 175368
rect 880 174280 239120 174560
rect 800 173472 239322 174280
rect 880 173192 239120 173472
rect 800 172520 239322 173192
rect 880 172240 239120 172520
rect 800 171432 239322 172240
rect 880 171152 239120 171432
rect 800 170344 239322 171152
rect 880 170064 239120 170344
rect 800 169256 239322 170064
rect 880 168976 239120 169256
rect 800 168304 239322 168976
rect 880 168024 239120 168304
rect 800 167216 239322 168024
rect 880 166936 239120 167216
rect 800 166128 239322 166936
rect 880 165848 239120 166128
rect 800 165176 239322 165848
rect 880 164896 239120 165176
rect 800 164088 239322 164896
rect 880 163808 239120 164088
rect 800 163000 239322 163808
rect 880 162720 239120 163000
rect 800 161912 239322 162720
rect 880 161632 239120 161912
rect 800 160960 239322 161632
rect 880 160680 239120 160960
rect 800 159872 239322 160680
rect 880 159592 239120 159872
rect 800 158784 239322 159592
rect 880 158504 239120 158784
rect 800 157832 239322 158504
rect 880 157552 239120 157832
rect 800 156744 239322 157552
rect 880 156464 239120 156744
rect 800 155656 239322 156464
rect 880 155376 239120 155656
rect 800 154568 239322 155376
rect 880 154288 239120 154568
rect 800 153616 239322 154288
rect 880 153336 239120 153616
rect 800 152528 239322 153336
rect 880 152248 239120 152528
rect 800 151440 239322 152248
rect 880 151160 239120 151440
rect 800 150488 239322 151160
rect 880 150208 239120 150488
rect 800 149400 239322 150208
rect 880 149120 239120 149400
rect 800 148312 239322 149120
rect 880 148032 239120 148312
rect 800 147360 239322 148032
rect 880 147080 239120 147360
rect 800 146272 239322 147080
rect 880 145992 239120 146272
rect 800 145184 239322 145992
rect 880 144904 239120 145184
rect 800 144096 239322 144904
rect 880 143816 239120 144096
rect 800 143144 239322 143816
rect 880 142864 239120 143144
rect 800 142056 239322 142864
rect 880 141776 239120 142056
rect 800 140968 239322 141776
rect 880 140688 239120 140968
rect 800 140016 239322 140688
rect 880 139736 239120 140016
rect 800 138928 239322 139736
rect 880 138648 239120 138928
rect 800 137840 239322 138648
rect 880 137560 239120 137840
rect 800 136752 239322 137560
rect 880 136472 239120 136752
rect 800 135800 239322 136472
rect 880 135520 239120 135800
rect 800 134712 239322 135520
rect 880 134432 239120 134712
rect 800 133624 239322 134432
rect 880 133344 239120 133624
rect 800 132672 239322 133344
rect 880 132392 239120 132672
rect 800 131584 239322 132392
rect 880 131304 239120 131584
rect 800 130496 239322 131304
rect 880 130216 239120 130496
rect 800 129544 239322 130216
rect 880 129264 239120 129544
rect 800 128456 239322 129264
rect 880 128176 239120 128456
rect 800 127368 239322 128176
rect 880 127088 239120 127368
rect 800 126280 239322 127088
rect 880 126000 239120 126280
rect 800 125328 239322 126000
rect 880 125048 239120 125328
rect 800 124240 239322 125048
rect 880 123960 239120 124240
rect 800 123152 239322 123960
rect 880 122872 239120 123152
rect 800 122200 239322 122872
rect 880 121920 239120 122200
rect 800 121112 239322 121920
rect 880 120832 239120 121112
rect 800 120024 239322 120832
rect 880 119744 239120 120024
rect 800 118936 239322 119744
rect 880 118656 239120 118936
rect 800 117984 239322 118656
rect 880 117704 239120 117984
rect 800 116896 239322 117704
rect 880 116616 239120 116896
rect 800 115808 239322 116616
rect 880 115528 239120 115808
rect 800 114856 239322 115528
rect 880 114576 239120 114856
rect 800 113768 239322 114576
rect 880 113488 239120 113768
rect 800 112680 239322 113488
rect 880 112400 239120 112680
rect 800 111592 239322 112400
rect 880 111312 239120 111592
rect 800 110640 239322 111312
rect 880 110360 239120 110640
rect 800 109552 239322 110360
rect 880 109272 239120 109552
rect 800 108464 239322 109272
rect 880 108184 239120 108464
rect 800 107512 239322 108184
rect 880 107232 239120 107512
rect 800 106424 239322 107232
rect 880 106144 239120 106424
rect 800 105336 239322 106144
rect 880 105056 239120 105336
rect 800 104384 239322 105056
rect 880 104104 239120 104384
rect 800 103296 239322 104104
rect 880 103016 239120 103296
rect 800 102208 239322 103016
rect 880 101928 239120 102208
rect 800 101120 239322 101928
rect 880 100840 239120 101120
rect 800 100168 239322 100840
rect 880 99888 239120 100168
rect 800 99080 239322 99888
rect 880 98800 239120 99080
rect 800 97992 239322 98800
rect 880 97712 239120 97992
rect 800 97040 239322 97712
rect 880 96760 239120 97040
rect 800 95952 239322 96760
rect 880 95672 239120 95952
rect 800 94864 239322 95672
rect 880 94584 239120 94864
rect 800 93776 239322 94584
rect 880 93496 239120 93776
rect 800 92824 239322 93496
rect 880 92544 239120 92824
rect 800 91736 239322 92544
rect 880 91456 239120 91736
rect 800 90648 239322 91456
rect 880 90368 239120 90648
rect 800 89696 239322 90368
rect 880 89416 239120 89696
rect 800 88608 239322 89416
rect 880 88328 239120 88608
rect 800 87520 239322 88328
rect 880 87240 239120 87520
rect 800 86568 239322 87240
rect 880 86288 239120 86568
rect 800 85480 239322 86288
rect 880 85200 239120 85480
rect 800 84392 239322 85200
rect 880 84112 239120 84392
rect 800 83304 239322 84112
rect 880 83024 239120 83304
rect 800 82352 239322 83024
rect 880 82072 239120 82352
rect 800 81264 239322 82072
rect 880 80984 239120 81264
rect 800 80176 239322 80984
rect 880 79896 239120 80176
rect 800 79224 239322 79896
rect 880 78944 239120 79224
rect 800 78136 239322 78944
rect 880 77856 239120 78136
rect 800 77048 239322 77856
rect 880 76768 239120 77048
rect 800 75960 239322 76768
rect 880 75680 239120 75960
rect 800 75008 239322 75680
rect 880 74728 239120 75008
rect 800 73920 239322 74728
rect 880 73640 239120 73920
rect 800 72832 239322 73640
rect 880 72552 239120 72832
rect 800 71880 239322 72552
rect 880 71600 239120 71880
rect 800 70792 239322 71600
rect 880 70512 239120 70792
rect 800 69704 239322 70512
rect 880 69424 239120 69704
rect 800 68616 239322 69424
rect 880 68336 239120 68616
rect 800 67664 239322 68336
rect 880 67384 239120 67664
rect 800 66576 239322 67384
rect 880 66296 239120 66576
rect 800 65488 239322 66296
rect 880 65208 239120 65488
rect 800 64536 239322 65208
rect 880 64256 239120 64536
rect 800 63448 239322 64256
rect 880 63168 239120 63448
rect 800 62360 239322 63168
rect 880 62080 239120 62360
rect 800 61408 239322 62080
rect 880 61128 239120 61408
rect 800 60320 239322 61128
rect 880 60040 239120 60320
rect 800 59232 239322 60040
rect 880 58952 239120 59232
rect 800 58144 239322 58952
rect 880 57864 239120 58144
rect 800 57192 239322 57864
rect 880 56912 239120 57192
rect 800 56104 239322 56912
rect 880 55824 239120 56104
rect 800 55016 239322 55824
rect 880 54736 239120 55016
rect 800 54064 239322 54736
rect 880 53784 239120 54064
rect 800 52976 239322 53784
rect 880 52696 239120 52976
rect 800 51888 239322 52696
rect 880 51608 239120 51888
rect 800 50800 239322 51608
rect 880 50520 239120 50800
rect 800 49848 239322 50520
rect 880 49568 239120 49848
rect 800 48760 239322 49568
rect 880 48480 239120 48760
rect 800 47672 239322 48480
rect 880 47392 239120 47672
rect 800 46720 239322 47392
rect 880 46440 239120 46720
rect 800 45632 239322 46440
rect 880 45352 239120 45632
rect 800 44544 239322 45352
rect 880 44264 239120 44544
rect 800 43592 239322 44264
rect 880 43312 239120 43592
rect 800 42504 239322 43312
rect 880 42224 239120 42504
rect 800 41416 239322 42224
rect 880 41136 239120 41416
rect 800 40328 239322 41136
rect 880 40048 239120 40328
rect 800 39376 239322 40048
rect 880 39096 239120 39376
rect 800 38288 239322 39096
rect 880 38008 239120 38288
rect 800 37200 239322 38008
rect 880 36920 239120 37200
rect 800 36248 239322 36920
rect 880 35968 239120 36248
rect 800 35160 239322 35968
rect 880 34880 239120 35160
rect 800 34072 239322 34880
rect 880 33792 239120 34072
rect 800 32984 239322 33792
rect 880 32704 239120 32984
rect 800 32032 239322 32704
rect 880 31752 239120 32032
rect 800 30944 239322 31752
rect 880 30664 239120 30944
rect 800 29856 239322 30664
rect 880 29576 239120 29856
rect 800 28904 239322 29576
rect 880 28624 239120 28904
rect 800 27816 239322 28624
rect 880 27536 239120 27816
rect 800 26728 239322 27536
rect 880 26448 239120 26728
rect 800 25640 239322 26448
rect 880 25360 239120 25640
rect 800 24688 239322 25360
rect 880 24408 239120 24688
rect 800 23600 239322 24408
rect 880 23320 239120 23600
rect 800 22512 239322 23320
rect 880 22232 239120 22512
rect 800 21560 239322 22232
rect 880 21280 239120 21560
rect 800 20472 239322 21280
rect 880 20192 239120 20472
rect 800 19384 239322 20192
rect 880 19104 239120 19384
rect 800 18432 239322 19104
rect 880 18152 239120 18432
rect 800 17344 239322 18152
rect 880 17064 239120 17344
rect 800 16256 239322 17064
rect 880 15976 239120 16256
rect 800 15168 239322 15976
rect 880 14888 239120 15168
rect 800 14216 239322 14888
rect 880 13936 239120 14216
rect 800 13128 239322 13936
rect 880 12848 239120 13128
rect 800 12040 239322 12848
rect 880 11760 239120 12040
rect 800 11088 239322 11760
rect 880 10808 239120 11088
rect 800 10000 239322 10808
rect 880 9720 239120 10000
rect 800 8912 239322 9720
rect 880 8632 239120 8912
rect 800 7824 239322 8632
rect 880 7544 239120 7824
rect 800 6872 239322 7544
rect 880 6592 239120 6872
rect 800 5784 239322 6592
rect 880 5504 239120 5784
rect 800 4696 239322 5504
rect 880 4416 239120 4696
rect 800 3744 239322 4416
rect 880 3464 239120 3744
rect 800 2656 239322 3464
rect 880 2376 239120 2656
rect 800 1568 239322 2376
rect 880 1288 239120 1568
rect 800 616 239322 1288
rect 880 443 239120 616
<< metal4 >>
rect 4208 2128 4528 237776
rect 9208 2128 9528 237776
rect 14208 2128 14528 237776
rect 19208 2128 19528 237776
rect 24208 2128 24528 237776
rect 29208 2128 29528 237776
rect 34208 2128 34528 237776
rect 39208 2128 39528 237776
rect 44208 2128 44528 237776
rect 49208 2128 49528 237776
rect 54208 2128 54528 237776
rect 59208 2128 59528 237776
rect 64208 2128 64528 237776
rect 69208 2128 69528 237776
rect 74208 2128 74528 237776
rect 79208 2128 79528 237776
rect 84208 2128 84528 237776
rect 89208 2128 89528 237776
rect 94208 2128 94528 237776
rect 99208 2128 99528 237776
rect 104208 2128 104528 237776
rect 109208 2128 109528 237776
rect 114208 2128 114528 237776
rect 119208 2128 119528 237776
rect 124208 2128 124528 237776
rect 129208 2128 129528 237776
rect 134208 2128 134528 237776
rect 139208 2128 139528 237776
rect 144208 2128 144528 237776
rect 149208 2128 149528 237776
rect 154208 2128 154528 237776
rect 159208 2128 159528 237776
rect 164208 2128 164528 237776
rect 169208 2128 169528 237776
rect 174208 2128 174528 237776
rect 179208 2128 179528 237776
rect 184208 2128 184528 237776
rect 189208 2128 189528 237776
rect 194208 2128 194528 237776
rect 199208 2128 199528 237776
rect 204208 2128 204528 237776
rect 209208 2128 209528 237776
rect 214208 2128 214528 237776
rect 219208 2128 219528 237776
rect 224208 2128 224528 237776
rect 229208 2128 229528 237776
rect 234208 2128 234528 237776
<< obsm4 >>
rect 28763 16491 29128 237421
rect 29608 16491 34128 237421
rect 34608 16491 39128 237421
rect 39608 16491 44128 237421
rect 44608 16491 49128 237421
rect 49608 16491 54128 237421
rect 54608 16491 59128 237421
rect 59608 16491 64128 237421
rect 64608 16491 69128 237421
rect 69608 16491 74128 237421
rect 74608 16491 79128 237421
rect 79608 16491 84128 237421
rect 84608 16491 89128 237421
rect 89608 16491 94128 237421
rect 94608 16491 99128 237421
rect 99608 16491 104128 237421
rect 104608 16491 109128 237421
rect 109608 16491 114128 237421
rect 114608 16491 119128 237421
rect 119608 16491 124128 237421
rect 124608 16491 129128 237421
rect 129608 16491 134128 237421
rect 134608 16491 139128 237421
rect 139608 16491 142173 237421
<< labels >>
rlabel metal3 s 0 416 800 536 6 alert_major_o
port 1 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 alert_minor_o
port 2 nsew signal output
rlabel metal3 s 239200 5584 240000 5704 6 boot_addr_i[0]
port 3 nsew signal input
rlabel metal3 s 239200 66376 240000 66496 6 boot_addr_i[10]
port 4 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 boot_addr_i[11]
port 5 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 boot_addr_i[12]
port 6 nsew signal input
rlabel metal2 s 85578 239200 85634 240000 6 boot_addr_i[13]
port 7 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 boot_addr_i[14]
port 8 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 boot_addr_i[15]
port 9 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 boot_addr_i[16]
port 10 nsew signal input
rlabel metal2 s 109130 239200 109186 240000 6 boot_addr_i[17]
port 11 nsew signal input
rlabel metal2 s 112258 239200 112314 240000 6 boot_addr_i[18]
port 12 nsew signal input
rlabel metal3 s 239200 117784 240000 117904 6 boot_addr_i[19]
port 13 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 boot_addr_i[1]
port 14 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 boot_addr_i[20]
port 15 nsew signal input
rlabel metal2 s 129646 239200 129702 240000 6 boot_addr_i[21]
port 16 nsew signal input
rlabel metal2 s 136822 239200 136878 240000 6 boot_addr_i[22]
port 17 nsew signal input
rlabel metal3 s 0 132472 800 132592 6 boot_addr_i[23]
port 18 nsew signal input
rlabel metal3 s 239200 137640 240000 137760 6 boot_addr_i[24]
port 19 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 boot_addr_i[25]
port 20 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 boot_addr_i[26]
port 21 nsew signal input
rlabel metal2 s 163502 239200 163558 240000 6 boot_addr_i[27]
port 22 nsew signal input
rlabel metal2 s 168654 239200 168710 240000 6 boot_addr_i[28]
port 23 nsew signal input
rlabel metal2 s 173806 239200 173862 240000 6 boot_addr_i[29]
port 24 nsew signal input
rlabel metal2 s 22006 239200 22062 240000 6 boot_addr_i[2]
port 25 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 boot_addr_i[30]
port 26 nsew signal input
rlabel metal3 s 0 173272 800 173392 6 boot_addr_i[31]
port 27 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 boot_addr_i[3]
port 28 nsew signal input
rlabel metal2 s 32218 239200 32274 240000 6 boot_addr_i[4]
port 29 nsew signal input
rlabel metal2 s 40406 239200 40462 240000 6 boot_addr_i[5]
port 30 nsew signal input
rlabel metal3 s 239200 45432 240000 45552 6 boot_addr_i[6]
port 31 nsew signal input
rlabel metal3 s 239200 50600 240000 50720 6 boot_addr_i[7]
port 32 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 boot_addr_i[8]
port 33 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 boot_addr_i[9]
port 34 nsew signal input
rlabel metal2 s 478 239200 534 240000 6 clk_i
port 35 nsew signal input
rlabel metal3 s 239200 416 240000 536 6 core_busy_o
port 36 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 crash_dump_o[0]
port 37 nsew signal output
rlabel metal3 s 239200 227808 240000 227928 6 crash_dump_o[100]
port 38 nsew signal output
rlabel metal2 s 223854 0 223910 800 6 crash_dump_o[101]
port 39 nsew signal output
rlabel metal3 s 239200 228896 240000 229016 6 crash_dump_o[102]
port 40 nsew signal output
rlabel metal2 s 229190 239200 229246 240000 6 crash_dump_o[103]
port 41 nsew signal output
rlabel metal2 s 230202 239200 230258 240000 6 crash_dump_o[104]
port 42 nsew signal output
rlabel metal3 s 0 226720 800 226840 6 crash_dump_o[105]
port 43 nsew signal output
rlabel metal3 s 0 227808 800 227928 6 crash_dump_o[106]
port 44 nsew signal output
rlabel metal2 s 227534 0 227590 800 6 crash_dump_o[107]
port 45 nsew signal output
rlabel metal3 s 0 229848 800 229968 6 crash_dump_o[108]
port 46 nsew signal output
rlabel metal3 s 239200 232024 240000 232144 6 crash_dump_o[109]
port 47 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 crash_dump_o[10]
port 48 nsew signal output
rlabel metal2 s 229374 0 229430 800 6 crash_dump_o[110]
port 49 nsew signal output
rlabel metal2 s 230294 0 230350 800 6 crash_dump_o[111]
port 50 nsew signal output
rlabel metal3 s 239200 233112 240000 233232 6 crash_dump_o[112]
port 51 nsew signal output
rlabel metal2 s 231214 0 231270 800 6 crash_dump_o[113]
port 52 nsew signal output
rlabel metal2 s 233238 239200 233294 240000 6 crash_dump_o[114]
port 53 nsew signal output
rlabel metal3 s 0 233112 800 233232 6 crash_dump_o[115]
port 54 nsew signal output
rlabel metal2 s 234342 239200 234398 240000 6 crash_dump_o[116]
port 55 nsew signal output
rlabel metal2 s 233054 0 233110 800 6 crash_dump_o[117]
port 56 nsew signal output
rlabel metal2 s 233974 0 234030 800 6 crash_dump_o[118]
port 57 nsew signal output
rlabel metal3 s 0 236240 800 236360 6 crash_dump_o[119]
port 58 nsew signal output
rlabel metal3 s 239200 72632 240000 72752 6 crash_dump_o[11]
port 59 nsew signal output
rlabel metal2 s 236366 239200 236422 240000 6 crash_dump_o[120]
port 60 nsew signal output
rlabel metal3 s 239200 237192 240000 237312 6 crash_dump_o[121]
port 61 nsew signal output
rlabel metal2 s 236734 0 236790 800 6 crash_dump_o[122]
port 62 nsew signal output
rlabel metal2 s 237378 239200 237434 240000 6 crash_dump_o[123]
port 63 nsew signal output
rlabel metal3 s 239200 238280 240000 238400 6 crash_dump_o[124]
port 64 nsew signal output
rlabel metal2 s 238390 239200 238446 240000 6 crash_dump_o[125]
port 65 nsew signal output
rlabel metal3 s 0 238280 800 238400 6 crash_dump_o[126]
port 66 nsew signal output
rlabel metal2 s 239494 0 239550 800 6 crash_dump_o[127]
port 67 nsew signal output
rlabel metal3 s 239200 79976 240000 80096 6 crash_dump_o[12]
port 68 nsew signal output
rlabel metal2 s 86590 239200 86646 240000 6 crash_dump_o[13]
port 69 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 crash_dump_o[14]
port 70 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 crash_dump_o[15]
port 71 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 crash_dump_o[16]
port 72 nsew signal output
rlabel metal3 s 239200 105136 240000 105256 6 crash_dump_o[17]
port 73 nsew signal output
rlabel metal2 s 113270 239200 113326 240000 6 crash_dump_o[18]
port 74 nsew signal output
rlabel metal2 s 118422 239200 118478 240000 6 crash_dump_o[19]
port 75 nsew signal output
rlabel metal2 s 14830 239200 14886 240000 6 crash_dump_o[1]
port 76 nsew signal output
rlabel metal2 s 124586 239200 124642 240000 6 crash_dump_o[20]
port 77 nsew signal output
rlabel metal2 s 130658 239200 130714 240000 6 crash_dump_o[21]
port 78 nsew signal output
rlabel metal3 s 239200 131384 240000 131504 6 crash_dump_o[22]
port 79 nsew signal output
rlabel metal2 s 138662 0 138718 800 6 crash_dump_o[23]
port 80 nsew signal output
rlabel metal2 s 144182 0 144238 800 6 crash_dump_o[24]
port 81 nsew signal output
rlabel metal2 s 153290 239200 153346 240000 6 crash_dump_o[25]
port 82 nsew signal output
rlabel metal2 s 157338 239200 157394 240000 6 crash_dump_o[26]
port 83 nsew signal output
rlabel metal3 s 0 150288 800 150408 6 crash_dump_o[27]
port 84 nsew signal output
rlabel metal3 s 239200 160760 240000 160880 6 crash_dump_o[28]
port 85 nsew signal output
rlabel metal3 s 239200 161712 240000 161832 6 crash_dump_o[29]
port 86 nsew signal output
rlabel metal3 s 239200 21360 240000 21480 6 crash_dump_o[2]
port 87 nsew signal output
rlabel metal2 s 177854 239200 177910 240000 6 crash_dump_o[30]
port 88 nsew signal output
rlabel metal2 s 180982 239200 181038 240000 6 crash_dump_o[31]
port 89 nsew signal output
rlabel metal2 s 186134 239200 186190 240000 6 crash_dump_o[32]
port 90 nsew signal output
rlabel metal3 s 239200 175448 240000 175568 6 crash_dump_o[33]
port 91 nsew signal output
rlabel metal3 s 0 178576 800 178696 6 crash_dump_o[34]
port 92 nsew signal output
rlabel metal3 s 239200 179528 240000 179648 6 crash_dump_o[35]
port 93 nsew signal output
rlabel metal2 s 185398 0 185454 800 6 crash_dump_o[36]
port 94 nsew signal output
rlabel metal3 s 0 182792 800 182912 6 crash_dump_o[37]
port 95 nsew signal output
rlabel metal2 s 187238 0 187294 800 6 crash_dump_o[38]
port 96 nsew signal output
rlabel metal2 s 194322 239200 194378 240000 6 crash_dump_o[39]
port 97 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 crash_dump_o[3]
port 98 nsew signal output
rlabel metal3 s 0 184832 800 184952 6 crash_dump_o[40]
port 99 nsew signal output
rlabel metal2 s 197358 239200 197414 240000 6 crash_dump_o[41]
port 100 nsew signal output
rlabel metal3 s 239200 184832 240000 184952 6 crash_dump_o[42]
port 101 nsew signal output
rlabel metal3 s 0 186872 800 186992 6 crash_dump_o[43]
port 102 nsew signal output
rlabel metal3 s 239200 189048 240000 189168 6 crash_dump_o[44]
port 103 nsew signal output
rlabel metal2 s 200486 239200 200542 240000 6 crash_dump_o[45]
port 104 nsew signal output
rlabel metal3 s 0 191088 800 191208 6 crash_dump_o[46]
port 105 nsew signal output
rlabel metal3 s 0 193264 800 193384 6 crash_dump_o[47]
port 106 nsew signal output
rlabel metal3 s 0 194216 800 194336 6 crash_dump_o[48]
port 107 nsew signal output
rlabel metal3 s 239200 195304 240000 195424 6 crash_dump_o[49]
port 108 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 crash_dump_o[4]
port 109 nsew signal output
rlabel metal2 s 202510 239200 202566 240000 6 crash_dump_o[50]
port 110 nsew signal output
rlabel metal2 s 196438 0 196494 800 6 crash_dump_o[51]
port 111 nsew signal output
rlabel metal3 s 0 195304 800 195424 6 crash_dump_o[52]
port 112 nsew signal output
rlabel metal3 s 0 196392 800 196512 6 crash_dump_o[53]
port 113 nsew signal output
rlabel metal2 s 199106 0 199162 800 6 crash_dump_o[54]
port 114 nsew signal output
rlabel metal2 s 206650 239200 206706 240000 6 crash_dump_o[55]
port 115 nsew signal output
rlabel metal2 s 207662 239200 207718 240000 6 crash_dump_o[56]
port 116 nsew signal output
rlabel metal3 s 239200 202648 240000 202768 6 crash_dump_o[57]
port 117 nsew signal output
rlabel metal3 s 0 200608 800 200728 6 crash_dump_o[58]
port 118 nsew signal output
rlabel metal2 s 200946 0 201002 800 6 crash_dump_o[59]
port 119 nsew signal output
rlabel metal3 s 239200 39176 240000 39296 6 crash_dump_o[5]
port 120 nsew signal output
rlabel metal3 s 0 203736 800 203856 6 crash_dump_o[60]
port 121 nsew signal output
rlabel metal3 s 0 204688 800 204808 6 crash_dump_o[61]
port 122 nsew signal output
rlabel metal2 s 201866 0 201922 800 6 crash_dump_o[62]
port 123 nsew signal output
rlabel metal2 s 213826 239200 213882 240000 6 crash_dump_o[63]
port 124 nsew signal output
rlabel metal3 s 0 208904 800 209024 6 crash_dump_o[64]
port 125 nsew signal output
rlabel metal2 s 214838 239200 214894 240000 6 crash_dump_o[65]
port 126 nsew signal output
rlabel metal2 s 216862 239200 216918 240000 6 crash_dump_o[66]
port 127 nsew signal output
rlabel metal2 s 203706 0 203762 800 6 crash_dump_o[67]
port 128 nsew signal output
rlabel metal3 s 0 209992 800 210112 6 crash_dump_o[68]
port 129 nsew signal output
rlabel metal2 s 205546 0 205602 800 6 crash_dump_o[69]
port 130 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 crash_dump_o[6]
port 131 nsew signal output
rlabel metal2 s 217874 239200 217930 240000 6 crash_dump_o[70]
port 132 nsew signal output
rlabel metal2 s 218886 239200 218942 240000 6 crash_dump_o[71]
port 133 nsew signal output
rlabel metal3 s 239200 209992 240000 210112 6 crash_dump_o[72]
port 134 nsew signal output
rlabel metal3 s 0 213120 800 213240 6 crash_dump_o[73]
port 135 nsew signal output
rlabel metal2 s 222014 239200 222070 240000 6 crash_dump_o[74]
port 136 nsew signal output
rlabel metal2 s 206466 0 206522 800 6 crash_dump_o[75]
port 137 nsew signal output
rlabel metal3 s 239200 211080 240000 211200 6 crash_dump_o[76]
port 138 nsew signal output
rlabel metal2 s 208306 0 208362 800 6 crash_dump_o[77]
port 139 nsew signal output
rlabel metal3 s 0 215296 800 215416 6 crash_dump_o[78]
port 140 nsew signal output
rlabel metal3 s 0 216248 800 216368 6 crash_dump_o[79]
port 141 nsew signal output
rlabel metal3 s 239200 51688 240000 51808 6 crash_dump_o[7]
port 142 nsew signal output
rlabel metal3 s 239200 213120 240000 213240 6 crash_dump_o[80]
port 143 nsew signal output
rlabel metal3 s 239200 214208 240000 214328 6 crash_dump_o[81]
port 144 nsew signal output
rlabel metal3 s 239200 215296 240000 215416 6 crash_dump_o[82]
port 145 nsew signal output
rlabel metal3 s 239200 216248 240000 216368 6 crash_dump_o[83]
port 146 nsew signal output
rlabel metal2 s 212906 0 212962 800 6 crash_dump_o[84]
port 147 nsew signal output
rlabel metal2 s 224038 239200 224094 240000 6 crash_dump_o[85]
port 148 nsew signal output
rlabel metal3 s 0 219376 800 219496 6 crash_dump_o[86]
port 149 nsew signal output
rlabel metal3 s 0 220464 800 220584 6 crash_dump_o[87]
port 150 nsew signal output
rlabel metal3 s 239200 217336 240000 217456 6 crash_dump_o[88]
port 151 nsew signal output
rlabel metal3 s 239200 218424 240000 218544 6 crash_dump_o[89]
port 152 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 crash_dump_o[8]
port 153 nsew signal output
rlabel metal2 s 215666 0 215722 800 6 crash_dump_o[90]
port 154 nsew signal output
rlabel metal2 s 217506 0 217562 800 6 crash_dump_o[91]
port 155 nsew signal output
rlabel metal2 s 218426 0 218482 800 6 crash_dump_o[92]
port 156 nsew signal output
rlabel metal3 s 239200 220464 240000 220584 6 crash_dump_o[93]
port 157 nsew signal output
rlabel metal3 s 0 223592 800 223712 6 crash_dump_o[94]
port 158 nsew signal output
rlabel metal2 s 221094 0 221150 800 6 crash_dump_o[95]
port 159 nsew signal output
rlabel metal2 s 222014 0 222070 800 6 crash_dump_o[96]
port 160 nsew signal output
rlabel metal3 s 239200 223592 240000 223712 6 crash_dump_o[97]
port 161 nsew signal output
rlabel metal3 s 239200 224680 240000 224800 6 crash_dump_o[98]
port 162 nsew signal output
rlabel metal3 s 239200 225768 240000 225888 6 crash_dump_o[99]
port 163 nsew signal output
rlabel metal2 s 68098 239200 68154 240000 6 crash_dump_o[9]
port 164 nsew signal output
rlabel metal2 s 5538 239200 5594 240000 6 data_addr_o[0]
port 165 nsew signal output
rlabel metal3 s 0 75760 800 75880 6 data_addr_o[10]
port 166 nsew signal output
rlabel metal3 s 0 79024 800 79144 6 data_addr_o[11]
port 167 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 data_addr_o[12]
port 168 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 data_addr_o[13]
port 169 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 data_addr_o[14]
port 170 nsew signal output
rlabel metal3 s 239200 89496 240000 89616 6 data_addr_o[15]
port 171 nsew signal output
rlabel metal2 s 104070 239200 104126 240000 6 data_addr_o[16]
port 172 nsew signal output
rlabel metal2 s 110234 239200 110290 240000 6 data_addr_o[17]
port 173 nsew signal output
rlabel metal3 s 239200 110440 240000 110560 6 data_addr_o[18]
port 174 nsew signal output
rlabel metal3 s 239200 118736 240000 118856 6 data_addr_o[19]
port 175 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 data_addr_o[1]
port 176 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 data_addr_o[20]
port 177 nsew signal output
rlabel metal2 s 131762 239200 131818 240000 6 data_addr_o[21]
port 178 nsew signal output
rlabel metal3 s 0 128256 800 128376 6 data_addr_o[22]
port 179 nsew signal output
rlabel metal3 s 0 133424 800 133544 6 data_addr_o[23]
port 180 nsew signal output
rlabel metal3 s 239200 138728 240000 138848 6 data_addr_o[24]
port 181 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 data_addr_o[25]
port 182 nsew signal output
rlabel metal3 s 239200 150288 240000 150408 6 data_addr_o[26]
port 183 nsew signal output
rlabel metal2 s 164514 239200 164570 240000 6 data_addr_o[27]
port 184 nsew signal output
rlabel metal3 s 0 153416 800 153536 6 data_addr_o[28]
port 185 nsew signal output
rlabel metal3 s 0 158584 800 158704 6 data_addr_o[29]
port 186 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 data_addr_o[2]
port 187 nsew signal output
rlabel metal3 s 0 167016 800 167136 6 data_addr_o[30]
port 188 nsew signal output
rlabel metal3 s 0 174360 800 174480 6 data_addr_o[31]
port 189 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 data_addr_o[3]
port 190 nsew signal output
rlabel metal2 s 33230 239200 33286 240000 6 data_addr_o[4]
port 191 nsew signal output
rlabel metal3 s 239200 40128 240000 40248 6 data_addr_o[5]
port 192 nsew signal output
rlabel metal3 s 239200 46520 240000 46640 6 data_addr_o[6]
port 193 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 data_addr_o[7]
port 194 nsew signal output
rlabel metal2 s 59910 239200 59966 240000 6 data_addr_o[8]
port 195 nsew signal output
rlabel metal2 s 69202 239200 69258 240000 6 data_addr_o[9]
port 196 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 data_be_o[0]
port 197 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 data_be_o[1]
port 198 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 data_be_o[2]
port 199 nsew signal output
rlabel metal3 s 239200 27616 240000 27736 6 data_be_o[3]
port 200 nsew signal output
rlabel metal2 s 1490 239200 1546 240000 6 data_err_i
port 201 nsew signal input
rlabel metal2 s 2502 239200 2558 240000 6 data_gnt_i
port 202 nsew signal input
rlabel metal2 s 6550 239200 6606 240000 6 data_rdata_i[0]
port 203 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 data_rdata_i[10]
port 204 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 data_rdata_i[11]
port 205 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 data_rdata_i[12]
port 206 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 data_rdata_i[13]
port 207 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 data_rdata_i[14]
port 208 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 data_rdata_i[15]
port 209 nsew signal input
rlabel metal2 s 105082 239200 105138 240000 6 data_rdata_i[16]
port 210 nsew signal input
rlabel metal3 s 239200 106224 240000 106344 6 data_rdata_i[17]
port 211 nsew signal input
rlabel metal2 s 114282 239200 114338 240000 6 data_rdata_i[18]
port 212 nsew signal input
rlabel metal3 s 239200 119824 240000 119944 6 data_rdata_i[19]
port 213 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 data_rdata_i[1]
port 214 nsew signal input
rlabel metal3 s 0 118736 800 118856 6 data_rdata_i[20]
port 215 nsew signal input
rlabel metal3 s 239200 127168 240000 127288 6 data_rdata_i[21]
port 216 nsew signal input
rlabel metal3 s 0 129344 800 129464 6 data_rdata_i[22]
port 217 nsew signal input
rlabel metal2 s 145102 239200 145158 240000 6 data_rdata_i[23]
port 218 nsew signal input
rlabel metal3 s 239200 139816 240000 139936 6 data_rdata_i[24]
port 219 nsew signal input
rlabel metal2 s 154302 239200 154358 240000 6 data_rdata_i[25]
port 220 nsew signal input
rlabel metal3 s 0 146072 800 146192 6 data_rdata_i[26]
port 221 nsew signal input
rlabel metal3 s 0 151240 800 151360 6 data_rdata_i[27]
port 222 nsew signal input
rlabel metal3 s 0 154368 800 154488 6 data_rdata_i[28]
port 223 nsew signal input
rlabel metal2 s 174818 239200 174874 240000 6 data_rdata_i[29]
port 224 nsew signal input
rlabel metal3 s 239200 22312 240000 22432 6 data_rdata_i[2]
port 225 nsew signal input
rlabel metal3 s 239200 164976 240000 165096 6 data_rdata_i[30]
port 226 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 data_rdata_i[31]
port 227 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 data_rdata_i[3]
port 228 nsew signal input
rlabel metal3 s 239200 32784 240000 32904 6 data_rdata_i[4]
port 229 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 data_rdata_i[5]
port 230 nsew signal input
rlabel metal3 s 239200 47472 240000 47592 6 data_rdata_i[6]
port 231 nsew signal input
rlabel metal2 s 52734 239200 52790 240000 6 data_rdata_i[7]
port 232 nsew signal input
rlabel metal3 s 239200 57944 240000 58064 6 data_rdata_i[8]
port 233 nsew signal input
rlabel metal3 s 239200 61208 240000 61328 6 data_rdata_i[9]
port 234 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 data_req_o
port 235 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 data_rvalid_i
port 236 nsew signal input
rlabel metal3 s 239200 6672 240000 6792 6 data_wdata_o[0]
port 237 nsew signal output
rlabel metal3 s 239200 67464 240000 67584 6 data_wdata_o[10]
port 238 nsew signal output
rlabel metal2 s 76378 239200 76434 240000 6 data_wdata_o[11]
port 239 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 data_wdata_o[12]
port 240 nsew signal output
rlabel metal2 s 87602 239200 87658 240000 6 data_wdata_o[13]
port 241 nsew signal output
rlabel metal2 s 93766 239200 93822 240000 6 data_wdata_o[14]
port 242 nsew signal output
rlabel metal3 s 239200 90448 240000 90568 6 data_wdata_o[15]
port 243 nsew signal output
rlabel metal3 s 239200 97792 240000 97912 6 data_wdata_o[16]
port 244 nsew signal output
rlabel metal2 s 111246 239200 111302 240000 6 data_wdata_o[17]
port 245 nsew signal output
rlabel metal2 s 115294 239200 115350 240000 6 data_wdata_o[18]
port 246 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 data_wdata_o[19]
port 247 nsew signal output
rlabel metal2 s 15842 239200 15898 240000 6 data_wdata_o[1]
port 248 nsew signal output
rlabel metal2 s 125598 239200 125654 240000 6 data_wdata_o[20]
port 249 nsew signal output
rlabel metal2 s 132774 239200 132830 240000 6 data_wdata_o[21]
port 250 nsew signal output
rlabel metal2 s 137926 239200 137982 240000 6 data_wdata_o[22]
port 251 nsew signal output
rlabel metal2 s 146114 239200 146170 240000 6 data_wdata_o[23]
port 252 nsew signal output
rlabel metal3 s 239200 140768 240000 140888 6 data_wdata_o[24]
port 253 nsew signal output
rlabel metal3 s 239200 146072 240000 146192 6 data_wdata_o[25]
port 254 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 data_wdata_o[26]
port 255 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 data_wdata_o[27]
port 256 nsew signal output
rlabel metal2 s 164330 0 164386 800 6 data_wdata_o[28]
port 257 nsew signal output
rlabel metal3 s 0 159672 800 159792 6 data_wdata_o[29]
port 258 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 data_wdata_o[2]
port 259 nsew signal output
rlabel metal3 s 0 168104 800 168224 6 data_wdata_o[30]
port 260 nsew signal output
rlabel metal3 s 0 175448 800 175568 6 data_wdata_o[31]
port 261 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 data_wdata_o[3]
port 262 nsew signal output
rlabel metal3 s 239200 33872 240000 33992 6 data_wdata_o[4]
port 263 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 data_wdata_o[5]
port 264 nsew signal output
rlabel metal2 s 46570 239200 46626 240000 6 data_wdata_o[6]
port 265 nsew signal output
rlabel metal2 s 53746 239200 53802 240000 6 data_wdata_o[7]
port 266 nsew signal output
rlabel metal2 s 60922 239200 60978 240000 6 data_wdata_o[8]
port 267 nsew signal output
rlabel metal3 s 0 68416 800 68536 6 data_wdata_o[9]
port 268 nsew signal output
rlabel metal3 s 239200 1368 240000 1488 6 data_we_o
port 269 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 debug_req_i
port 270 nsew signal input
rlabel metal3 s 239200 2456 240000 2576 6 dummy_instr_id_o
port 271 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 eFPGA_delay_o[0]
port 272 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 eFPGA_delay_o[1]
port 273 nsew signal output
rlabel metal2 s 23018 239200 23074 240000 6 eFPGA_delay_o[2]
port 274 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 eFPGA_delay_o[3]
port 275 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 eFPGA_en_o
port 276 nsew signal output
rlabel metal3 s 239200 3544 240000 3664 6 eFPGA_fpga_done_i
port 277 nsew signal input
rlabel metal2 s 7654 239200 7710 240000 6 eFPGA_operand_a_o[0]
port 278 nsew signal output
rlabel metal3 s 239200 68416 240000 68536 6 eFPGA_operand_a_o[10]
port 279 nsew signal output
rlabel metal3 s 239200 73720 240000 73840 6 eFPGA_operand_a_o[11]
port 280 nsew signal output
rlabel metal3 s 239200 81064 240000 81184 6 eFPGA_operand_a_o[12]
port 281 nsew signal output
rlabel metal2 s 88614 239200 88670 240000 6 eFPGA_operand_a_o[13]
port 282 nsew signal output
rlabel metal3 s 239200 87320 240000 87440 6 eFPGA_operand_a_o[14]
port 283 nsew signal output
rlabel metal2 s 99930 239200 99986 240000 6 eFPGA_operand_a_o[15]
port 284 nsew signal output
rlabel metal3 s 239200 98880 240000 99000 6 eFPGA_operand_a_o[16]
port 285 nsew signal output
rlabel metal2 s 110234 0 110290 800 6 eFPGA_operand_a_o[17]
port 286 nsew signal output
rlabel metal3 s 239200 111392 240000 111512 6 eFPGA_operand_a_o[18]
port 287 nsew signal output
rlabel metal2 s 119434 239200 119490 240000 6 eFPGA_operand_a_o[19]
port 288 nsew signal output
rlabel metal3 s 0 19184 800 19304 6 eFPGA_operand_a_o[1]
port 289 nsew signal output
rlabel metal2 s 126794 0 126850 800 6 eFPGA_operand_a_o[20]
port 290 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 eFPGA_operand_a_o[21]
port 291 nsew signal output
rlabel metal2 s 138938 239200 138994 240000 6 eFPGA_operand_a_o[22]
port 292 nsew signal output
rlabel metal2 s 147126 239200 147182 240000 6 eFPGA_operand_a_o[23]
port 293 nsew signal output
rlabel metal3 s 0 139816 800 139936 6 eFPGA_operand_a_o[24]
port 294 nsew signal output
rlabel metal2 s 155314 239200 155370 240000 6 eFPGA_operand_a_o[25]
port 295 nsew signal output
rlabel metal3 s 239200 151240 240000 151360 6 eFPGA_operand_a_o[26]
port 296 nsew signal output
rlabel metal2 s 157890 0 157946 800 6 eFPGA_operand_a_o[27]
port 297 nsew signal output
rlabel metal2 s 169666 239200 169722 240000 6 eFPGA_operand_a_o[28]
port 298 nsew signal output
rlabel metal3 s 239200 162800 240000 162920 6 eFPGA_operand_a_o[29]
port 299 nsew signal output
rlabel metal3 s 239200 23400 240000 23520 6 eFPGA_operand_a_o[2]
port 300 nsew signal output
rlabel metal3 s 0 169056 800 169176 6 eFPGA_operand_a_o[30]
port 301 nsew signal output
rlabel metal2 s 180798 0 180854 800 6 eFPGA_operand_a_o[31]
port 302 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 eFPGA_operand_a_o[3]
port 303 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 eFPGA_operand_a_o[4]
port 304 nsew signal output
rlabel metal2 s 41418 239200 41474 240000 6 eFPGA_operand_a_o[5]
port 305 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 eFPGA_operand_a_o[6]
port 306 nsew signal output
rlabel metal2 s 54758 239200 54814 240000 6 eFPGA_operand_a_o[7]
port 307 nsew signal output
rlabel metal2 s 61934 239200 61990 240000 6 eFPGA_operand_a_o[8]
port 308 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 eFPGA_operand_a_o[9]
port 309 nsew signal output
rlabel metal3 s 239200 7624 240000 7744 6 eFPGA_operand_b_o[0]
port 310 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 eFPGA_operand_b_o[10]
port 311 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 eFPGA_operand_b_o[11]
port 312 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 eFPGA_operand_b_o[12]
port 313 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 eFPGA_operand_b_o[13]
port 314 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 eFPGA_operand_b_o[14]
port 315 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 eFPGA_operand_b_o[15]
port 316 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 eFPGA_operand_b_o[16]
port 317 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 eFPGA_operand_b_o[17]
port 318 nsew signal output
rlabel metal3 s 239200 112480 240000 112600 6 eFPGA_operand_b_o[18]
port 319 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 eFPGA_operand_b_o[19]
port 320 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 eFPGA_operand_b_o[1]
port 321 nsew signal output
rlabel metal3 s 0 119824 800 119944 6 eFPGA_operand_b_o[20]
port 322 nsew signal output
rlabel metal2 s 133786 239200 133842 240000 6 eFPGA_operand_b_o[21]
port 323 nsew signal output
rlabel metal3 s 0 130296 800 130416 6 eFPGA_operand_b_o[22]
port 324 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 eFPGA_operand_b_o[23]
port 325 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 eFPGA_operand_b_o[24]
port 326 nsew signal output
rlabel metal3 s 0 141856 800 141976 6 eFPGA_operand_b_o[25]
port 327 nsew signal output
rlabel metal3 s 239200 152328 240000 152448 6 eFPGA_operand_b_o[26]
port 328 nsew signal output
rlabel metal3 s 239200 157632 240000 157752 6 eFPGA_operand_b_o[27]
port 329 nsew signal output
rlabel metal3 s 0 155456 800 155576 6 eFPGA_operand_b_o[28]
port 330 nsew signal output
rlabel metal3 s 0 160760 800 160880 6 eFPGA_operand_b_o[29]
port 331 nsew signal output
rlabel metal2 s 24030 239200 24086 240000 6 eFPGA_operand_b_o[2]
port 332 nsew signal output
rlabel metal3 s 239200 165928 240000 166048 6 eFPGA_operand_b_o[30]
port 333 nsew signal output
rlabel metal3 s 0 176400 800 176520 6 eFPGA_operand_b_o[31]
port 334 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 eFPGA_operand_b_o[3]
port 335 nsew signal output
rlabel metal2 s 34242 239200 34298 240000 6 eFPGA_operand_b_o[4]
port 336 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 eFPGA_operand_b_o[5]
port 337 nsew signal output
rlabel metal3 s 0 54816 800 54936 6 eFPGA_operand_b_o[6]
port 338 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 eFPGA_operand_b_o[7]
port 339 nsew signal output
rlabel metal2 s 63038 239200 63094 240000 6 eFPGA_operand_b_o[8]
port 340 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 eFPGA_operand_b_o[9]
port 341 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 eFPGA_operator_o[0]
port 342 nsew signal output
rlabel metal3 s 239200 16056 240000 16176 6 eFPGA_operator_o[1]
port 343 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 eFPGA_result_a_i[0]
port 344 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 eFPGA_result_a_i[10]
port 345 nsew signal input
rlabel metal3 s 239200 74808 240000 74928 6 eFPGA_result_a_i[11]
port 346 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 eFPGA_result_a_i[12]
port 347 nsew signal input
rlabel metal2 s 89718 239200 89774 240000 6 eFPGA_result_a_i[13]
port 348 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 eFPGA_result_a_i[14]
port 349 nsew signal input
rlabel metal2 s 100942 239200 100998 240000 6 eFPGA_result_a_i[15]
port 350 nsew signal input
rlabel metal2 s 106094 239200 106150 240000 6 eFPGA_result_a_i[16]
port 351 nsew signal input
rlabel metal3 s 0 107312 800 107432 6 eFPGA_result_a_i[17]
port 352 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 eFPGA_result_a_i[18]
port 353 nsew signal input
rlabel metal2 s 120446 239200 120502 240000 6 eFPGA_result_a_i[19]
port 354 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 eFPGA_result_a_i[1]
port 355 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 eFPGA_result_a_i[20]
port 356 nsew signal input
rlabel metal3 s 0 124040 800 124160 6 eFPGA_result_a_i[21]
port 357 nsew signal input
rlabel metal2 s 139950 239200 140006 240000 6 eFPGA_result_a_i[22]
port 358 nsew signal input
rlabel metal3 s 239200 135600 240000 135720 6 eFPGA_result_a_i[23]
port 359 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 eFPGA_result_a_i[24]
port 360 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 eFPGA_result_a_i[25]
port 361 nsew signal input
rlabel metal3 s 239200 153416 240000 153536 6 eFPGA_result_a_i[26]
port 362 nsew signal input
rlabel metal3 s 239200 158584 240000 158704 6 eFPGA_result_a_i[27]
port 363 nsew signal input
rlabel metal3 s 0 156544 800 156664 6 eFPGA_result_a_i[28]
port 364 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 eFPGA_result_a_i[29]
port 365 nsew signal input
rlabel metal3 s 239200 24488 240000 24608 6 eFPGA_result_a_i[2]
port 366 nsew signal input
rlabel metal3 s 0 170144 800 170264 6 eFPGA_result_a_i[30]
port 367 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 eFPGA_result_a_i[31]
port 368 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 eFPGA_result_a_i[3]
port 369 nsew signal input
rlabel metal2 s 35346 239200 35402 240000 6 eFPGA_result_a_i[4]
port 370 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 eFPGA_result_a_i[5]
port 371 nsew signal input
rlabel metal3 s 239200 48560 240000 48680 6 eFPGA_result_a_i[6]
port 372 nsew signal input
rlabel metal2 s 55862 239200 55918 240000 6 eFPGA_result_a_i[7]
port 373 nsew signal input
rlabel metal3 s 239200 59032 240000 59152 6 eFPGA_result_a_i[8]
port 374 nsew signal input
rlabel metal2 s 70214 239200 70270 240000 6 eFPGA_result_a_i[9]
port 375 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 eFPGA_result_b_i[0]
port 376 nsew signal input
rlabel metal2 s 72238 239200 72294 240000 6 eFPGA_result_b_i[10]
port 377 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 eFPGA_result_b_i[11]
port 378 nsew signal input
rlabel metal2 s 80426 239200 80482 240000 6 eFPGA_result_b_i[12]
port 379 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 eFPGA_result_b_i[13]
port 380 nsew signal input
rlabel metal3 s 0 97792 800 97912 6 eFPGA_result_b_i[14]
port 381 nsew signal input
rlabel metal3 s 239200 91536 240000 91656 6 eFPGA_result_b_i[15]
port 382 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 eFPGA_result_b_i[16]
port 383 nsew signal input
rlabel metal3 s 239200 107312 240000 107432 6 eFPGA_result_b_i[17]
port 384 nsew signal input
rlabel metal3 s 0 114656 800 114776 6 eFPGA_result_b_i[18]
port 385 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 eFPGA_result_b_i[19]
port 386 nsew signal input
rlabel metal3 s 239200 17144 240000 17264 6 eFPGA_result_b_i[1]
port 387 nsew signal input
rlabel metal3 s 239200 124040 240000 124160 6 eFPGA_result_b_i[20]
port 388 nsew signal input
rlabel metal3 s 239200 128256 240000 128376 6 eFPGA_result_b_i[21]
port 389 nsew signal input
rlabel metal3 s 239200 132472 240000 132592 6 eFPGA_result_b_i[22]
port 390 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 eFPGA_result_b_i[23]
port 391 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 eFPGA_result_b_i[24]
port 392 nsew signal input
rlabel metal3 s 239200 147160 240000 147280 6 eFPGA_result_b_i[25]
port 393 nsew signal input
rlabel metal2 s 158442 239200 158498 240000 6 eFPGA_result_b_i[26]
port 394 nsew signal input
rlabel metal3 s 0 152328 800 152448 6 eFPGA_result_b_i[27]
port 395 nsew signal input
rlabel metal2 s 170678 239200 170734 240000 6 eFPGA_result_b_i[28]
port 396 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 eFPGA_result_b_i[29]
port 397 nsew signal input
rlabel metal2 s 25042 239200 25098 240000 6 eFPGA_result_b_i[2]
port 398 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 eFPGA_result_b_i[30]
port 399 nsew signal input
rlabel metal3 s 239200 170144 240000 170264 6 eFPGA_result_b_i[31]
port 400 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 eFPGA_result_b_i[3]
port 401 nsew signal input
rlabel metal3 s 239200 34960 240000 35080 6 eFPGA_result_b_i[4]
port 402 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 eFPGA_result_b_i[5]
port 403 nsew signal input
rlabel metal3 s 0 55904 800 56024 6 eFPGA_result_b_i[6]
port 404 nsew signal input
rlabel metal3 s 239200 52776 240000 52896 6 eFPGA_result_b_i[7]
port 405 nsew signal input
rlabel metal2 s 64050 239200 64106 240000 6 eFPGA_result_b_i[8]
port 406 nsew signal input
rlabel metal3 s 0 69504 800 69624 6 eFPGA_result_b_i[9]
port 407 nsew signal input
rlabel metal3 s 239200 8712 240000 8832 6 eFPGA_result_c_i[0]
port 408 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 eFPGA_result_c_i[10]
port 409 nsew signal input
rlabel metal3 s 239200 75760 240000 75880 6 eFPGA_result_c_i[11]
port 410 nsew signal input
rlabel metal2 s 81438 239200 81494 240000 6 eFPGA_result_c_i[12]
port 411 nsew signal input
rlabel metal3 s 239200 84192 240000 84312 6 eFPGA_result_c_i[13]
port 412 nsew signal input
rlabel metal3 s 0 98880 800 99000 6 eFPGA_result_c_i[14]
port 413 nsew signal input
rlabel metal2 s 101954 239200 102010 240000 6 eFPGA_result_c_i[15]
port 414 nsew signal input
rlabel metal3 s 0 105136 800 105256 6 eFPGA_result_c_i[16]
port 415 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 eFPGA_result_c_i[17]
port 416 nsew signal input
rlabel metal3 s 239200 113568 240000 113688 6 eFPGA_result_c_i[18]
port 417 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 eFPGA_result_c_i[19]
port 418 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 eFPGA_result_c_i[1]
port 419 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 eFPGA_result_c_i[20]
port 420 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 eFPGA_result_c_i[21]
port 421 nsew signal input
rlabel metal2 s 140962 239200 141018 240000 6 eFPGA_result_c_i[22]
port 422 nsew signal input
rlabel metal3 s 239200 136552 240000 136672 6 eFPGA_result_c_i[23]
port 423 nsew signal input
rlabel metal2 s 149150 239200 149206 240000 6 eFPGA_result_c_i[24]
port 424 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 eFPGA_result_c_i[25]
port 425 nsew signal input
rlabel metal3 s 239200 154368 240000 154488 6 eFPGA_result_c_i[26]
port 426 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 eFPGA_result_c_i[27]
port 427 nsew signal input
rlabel metal2 s 171690 239200 171746 240000 6 eFPGA_result_c_i[28]
port 428 nsew signal input
rlabel metal3 s 239200 163888 240000 164008 6 eFPGA_result_c_i[29]
port 429 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 eFPGA_result_c_i[2]
port 430 nsew signal input
rlabel metal3 s 239200 167016 240000 167136 6 eFPGA_result_c_i[30]
port 431 nsew signal input
rlabel metal3 s 0 177488 800 177608 6 eFPGA_result_c_i[31]
port 432 nsew signal input
rlabel metal3 s 239200 28704 240000 28824 6 eFPGA_result_c_i[3]
port 433 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 eFPGA_result_c_i[4]
port 434 nsew signal input
rlabel metal3 s 0 52776 800 52896 6 eFPGA_result_c_i[5]
port 435 nsew signal input
rlabel metal2 s 47582 239200 47638 240000 6 eFPGA_result_c_i[6]
port 436 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 eFPGA_result_c_i[7]
port 437 nsew signal input
rlabel metal3 s 0 62160 800 62280 6 eFPGA_result_c_i[8]
port 438 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 eFPGA_result_c_i[9]
port 439 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 eFPGA_write_strobe_o
port 440 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 fetch_enable_i
port 441 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 hart_id_i[0]
port 442 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 hart_id_i[10]
port 443 nsew signal input
rlabel metal2 s 77390 239200 77446 240000 6 hart_id_i[11]
port 444 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 hart_id_i[12]
port 445 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 hart_id_i[13]
port 446 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 hart_id_i[14]
port 447 nsew signal input
rlabel metal2 s 102966 239200 103022 240000 6 hart_id_i[15]
port 448 nsew signal input
rlabel metal3 s 239200 99968 240000 100088 6 hart_id_i[16]
port 449 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 hart_id_i[17]
port 450 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 hart_id_i[18]
port 451 nsew signal input
rlabel metal3 s 239200 120912 240000 121032 6 hart_id_i[19]
port 452 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 hart_id_i[1]
port 453 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 hart_id_i[20]
port 454 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 hart_id_i[21]
port 455 nsew signal input
rlabel metal3 s 0 131384 800 131504 6 hart_id_i[22]
port 456 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 hart_id_i[23]
port 457 nsew signal input
rlabel metal3 s 239200 141856 240000 141976 6 hart_id_i[24]
port 458 nsew signal input
rlabel metal3 s 239200 148112 240000 148232 6 hart_id_i[25]
port 459 nsew signal input
rlabel metal3 s 239200 155456 240000 155576 6 hart_id_i[26]
port 460 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 hart_id_i[27]
port 461 nsew signal input
rlabel metal2 s 172794 239200 172850 240000 6 hart_id_i[28]
port 462 nsew signal input
rlabel metal3 s 0 161712 800 161832 6 hart_id_i[29]
port 463 nsew signal input
rlabel metal3 s 239200 25440 240000 25560 6 hart_id_i[2]
port 464 nsew signal input
rlabel metal3 s 239200 168104 240000 168224 6 hart_id_i[30]
port 465 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 hart_id_i[31]
port 466 nsew signal input
rlabel metal3 s 239200 29656 240000 29776 6 hart_id_i[3]
port 467 nsew signal input
rlabel metal2 s 36358 239200 36414 240000 6 hart_id_i[4]
port 468 nsew signal input
rlabel metal3 s 239200 41216 240000 41336 6 hart_id_i[5]
port 469 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 hart_id_i[6]
port 470 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 hart_id_i[7]
port 471 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 hart_id_i[8]
port 472 nsew signal input
rlabel metal3 s 239200 62160 240000 62280 6 hart_id_i[9]
port 473 nsew signal input
rlabel metal3 s 0 14016 800 14136 6 ic_data_addr_o[0]
port 474 nsew signal output
rlabel metal2 s 16854 239200 16910 240000 6 ic_data_addr_o[1]
port 475 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 ic_data_addr_o[2]
port 476 nsew signal output
rlabel metal2 s 29182 239200 29238 240000 6 ic_data_addr_o[3]
port 477 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 ic_data_addr_o[4]
port 478 nsew signal output
rlabel metal3 s 239200 42304 240000 42424 6 ic_data_addr_o[5]
port 479 nsew signal output
rlabel metal2 s 48686 239200 48742 240000 6 ic_data_addr_o[6]
port 480 nsew signal output
rlabel metal3 s 239200 53864 240000 53984 6 ic_data_addr_o[7]
port 481 nsew signal output
rlabel metal2 s 8666 239200 8722 240000 6 ic_data_rdata_i[0]
port 482 nsew signal input
rlabel metal2 s 222934 0 222990 800 6 ic_data_rdata_i[100]
port 483 nsew signal input
rlabel metal2 s 228178 239200 228234 240000 6 ic_data_rdata_i[101]
port 484 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 ic_data_rdata_i[102]
port 485 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 ic_data_rdata_i[103]
port 486 nsew signal input
rlabel metal3 s 239200 229848 240000 229968 6 ic_data_rdata_i[104]
port 487 nsew signal input
rlabel metal2 s 226614 0 226670 800 6 ic_data_rdata_i[105]
port 488 nsew signal input
rlabel metal3 s 239200 230936 240000 231056 6 ic_data_rdata_i[106]
port 489 nsew signal input
rlabel metal3 s 0 228896 800 229016 6 ic_data_rdata_i[107]
port 490 nsew signal input
rlabel metal3 s 0 230936 800 231056 6 ic_data_rdata_i[108]
port 491 nsew signal input
rlabel metal2 s 228454 0 228510 800 6 ic_data_rdata_i[109]
port 492 nsew signal input
rlabel metal3 s 239200 69504 240000 69624 6 ic_data_rdata_i[10]
port 493 nsew signal input
rlabel metal2 s 231214 239200 231270 240000 6 ic_data_rdata_i[110]
port 494 nsew signal input
rlabel metal2 s 232226 239200 232282 240000 6 ic_data_rdata_i[111]
port 495 nsew signal input
rlabel metal3 s 0 232024 800 232144 6 ic_data_rdata_i[112]
port 496 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 ic_data_rdata_i[113]
port 497 nsew signal input
rlabel metal3 s 239200 234064 240000 234184 6 ic_data_rdata_i[114]
port 498 nsew signal input
rlabel metal3 s 0 234064 800 234184 6 ic_data_rdata_i[115]
port 499 nsew signal input
rlabel metal3 s 0 235152 800 235272 6 ic_data_rdata_i[116]
port 500 nsew signal input
rlabel metal3 s 239200 235152 240000 235272 6 ic_data_rdata_i[117]
port 501 nsew signal input
rlabel metal2 s 234894 0 234950 800 6 ic_data_rdata_i[118]
port 502 nsew signal input
rlabel metal2 s 235354 239200 235410 240000 6 ic_data_rdata_i[119]
port 503 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 ic_data_rdata_i[11]
port 504 nsew signal input
rlabel metal3 s 239200 236240 240000 236360 6 ic_data_rdata_i[120]
port 505 nsew signal input
rlabel metal2 s 235814 0 235870 800 6 ic_data_rdata_i[121]
port 506 nsew signal input
rlabel metal2 s 237654 0 237710 800 6 ic_data_rdata_i[122]
port 507 nsew signal input
rlabel metal2 s 238574 0 238630 800 6 ic_data_rdata_i[123]
port 508 nsew signal input
rlabel metal3 s 0 237192 800 237312 6 ic_data_rdata_i[124]
port 509 nsew signal input
rlabel metal3 s 239200 239368 240000 239488 6 ic_data_rdata_i[125]
port 510 nsew signal input
rlabel metal3 s 0 239368 800 239488 6 ic_data_rdata_i[126]
port 511 nsew signal input
rlabel metal2 s 239402 239200 239458 240000 6 ic_data_rdata_i[127]
port 512 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 ic_data_rdata_i[12]
port 513 nsew signal input
rlabel metal2 s 90730 239200 90786 240000 6 ic_data_rdata_i[13]
port 514 nsew signal input
rlabel metal2 s 94778 239200 94834 240000 6 ic_data_rdata_i[14]
port 515 nsew signal input
rlabel metal3 s 239200 92624 240000 92744 6 ic_data_rdata_i[15]
port 516 nsew signal input
rlabel metal2 s 107106 239200 107162 240000 6 ic_data_rdata_i[16]
port 517 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 ic_data_rdata_i[17]
port 518 nsew signal input
rlabel metal3 s 239200 114656 240000 114776 6 ic_data_rdata_i[18]
port 519 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 ic_data_rdata_i[19]
port 520 nsew signal input
rlabel metal2 s 17866 239200 17922 240000 6 ic_data_rdata_i[1]
port 521 nsew signal input
rlabel metal2 s 126610 239200 126666 240000 6 ic_data_rdata_i[20]
port 522 nsew signal input
rlabel metal2 s 134798 239200 134854 240000 6 ic_data_rdata_i[21]
port 523 nsew signal input
rlabel metal2 s 141974 239200 142030 240000 6 ic_data_rdata_i[22]
port 524 nsew signal input
rlabel metal2 s 148138 239200 148194 240000 6 ic_data_rdata_i[23]
port 525 nsew signal input
rlabel metal2 s 150162 239200 150218 240000 6 ic_data_rdata_i[24]
port 526 nsew signal input
rlabel metal3 s 0 142944 800 143064 6 ic_data_rdata_i[25]
port 527 nsew signal input
rlabel metal3 s 0 147160 800 147280 6 ic_data_rdata_i[26]
port 528 nsew signal input
rlabel metal2 s 165618 239200 165674 240000 6 ic_data_rdata_i[27]
port 529 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 ic_data_rdata_i[28]
port 530 nsew signal input
rlabel metal3 s 0 162800 800 162920 6 ic_data_rdata_i[29]
port 531 nsew signal input
rlabel metal3 s 239200 26528 240000 26648 6 ic_data_rdata_i[2]
port 532 nsew signal input
rlabel metal3 s 0 171232 800 171352 6 ic_data_rdata_i[30]
port 533 nsew signal input
rlabel metal3 s 239200 171232 240000 171352 6 ic_data_rdata_i[31]
port 534 nsew signal input
rlabel metal3 s 239200 174360 240000 174480 6 ic_data_rdata_i[32]
port 535 nsew signal input
rlabel metal2 s 188158 239200 188214 240000 6 ic_data_rdata_i[33]
port 536 nsew signal input
rlabel metal2 s 190182 239200 190238 240000 6 ic_data_rdata_i[34]
port 537 nsew signal input
rlabel metal3 s 239200 180616 240000 180736 6 ic_data_rdata_i[35]
port 538 nsew signal input
rlabel metal3 s 0 179528 800 179648 6 ic_data_rdata_i[36]
port 539 nsew signal input
rlabel metal2 s 192206 239200 192262 240000 6 ic_data_rdata_i[37]
port 540 nsew signal input
rlabel metal3 s 0 183744 800 183864 6 ic_data_rdata_i[38]
port 541 nsew signal input
rlabel metal3 s 239200 182792 240000 182912 6 ic_data_rdata_i[39]
port 542 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 ic_data_rdata_i[3]
port 543 nsew signal input
rlabel metal2 s 195334 239200 195390 240000 6 ic_data_rdata_i[40]
port 544 nsew signal input
rlabel metal2 s 191838 0 191894 800 6 ic_data_rdata_i[41]
port 545 nsew signal input
rlabel metal3 s 239200 185920 240000 186040 6 ic_data_rdata_i[42]
port 546 nsew signal input
rlabel metal2 s 193678 0 193734 800 6 ic_data_rdata_i[43]
port 547 nsew signal input
rlabel metal3 s 0 187960 800 188080 6 ic_data_rdata_i[44]
port 548 nsew signal input
rlabel metal3 s 0 190136 800 190256 6 ic_data_rdata_i[45]
port 549 nsew signal input
rlabel metal3 s 0 192176 800 192296 6 ic_data_rdata_i[46]
port 550 nsew signal input
rlabel metal3 s 239200 192176 240000 192296 6 ic_data_rdata_i[47]
port 551 nsew signal input
rlabel metal3 s 239200 193264 240000 193384 6 ic_data_rdata_i[48]
port 552 nsew signal input
rlabel metal3 s 239200 196392 240000 196512 6 ic_data_rdata_i[49]
port 553 nsew signal input
rlabel metal3 s 239200 36048 240000 36168 6 ic_data_rdata_i[4]
port 554 nsew signal input
rlabel metal3 s 239200 197344 240000 197464 6 ic_data_rdata_i[50]
port 555 nsew signal input
rlabel metal2 s 203522 239200 203578 240000 6 ic_data_rdata_i[51]
port 556 nsew signal input
rlabel metal2 s 197266 0 197322 800 6 ic_data_rdata_i[52]
port 557 nsew signal input
rlabel metal3 s 0 197344 800 197464 6 ic_data_rdata_i[53]
port 558 nsew signal input
rlabel metal3 s 239200 198432 240000 198552 6 ic_data_rdata_i[54]
port 559 nsew signal input
rlabel metal3 s 239200 200608 240000 200728 6 ic_data_rdata_i[55]
port 560 nsew signal input
rlabel metal3 s 0 198432 800 198552 6 ic_data_rdata_i[56]
port 561 nsew signal input
rlabel metal3 s 0 199520 800 199640 6 ic_data_rdata_i[57]
port 562 nsew signal input
rlabel metal3 s 0 201560 800 201680 6 ic_data_rdata_i[58]
port 563 nsew signal input
rlabel metal2 s 209686 239200 209742 240000 6 ic_data_rdata_i[59]
port 564 nsew signal input
rlabel metal3 s 239200 43392 240000 43512 6 ic_data_rdata_i[5]
port 565 nsew signal input
rlabel metal2 s 210698 239200 210754 240000 6 ic_data_rdata_i[60]
port 566 nsew signal input
rlabel metal3 s 0 205776 800 205896 6 ic_data_rdata_i[61]
port 567 nsew signal input
rlabel metal3 s 239200 204688 240000 204808 6 ic_data_rdata_i[62]
port 568 nsew signal input
rlabel metal3 s 0 206864 800 206984 6 ic_data_rdata_i[63]
port 569 nsew signal input
rlabel metal2 s 202786 0 202842 800 6 ic_data_rdata_i[64]
port 570 nsew signal input
rlabel metal2 s 215850 239200 215906 240000 6 ic_data_rdata_i[65]
port 571 nsew signal input
rlabel metal3 s 239200 206864 240000 206984 6 ic_data_rdata_i[66]
port 572 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 ic_data_rdata_i[67]
port 573 nsew signal input
rlabel metal3 s 0 211080 800 211200 6 ic_data_rdata_i[68]
port 574 nsew signal input
rlabel metal3 s 239200 207952 240000 208072 6 ic_data_rdata_i[69]
port 575 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 ic_data_rdata_i[6]
port 576 nsew signal input
rlabel metal3 s 239200 208904 240000 209024 6 ic_data_rdata_i[70]
port 577 nsew signal input
rlabel metal2 s 219990 239200 220046 240000 6 ic_data_rdata_i[71]
port 578 nsew signal input
rlabel metal3 s 0 212032 800 212152 6 ic_data_rdata_i[72]
port 579 nsew signal input
rlabel metal2 s 221002 239200 221058 240000 6 ic_data_rdata_i[73]
port 580 nsew signal input
rlabel metal3 s 0 214208 800 214328 6 ic_data_rdata_i[74]
port 581 nsew signal input
rlabel metal2 s 207386 0 207442 800 6 ic_data_rdata_i[75]
port 582 nsew signal input
rlabel metal3 s 239200 212032 240000 212152 6 ic_data_rdata_i[76]
port 583 nsew signal input
rlabel metal2 s 209226 0 209282 800 6 ic_data_rdata_i[77]
port 584 nsew signal input
rlabel metal2 s 210146 0 210202 800 6 ic_data_rdata_i[78]
port 585 nsew signal input
rlabel metal3 s 0 217336 800 217456 6 ic_data_rdata_i[79]
port 586 nsew signal input
rlabel metal3 s 239200 54816 240000 54936 6 ic_data_rdata_i[7]
port 587 nsew signal input
rlabel metal3 s 0 218424 800 218544 6 ic_data_rdata_i[80]
port 588 nsew signal input
rlabel metal2 s 211066 0 211122 800 6 ic_data_rdata_i[81]
port 589 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 ic_data_rdata_i[82]
port 590 nsew signal input
rlabel metal2 s 223026 239200 223082 240000 6 ic_data_rdata_i[83]
port 591 nsew signal input
rlabel metal2 s 213826 0 213882 800 6 ic_data_rdata_i[84]
port 592 nsew signal input
rlabel metal2 s 214746 0 214802 800 6 ic_data_rdata_i[85]
port 593 nsew signal input
rlabel metal2 s 225050 239200 225106 240000 6 ic_data_rdata_i[86]
port 594 nsew signal input
rlabel metal3 s 0 221552 800 221672 6 ic_data_rdata_i[87]
port 595 nsew signal input
rlabel metal3 s 0 222504 800 222624 6 ic_data_rdata_i[88]
port 596 nsew signal input
rlabel metal3 s 239200 219376 240000 219496 6 ic_data_rdata_i[89]
port 597 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 ic_data_rdata_i[8]
port 598 nsew signal input
rlabel metal2 s 216586 0 216642 800 6 ic_data_rdata_i[90]
port 599 nsew signal input
rlabel metal2 s 226062 239200 226118 240000 6 ic_data_rdata_i[91]
port 600 nsew signal input
rlabel metal2 s 219254 0 219310 800 6 ic_data_rdata_i[92]
port 601 nsew signal input
rlabel metal2 s 220174 0 220230 800 6 ic_data_rdata_i[93]
port 602 nsew signal input
rlabel metal2 s 227166 239200 227222 240000 6 ic_data_rdata_i[94]
port 603 nsew signal input
rlabel metal3 s 239200 221552 240000 221672 6 ic_data_rdata_i[95]
port 604 nsew signal input
rlabel metal3 s 239200 222504 240000 222624 6 ic_data_rdata_i[96]
port 605 nsew signal input
rlabel metal3 s 0 224680 800 224800 6 ic_data_rdata_i[97]
port 606 nsew signal input
rlabel metal3 s 0 225768 800 225888 6 ic_data_rdata_i[98]
port 607 nsew signal input
rlabel metal3 s 239200 226720 240000 226840 6 ic_data_rdata_i[99]
port 608 nsew signal input
rlabel metal2 s 71226 239200 71282 240000 6 ic_data_rdata_i[9]
port 609 nsew signal input
rlabel metal3 s 239200 9800 240000 9920 6 ic_data_req_o[0]
port 610 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 ic_data_req_o[1]
port 611 nsew signal output
rlabel metal3 s 239200 10888 240000 11008 6 ic_data_wdata_o[0]
port 612 nsew signal output
rlabel metal3 s 239200 70592 240000 70712 6 ic_data_wdata_o[10]
port 613 nsew signal output
rlabel metal3 s 239200 76848 240000 76968 6 ic_data_wdata_o[11]
port 614 nsew signal output
rlabel metal3 s 239200 82152 240000 82272 6 ic_data_wdata_o[12]
port 615 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 ic_data_wdata_o[13]
port 616 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 ic_data_wdata_o[14]
port 617 nsew signal output
rlabel metal3 s 239200 93576 240000 93696 6 ic_data_wdata_o[15]
port 618 nsew signal output
rlabel metal3 s 239200 100920 240000 101040 6 ic_data_wdata_o[16]
port 619 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 ic_data_wdata_o[17]
port 620 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 ic_data_wdata_o[18]
port 621 nsew signal output
rlabel metal3 s 239200 122000 240000 122120 6 ic_data_wdata_o[19]
port 622 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 ic_data_wdata_o[1]
port 623 nsew signal output
rlabel metal3 s 239200 125128 240000 125248 6 ic_data_wdata_o[20]
port 624 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 ic_data_wdata_o[21]
port 625 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 ic_data_wdata_o[22]
port 626 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 ic_data_wdata_o[23]
port 627 nsew signal output
rlabel metal3 s 239200 142944 240000 143064 6 ic_data_wdata_o[24]
port 628 nsew signal output
rlabel metal3 s 239200 149200 240000 149320 6 ic_data_wdata_o[25]
port 629 nsew signal output
rlabel metal2 s 159454 239200 159510 240000 6 ic_data_wdata_o[26]
port 630 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 ic_data_wdata_o[27]
port 631 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 ic_data_wdata_o[28]
port 632 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 ic_data_wdata_o[29]
port 633 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 ic_data_wdata_o[2]
port 634 nsew signal output
rlabel metal2 s 177118 0 177174 800 6 ic_data_wdata_o[30]
port 635 nsew signal output
rlabel metal2 s 183558 0 183614 800 6 ic_data_wdata_o[31]
port 636 nsew signal output
rlabel metal2 s 187146 239200 187202 240000 6 ic_data_wdata_o[32]
port 637 nsew signal output
rlabel metal2 s 189170 239200 189226 240000 6 ic_data_wdata_o[33]
port 638 nsew signal output
rlabel metal3 s 239200 177488 240000 177608 6 ic_data_wdata_o[34]
port 639 nsew signal output
rlabel metal2 s 191194 239200 191250 240000 6 ic_data_wdata_o[35]
port 640 nsew signal output
rlabel metal3 s 0 180616 800 180736 6 ic_data_wdata_o[36]
port 641 nsew signal output
rlabel metal2 s 186318 0 186374 800 6 ic_data_wdata_o[37]
port 642 nsew signal output
rlabel metal2 s 188158 0 188214 800 6 ic_data_wdata_o[38]
port 643 nsew signal output
rlabel metal3 s 239200 183744 240000 183864 6 ic_data_wdata_o[39]
port 644 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 ic_data_wdata_o[3]
port 645 nsew signal output
rlabel metal2 s 196346 239200 196402 240000 6 ic_data_wdata_o[40]
port 646 nsew signal output
rlabel metal2 s 198370 239200 198426 240000 6 ic_data_wdata_o[41]
port 647 nsew signal output
rlabel metal2 s 192758 0 192814 800 6 ic_data_wdata_o[42]
port 648 nsew signal output
rlabel metal3 s 239200 186872 240000 186992 6 ic_data_wdata_o[43]
port 649 nsew signal output
rlabel metal3 s 0 189048 800 189168 6 ic_data_wdata_o[44]
port 650 nsew signal output
rlabel metal3 s 239200 190136 240000 190256 6 ic_data_wdata_o[45]
port 651 nsew signal output
rlabel metal3 s 239200 191088 240000 191208 6 ic_data_wdata_o[46]
port 652 nsew signal output
rlabel metal2 s 201498 239200 201554 240000 6 ic_data_wdata_o[47]
port 653 nsew signal output
rlabel metal3 s 239200 194216 240000 194336 6 ic_data_wdata_o[48]
port 654 nsew signal output
rlabel metal2 s 194598 0 194654 800 6 ic_data_wdata_o[49]
port 655 nsew signal output
rlabel metal3 s 239200 37000 240000 37120 6 ic_data_wdata_o[4]
port 656 nsew signal output
rlabel metal2 s 195518 0 195574 800 6 ic_data_wdata_o[50]
port 657 nsew signal output
rlabel metal2 s 204534 239200 204590 240000 6 ic_data_wdata_o[51]
port 658 nsew signal output
rlabel metal2 s 205546 239200 205602 240000 6 ic_data_wdata_o[52]
port 659 nsew signal output
rlabel metal2 s 198186 0 198242 800 6 ic_data_wdata_o[53]
port 660 nsew signal output
rlabel metal3 s 239200 199520 240000 199640 6 ic_data_wdata_o[54]
port 661 nsew signal output
rlabel metal2 s 200026 0 200082 800 6 ic_data_wdata_o[55]
port 662 nsew signal output
rlabel metal3 s 239200 201560 240000 201680 6 ic_data_wdata_o[56]
port 663 nsew signal output
rlabel metal2 s 208674 239200 208730 240000 6 ic_data_wdata_o[57]
port 664 nsew signal output
rlabel metal3 s 239200 203736 240000 203856 6 ic_data_wdata_o[58]
port 665 nsew signal output
rlabel metal3 s 0 202648 800 202768 6 ic_data_wdata_o[59]
port 666 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 ic_data_wdata_o[5]
port 667 nsew signal output
rlabel metal2 s 211710 239200 211766 240000 6 ic_data_wdata_o[60]
port 668 nsew signal output
rlabel metal2 s 212722 239200 212778 240000 6 ic_data_wdata_o[61]
port 669 nsew signal output
rlabel metal3 s 239200 205776 240000 205896 6 ic_data_wdata_o[62]
port 670 nsew signal output
rlabel metal3 s 0 207952 800 208072 6 ic_data_wdata_o[63]
port 671 nsew signal output
rlabel metal2 s 49698 239200 49754 240000 6 ic_data_wdata_o[6]
port 672 nsew signal output
rlabel metal3 s 239200 55904 240000 56024 6 ic_data_wdata_o[7]
port 673 nsew signal output
rlabel metal2 s 65062 239200 65118 240000 6 ic_data_wdata_o[8]
port 674 nsew signal output
rlabel metal3 s 0 71680 800 71800 6 ic_data_wdata_o[9]
port 675 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 ic_data_write_o
port 676 nsew signal output
rlabel metal2 s 9678 239200 9734 240000 6 ic_tag_addr_o[0]
port 677 nsew signal output
rlabel metal3 s 239200 18232 240000 18352 6 ic_tag_addr_o[1]
port 678 nsew signal output
rlabel metal2 s 26054 239200 26110 240000 6 ic_tag_addr_o[2]
port 679 nsew signal output
rlabel metal3 s 0 42304 800 42424 6 ic_tag_addr_o[3]
port 680 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 ic_tag_addr_o[4]
port 681 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 ic_tag_addr_o[5]
port 682 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 ic_tag_addr_o[6]
port 683 nsew signal output
rlabel metal2 s 56874 239200 56930 240000 6 ic_tag_addr_o[7]
port 684 nsew signal output
rlabel metal2 s 10690 239200 10746 240000 6 ic_tag_rdata_i[0]
port 685 nsew signal input
rlabel metal2 s 73250 239200 73306 240000 6 ic_tag_rdata_i[10]
port 686 nsew signal input
rlabel metal2 s 78402 239200 78458 240000 6 ic_tag_rdata_i[11]
port 687 nsew signal input
rlabel metal2 s 82450 239200 82506 240000 6 ic_tag_rdata_i[12]
port 688 nsew signal input
rlabel metal3 s 239200 85280 240000 85400 6 ic_tag_rdata_i[13]
port 689 nsew signal input
rlabel metal2 s 95790 239200 95846 240000 6 ic_tag_rdata_i[14]
port 690 nsew signal input
rlabel metal3 s 239200 94664 240000 94784 6 ic_tag_rdata_i[15]
port 691 nsew signal input
rlabel metal3 s 239200 102008 240000 102128 6 ic_tag_rdata_i[16]
port 692 nsew signal input
rlabel metal3 s 239200 108264 240000 108384 6 ic_tag_rdata_i[17]
port 693 nsew signal input
rlabel metal3 s 239200 115608 240000 115728 6 ic_tag_rdata_i[18]
port 694 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 ic_tag_rdata_i[19]
port 695 nsew signal input
rlabel metal2 s 18878 239200 18934 240000 6 ic_tag_rdata_i[1]
port 696 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 ic_tag_rdata_i[20]
port 697 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 ic_tag_rdata_i[21]
port 698 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 ic_tag_rdata_i[22]
port 699 nsew signal input
rlabel metal3 s 0 134512 800 134632 6 ic_tag_rdata_i[23]
port 700 nsew signal input
rlabel metal3 s 239200 143896 240000 144016 6 ic_tag_rdata_i[24]
port 701 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 ic_tag_rdata_i[25]
port 702 nsew signal input
rlabel metal2 s 160466 239200 160522 240000 6 ic_tag_rdata_i[26]
port 703 nsew signal input
rlabel metal2 s 166630 239200 166686 240000 6 ic_tag_rdata_i[27]
port 704 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 ic_tag_rdata_i[28]
port 705 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 ic_tag_rdata_i[29]
port 706 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 ic_tag_rdata_i[2]
port 707 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 ic_tag_rdata_i[30]
port 708 nsew signal input
rlabel metal2 s 181994 239200 182050 240000 6 ic_tag_rdata_i[31]
port 709 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 ic_tag_rdata_i[32]
port 710 nsew signal input
rlabel metal3 s 239200 176400 240000 176520 6 ic_tag_rdata_i[33]
port 711 nsew signal input
rlabel metal3 s 239200 178576 240000 178696 6 ic_tag_rdata_i[34]
port 712 nsew signal input
rlabel metal3 s 239200 181704 240000 181824 6 ic_tag_rdata_i[35]
port 713 nsew signal input
rlabel metal3 s 0 181704 800 181824 6 ic_tag_rdata_i[36]
port 714 nsew signal input
rlabel metal2 s 193310 239200 193366 240000 6 ic_tag_rdata_i[37]
port 715 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 ic_tag_rdata_i[38]
port 716 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 ic_tag_rdata_i[39]
port 717 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 ic_tag_rdata_i[3]
port 718 nsew signal input
rlabel metal2 s 190918 0 190974 800 6 ic_tag_rdata_i[40]
port 719 nsew signal input
rlabel metal3 s 0 185920 800 186040 6 ic_tag_rdata_i[41]
port 720 nsew signal input
rlabel metal2 s 199474 239200 199530 240000 6 ic_tag_rdata_i[42]
port 721 nsew signal input
rlabel metal3 s 239200 187960 240000 188080 6 ic_tag_rdata_i[43]
port 722 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 ic_tag_rdata_i[4]
port 723 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 ic_tag_rdata_i[5]
port 724 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 ic_tag_rdata_i[6]
port 725 nsew signal input
rlabel metal2 s 57886 239200 57942 240000 6 ic_tag_rdata_i[7]
port 726 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 ic_tag_rdata_i[8]
port 727 nsew signal input
rlabel metal3 s 239200 63248 240000 63368 6 ic_tag_rdata_i[9]
port 728 nsew signal input
rlabel metal2 s 11702 239200 11758 240000 6 ic_tag_req_o[0]
port 729 nsew signal output
rlabel metal3 s 239200 19184 240000 19304 6 ic_tag_req_o[1]
port 730 nsew signal output
rlabel metal2 s 12714 239200 12770 240000 6 ic_tag_wdata_o[0]
port 731 nsew signal output
rlabel metal3 s 239200 71680 240000 71800 6 ic_tag_wdata_o[10]
port 732 nsew signal output
rlabel metal3 s 0 83104 800 83224 6 ic_tag_wdata_o[11]
port 733 nsew signal output
rlabel metal2 s 83554 239200 83610 240000 6 ic_tag_wdata_o[12]
port 734 nsew signal output
rlabel metal3 s 0 92624 800 92744 6 ic_tag_wdata_o[13]
port 735 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 ic_tag_wdata_o[14]
port 736 nsew signal output
rlabel metal3 s 239200 95752 240000 95872 6 ic_tag_wdata_o[15]
port 737 nsew signal output
rlabel metal3 s 0 106224 800 106344 6 ic_tag_wdata_o[16]
port 738 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 ic_tag_wdata_o[17]
port 739 nsew signal output
rlabel metal2 s 116306 239200 116362 240000 6 ic_tag_wdata_o[18]
port 740 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 ic_tag_wdata_o[19]
port 741 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 ic_tag_wdata_o[1]
port 742 nsew signal output
rlabel metal2 s 127622 239200 127678 240000 6 ic_tag_wdata_o[20]
port 743 nsew signal output
rlabel metal3 s 0 126080 800 126200 6 ic_tag_wdata_o[21]
port 744 nsew signal output
rlabel metal2 s 27066 239200 27122 240000 6 ic_tag_wdata_o[2]
port 745 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 ic_tag_wdata_o[3]
port 746 nsew signal output
rlabel metal3 s 239200 38088 240000 38208 6 ic_tag_wdata_o[4]
port 747 nsew signal output
rlabel metal2 s 42522 239200 42578 240000 6 ic_tag_wdata_o[5]
port 748 nsew signal output
rlabel metal2 s 50710 239200 50766 240000 6 ic_tag_wdata_o[6]
port 749 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 ic_tag_wdata_o[7]
port 750 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 ic_tag_wdata_o[8]
port 751 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 ic_tag_wdata_o[9]
port 752 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 ic_tag_write_o
port 753 nsew signal output
rlabel metal3 s 239200 11840 240000 11960 6 instr_addr_o[0]
port 754 nsew signal output
rlabel metal2 s 74262 239200 74318 240000 6 instr_addr_o[10]
port 755 nsew signal output
rlabel metal3 s 0 84192 800 84312 6 instr_addr_o[11]
port 756 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 instr_addr_o[12]
port 757 nsew signal output
rlabel metal2 s 91742 239200 91798 240000 6 instr_addr_o[13]
port 758 nsew signal output
rlabel metal2 s 96894 239200 96950 240000 6 instr_addr_o[14]
port 759 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 instr_addr_o[15]
port 760 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 instr_addr_o[16]
port 761 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 instr_addr_o[17]
port 762 nsew signal output
rlabel metal2 s 117410 239200 117466 240000 6 instr_addr_o[18]
port 763 nsew signal output
rlabel metal2 s 121458 239200 121514 240000 6 instr_addr_o[19]
port 764 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 instr_addr_o[1]
port 765 nsew signal output
rlabel metal2 s 128634 239200 128690 240000 6 instr_addr_o[20]
port 766 nsew signal output
rlabel metal3 s 0 127168 800 127288 6 instr_addr_o[21]
port 767 nsew signal output
rlabel metal2 s 142986 239200 143042 240000 6 instr_addr_o[22]
port 768 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 instr_addr_o[23]
port 769 nsew signal output
rlabel metal2 s 151174 239200 151230 240000 6 instr_addr_o[24]
port 770 nsew signal output
rlabel metal3 s 0 143896 800 144016 6 instr_addr_o[25]
port 771 nsew signal output
rlabel metal3 s 239200 156544 240000 156664 6 instr_addr_o[26]
port 772 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 instr_addr_o[27]
port 773 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 instr_addr_o[28]
port 774 nsew signal output
rlabel metal3 s 0 163888 800 164008 6 instr_addr_o[29]
port 775 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 instr_addr_o[2]
port 776 nsew signal output
rlabel metal2 s 178958 239200 179014 240000 6 instr_addr_o[30]
port 777 nsew signal output
rlabel metal2 s 183006 239200 183062 240000 6 instr_addr_o[31]
port 778 nsew signal output
rlabel metal2 s 30194 239200 30250 240000 6 instr_addr_o[3]
port 779 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 instr_addr_o[4]
port 780 nsew signal output
rlabel metal2 s 43534 239200 43590 240000 6 instr_addr_o[5]
port 781 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 instr_addr_o[6]
port 782 nsew signal output
rlabel metal3 s 239200 56992 240000 57112 6 instr_addr_o[7]
port 783 nsew signal output
rlabel metal3 s 239200 60120 240000 60240 6 instr_addr_o[8]
port 784 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 instr_addr_o[9]
port 785 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 instr_err_i
port 786 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 instr_gnt_i
port 787 nsew signal input
rlabel metal3 s 239200 12928 240000 13048 6 instr_rdata_i[0]
port 788 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 instr_rdata_i[10]
port 789 nsew signal input
rlabel metal2 s 79414 239200 79470 240000 6 instr_rdata_i[11]
port 790 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 instr_rdata_i[12]
port 791 nsew signal input
rlabel metal3 s 239200 86368 240000 86488 6 instr_rdata_i[13]
port 792 nsew signal input
rlabel metal2 s 97906 239200 97962 240000 6 instr_rdata_i[14]
port 793 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 instr_rdata_i[15]
port 794 nsew signal input
rlabel metal3 s 239200 103096 240000 103216 6 instr_rdata_i[16]
port 795 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 instr_rdata_i[17]
port 796 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 instr_rdata_i[18]
port 797 nsew signal input
rlabel metal2 s 122470 239200 122526 240000 6 instr_rdata_i[19]
port 798 nsew signal input
rlabel metal2 s 19890 239200 19946 240000 6 instr_rdata_i[1]
port 799 nsew signal input
rlabel metal3 s 0 122000 800 122120 6 instr_rdata_i[20]
port 800 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 instr_rdata_i[21]
port 801 nsew signal input
rlabel metal2 s 143998 239200 144054 240000 6 instr_rdata_i[22]
port 802 nsew signal input
rlabel metal3 s 0 136552 800 136672 6 instr_rdata_i[23]
port 803 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 instr_rdata_i[24]
port 804 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 instr_rdata_i[25]
port 805 nsew signal input
rlabel metal2 s 161478 239200 161534 240000 6 instr_rdata_i[26]
port 806 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 instr_rdata_i[27]
port 807 nsew signal input
rlabel metal3 s 0 157632 800 157752 6 instr_rdata_i[28]
port 808 nsew signal input
rlabel metal2 s 175830 239200 175886 240000 6 instr_rdata_i[29]
port 809 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 instr_rdata_i[2]
port 810 nsew signal input
rlabel metal2 s 179970 239200 180026 240000 6 instr_rdata_i[30]
port 811 nsew signal input
rlabel metal2 s 184018 239200 184074 240000 6 instr_rdata_i[31]
port 812 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 instr_rdata_i[3]
port 813 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 instr_rdata_i[4]
port 814 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 instr_rdata_i[5]
port 815 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 instr_rdata_i[6]
port 816 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 instr_rdata_i[7]
port 817 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 instr_rdata_i[8]
port 818 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 instr_rdata_i[9]
port 819 nsew signal input
rlabel metal2 s 3514 239200 3570 240000 6 instr_req_o
port 820 nsew signal output
rlabel metal2 s 4526 239200 4582 240000 6 instr_rvalid_i
port 821 nsew signal input
rlabel metal2 s 386 0 442 800 6 irq_external_i
port 822 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 irq_fast_i[0]
port 823 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 irq_fast_i[10]
port 824 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 irq_fast_i[11]
port 825 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 irq_fast_i[12]
port 826 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 irq_fast_i[13]
port 827 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 irq_fast_i[14]
port 828 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 irq_fast_i[1]
port 829 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 irq_fast_i[2]
port 830 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 irq_fast_i[3]
port 831 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 irq_fast_i[4]
port 832 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 irq_fast_i[5]
port 833 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 irq_fast_i[6]
port 834 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 irq_fast_i[7]
port 835 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 irq_fast_i[8]
port 836 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 irq_fast_i[9]
port 837 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 irq_nm_i
port 838 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 irq_pending_o
port 839 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 irq_software_i
port 840 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 irq_timer_i
port 841 nsew signal input
rlabel metal3 s 239200 14016 240000 14136 6 rf_raddr_a_o[0]
port 842 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 rf_raddr_a_o[1]
port 843 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 rf_raddr_a_o[2]
port 844 nsew signal output
rlabel metal3 s 239200 30744 240000 30864 6 rf_raddr_a_o[3]
port 845 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 rf_raddr_a_o[4]
port 846 nsew signal output
rlabel metal3 s 239200 14968 240000 15088 6 rf_raddr_b_o[0]
port 847 nsew signal output
rlabel metal3 s 239200 20272 240000 20392 6 rf_raddr_b_o[1]
port 848 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 rf_raddr_b_o[2]
port 849 nsew signal output
rlabel metal3 s 239200 31832 240000 31952 6 rf_raddr_b_o[3]
port 850 nsew signal output
rlabel metal2 s 37370 239200 37426 240000 6 rf_raddr_b_o[4]
port 851 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 rf_rdata_a_ecc_i[0]
port 852 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 rf_rdata_a_ecc_i[10]
port 853 nsew signal input
rlabel metal3 s 0 85280 800 85400 6 rf_rdata_a_ecc_i[11]
port 854 nsew signal input
rlabel metal3 s 239200 83104 240000 83224 6 rf_rdata_a_ecc_i[12]
port 855 nsew signal input
rlabel metal2 s 92754 239200 92810 240000 6 rf_rdata_a_ecc_i[13]
port 856 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 rf_rdata_a_ecc_i[14]
port 857 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 rf_rdata_a_ecc_i[15]
port 858 nsew signal input
rlabel metal2 s 108118 239200 108174 240000 6 rf_rdata_a_ecc_i[16]
port 859 nsew signal input
rlabel metal3 s 0 111392 800 111512 6 rf_rdata_a_ecc_i[17]
port 860 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 rf_rdata_a_ecc_i[18]
port 861 nsew signal input
rlabel metal3 s 0 117784 800 117904 6 rf_rdata_a_ecc_i[19]
port 862 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 rf_rdata_a_ecc_i[1]
port 863 nsew signal input
rlabel metal3 s 239200 126080 240000 126200 6 rf_rdata_a_ecc_i[20]
port 864 nsew signal input
rlabel metal2 s 135810 239200 135866 240000 6 rf_rdata_a_ecc_i[21]
port 865 nsew signal input
rlabel metal3 s 239200 133424 240000 133544 6 rf_rdata_a_ecc_i[22]
port 866 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 rf_rdata_a_ecc_i[23]
port 867 nsew signal input
rlabel metal2 s 152278 239200 152334 240000 6 rf_rdata_a_ecc_i[24]
port 868 nsew signal input
rlabel metal2 s 156326 239200 156382 240000 6 rf_rdata_a_ecc_i[25]
port 869 nsew signal input
rlabel metal2 s 162490 239200 162546 240000 6 rf_rdata_a_ecc_i[26]
port 870 nsew signal input
rlabel metal2 s 167642 239200 167698 240000 6 rf_rdata_a_ecc_i[27]
port 871 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 rf_rdata_a_ecc_i[28]
port 872 nsew signal input
rlabel metal2 s 176842 239200 176898 240000 6 rf_rdata_a_ecc_i[29]
port 873 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 rf_rdata_a_ecc_i[2]
port 874 nsew signal input
rlabel metal3 s 0 172320 800 172440 6 rf_rdata_a_ecc_i[30]
port 875 nsew signal input
rlabel metal3 s 239200 172320 240000 172440 6 rf_rdata_a_ecc_i[31]
port 876 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 rf_rdata_a_ecc_i[3]
port 877 nsew signal input
rlabel metal2 s 38382 239200 38438 240000 6 rf_rdata_a_ecc_i[4]
port 878 nsew signal input
rlabel metal2 s 44546 239200 44602 240000 6 rf_rdata_a_ecc_i[5]
port 879 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 rf_rdata_a_ecc_i[6]
port 880 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 rf_rdata_a_ecc_i[7]
port 881 nsew signal input
rlabel metal2 s 66074 239200 66130 240000 6 rf_rdata_a_ecc_i[8]
port 882 nsew signal input
rlabel metal3 s 239200 64336 240000 64456 6 rf_rdata_a_ecc_i[9]
port 883 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 rf_rdata_b_ecc_i[0]
port 884 nsew signal input
rlabel metal2 s 75274 239200 75330 240000 6 rf_rdata_b_ecc_i[10]
port 885 nsew signal input
rlabel metal3 s 239200 77936 240000 78056 6 rf_rdata_b_ecc_i[11]
port 886 nsew signal input
rlabel metal2 s 84566 239200 84622 240000 6 rf_rdata_b_ecc_i[12]
port 887 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 rf_rdata_b_ecc_i[13]
port 888 nsew signal input
rlabel metal3 s 239200 88408 240000 88528 6 rf_rdata_b_ecc_i[14]
port 889 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 rf_rdata_b_ecc_i[15]
port 890 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 rf_rdata_b_ecc_i[16]
port 891 nsew signal input
rlabel metal3 s 0 112480 800 112600 6 rf_rdata_b_ecc_i[17]
port 892 nsew signal input
rlabel metal3 s 239200 116696 240000 116816 6 rf_rdata_b_ecc_i[18]
port 893 nsew signal input
rlabel metal2 s 123482 239200 123538 240000 6 rf_rdata_b_ecc_i[19]
port 894 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 rf_rdata_b_ecc_i[1]
port 895 nsew signal input
rlabel metal3 s 0 122952 800 123072 6 rf_rdata_b_ecc_i[20]
port 896 nsew signal input
rlabel metal3 s 239200 129344 240000 129464 6 rf_rdata_b_ecc_i[21]
port 897 nsew signal input
rlabel metal3 s 239200 134512 240000 134632 6 rf_rdata_b_ecc_i[22]
port 898 nsew signal input
rlabel metal3 s 0 137640 800 137760 6 rf_rdata_b_ecc_i[23]
port 899 nsew signal input
rlabel metal3 s 239200 144984 240000 145104 6 rf_rdata_b_ecc_i[24]
port 900 nsew signal input
rlabel metal3 s 0 144984 800 145104 6 rf_rdata_b_ecc_i[25]
port 901 nsew signal input
rlabel metal3 s 0 148112 800 148232 6 rf_rdata_b_ecc_i[26]
port 902 nsew signal input
rlabel metal3 s 239200 159672 240000 159792 6 rf_rdata_b_ecc_i[27]
port 903 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 rf_rdata_b_ecc_i[28]
port 904 nsew signal input
rlabel metal3 s 0 164976 800 165096 6 rf_rdata_b_ecc_i[29]
port 905 nsew signal input
rlabel metal2 s 28170 239200 28226 240000 6 rf_rdata_b_ecc_i[2]
port 906 nsew signal input
rlabel metal3 s 239200 169056 240000 169176 6 rf_rdata_b_ecc_i[30]
port 907 nsew signal input
rlabel metal2 s 185030 239200 185086 240000 6 rf_rdata_b_ecc_i[31]
port 908 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 rf_rdata_b_ecc_i[3]
port 909 nsew signal input
rlabel metal2 s 39394 239200 39450 240000 6 rf_rdata_b_ecc_i[4]
port 910 nsew signal input
rlabel metal3 s 239200 44344 240000 44464 6 rf_rdata_b_ecc_i[5]
port 911 nsew signal input
rlabel metal2 s 51722 239200 51778 240000 6 rf_rdata_b_ecc_i[6]
port 912 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 rf_rdata_b_ecc_i[7]
port 913 nsew signal input
rlabel metal2 s 67086 239200 67142 240000 6 rf_rdata_b_ecc_i[8]
port 914 nsew signal input
rlabel metal3 s 239200 65288 240000 65408 6 rf_rdata_b_ecc_i[9]
port 915 nsew signal input
rlabel metal2 s 13726 239200 13782 240000 6 rf_waddr_wb_o[0]
port 916 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 rf_waddr_wb_o[1]
port 917 nsew signal output
rlabel metal3 s 0 33872 800 33992 6 rf_waddr_wb_o[2]
port 918 nsew signal output
rlabel metal2 s 31206 239200 31262 240000 6 rf_waddr_wb_o[3]
port 919 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 rf_waddr_wb_o[4]
port 920 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 rf_wdata_wb_ecc_o[0]
port 921 nsew signal output
rlabel metal3 s 0 77936 800 78056 6 rf_wdata_wb_ecc_o[10]
port 922 nsew signal output
rlabel metal3 s 239200 79024 240000 79144 6 rf_wdata_wb_ecc_o[11]
port 923 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 rf_wdata_wb_ecc_o[12]
port 924 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 rf_wdata_wb_ecc_o[13]
port 925 nsew signal output
rlabel metal2 s 98918 239200 98974 240000 6 rf_wdata_wb_ecc_o[14]
port 926 nsew signal output
rlabel metal3 s 239200 96840 240000 96960 6 rf_wdata_wb_ecc_o[15]
port 927 nsew signal output
rlabel metal3 s 239200 104184 240000 104304 6 rf_wdata_wb_ecc_o[16]
port 928 nsew signal output
rlabel metal3 s 239200 109352 240000 109472 6 rf_wdata_wb_ecc_o[17]
port 929 nsew signal output
rlabel metal3 s 0 116696 800 116816 6 rf_wdata_wb_ecc_o[18]
port 930 nsew signal output
rlabel metal3 s 239200 122952 240000 123072 6 rf_wdata_wb_ecc_o[19]
port 931 nsew signal output
rlabel metal2 s 20902 239200 20958 240000 6 rf_wdata_wb_ecc_o[1]
port 932 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 rf_wdata_wb_ecc_o[20]
port 933 nsew signal output
rlabel metal3 s 239200 130296 240000 130416 6 rf_wdata_wb_ecc_o[21]
port 934 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 rf_wdata_wb_ecc_o[22]
port 935 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 rf_wdata_wb_ecc_o[23]
port 936 nsew signal output
rlabel metal2 s 147862 0 147918 800 6 rf_wdata_wb_ecc_o[24]
port 937 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 rf_wdata_wb_ecc_o[25]
port 938 nsew signal output
rlabel metal3 s 0 149200 800 149320 6 rf_wdata_wb_ecc_o[26]
port 939 nsew signal output
rlabel metal2 s 163410 0 163466 800 6 rf_wdata_wb_ecc_o[27]
port 940 nsew signal output
rlabel metal2 s 170770 0 170826 800 6 rf_wdata_wb_ecc_o[28]
port 941 nsew signal output
rlabel metal2 s 175278 0 175334 800 6 rf_wdata_wb_ecc_o[29]
port 942 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 rf_wdata_wb_ecc_o[2]
port 943 nsew signal output
rlabel metal2 s 178958 0 179014 800 6 rf_wdata_wb_ecc_o[30]
port 944 nsew signal output
rlabel metal3 s 239200 173272 240000 173392 6 rf_wdata_wb_ecc_o[31]
port 945 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 rf_wdata_wb_ecc_o[3]
port 946 nsew signal output
rlabel metal3 s 0 50600 800 50720 6 rf_wdata_wb_ecc_o[4]
port 947 nsew signal output
rlabel metal2 s 45558 239200 45614 240000 6 rf_wdata_wb_ecc_o[5]
port 948 nsew signal output
rlabel metal3 s 239200 49648 240000 49768 6 rf_wdata_wb_ecc_o[6]
port 949 nsew signal output
rlabel metal2 s 58898 239200 58954 240000 6 rf_wdata_wb_ecc_o[7]
port 950 nsew signal output
rlabel metal3 s 0 67464 800 67584 6 rf_wdata_wb_ecc_o[8]
port 951 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 rf_wdata_wb_ecc_o[9]
port 952 nsew signal output
rlabel metal3 s 239200 4496 240000 4616 6 rf_we_wb_o
port 953 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 rst_ni
port 954 nsew signal input
rlabel metal4 s 4208 2128 4528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 14208 2128 14528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 24208 2128 24528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 34208 2128 34528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 44208 2128 44528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 54208 2128 54528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 64208 2128 64528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 74208 2128 74528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 84208 2128 84528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 94208 2128 94528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 104208 2128 104528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 114208 2128 114528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 124208 2128 124528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 134208 2128 134528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 144208 2128 144528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 154208 2128 154528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 164208 2128 164528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 174208 2128 174528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 184208 2128 184528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 194208 2128 194528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 204208 2128 204528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 214208 2128 214528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 224208 2128 224528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 234208 2128 234528 237776 6 vccd1
port 955 nsew power input
rlabel metal4 s 9208 2128 9528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 19208 2128 19528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 29208 2128 29528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 39208 2128 39528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 49208 2128 49528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 59208 2128 59528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 69208 2128 69528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 79208 2128 79528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 89208 2128 89528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 99208 2128 99528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 109208 2128 109528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 119208 2128 119528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 129208 2128 129528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 139208 2128 139528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 149208 2128 149528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 159208 2128 159528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 169208 2128 169528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 179208 2128 179528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 189208 2128 189528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 199208 2128 199528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 209208 2128 209528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 219208 2128 219528 237776 6 vssd1
port 956 nsew ground input
rlabel metal4 s 229208 2128 229528 237776 6 vssd1
port 956 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 240000 240000
string LEFview TRUE
string GDS_FILE /project/openlane/ibex_core/runs/ibex_core/results/magic/ibex_core.gds
string GDS_END 58354090
string GDS_START 671490
<< end >>

