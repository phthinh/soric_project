* NGSPICE file created from uart_to_mem.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

.subckt uart_to_mem clk_i data_addr_o[0] data_addr_o[10] data_addr_o[11] data_addr_o[1]
+ data_addr_o[2] data_addr_o[3] data_addr_o[4] data_addr_o[5] data_addr_o[6] data_addr_o[7]
+ data_addr_o[8] data_addr_o[9] data_be_o[0] data_be_o[1] data_be_o[2] data_be_o[3]
+ data_gnt_i data_rdata_i[0] data_rdata_i[10] data_rdata_i[11] data_rdata_i[12] data_rdata_i[13]
+ data_rdata_i[14] data_rdata_i[15] data_rdata_i[16] data_rdata_i[17] data_rdata_i[18]
+ data_rdata_i[19] data_rdata_i[1] data_rdata_i[20] data_rdata_i[21] data_rdata_i[22]
+ data_rdata_i[23] data_rdata_i[24] data_rdata_i[25] data_rdata_i[26] data_rdata_i[27]
+ data_rdata_i[28] data_rdata_i[29] data_rdata_i[2] data_rdata_i[30] data_rdata_i[31]
+ data_rdata_i[3] data_rdata_i[4] data_rdata_i[5] data_rdata_i[6] data_rdata_i[7]
+ data_rdata_i[8] data_rdata_i[9] data_req_o data_rvalid_i data_wdata_o[0] data_wdata_o[10]
+ data_wdata_o[11] data_wdata_o[12] data_wdata_o[13] data_wdata_o[14] data_wdata_o[15]
+ data_wdata_o[16] data_wdata_o[17] data_wdata_o[18] data_wdata_o[19] data_wdata_o[1]
+ data_wdata_o[20] data_wdata_o[21] data_wdata_o[22] data_wdata_o[23] data_wdata_o[24]
+ data_wdata_o[25] data_wdata_o[26] data_wdata_o[27] data_wdata_o[28] data_wdata_o[29]
+ data_wdata_o[2] data_wdata_o[30] data_wdata_o[31] data_wdata_o[3] data_wdata_o[4]
+ data_wdata_o[5] data_wdata_o[6] data_wdata_o[7] data_wdata_o[8] data_wdata_o[9]
+ data_we_o rst_i rx_i tx_o uart_error vccd1 vssd1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0965__B1 _1780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1142__B1 data_rdata_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1874__CLK _1875_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1270_ _1270_/A vssd1 vssd1 vccd1 vccd1 _1414_/A sky130_fd_sc_hd__inv_2
XFILLER_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0985_ _0985_/A _1777_/Q _1778_/Q vssd1 vssd1 vccd1 vccd1 _1023_/C sky130_fd_sc_hd__or3b_2
X_1606_ _1691_/X _1592_/X _1232_/B _1605_/X vssd1 vssd1 vccd1 vccd1 _1606_/Y sky130_fd_sc_hd__o22ai_2
X_1399_ _1710_/X _1186_/X _1790_/Q _1397_/X vssd1 vssd1 vccd1 vccd1 _1790_/D sky130_fd_sc_hd__o22a_2
X_1468_ _1468_/A _1468_/B vssd1 vssd1 vccd1 vccd1 _1468_/Y sky130_fd_sc_hd__nor2_2
X_1537_ _1537_/A vssd1 vssd1 vccd1 vccd1 _1538_/B sky130_fd_sc_hd__buf_1
XFILLER_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0938__B1 _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1418__A1 _1777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1322_ _1325_/A vssd1 vssd1 vccd1 vccd1 _1323_/A sky130_fd_sc_hd__buf_1
X_1253_ _1689_/X _1253_/B _1253_/C _1253_/D vssd1 vssd1 vccd1 vccd1 _1254_/A sky130_fd_sc_hd__or4_2
XANTENNA__1106__B1 data_rdata_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1184_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1195_/A sky130_fd_sc_hd__inv_2
XANTENNA__1409__A1 _1784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0968_ _0968_/A vssd1 vssd1 vccd1 vccd1 _0968_/X sky130_fd_sc_hd__buf_1
X_0899_ data_wdata_o[18] _0893_/X _1779_/Q _0894_/X vssd1 vssd1 vccd1 vccd1 _1903_/D
+ sky130_fd_sc_hd__a22o_2
XANTENNA__1345__B1 _1784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1336__B1 _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1871_ _1904_/CLK _1871_/D vssd1 vssd1 vccd1 vccd1 _1871_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1305_ data_addr_o[8] _1292_/X _1777_/Q _1294_/A vssd1 vssd1 vccd1 vccd1 _1821_/D
+ sky130_fd_sc_hd__a22o_2
X_1236_ _1688_/X vssd1 vssd1 vccd1 vccd1 _1238_/B sky130_fd_sc_hd__inv_2
XFILLER_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1098_ _1867_/Q _1095_/X data_rdata_i[26] _1096_/X _1093_/X vssd1 vssd1 vccd1 vccd1
+ _1867_/D sky130_fd_sc_hd__o221a_2
X_1167_ _1755_/Q _1756_/Q vssd1 vssd1 vccd1 vccd1 _1530_/B sky130_fd_sc_hd__or2_2
XANTENNA__1318__B1 _1783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1021_ _1021_/A uart_error vssd1 vssd1 vccd1 vccd1 _1021_/X sky130_fd_sc_hd__or2_2
X_1785_ _1835_/CLK _1785_/D vssd1 vssd1 vccd1 vccd1 tx_o sky130_fd_sc_hd__dfxtp_2
X_1854_ _1903_/CLK _1854_/D vssd1 vssd1 vccd1 vccd1 _1854_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1219_ _1219_/A vssd1 vssd1 vccd1 vccd1 _1258_/B sky130_fd_sc_hd__inv_2
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _1570_/A vssd1 vssd1 vccd1 vccd1 _1570_/X sky130_fd_sc_hd__buf_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1004_ data_req_o _1837_/Q _1021_/A _1004_/D vssd1 vssd1 vccd1 vccd1 _1428_/C sky130_fd_sc_hd__or4_2
X_1906_ _1908_/CLK _1906_/D _0886_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[21] sky130_fd_sc_hd__dfrtp_2
X_1768_ _1888_/CLK _1768_/D vssd1 vssd1 vccd1 vccd1 _1768_/Q sky130_fd_sc_hd__dfxtp_2
X_1837_ _1840_/CLK _1837_/D vssd1 vssd1 vccd1 vccd1 _1837_/Q sky130_fd_sc_hd__dfxtp_2
X_1699_ _1842_/Q _1850_/Q _1796_/Q vssd1 vssd1 vccd1 vccd1 _1699_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1622_ _1657_/X _1714_/S _1725_/S _1621_/X vssd1 vssd1 vccd1 vccd1 _1622_/X sky130_fd_sc_hd__a22o_2
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1553_ _1553_/A vssd1 vssd1 vccd1 vccd1 _1554_/B sky130_fd_sc_hd__buf_1
X_1484_ _1600_/A _1484_/B vssd1 vssd1 vccd1 vccd1 _1485_/A sky130_fd_sc_hd__or2_2
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_12_0_clk_i clkbuf_3_6_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1859_/CLK sky130_fd_sc_hd__clkbuf_2
X_0984_ _1778_/Q _0985_/A _1777_/Q vssd1 vssd1 vccd1 vccd1 _1468_/A sky130_fd_sc_hd__or3b_2
X_1536_ _1758_/Q _1530_/X _1540_/B vssd1 vssd1 vccd1 vccd1 _1537_/A sky130_fd_sc_hd__a21bo_2
XFILLER_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1605_ _1605_/A _1646_/X vssd1 vssd1 vccd1 vccd1 _1605_/X sky130_fd_sc_hd__and2_2
X_1398_ _1709_/X _1186_/X _1791_/Q _1397_/X vssd1 vssd1 vccd1 vccd1 _1791_/D sky130_fd_sc_hd__o22a_2
XFILLER_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1467_ _1278_/A _1358_/A _0871_/A _0946_/B vssd1 vssd1 vccd1 vccd1 _1803_/D sky130_fd_sc_hd__o22ai_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0938__A1 data_wdata_o[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1321_ data_wdata_o[29] _1310_/X _1782_/Q _1312_/X vssd1 vssd1 vccd1 vccd1 _1818_/D
+ sky130_fd_sc_hd__a22o_2
X_1252_ _1589_/B vssd1 vssd1 vccd1 vccd1 _1253_/D sky130_fd_sc_hd__inv_2
X_1183_ _1613_/A _1196_/A _1613_/B _1405_/B vssd1 vssd1 vccd1 vccd1 _1397_/A sky130_fd_sc_hd__o211a_2
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1042__B1 _1781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0967_ _0976_/A vssd1 vssd1 vccd1 vccd1 _0968_/A sky130_fd_sc_hd__buf_1
X_0898_ _0898_/A vssd1 vssd1 vccd1 vccd1 _0898_/X sky130_fd_sc_hd__buf_1
X_1519_ _1775_/Q _1514_/X _1243_/Y vssd1 vssd1 vccd1 vccd1 _1521_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__1345__A1 data_addr_o[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1336__A1 data_wdata_o[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1870_ _1904_/CLK _1870_/D vssd1 vssd1 vccd1 vccd1 _1870_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1304_ _1304_/A vssd1 vssd1 vccd1 vccd1 _1304_/X sky130_fd_sc_hd__buf_1
X_1235_ _1692_/X vssd1 vssd1 vccd1 vccd1 _1600_/B sky130_fd_sc_hd__inv_4
X_1166_ _1738_/Q vssd1 vssd1 vccd1 vccd1 _1166_/Y sky130_fd_sc_hd__inv_2
X_1097_ _1868_/Q _1095_/X data_rdata_i[27] _1096_/X _1093_/X vssd1 vssd1 vccd1 vccd1
+ _1868_/D sky130_fd_sc_hd__o221a_2
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1318__A1 data_wdata_o[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1020_ _1784_/Q _1020_/B _1782_/Q vssd1 vssd1 vccd1 vccd1 _1469_/B sky130_fd_sc_hd__or3b_2
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1784_ _1895_/CLK _1784_/D vssd1 vssd1 vccd1 vccd1 _1784_/Q sky130_fd_sc_hd__dfxtp_2
X_1853_ _1895_/CLK _1853_/D vssd1 vssd1 vccd1 vccd1 _1853_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1218_ _1828_/Q _1827_/Q vssd1 vssd1 vccd1 vccd1 _1219_/A sky130_fd_sc_hd__or2_2
X_1149_ _1831_/Q vssd1 vssd1 vccd1 vccd1 _1149_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1003_ _1825_/Q data_rvalid_i data_gnt_i vssd1 vssd1 vccd1 vccd1 _1004_/D sky130_fd_sc_hd__or3_2
X_1905_ _1908_/CLK _1905_/D _0889_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[20] sky130_fd_sc_hd__dfrtp_2
X_1698_ _1697_/X _1871_/Q _1794_/Q vssd1 vssd1 vccd1 vccd1 _1698_/X sky130_fd_sc_hd__mux2_1
X_1836_ _1881_/CLK _1836_/D vssd1 vssd1 vccd1 vccd1 _1836_/Q sky130_fd_sc_hd__dfxtp_2
X_1767_ _1830_/CLK _1767_/D vssd1 vssd1 vccd1 vccd1 _1767_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1621_ _1837_/Q _1652_/X vssd1 vssd1 vccd1 vccd1 _1621_/X sky130_fd_sc_hd__or2_2
X_1552_ _1761_/Q _1545_/X _1551_/X vssd1 vssd1 vccd1 vccd1 _1553_/A sky130_fd_sc_hd__a21bo_2
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1483_ _1595_/A vssd1 vssd1 vccd1 vccd1 _1600_/A sky130_fd_sc_hd__buf_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1819_ _1908_/CLK _1819_/D _1317_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[30] sky130_fd_sc_hd__dfrtp_2
XFILLER_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0983_ _1784_/Q _1020_/B _0983_/C vssd1 vssd1 vccd1 vccd1 _0985_/A sky130_fd_sc_hd__or3_2
XFILLER_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1604_ _1604_/A vssd1 vssd1 vccd1 vccd1 _1604_/X sky130_fd_sc_hd__buf_1
X_1535_ _1535_/A vssd1 vssd1 vccd1 vccd1 _1535_/X sky130_fd_sc_hd__buf_1
X_1397_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1397_/X sky130_fd_sc_hd__buf_1
X_1466_ _1743_/Q _1463_/A _1465_/Y _1463_/Y vssd1 vssd1 vccd1 vccd1 _1466_/X sky130_fd_sc_hd__a22o_2
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1320_ _1320_/A vssd1 vssd1 vccd1 vccd1 _1320_/X sky130_fd_sc_hd__buf_1
X_1182_ _1189_/A _1674_/S _1837_/Q _1181_/Y vssd1 vssd1 vccd1 vccd1 _1405_/B sky130_fd_sc_hd__o2bb2a_2
X_1251_ _1251_/A vssd1 vssd1 vccd1 vccd1 _1589_/B sky130_fd_sc_hd__buf_1
XFILLER_32_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0897_ _0906_/A vssd1 vssd1 vccd1 vccd1 _0898_/A sky130_fd_sc_hd__buf_1
X_0966_ _0966_/A vssd1 vssd1 vccd1 vccd1 _0976_/A sky130_fd_sc_hd__buf_1
X_1518_ _1518_/A vssd1 vssd1 vccd1 vccd1 _1518_/X sky130_fd_sc_hd__buf_1
X_1449_ _1749_/Q _1447_/B _1448_/Y vssd1 vssd1 vccd1 vccd1 _1449_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1303_ _1306_/A vssd1 vssd1 vccd1 vccd1 _1304_/A sky130_fd_sc_hd__buf_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1096_ _1111_/A vssd1 vssd1 vccd1 vccd1 _1096_/X sky130_fd_sc_hd__buf_1
X_1234_ _1691_/X vssd1 vssd1 vccd1 vccd1 _1253_/B sky130_fd_sc_hd__inv_2
X_1165_ _1652_/X _1648_/X _1647_/X vssd1 vssd1 vccd1 vccd1 _1179_/C sky130_fd_sc_hd__or3_2
X_0949_ _0964_/A vssd1 vssd1 vccd1 vccd1 _0949_/X sky130_fd_sc_hd__buf_1
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1852_ _1852_/CLK _1852_/D vssd1 vssd1 vccd1 vccd1 _1852_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1783_ _1895_/CLK _1783_/D vssd1 vssd1 vccd1 vccd1 _1783_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1079_ _1873_/Q vssd1 vssd1 vccd1 vccd1 _1079_/Y sky130_fd_sc_hd__inv_2
X_1217_ _1829_/Q vssd1 vssd1 vccd1 vccd1 _1258_/A sky130_fd_sc_hd__inv_2
X_1148_ data_we_o _1737_/X _1147_/Y _1737_/S _1145_/X vssd1 vssd1 vccd1 vccd1 _1840_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_20_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ _1002_/A vssd1 vssd1 vccd1 vccd1 _1605_/A sky130_fd_sc_hd__buf_1
X_1904_ _1904_/CLK _1904_/D _0892_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[19] sky130_fd_sc_hd__dfrtp_2
X_1835_ _1835_/CLK _1835_/D vssd1 vssd1 vccd1 vccd1 _1835_/Q sky130_fd_sc_hd__dfxtp_2
X_1697_ _1696_/X _1863_/Q _1798_/Q vssd1 vssd1 vccd1 vccd1 _1697_/X sky130_fd_sc_hd__mux2_1
X_1766_ _1851_/CLK _1766_/D vssd1 vssd1 vccd1 vccd1 _1766_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1551_ _1760_/Q _1761_/Q _1551_/C vssd1 vssd1 vccd1 vccd1 _1551_/X sky130_fd_sc_hd__or3_2
XANTENNA__1474__A rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1482_ _1482_/A vssd1 vssd1 vccd1 vccd1 _1484_/B sky130_fd_sc_hd__buf_1
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1620_ _1620_/A vssd1 vssd1 vccd1 vccd1 _1620_/X sky130_fd_sc_hd__buf_1
XFILLER_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1687__A1 rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1136__B1 data_rdata_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1818_ _1908_/CLK _1818_/D _1320_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[29] sky130_fd_sc_hd__dfrtp_2
X_1749_ _1830_/CLK _1749_/D vssd1 vssd1 vccd1 vccd1 _1749_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_4_6_0_clk_i clkbuf_4_7_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1852_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_26_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0982_ _1782_/Q _1781_/Q _1780_/Q _1779_/Q vssd1 vssd1 vccd1 vccd1 _0983_/C sky130_fd_sc_hd__or4_2
XANTENNA__1109__B1 data_rdata_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1534_ _1543_/A _1534_/B vssd1 vssd1 vccd1 vccd1 _1535_/A sky130_fd_sc_hd__and2_2
X_1603_ _1610_/A _1691_/X vssd1 vssd1 vccd1 vccd1 _1604_/A sky130_fd_sc_hd__or2_2
X_1465_ _1743_/Q vssd1 vssd1 vccd1 vccd1 _1465_/Y sky130_fd_sc_hd__inv_2
X_1396_ _1708_/X _1186_/X _1792_/Q _1187_/X vssd1 vssd1 vccd1 vccd1 _1792_/D sky130_fd_sc_hd__o22a_2
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1339__B1 _1777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1181_ _1613_/A vssd1 vssd1 vccd1 vccd1 _1181_/Y sky130_fd_sc_hd__inv_2
X_1250_ _1746_/Q _1692_/S _1746_/Q _1692_/S vssd1 vssd1 vccd1 vccd1 _1251_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0896_ _1145_/A vssd1 vssd1 vccd1 vccd1 _0906_/A sky130_fd_sc_hd__buf_1
X_0965_ data_wdata_o[3] _0963_/X _1780_/Q _0964_/X vssd1 vssd1 vccd1 vccd1 _1888_/D
+ sky130_fd_sc_hd__a22o_2
X_1517_ rx_i _1517_/B vssd1 vssd1 vccd1 vccd1 _1518_/A sky130_fd_sc_hd__and2_2
X_1448_ _1451_/B vssd1 vssd1 vccd1 vccd1 _1448_/Y sky130_fd_sc_hd__inv_2
X_1379_ _1379_/A vssd1 vssd1 vccd1 vccd1 _1379_/X sky130_fd_sc_hd__buf_1
XFILLER_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1024__A2 _1006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1302_ data_addr_o[9] _1292_/X _1778_/Q _1294_/X vssd1 vssd1 vccd1 vccd1 _1822_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1233_ rx_i _1580_/A vssd1 vssd1 vccd1 vccd1 _1233_/Y sky130_fd_sc_hd__nor2_2
X_1095_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1095_/X sky130_fd_sc_hd__buf_1
X_1164_ _1164_/A vssd1 vssd1 vccd1 vccd1 _1189_/A sky130_fd_sc_hd__inv_2
X_0948_ _0963_/A vssd1 vssd1 vccd1 vccd1 _0964_/A sky130_fd_sc_hd__inv_2
XFILLER_20_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0879_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1154_/A sky130_fd_sc_hd__buf_1
XFILLER_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1851_ _1851_/CLK _1851_/D vssd1 vssd1 vccd1 vccd1 _1851_/Q sky130_fd_sc_hd__dfxtp_2
X_1782_ _1895_/CLK _1782_/D vssd1 vssd1 vccd1 vccd1 _1782_/Q sky130_fd_sc_hd__dfxtp_2
X_1216_ _1830_/Q vssd1 vssd1 vccd1 vccd1 _1216_/Y sky130_fd_sc_hd__inv_2
X_1078_ _1065_/Y _1737_/S _1072_/B _0891_/A _1077_/Y vssd1 vssd1 vccd1 vccd1 _1874_/D
+ sky130_fd_sc_hd__o311a_2
X_1147_ _1737_/X vssd1 vssd1 vccd1 vccd1 _1147_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _1752_/Q vssd1 vssd1 vccd1 vccd1 _1220_/B sky130_fd_sc_hd__inv_2
X_1834_ _1881_/CLK _1834_/D vssd1 vssd1 vccd1 vccd1 _1834_/Q sky130_fd_sc_hd__dfxtp_2
X_1903_ _1903_/CLK _1903_/D _0898_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[18] sky130_fd_sc_hd__dfrtp_2
X_1765_ _1840_/CLK _1765_/D vssd1 vssd1 vccd1 vccd1 _1765_/Q sky130_fd_sc_hd__dfxtp_2
X_1696_ _1847_/Q _1855_/Q _1796_/Q vssd1 vssd1 vccd1 vccd1 _1696_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1090__B1 data_rdata_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_2_0_clk_i clkbuf_4_3_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1840_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1550_ _1550_/A vssd1 vssd1 vccd1 vccd1 _1550_/X sky130_fd_sc_hd__buf_1
X_1481_ _1692_/S _1481_/B vssd1 vssd1 vccd1 vccd1 _1482_/A sky130_fd_sc_hd__or2_2
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0895__B1 _1780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1817_ _1908_/CLK _1817_/D _1323_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[28] sky130_fd_sc_hd__dfrtp_2
X_1748_ _1830_/CLK _1748_/D vssd1 vssd1 vccd1 vccd1 _1748_/Q sky130_fd_sc_hd__dfxtp_2
X_1679_ _1678_/X _1859_/Q _1798_/Q vssd1 vssd1 vccd1 vccd1 _1679_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0877__B1 _1784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0981_ _1783_/Q vssd1 vssd1 vccd1 vccd1 _1020_/B sky130_fd_sc_hd__inv_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1602_ _1692_/X _1592_/B _1695_/X _1584_/A _1601_/Y vssd1 vssd1 vccd1 vccd1 _1602_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1533_ _1548_/A vssd1 vssd1 vccd1 vccd1 _1543_/A sky130_fd_sc_hd__buf_1
X_1395_ rst_i _1395_/B vssd1 vssd1 vccd1 vccd1 _1793_/D sky130_fd_sc_hd__nor2_2
X_1464_ _1742_/Q _1462_/B _1463_/Y vssd1 vssd1 vccd1 vccd1 _1464_/X sky130_fd_sc_hd__a21o_2
XFILLER_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1395__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1180_ _1180_/A vssd1 vssd1 vccd1 vccd1 _1674_/S sky130_fd_sc_hd__buf_1
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0964_ _0964_/A vssd1 vssd1 vccd1 vccd1 _0964_/X sky130_fd_sc_hd__buf_1
X_0895_ data_wdata_o[19] _0893_/X _1780_/Q _0894_/X vssd1 vssd1 vccd1 vccd1 _1904_/D
+ sky130_fd_sc_hd__a22o_2
X_1516_ _1516_/A vssd1 vssd1 vccd1 vccd1 _1517_/B sky130_fd_sc_hd__buf_1
X_1378_ _1382_/A vssd1 vssd1 vccd1 vccd1 _1379_/A sky130_fd_sc_hd__buf_1
X_1447_ _1749_/Q _1447_/B vssd1 vssd1 vccd1 vccd1 _1451_/B sky130_fd_sc_hd__or2_2
XFILLER_14_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1301_ _1301_/A vssd1 vssd1 vccd1 vccd1 _1301_/X sky130_fd_sc_hd__buf_1
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1232_ _1754_/Q _1232_/B vssd1 vssd1 vccd1 vccd1 _1580_/A sky130_fd_sc_hd__or2_2
X_1094_ _1869_/Q _1086_/X data_rdata_i[28] _1088_/X _1093_/X vssd1 vssd1 vccd1 vccd1
+ _1869_/D sky130_fd_sc_hd__o221a_2
X_1163_ _1163_/A vssd1 vssd1 vccd1 vccd1 _1196_/A sky130_fd_sc_hd__buf_1
X_0947_ _0963_/A vssd1 vssd1 vccd1 vccd1 _0947_/X sky130_fd_sc_hd__buf_1
X_0878_ rst_i vssd1 vssd1 vccd1 vccd1 _1155_/A sky130_fd_sc_hd__inv_2
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1411__B1 _1783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1850_ _1852_/CLK _1850_/D vssd1 vssd1 vccd1 vccd1 _1850_/Q sky130_fd_sc_hd__dfxtp_2
X_1781_ _1895_/CLK _1781_/D vssd1 vssd1 vccd1 vccd1 _1781_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1493__A rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1146_ _1841_/Q _1140_/X data_rdata_i[0] _1141_/X _1145_/X vssd1 vssd1 vccd1 vccd1
+ _1841_/D sky130_fd_sc_hd__o221a_2
X_1215_ rst_i _1215_/B vssd1 vssd1 vccd1 vccd1 _1831_/D sky130_fd_sc_hd__nor2_2
X_1077_ _1065_/Y _1737_/S _1067_/A vssd1 vssd1 vccd1 vccd1 _1077_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1000_ _1000_/A vssd1 vssd1 vccd1 vccd1 _1000_/X sky130_fd_sc_hd__buf_1
X_1902_ _1908_/CLK _1902_/D _0901_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[17] sky130_fd_sc_hd__dfrtp_2
XANTENNA__1488__A rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1833_ _1881_/CLK _1833_/D vssd1 vssd1 vccd1 vccd1 _1833_/Q sky130_fd_sc_hd__dfxtp_2
X_1764_ _1771_/CLK _1764_/D vssd1 vssd1 vccd1 vccd1 _1764_/Q sky130_fd_sc_hd__dfxtp_2
X_1695_ _1692_/X _1600_/Y _1695_/S vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1129_ _1851_/Q _1126_/X data_rdata_i[10] _1127_/X _1124_/X vssd1 vssd1 vccd1 vccd1
+ _1851_/D sky130_fd_sc_hd__o221a_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1247_/C _1767_/Q _1766_/Q _1479_/Y vssd1 vssd1 vccd1 vccd1 _1481_/B sky130_fd_sc_hd__o22a_2
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1816_ _1908_/CLK _1816_/D _1326_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[27] sky130_fd_sc_hd__dfrtp_2
X_1747_ _1830_/CLK _1747_/D vssd1 vssd1 vccd1 vccd1 _1747_/Q sky130_fd_sc_hd__dfxtp_2
X_1678_ _1843_/Q _1851_/Q _1796_/Q vssd1 vssd1 vccd1 vccd1 _1678_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0980_ _1371_/B vssd1 vssd1 vccd1 vccd1 _0980_/X sky130_fd_sc_hd__buf_1
X_1532_ _1532_/A vssd1 vssd1 vccd1 vccd1 _1534_/B sky130_fd_sc_hd__buf_1
X_1601_ _1600_/B _1695_/S _1229_/Y vssd1 vssd1 vccd1 vccd1 _1601_/Y sky130_fd_sc_hd__o21ai_2
X_1394_ _1394_/A vssd1 vssd1 vccd1 vccd1 _1394_/X sky130_fd_sc_hd__buf_1
X_1463_ _1463_/A vssd1 vssd1 vccd1 vccd1 _1463_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0894_ _0894_/A vssd1 vssd1 vccd1 vccd1 _0894_/X sky130_fd_sc_hd__buf_1
XFILLER_32_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0963_ _0963_/A vssd1 vssd1 vccd1 vccd1 _0963_/X sky130_fd_sc_hd__buf_1
X_1515_ _1774_/Q _1514_/B _1514_/X vssd1 vssd1 vccd1 vccd1 _1516_/A sky130_fd_sc_hd__a21bo_2
X_1377_ _1377_/A vssd1 vssd1 vccd1 vccd1 _1377_/X sky130_fd_sc_hd__buf_1
X_1446_ _1749_/Q vssd1 vssd1 vccd1 vccd1 _1446_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1300_ _1306_/A vssd1 vssd1 vccd1 vccd1 _1301_/A sky130_fd_sc_hd__buf_1
X_1162_ _1835_/Q _1201_/A _1836_/Q vssd1 vssd1 vccd1 vccd1 _1163_/A sky130_fd_sc_hd__or3_2
X_1231_ _1576_/A _1581_/B vssd1 vssd1 vccd1 vccd1 _1232_/B sky130_fd_sc_hd__or2_2
X_1093_ _1628_/A vssd1 vssd1 vccd1 vccd1 _1093_/X sky130_fd_sc_hd__buf_1
XFILLER_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1003__B data_rvalid_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0877_ data_wdata_o[23] _0874_/X _1784_/Q _0876_/X vssd1 vssd1 vccd1 vccd1 _1908_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0946_ _1803_/Q _0946_/B vssd1 vssd1 vccd1 vccd1 _0963_/A sky130_fd_sc_hd__nand2_2
X_1429_ _1275_/X _1420_/X _1800_/Q _1428_/X vssd1 vssd1 vccd1 vccd1 _1800_/D sky130_fd_sc_hd__a2bb2o_2
XANTENNA__0931__B1 _1780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1411__A1 _1782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1780_ _1895_/CLK _1780_/D vssd1 vssd1 vccd1 vccd1 _1780_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1145_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1145_/X sky130_fd_sc_hd__buf_1
X_1214_ _1831_/Q _1069_/A _1149_/Y _1150_/X vssd1 vssd1 vccd1 vccd1 _1215_/B sky130_fd_sc_hd__o22a_2
X_1076_ _1076_/A vssd1 vssd1 vccd1 vccd1 _1737_/S sky130_fd_sc_hd__buf_1
X_0929_ _0929_/A vssd1 vssd1 vccd1 vccd1 _0929_/X sky130_fd_sc_hd__buf_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1901_ _1903_/CLK _1901_/D _0904_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[16] sky130_fd_sc_hd__dfrtp_2
X_1832_ _1835_/CLK _1832_/D _1212_/X vssd1 vssd1 vccd1 vccd1 _1832_/Q sky130_fd_sc_hd__dfrtp_2
X_1694_ _1581_/A rx_i _1695_/S vssd1 vssd1 vccd1 vccd1 _1694_/X sky130_fd_sc_hd__mux2_1
X_1763_ _1771_/CLK _1763_/D vssd1 vssd1 vccd1 vccd1 _1763_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_clkbuf_3_4_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1139__B1 data_rdata_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1059_ _1059_/A vssd1 vssd1 vccd1 vccd1 _1059_/X sky130_fd_sc_hd__buf_1
X_1128_ _1852_/Q _1126_/X data_rdata_i[11] _1127_/X _1124_/X vssd1 vssd1 vccd1 vccd1
+ _1852_/D sky130_fd_sc_hd__o221a_2
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1614__B2 _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1075__C1 rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1302__B1 _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1815_ _1908_/CLK _1815_/D _1332_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[26] sky130_fd_sc_hd__dfrtp_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1677_ _1676_/X _1870_/Q _1794_/Q vssd1 vssd1 vccd1 vccd1 _1677_/X sky130_fd_sc_hd__mux2_1
X_1746_ _1830_/CLK _1746_/D vssd1 vssd1 vccd1 vccd1 _1746_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1600_ _1600_/A _1600_/B vssd1 vssd1 vccd1 vccd1 _1600_/Y sky130_fd_sc_hd__nor2_2
X_1531_ _1757_/Q _1530_/B _1530_/X vssd1 vssd1 vccd1 vccd1 _1532_/A sky130_fd_sc_hd__a21bo_2
X_1462_ _1742_/Q _1462_/B vssd1 vssd1 vccd1 vccd1 _1463_/A sky130_fd_sc_hd__or2_2
X_1393_ _1628_/A vssd1 vssd1 vccd1 vccd1 _1394_/A sky130_fd_sc_hd__buf_1
XANTENNA__1721__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1729_ _1512_/B _1513_/X _1736_/S vssd1 vssd1 vccd1 vccd1 _1773_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0893_ _0893_/A vssd1 vssd1 vccd1 vccd1 _0893_/X sky130_fd_sc_hd__buf_1
X_0962_ _0962_/A vssd1 vssd1 vccd1 vccd1 _0962_/X sky130_fd_sc_hd__buf_1
X_1514_ _1774_/Q _1514_/B vssd1 vssd1 vccd1 vccd1 _1514_/X sky130_fd_sc_hd__or2_2
X_1445_ _1443_/Y _1441_/Y _1447_/B vssd1 vssd1 vccd1 vccd1 _1445_/X sky130_fd_sc_hd__o21a_2
XANTENNA__1716__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1376_ _1382_/A vssd1 vssd1 vccd1 vccd1 _1377_/A sky130_fd_sc_hd__buf_1
XANTENNA__1801__CLK _1875_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1092_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1628_/A sky130_fd_sc_hd__buf_1
X_1161_ _1834_/Q _1833_/Q vssd1 vssd1 vccd1 vccd1 _1201_/A sky130_fd_sc_hd__or2_2
X_1230_ _1581_/A vssd1 vssd1 vccd1 vccd1 _1576_/A sky130_fd_sc_hd__inv_2
XANTENNA__1824__CLK _1875_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1003__C data_gnt_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0876_ _0894_/A vssd1 vssd1 vccd1 vccd1 _0876_/X sky130_fd_sc_hd__buf_1
X_0945_ _1013_/C _0945_/B _1797_/Q _1276_/A vssd1 vssd1 vccd1 vccd1 _0946_/B sky130_fd_sc_hd__and4b_2
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1428_ _1428_/A _1428_/B _1428_/C vssd1 vssd1 vccd1 vccd1 _1428_/X sky130_fd_sc_hd__or3_2
X_1359_ _1434_/B vssd1 vssd1 vccd1 vccd1 _1359_/X sky130_fd_sc_hd__buf_1
XFILLER_18_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1213_ _0980_/X _0991_/X _1832_/Q _0995_/B vssd1 vssd1 vccd1 vccd1 _1832_/D sky130_fd_sc_hd__a2bb2o_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1144_ _1842_/Q _1140_/X data_rdata_i[1] _1141_/X _1138_/X vssd1 vssd1 vccd1 vccd1
+ _1842_/D sky130_fd_sc_hd__o221a_2
X_1075_ _1083_/A _1073_/Y _1420_/C _1073_/A rst_i vssd1 vssd1 vccd1 vccd1 _1875_/D
+ sky130_fd_sc_hd__a221oi_2
X_0928_ _0928_/A vssd1 vssd1 vccd1 vccd1 _0928_/X sky130_fd_sc_hd__buf_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1148__A1 data_we_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1900_ _1903_/CLK _1900_/D _0907_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[15] sky130_fd_sc_hd__dfrtp_2
XANTENNA__1623__A2 _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1831_ _1840_/CLK _1831_/D vssd1 vssd1 vccd1 vccd1 _1831_/Q sky130_fd_sc_hd__dfxtp_2
X_1762_ _1771_/CLK _1762_/D vssd1 vssd1 vccd1 vccd1 _1762_/Q sky130_fd_sc_hd__dfxtp_2
X_1693_ _1581_/A _1521_/A _1695_/S vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1724__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1058_ _1058_/A vssd1 vssd1 vccd1 vccd1 _1059_/A sky130_fd_sc_hd__buf_1
X_1127_ _1141_/A vssd1 vssd1 vccd1 vccd1 _1127_/X sky130_fd_sc_hd__buf_1
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1814_ _1908_/CLK _1814_/D _1335_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[25] sky130_fd_sc_hd__dfrtp_2
X_1745_ _1835_/CLK _1745_/D vssd1 vssd1 vccd1 vccd1 _1745_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1719__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1676_ _1675_/X _1862_/Q _1798_/Q vssd1 vssd1 vccd1 vccd1 _1676_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1048__B1 _1780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1599__A1 rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1530_ _1757_/Q _1530_/B vssd1 vssd1 vccd1 vccd1 _1530_/X sky130_fd_sc_hd__or2_2
X_1392_ _1392_/A vssd1 vssd1 vccd1 vccd1 _1392_/X sky130_fd_sc_hd__buf_1
X_1461_ _1741_/Q _1460_/B _1462_/B vssd1 vssd1 vccd1 vccd1 _1461_/X sky130_fd_sc_hd__a21bo_2
XFILLER_50_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1728_ _1517_/B _1518_/X _1736_/S vssd1 vssd1 vccd1 vccd1 _1774_/D sky130_fd_sc_hd__mux2_1
X_1659_ _1599_/Y _1689_/X _1681_/X vssd1 vssd1 vccd1 vccd1 _1747_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0961_ _0961_/A vssd1 vssd1 vccd1 vccd1 _0962_/A sky130_fd_sc_hd__buf_1
X_0892_ _0892_/A vssd1 vssd1 vccd1 vccd1 _0892_/X sky130_fd_sc_hd__buf_1
X_1375_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1382_/A sky130_fd_sc_hd__buf_1
X_1513_ _1513_/A vssd1 vssd1 vccd1 vccd1 _1513_/X sky130_fd_sc_hd__buf_1
X_1444_ _1748_/Q _1444_/B vssd1 vssd1 vccd1 vccd1 _1447_/B sky130_fd_sc_hd__or2_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1091_ _1870_/Q _1086_/X data_rdata_i[29] _1088_/X _0881_/X vssd1 vssd1 vccd1 vccd1
+ _1870_/D sky130_fd_sc_hd__o221a_2
X_1160_ _1160_/A vssd1 vssd1 vccd1 vccd1 _1613_/A sky130_fd_sc_hd__buf_1
X_0944_ _1017_/A vssd1 vssd1 vccd1 vccd1 _1276_/A sky130_fd_sc_hd__inv_2
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0875_ _0893_/A vssd1 vssd1 vccd1 vccd1 _0894_/A sky130_fd_sc_hd__inv_2
X_1358_ _1358_/A vssd1 vssd1 vccd1 vccd1 _1358_/X sky130_fd_sc_hd__buf_1
X_1427_ _1795_/Q vssd1 vssd1 vccd1 vccd1 _1428_/A sky130_fd_sc_hd__inv_2
X_1289_ _1289_/A vssd1 vssd1 vccd1 vccd1 _1290_/A sky130_fd_sc_hd__buf_1
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1212_ _1212_/A vssd1 vssd1 vccd1 vccd1 _1212_/X sky130_fd_sc_hd__buf_1
X_1074_ _1875_/Q vssd1 vssd1 vccd1 vccd1 _1420_/C sky130_fd_sc_hd__inv_2
X_1143_ _1843_/Q _1140_/X data_rdata_i[2] _1141_/X _1138_/X vssd1 vssd1 vccd1 vccd1
+ _1843_/D sky130_fd_sc_hd__o221a_2
X_0927_ _0927_/A vssd1 vssd1 vccd1 vccd1 _0928_/A sky130_fd_sc_hd__buf_1
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1761_ _1771_/CLK _1761_/D vssd1 vssd1 vccd1 vccd1 _1761_/Q sky130_fd_sc_hd__dfxtp_2
X_1830_ _1830_/CLK _1830_/D vssd1 vssd1 vccd1 vccd1 _1830_/Q sky130_fd_sc_hd__dfxtp_2
X_1692_ _1443_/Y _1445_/X _1692_/S vssd1 vssd1 vccd1 vccd1 _1692_/X sky130_fd_sc_hd__mux2_1
X_1126_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1126_/X sky130_fd_sc_hd__buf_1
X_1057_ _1057_/A vssd1 vssd1 vccd1 vccd1 _1877_/D sky130_fd_sc_hd__buf_1
XFILLER_40_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1813_ _1908_/CLK _1813_/D _1338_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[24] sky130_fd_sc_hd__dfrtp_2
X_1744_ _1835_/CLK _1744_/D vssd1 vssd1 vccd1 vccd1 _1744_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1675_ _1846_/Q _1854_/Q _1796_/Q vssd1 vssd1 vccd1 vccd1 _1675_/X sky130_fd_sc_hd__mux2_1
X_1109_ _1861_/Q _1102_/X data_rdata_i[20] _1103_/X _1108_/X vssd1 vssd1 vccd1 vccd1
+ _1861_/D sky130_fd_sc_hd__o221a_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1391_ _1391_/A vssd1 vssd1 vccd1 vccd1 _1392_/A sky130_fd_sc_hd__buf_1
X_1460_ _1741_/Q _1460_/B vssd1 vssd1 vccd1 vccd1 _1462_/B sky130_fd_sc_hd__or2_2
X_1658_ _1593_/Y _1253_/D _1681_/X vssd1 vssd1 vccd1 vccd1 _1746_/D sky130_fd_sc_hd__mux2_1
X_1727_ _1520_/Y _1521_/Y _1736_/S vssd1 vssd1 vccd1 vccd1 _1775_/D sky130_fd_sc_hd__mux2_1
X_1589_ _1600_/A _1589_/B vssd1 vssd1 vccd1 vccd1 _1590_/A sky130_fd_sc_hd__or2_2
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0960_ data_wdata_o[4] _0947_/X _1781_/Q _0949_/X vssd1 vssd1 vccd1 vccd1 _1889_/D
+ sky130_fd_sc_hd__a22o_2
X_0891_ _0891_/A vssd1 vssd1 vccd1 vccd1 _0892_/A sky130_fd_sc_hd__buf_1
X_1512_ rx_i _1512_/B vssd1 vssd1 vccd1 vccd1 _1513_/A sky130_fd_sc_hd__and2_2
XFILLER_4_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1443_ _1748_/Q vssd1 vssd1 vccd1 vccd1 _1443_/Y sky130_fd_sc_hd__inv_2
X_1374_ _1374_/A vssd1 vssd1 vccd1 vccd1 _1374_/X sky130_fd_sc_hd__buf_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1090_ _1871_/Q _1086_/X data_rdata_i[30] _1088_/X _0881_/X vssd1 vssd1 vccd1 vccd1
+ _1871_/D sky130_fd_sc_hd__o221a_2
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0874_ _0893_/A vssd1 vssd1 vccd1 vccd1 _0874_/X sky130_fd_sc_hd__buf_1
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0943_ _0943_/A vssd1 vssd1 vccd1 vccd1 _0943_/X sky130_fd_sc_hd__buf_1
X_1288_ _1288_/A vssd1 vssd1 vccd1 vccd1 _1825_/D sky130_fd_sc_hd__buf_1
X_1426_ _0873_/B _1423_/X _0945_/B _1425_/X vssd1 vssd1 vccd1 vccd1 _1796_/D sky130_fd_sc_hd__o22ai_2
X_1357_ _1357_/A vssd1 vssd1 vccd1 vccd1 _1357_/X sky130_fd_sc_hd__buf_1
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1571__B1 _1777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1211_ _1289_/A vssd1 vssd1 vccd1 vccd1 _1212_/A sky130_fd_sc_hd__buf_1
X_1142_ _1844_/Q _1140_/X data_rdata_i[3] _1141_/X _1138_/X vssd1 vssd1 vccd1 vccd1
+ _1844_/D sky130_fd_sc_hd__o221a_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1073_ _1073_/A vssd1 vssd1 vccd1 vccd1 _1073_/Y sky130_fd_sc_hd__inv_2
X_0926_ data_wdata_o[12] _0911_/X _1781_/Q _0913_/X vssd1 vssd1 vccd1 vccd1 _1897_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0878__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1409_ _1784_/Q _1407_/X rx_i _1408_/X vssd1 vssd1 vccd1 vccd1 _1784_/D sky130_fd_sc_hd__a22o_2
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1305__B1 _1777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1760_ _1771_/CLK _1760_/D vssd1 vssd1 vccd1 vccd1 _1760_/Q sky130_fd_sc_hd__dfxtp_2
X_1691_ _1446_/Y _1449_/Y _1692_/S vssd1 vssd1 vccd1 vccd1 _1691_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1125_ _1853_/Q _1118_/X data_rdata_i[12] _1120_/X _1124_/X vssd1 vssd1 vccd1 vccd1
+ _1853_/D sky130_fd_sc_hd__o221a_2
X_1056_ _1641_/X _1877_/Q _1060_/S vssd1 vssd1 vccd1 vccd1 _1057_/A sky130_fd_sc_hd__mux2_2
X_0909_ _1794_/Q _1798_/Q vssd1 vssd1 vccd1 vccd1 _1013_/C sky130_fd_sc_hd__or2_2
X_1889_ _1892_/CLK _1889_/D _0959_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[4] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1066__A2 data_gnt_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0981__A _1783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1674_ _1404_/B _1672_/S _1674_/S vssd1 vssd1 vccd1 vccd1 _1674_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1812_ _1852_/CLK _1812_/D _1341_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[7] sky130_fd_sc_hd__dfrtp_2
X_1743_ _1840_/CLK _1743_/D vssd1 vssd1 vccd1 vccd1 _1743_/Q sky130_fd_sc_hd__dfxtp_2
X_1039_ _1039_/A vssd1 vssd1 vccd1 vccd1 _1881_/D sky130_fd_sc_hd__buf_1
XANTENNA__0891__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1108_ _1131_/A vssd1 vssd1 vccd1 vccd1 _1108_/X sky130_fd_sc_hd__buf_1
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1390_ _1390_/A vssd1 vssd1 vccd1 vccd1 _1390_/X sky130_fd_sc_hd__buf_1
X_1657_ _1196_/A _1652_/X _1674_/S vssd1 vssd1 vccd1 vccd1 _1657_/X sky130_fd_sc_hd__mux2_1
X_1726_ _1249_/A _1522_/Y _1736_/S vssd1 vssd1 vccd1 vccd1 _1776_/D sky130_fd_sc_hd__mux2_1
X_1588_ _1683_/S _1581_/X _1232_/B _1586_/X _1587_/X vssd1 vssd1 vccd1 vccd1 _1588_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_26_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0890_ data_wdata_o[20] _0874_/X _1781_/Q _0876_/X vssd1 vssd1 vccd1 vccd1 _1905_/D
+ sky130_fd_sc_hd__a22o_2
X_1511_ _1509_/Y _1505_/Y _1514_/B vssd1 vssd1 vccd1 vccd1 _1512_/B sky130_fd_sc_hd__o21ai_2
XFILLER_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1442_ _1746_/Q _1747_/Q _1441_/Y vssd1 vssd1 vccd1 vccd1 _1442_/X sky130_fd_sc_hd__a21o_2
X_1373_ _1373_/A vssd1 vssd1 vccd1 vccd1 _1374_/A sky130_fd_sc_hd__buf_1
XANTENNA__1330__A _1361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk_i clkbuf_3_7_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1908_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1709_ _1881_/Q _1792_/Q _1714_/S vssd1 vssd1 vccd1 vccd1 _1709_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1150__A data_gnt_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0873_ _1794_/Q _0873_/B _1471_/B vssd1 vssd1 vccd1 vccd1 _0893_/A sky130_fd_sc_hd__or3_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0942_ _0942_/A vssd1 vssd1 vccd1 vccd1 _0943_/A sky130_fd_sc_hd__buf_1
X_1425_ _1422_/A _1016_/B _1275_/X _1420_/B _1424_/X vssd1 vssd1 vccd1 vccd1 _1425_/X
+ sky130_fd_sc_hd__o221a_2
X_1287_ _1825_/Q _1649_/X _1287_/S vssd1 vssd1 vccd1 vccd1 _1288_/A sky130_fd_sc_hd__mux2_2
X_1356_ _1356_/A vssd1 vssd1 vccd1 vccd1 _1357_/A sky130_fd_sc_hd__buf_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0984__A _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1210_ _1296_/A vssd1 vssd1 vccd1 vccd1 _1289_/A sky130_fd_sc_hd__buf_1
XFILLER_1_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1141_ _1141_/A vssd1 vssd1 vccd1 vccd1 _1141_/X sky130_fd_sc_hd__buf_1
X_1072_ _1076_/A _1072_/B vssd1 vssd1 vccd1 vccd1 _1073_/A sky130_fd_sc_hd__or2_2
X_0925_ _0925_/A vssd1 vssd1 vccd1 vccd1 _0925_/X sky130_fd_sc_hd__buf_1
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1408_ _1414_/A vssd1 vssd1 vccd1 vccd1 _1408_/X sky130_fd_sc_hd__buf_1
X_1339_ data_wdata_o[24] _1327_/X _1777_/Q _1328_/X vssd1 vssd1 vccd1 vccd1 _1813_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1078__B1 _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1305__A1 data_addr_o[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1690_ _1450_/Y _1452_/X _1692_/S vssd1 vssd1 vccd1 vccd1 _1690_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1055_ _1055_/A vssd1 vssd1 vccd1 vccd1 _1055_/X sky130_fd_sc_hd__buf_1
X_1124_ _1131_/A vssd1 vssd1 vccd1 vccd1 _1124_/X sky130_fd_sc_hd__buf_1
X_0908_ _1796_/Q vssd1 vssd1 vccd1 vccd1 _0945_/B sky130_fd_sc_hd__inv_2
X_1888_ _1888_/CLK _1888_/D _0962_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[3] sky130_fd_sc_hd__dfrtp_2
XANTENNA__1299__B1 _1779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1811_ _1892_/CLK _1811_/D _1348_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[6] sky130_fd_sc_hd__dfrtp_2
XFILLER_7_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1673_ _1690_/X _1608_/X _1695_/S vssd1 vssd1 vccd1 vccd1 _1673_/X sky130_fd_sc_hd__mux2_1
X_1742_ _1840_/CLK _1742_/D vssd1 vssd1 vccd1 vccd1 _1742_/Q sky130_fd_sc_hd__dfxtp_2
X_1038_ _1642_/X _1881_/Q _1047_/A vssd1 vssd1 vccd1 vccd1 _1039_/A sky130_fd_sc_hd__mux2_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1107_ _1314_/A vssd1 vssd1 vccd1 vccd1 _1131_/A sky130_fd_sc_hd__buf_1
XFILLER_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1725_ _1176_/A _1523_/Y _1725_/S vssd1 vssd1 vccd1 vccd1 _1755_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_4_11_0_clk_i clkbuf_3_5_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1883_/CLK sky130_fd_sc_hd__clkbuf_2
X_1587_ _1752_/Q _1753_/Q _1587_/C _1695_/S vssd1 vssd1 vccd1 vccd1 _1587_/X sky130_fd_sc_hd__or4_2
X_1656_ _1588_/Y _1598_/B _1656_/S vssd1 vssd1 vccd1 vccd1 _1754_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1063__A data_rvalid_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1417__B1 _1779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1510_ _1510_/A _1510_/B vssd1 vssd1 vccd1 vccd1 _1514_/B sky130_fd_sc_hd__or2_2
XFILLER_4_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1441_ _1444_/B vssd1 vssd1 vccd1 vccd1 _1441_/Y sky130_fd_sc_hd__inv_2
X_1372_ _1455_/A vssd1 vssd1 vccd1 vccd1 _1804_/D sky130_fd_sc_hd__inv_2
X_1708_ _1882_/Q _1838_/Q _1714_/S vssd1 vssd1 vccd1 vccd1 _1708_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1639_ _1581_/B _1521_/A _1695_/S vssd1 vssd1 vccd1 vccd1 _1639_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0941_ data_wdata_o[8] _0929_/X _1777_/Q _0930_/X vssd1 vssd1 vccd1 vccd1 _1893_/D
+ sky130_fd_sc_hd__a22o_2
X_0872_ _0910_/C vssd1 vssd1 vccd1 vccd1 _1471_/B sky130_fd_sc_hd__buf_1
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1424_ _1800_/Q _1803_/Q _1280_/X _0871_/A _1419_/A vssd1 vssd1 vccd1 vccd1 _1424_/X
+ sky130_fd_sc_hd__o32a_2
X_1355_ data_addr_o[4] _1342_/X _1781_/Q _1344_/X vssd1 vssd1 vccd1 vccd1 _1809_/D
+ sky130_fd_sc_hd__a22o_2
X_1286_ _1275_/A _1419_/A _1285_/Y _1015_/X _1025_/Y vssd1 vssd1 vccd1 vccd1 _1287_/S
+ sky130_fd_sc_hd__o311a_2
XFILLER_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1140_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1140_/X sky130_fd_sc_hd__buf_1
X_1071_ _1874_/Q _1067_/B _1080_/A _1873_/Q data_gnt_i vssd1 vssd1 vccd1 vccd1 _1072_/B
+ sky130_fd_sc_hd__a32o_2
X_0924_ _0927_/A vssd1 vssd1 vccd1 vccd1 _0925_/A sky130_fd_sc_hd__buf_1
X_1338_ _1338_/A vssd1 vssd1 vccd1 vccd1 _1338_/X sky130_fd_sc_hd__buf_1
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1407_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1407_/X sky130_fd_sc_hd__buf_1
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1269_ _1266_/Y _1258_/C _1413_/A _1268_/X vssd1 vssd1 vccd1 vccd1 _1828_/D sky130_fd_sc_hd__o22ai_2
XFILLER_3_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1054_ _1058_/A vssd1 vssd1 vccd1 vccd1 _1055_/A sky130_fd_sc_hd__buf_1
X_1123_ _1854_/Q _1118_/X data_rdata_i[13] _1120_/X _1115_/X vssd1 vssd1 vccd1 vccd1
+ _1854_/D sky130_fd_sc_hd__o221a_2
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0907_ _0907_/A vssd1 vssd1 vccd1 vccd1 _0907_/X sky130_fd_sc_hd__buf_1
X_1887_ _1888_/CLK _1887_/D _0968_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[2] sky130_fd_sc_hd__dfrtp_2
XFILLER_16_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1741_ _1875_/CLK _1741_/D vssd1 vssd1 vccd1 vccd1 _1741_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1810_ _1892_/CLK _1810_/D _1351_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[5] sky130_fd_sc_hd__dfrtp_2
X_1672_ _1627_/X _1648_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1743_/D sky130_fd_sc_hd__mux2_1
X_1106_ _1862_/Q _1102_/X data_rdata_i[21] _1103_/X _1100_/X vssd1 vssd1 vccd1 vccd1
+ _1862_/D sky130_fd_sc_hd__o221a_2
X_1037_ _1037_/A vssd1 vssd1 vccd1 vccd1 _1037_/X sky130_fd_sc_hd__buf_1
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1132__B1 data_rdata_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1873__CLK _1875_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1724_ _1528_/B _1529_/X _1725_/S vssd1 vssd1 vccd1 vccd1 _1756_/D sky130_fd_sc_hd__mux2_1
X_1655_ _1585_/Y _1576_/A _1656_/S vssd1 vssd1 vccd1 vccd1 _1753_/D sky130_fd_sc_hd__mux2_1
X_1586_ _1605_/A _1664_/X vssd1 vssd1 vccd1 vccd1 _1586_/X sky130_fd_sc_hd__and2_2
XANTENNA__1123__B1 data_rdata_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1114__B1 data_rdata_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1417__A1 _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1371_ rst_i _1371_/B vssd1 vssd1 vccd1 vccd1 _1455_/A sky130_fd_sc_hd__or2_2
XFILLER_4_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1440_ _1746_/Q _1747_/Q vssd1 vssd1 vccd1 vccd1 _1444_/B sky130_fd_sc_hd__or2_2
XANTENNA__1105__B1 data_rdata_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1707_ _1706_/X _1868_/Q _1794_/Q vssd1 vssd1 vccd1 vccd1 _1707_/X sky130_fd_sc_hd__mux2_1
X_1638_ _1581_/B _1579_/X _1695_/S vssd1 vssd1 vccd1 vccd1 _1638_/X sky130_fd_sc_hd__mux2_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _1569_/A vssd1 vssd1 vccd1 vccd1 _1649_/S sky130_fd_sc_hd__inv_2
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clk_i clkbuf_4_9_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1875_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0940_ _0940_/A vssd1 vssd1 vccd1 vccd1 _0940_/X sky130_fd_sc_hd__buf_1
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1574__B1 _1783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0871_ _0871_/A _1017_/A vssd1 vssd1 vccd1 vccd1 _0910_/C sky130_fd_sc_hd__or2_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1423_ _1471_/A _1428_/C _1471_/B vssd1 vssd1 vccd1 vccd1 _1423_/X sky130_fd_sc_hd__o21a_2
X_1285_ _1875_/Q _1873_/Q vssd1 vssd1 vccd1 vccd1 _1285_/Y sky130_fd_sc_hd__nor2_2
X_1354_ _1354_/A vssd1 vssd1 vccd1 vccd1 _1354_/X sky130_fd_sc_hd__buf_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1070_ _1150_/B vssd1 vssd1 vccd1 vccd1 _1076_/A sky130_fd_sc_hd__buf_1
X_0923_ data_wdata_o[13] _0911_/X _1782_/Q _0913_/X vssd1 vssd1 vccd1 vccd1 _1898_/D
+ sky130_fd_sc_hd__a22o_2
X_1337_ _1340_/A vssd1 vssd1 vccd1 vccd1 _1338_/A sky130_fd_sc_hd__buf_1
X_1406_ _1190_/A _1404_/X _1405_/B tx_o _1405_/Y vssd1 vssd1 vccd1 vccd1 _1785_/D
+ sky130_fd_sc_hd__a32o_2
X_1268_ _1266_/Y _1827_/Q _1828_/Q _1578_/B vssd1 vssd1 vccd1 vccd1 _1268_/X sky130_fd_sc_hd__a22o_2
X_1199_ _1836_/Q _1195_/X _1187_/X _1198_/X vssd1 vssd1 vccd1 vccd1 _1836_/D sky130_fd_sc_hd__a22o_2
XFILLER_10_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_6_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1122_ _1855_/Q _1118_/X data_rdata_i[14] _1120_/X _1115_/X vssd1 vssd1 vccd1 vccd1
+ _1855_/D sky130_fd_sc_hd__o221a_2
X_1053_ _1878_/Q _1047_/X _1047_/X _1052_/Y vssd1 vssd1 vccd1 vccd1 _1878_/D sky130_fd_sc_hd__o2bb2ai_2
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0906_ _0906_/A vssd1 vssd1 vccd1 vccd1 _0907_/A sky130_fd_sc_hd__buf_1
X_1886_ _1888_/CLK _1886_/D _0971_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[1] sky130_fd_sc_hd__dfrtp_2
XANTENNA__1082__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1740_ _1835_/CLK _1740_/D vssd1 vssd1 vccd1 vccd1 _1740_/Q sky130_fd_sc_hd__dfxtp_2
X_1671_ _1625_/X _1647_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1742_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1105_ _1863_/Q _1102_/X data_rdata_i[22] _1103_/X _1100_/X vssd1 vssd1 vccd1 vccd1
+ _1863_/D sky130_fd_sc_hd__o221a_2
X_1036_ _1040_/A vssd1 vssd1 vccd1 vccd1 _1037_/A sky130_fd_sc_hd__buf_1
X_1869_ _1904_/CLK _1869_/D vssd1 vssd1 vccd1 vccd1 _1869_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1723_ _1534_/B _1535_/X _1725_/S vssd1 vssd1 vccd1 vccd1 _1757_/D sky130_fd_sc_hd__mux2_1
X_1654_ _1583_/Y _1681_/S _1656_/S vssd1 vssd1 vccd1 vccd1 _1752_/D sky130_fd_sc_hd__mux2_1
X_1585_ _1694_/X _1584_/X _1693_/X _1581_/X _1592_/A vssd1 vssd1 vccd1 vccd1 _1585_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_41_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0882__B1 _1783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1019_ _1800_/Q _1016_/Y _1469_/A _1570_/A vssd1 vssd1 vccd1 vccd1 _1019_/Y sky130_fd_sc_hd__a22oi_2
Xclkbuf_4_5_0_clk_i clkbuf_4_5_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1830_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1370_ data_addr_o[0] _1358_/X _1777_/Q _1359_/X vssd1 vssd1 vccd1 vccd1 _1805_/D
+ sky130_fd_sc_hd__a22o_2
X_1637_ _1636_/X _1865_/Q _1794_/Q vssd1 vssd1 vccd1 vccd1 _1637_/X sky130_fd_sc_hd__mux2_1
X_1706_ _1705_/X _1860_/Q _1798_/Q vssd1 vssd1 vccd1 vccd1 _1706_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1499_/A vssd1 vssd1 vccd1 vccd1 _1499_/X sky130_fd_sc_hd__buf_1
X_1568_ _1837_/Q _1568_/B vssd1 vssd1 vccd1 vccd1 _1568_/Y sky130_fd_sc_hd__nor2_2
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1099__B1 data_rdata_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0870_ _1752_/Q _1226_/B _1002_/A vssd1 vssd1 vccd1 vccd1 _1017_/A sky130_fd_sc_hd__or3_2
X_1422_ _1422_/A vssd1 vssd1 vccd1 vccd1 _1471_/A sky130_fd_sc_hd__buf_1
X_1284_ _1284_/A vssd1 vssd1 vccd1 vccd1 _1284_/X sky130_fd_sc_hd__buf_1
X_1353_ _1356_/A vssd1 vssd1 vccd1 vccd1 _1354_/A sky130_fd_sc_hd__buf_1
Xclkbuf_0_clk_i clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_0999_ _1040_/A vssd1 vssd1 vccd1 vccd1 _1000_/A sky130_fd_sc_hd__buf_1
XFILLER_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_2_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0922_ _0922_/A vssd1 vssd1 vccd1 vccd1 _0922_/X sky130_fd_sc_hd__buf_1
X_1405_ _1613_/B _1405_/B vssd1 vssd1 vccd1 vccd1 _1405_/Y sky130_fd_sc_hd__nand2_2
X_1336_ data_wdata_o[25] _1327_/X _1778_/Q _1328_/X vssd1 vssd1 vccd1 vccd1 _1814_/D
+ sky130_fd_sc_hd__a22o_2
X_1198_ _1208_/B _1404_/B _1198_/C vssd1 vssd1 vccd1 vccd1 _1198_/X sky130_fd_sc_hd__or3_2
X_1267_ _1827_/Q vssd1 vssd1 vccd1 vccd1 _1578_/B sky130_fd_sc_hd__inv_2
XFILLER_10_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1052_ _1800_/Q _1680_/X _1779_/Q _1570_/A vssd1 vssd1 vccd1 vccd1 _1052_/Y sky130_fd_sc_hd__a22oi_2
X_1121_ _1856_/Q _1118_/X data_rdata_i[15] _1120_/X _1115_/X vssd1 vssd1 vccd1 vccd1
+ _1856_/D sky130_fd_sc_hd__o221a_2
X_0905_ data_wdata_o[16] _0893_/X _1777_/Q _0894_/X vssd1 vssd1 vccd1 vccd1 _1901_/D
+ sky130_fd_sc_hd__a22o_2
X_1885_ _1888_/CLK _1885_/D _0974_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[0] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1319_ _1325_/A vssd1 vssd1 vccd1 vccd1 _1320_/A sky130_fd_sc_hd__buf_1
XFILLER_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1670_ _1623_/X _1651_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1741_/D sky130_fd_sc_hd__mux2_1
X_1035_ _1035_/A vssd1 vssd1 vccd1 vccd1 _1882_/D sky130_fd_sc_hd__buf_1
X_1104_ _1864_/Q _1102_/X data_rdata_i[23] _1103_/X _1100_/X vssd1 vssd1 vccd1 vccd1
+ _1864_/D sky130_fd_sc_hd__o221a_2
XFILLER_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1868_ _1904_/CLK _1868_/D vssd1 vssd1 vccd1 vccd1 _1868_/Q sky130_fd_sc_hd__dfxtp_2
X_1799_ _1883_/CLK _1799_/D _1383_/X vssd1 vssd1 vccd1 vccd1 _1799_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_1_0_clk_i clkbuf_4_1_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1888_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1653_ _1404_/B _1651_/X _1674_/S vssd1 vssd1 vccd1 vccd1 _1653_/X sky130_fd_sc_hd__mux2_1
X_1722_ _1538_/B _1539_/X _1725_/S vssd1 vssd1 vccd1 vccd1 _1758_/D sky130_fd_sc_hd__mux2_1
X_1584_ _1584_/A vssd1 vssd1 vccd1 vccd1 _1584_/X sky130_fd_sc_hd__buf_1
XANTENNA__0882__A1 data_wdata_o[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1018_ _1018_/A vssd1 vssd1 vccd1 vccd1 _1570_/A sky130_fd_sc_hd__buf_1
XFILLER_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1705_ _1844_/Q _1852_/Q _1796_/Q vssd1 vssd1 vccd1 vccd1 _1705_/X sky130_fd_sc_hd__mux2_1
X_1636_ _1635_/X _1857_/Q _1798_/Q vssd1 vssd1 vccd1 vccd1 _1636_/X sky130_fd_sc_hd__mux2_1
X_1567_ _1567_/A vssd1 vssd1 vccd1 vccd1 _1567_/X sky130_fd_sc_hd__buf_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ rx_i _1498_/B vssd1 vssd1 vccd1 vccd1 _1499_/A sky130_fd_sc_hd__and2_2
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1421_ _1801_/Q _1278_/X _1420_/X _1294_/X vssd1 vssd1 vccd1 vccd1 _1801_/D sky130_fd_sc_hd__a31o_2
X_1283_ _1289_/A vssd1 vssd1 vccd1 vccd1 _1284_/A sky130_fd_sc_hd__buf_1
X_1352_ data_addr_o[5] _1342_/X _1782_/Q _1344_/X vssd1 vssd1 vccd1 vccd1 _1810_/D
+ sky130_fd_sc_hd__a22o_2
X_0998_ _1296_/A vssd1 vssd1 vccd1 vccd1 _1040_/A sky130_fd_sc_hd__buf_1
X_1619_ _1616_/X _1645_/X vssd1 vssd1 vccd1 vccd1 _1620_/A sky130_fd_sc_hd__and2b_2
XFILLER_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0921_ _0927_/A vssd1 vssd1 vccd1 vccd1 _0922_/A sky130_fd_sc_hd__buf_1
X_1335_ _1335_/A vssd1 vssd1 vccd1 vccd1 _1335_/X sky130_fd_sc_hd__buf_1
X_1404_ _1786_/Q _1404_/B vssd1 vssd1 vccd1 vccd1 _1404_/X sky130_fd_sc_hd__or2_2
X_1197_ _1835_/Q _1201_/A _1836_/Q vssd1 vssd1 vccd1 vccd1 _1198_/C sky130_fd_sc_hd__o21a_2
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1266_ _1828_/Q vssd1 vssd1 vccd1 vccd1 _1266_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1051_ _1051_/A vssd1 vssd1 vccd1 vccd1 _1051_/X sky130_fd_sc_hd__buf_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1120_ _1141_/A vssd1 vssd1 vccd1 vccd1 _1120_/X sky130_fd_sc_hd__buf_1
X_0904_ _0904_/A vssd1 vssd1 vccd1 vccd1 _0904_/X sky130_fd_sc_hd__buf_1
X_1884_ _1892_/CLK _1884_/D _0977_/X vssd1 vssd1 vccd1 vccd1 _1884_/Q sky130_fd_sc_hd__dfrtp_2
X_1318_ data_wdata_o[30] _1310_/X _1783_/Q _1312_/X vssd1 vssd1 vccd1 vccd1 _1819_/D
+ sky130_fd_sc_hd__a22o_2
X_1249_ _1249_/A _1249_/B vssd1 vssd1 vccd1 vccd1 _1692_/S sky130_fd_sc_hd__nor2_2
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1144__B1 data_rdata_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1135__B1 data_rdata_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1034_ _1643_/X _1882_/Q _1047_/A vssd1 vssd1 vccd1 vccd1 _1035_/A sky130_fd_sc_hd__mux2_2
X_1103_ _1111_/A vssd1 vssd1 vccd1 vccd1 _1103_/X sky130_fd_sc_hd__buf_1
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1867_ _1904_/CLK _1867_/D vssd1 vssd1 vccd1 vccd1 _1867_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1798_ _1859_/CLK _1798_/D _1386_/X vssd1 vssd1 vccd1 vccd1 _1798_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1721_ _1543_/B _1544_/X _1725_/S vssd1 vssd1 vccd1 vccd1 _1759_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1583_ _1638_/X _1592_/A _1639_/X _1584_/A _1582_/X vssd1 vssd1 vccd1 vccd1 _1583_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1652_ _1740_/Q _1459_/X _1652_/S vssd1 vssd1 vccd1 vccd1 _1652_/X sky130_fd_sc_hd__mux2_1
X_1017_ _1017_/A vssd1 vssd1 vccd1 vccd1 _1469_/A sky130_fd_sc_hd__buf_1
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1704_ _1703_/X _1869_/Q _1794_/Q vssd1 vssd1 vccd1 vccd1 _1704_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1329__B1 _1780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _1497_/A vssd1 vssd1 vccd1 vccd1 _1498_/B sky130_fd_sc_hd__buf_1
X_1566_ _1566_/A _1566_/B vssd1 vssd1 vccd1 vccd1 _1567_/A sky130_fd_sc_hd__and2_2
X_1635_ _1841_/Q _1849_/Q _1796_/Q vssd1 vssd1 vccd1 vccd1 _1635_/X sky130_fd_sc_hd__mux2_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1420_ _1873_/Q _1420_/B _1420_/C vssd1 vssd1 vccd1 vccd1 _1420_/X sky130_fd_sc_hd__or3_2
X_1351_ _1351_/A vssd1 vssd1 vccd1 vccd1 _1351_/X sky130_fd_sc_hd__buf_1
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1282_ _1884_/Q _1358_/A _1065_/B _1281_/X vssd1 vssd1 vccd1 vccd1 _1826_/D sky130_fd_sc_hd__o22ai_2
X_0997_ _1314_/A vssd1 vssd1 vccd1 vccd1 _1296_/A sky130_fd_sc_hd__buf_1
X_1618_ _1618_/A vssd1 vssd1 vccd1 vccd1 _1618_/X sky130_fd_sc_hd__buf_1
XFILLER_5_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1549_ _1566_/A _1549_/B vssd1 vssd1 vccd1 vccd1 _1550_/A sky130_fd_sc_hd__and2_2
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_3_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0920_ data_wdata_o[14] _0911_/X _1783_/Q _0913_/X vssd1 vssd1 vccd1 vccd1 _1899_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1334_ _1340_/A vssd1 vssd1 vccd1 vccd1 _1335_/A sky130_fd_sc_hd__buf_1
X_1403_ _1786_/Q _1186_/A _1714_/X _1203_/X vssd1 vssd1 vccd1 vccd1 _1786_/D sky130_fd_sc_hd__a22o_2
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1265_ _1258_/A _1258_/C _1413_/A _1264_/X vssd1 vssd1 vccd1 vccd1 _1829_/D sky130_fd_sc_hd__o22ai_2
XFILLER_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1196_ _1196_/A vssd1 vssd1 vccd1 vccd1 _1404_/B sky130_fd_sc_hd__inv_2
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1050_ _1058_/A vssd1 vssd1 vccd1 vccd1 _1051_/A sky130_fd_sc_hd__buf_1
XFILLER_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1883_ _1883_/CLK _1883_/D _1000_/X vssd1 vssd1 vccd1 vccd1 _1883_/Q sky130_fd_sc_hd__dfrtp_2
X_0903_ _0906_/A vssd1 vssd1 vccd1 vccd1 _0904_/A sky130_fd_sc_hd__buf_1
XFILLER_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1317_ _1317_/A vssd1 vssd1 vccd1 vccd1 _1317_/X sky130_fd_sc_hd__buf_1
X_1248_ _1774_/Q _1775_/Q _1510_/B _1248_/D vssd1 vssd1 vccd1 vccd1 _1249_/B sky130_fd_sc_hd__or4_2
XANTENNA__1153__A1 data_req_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1179_ _1645_/X _1651_/X _1179_/C _1617_/B vssd1 vssd1 vccd1 vccd1 _1180_/A sky130_fd_sc_hd__or4_2
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1102_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1102_/X sky130_fd_sc_hd__buf_1
X_1033_ _1033_/A vssd1 vssd1 vccd1 vccd1 _1033_/X sky130_fd_sc_hd__buf_1
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1866_ _1904_/CLK _1866_/D vssd1 vssd1 vccd1 vccd1 _1866_/Q sky130_fd_sc_hd__dfxtp_2
X_1797_ _1859_/CLK _1797_/D _1388_/X vssd1 vssd1 vccd1 vccd1 _1797_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1720_ _1549_/B _1550_/X _1725_/S vssd1 vssd1 vccd1 vccd1 _1760_/D sky130_fd_sc_hd__mux2_1
X_1651_ _1741_/Q _1461_/X _1652_/S vssd1 vssd1 vccd1 vccd1 _1651_/X sky130_fd_sc_hd__mux2_1
X_1582_ _1687_/X _1581_/X rx_i _1591_/B vssd1 vssd1 vccd1 vccd1 _1582_/X sky130_fd_sc_hd__o22a_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1016_ _1794_/Q _1016_/B vssd1 vssd1 vccd1 vccd1 _1016_/Y sky130_fd_sc_hd__nor2_2
X_1849_ _1852_/CLK _1849_/D vssd1 vssd1 vccd1 vccd1 _1849_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1703_ _1702_/X _1861_/Q _1798_/Q vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__mux2_1
X_1634_ tx_o vssd1 vssd1 vccd1 vccd1 _1634_/X sky130_fd_sc_hd__buf_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _1770_/Q _1510_/A _1500_/B vssd1 vssd1 vccd1 vccd1 _1497_/A sky130_fd_sc_hd__a21bo_2
X_1565_ _1564_/Y _1560_/Y _1171_/X vssd1 vssd1 vccd1 vccd1 _1566_/B sky130_fd_sc_hd__o21ai_2
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1281_ _1275_/X _1279_/X _1280_/X vssd1 vssd1 vccd1 vccd1 _1281_/X sky130_fd_sc_hd__o21a_2
XFILLER_0_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1350_ _1356_/A vssd1 vssd1 vccd1 vccd1 _1351_/A sky130_fd_sc_hd__buf_1
XFILLER_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0996_ _0980_/X _0993_/Y _1022_/A _1884_/Q _0995_/X vssd1 vssd1 vccd1 vccd1 _1884_/D
+ sky130_fd_sc_hd__a32o_2
X_1617_ _1616_/X _1617_/B vssd1 vssd1 vccd1 vccd1 _1618_/A sky130_fd_sc_hd__and2b_2
X_1479_ _1767_/Q vssd1 vssd1 vccd1 vccd1 _1479_/Y sky130_fd_sc_hd__inv_2
X_1548_ _1548_/A vssd1 vssd1 vccd1 vccd1 _1566_/A sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_3_7_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1410__B1 _1784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1402_ _1713_/X _1195_/X _1787_/Q _1203_/X vssd1 vssd1 vccd1 vccd1 _1787_/D sky130_fd_sc_hd__o22a_2
X_1333_ data_wdata_o[26] _1327_/X _1779_/Q _1328_/X vssd1 vssd1 vccd1 vccd1 _1815_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1264_ _1829_/Q _1219_/A _1258_/A _1258_/B vssd1 vssd1 vccd1 vccd1 _1264_/X sky130_fd_sc_hd__o22a_2
XFILLER_51_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1195_ _1195_/A vssd1 vssd1 vccd1 vccd1 _1195_/X sky130_fd_sc_hd__buf_1
X_0979_ _1021_/A vssd1 vssd1 vccd1 vccd1 _1371_/B sky130_fd_sc_hd__inv_2
XFILLER_35_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1882_ _1883_/CLK _1882_/D _1033_/X vssd1 vssd1 vccd1 vccd1 _1882_/Q sky130_fd_sc_hd__dfrtp_2
X_0902_ data_wdata_o[17] _0893_/X _1778_/Q _0894_/X vssd1 vssd1 vccd1 vccd1 _1902_/D
+ sky130_fd_sc_hd__a22o_2
XANTENNA__1622__B1 _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1316_ _1325_/A vssd1 vssd1 vccd1 vccd1 _1317_/A sky130_fd_sc_hd__buf_1
X_1247_ _1768_/Q _1769_/Q _1247_/C _1767_/Q vssd1 vssd1 vccd1 vccd1 _1248_/D sky130_fd_sc_hd__or4_2
XFILLER_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1178_ _1166_/Y _1652_/S _1166_/Y _1652_/S vssd1 vssd1 vccd1 vccd1 _1617_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1032_ _1040_/A vssd1 vssd1 vccd1 vccd1 _1033_/A sky130_fd_sc_hd__buf_1
X_1101_ _1865_/Q _1095_/X data_rdata_i[24] _1096_/X _1100_/X vssd1 vssd1 vccd1 vccd1
+ _1865_/D sky130_fd_sc_hd__o221a_2
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1865_ _1908_/CLK _1865_/D vssd1 vssd1 vccd1 vccd1 _1865_/Q sky130_fd_sc_hd__dfxtp_2
X_1796_ _1859_/CLK _1796_/D _1390_/X vssd1 vssd1 vccd1 vccd1 _1796_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1071__B2 data_gnt_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1650_ _1611_/X _1688_/X _1683_/S vssd1 vssd1 vccd1 vccd1 _1650_/X sky130_fd_sc_hd__mux2_1
X_1581_ _1581_/A _1581_/B _1754_/Q vssd1 vssd1 vccd1 vccd1 _1581_/X sky130_fd_sc_hd__or3_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1015_ _1799_/Q _1569_/A _1884_/Q _1343_/A _1014_/X vssd1 vssd1 vccd1 vccd1 _1015_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1779_ _1895_/CLK _1779_/D vssd1 vssd1 vccd1 vccd1 _1779_/Q sky130_fd_sc_hd__dfxtp_2
X_1848_ _1852_/CLK _1848_/D vssd1 vssd1 vccd1 vccd1 _1848_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1633_ vssd1 vssd1 vccd1 vccd1 data_be_o[3] _1633_/LO sky130_fd_sc_hd__conb_1
X_1564_ _1764_/Q vssd1 vssd1 vccd1 vccd1 _1564_/Y sky130_fd_sc_hd__inv_2
X_1702_ _1845_/Q _1853_/Q _1796_/Q vssd1 vssd1 vccd1 vccd1 _1702_/X sky130_fd_sc_hd__mux2_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1770_/Q _1510_/A vssd1 vssd1 vccd1 vccd1 _1500_/B sky130_fd_sc_hd__or2_2
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1280_ _1801_/Q _1799_/Q vssd1 vssd1 vccd1 vccd1 _1280_/X sky130_fd_sc_hd__or2_2
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0995_ _1021_/A _0995_/B vssd1 vssd1 vccd1 vccd1 _0995_/X sky130_fd_sc_hd__or2_2
X_1547_ _1547_/A vssd1 vssd1 vccd1 vccd1 _1549_/B sky130_fd_sc_hd__buf_1
X_1616_ _1837_/Q _1804_/D _1164_/A vssd1 vssd1 vccd1 vccd1 _1616_/X sky130_fd_sc_hd__o21a_2
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1478_ _1591_/B vssd1 vssd1 vccd1 vccd1 _1736_/S sky130_fd_sc_hd__inv_2
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1410__A1 _1783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1401_ _1712_/X _1195_/X _1788_/Q _1397_/X vssd1 vssd1 vccd1 vccd1 _1788_/D sky130_fd_sc_hd__o22a_2
X_1332_ _1332_/A vssd1 vssd1 vccd1 vccd1 _1332_/X sky130_fd_sc_hd__buf_1
X_1263_ _1270_/A vssd1 vssd1 vccd1 vccd1 _1413_/A sky130_fd_sc_hd__buf_1
X_1194_ _1837_/Q _1825_/Q _1145_/X _1193_/X vssd1 vssd1 vccd1 vccd1 _1837_/D sky130_fd_sc_hd__o211a_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1004__A data_req_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0978_ _1745_/Q _1744_/Q vssd1 vssd1 vccd1 vccd1 _1021_/A sky130_fd_sc_hd__or2_2
XFILLER_10_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1881_ _1881_/CLK _1881_/D _1037_/X vssd1 vssd1 vccd1 vccd1 _1881_/Q sky130_fd_sc_hd__dfrtp_2
X_0901_ _0901_/A vssd1 vssd1 vccd1 vccd1 _0901_/X sky130_fd_sc_hd__buf_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1315_ _1361_/A vssd1 vssd1 vccd1 vccd1 _1325_/A sky130_fd_sc_hd__buf_1
X_1246_ _1766_/Q vssd1 vssd1 vccd1 vccd1 _1247_/C sky130_fd_sc_hd__inv_2
X_1177_ _1177_/A _1177_/B vssd1 vssd1 vccd1 vccd1 _1652_/S sky130_fd_sc_hd__nor2_2
XFILLER_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1129__B1 data_rdata_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1031_ _1883_/Q _1028_/X _1028_/X _1030_/Y vssd1 vssd1 vccd1 vccd1 _1883_/D sky130_fd_sc_hd__o2bb2ai_2
X_1100_ _1628_/A vssd1 vssd1 vccd1 vccd1 _1100_/X sky130_fd_sc_hd__buf_1
XFILLER_38_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1864_ _1904_/CLK _1864_/D vssd1 vssd1 vccd1 vccd1 _1864_/Q sky130_fd_sc_hd__dfxtp_2
X_1795_ _1859_/CLK _1795_/D _1392_/X vssd1 vssd1 vccd1 vccd1 _1795_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1229_ _1261_/A vssd1 vssd1 vccd1 vccd1 _1229_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1580_ _1580_/A vssd1 vssd1 vccd1 vccd1 _1584_/A sky130_fd_sc_hd__buf_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1014_ _1422_/A _1428_/C _1428_/B vssd1 vssd1 vccd1 vccd1 _1014_/X sky130_fd_sc_hd__or3_2
XFILLER_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1847_ _1895_/CLK _1847_/D vssd1 vssd1 vccd1 vccd1 _1847_/Q sky130_fd_sc_hd__dfxtp_2
X_1778_ _1895_/CLK _1778_/D vssd1 vssd1 vccd1 vccd1 _1778_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_40_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1701_ _1700_/X _1866_/Q _1794_/Q vssd1 vssd1 vccd1 vccd1 _1701_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1632_ vssd1 vssd1 vccd1 vccd1 data_be_o[2] _1632_/LO sky130_fd_sc_hd__conb_1
X_1494_ _1494_/A vssd1 vssd1 vccd1 vccd1 _1494_/X sky130_fd_sc_hd__buf_1
X_1563_ _1837_/Q _1563_/B vssd1 vssd1 vccd1 vccd1 _1563_/Y sky130_fd_sc_hd__nor2_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1800__CLK _1875_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0994_ _1468_/A vssd1 vssd1 vccd1 vccd1 _1022_/A sky130_fd_sc_hd__inv_2
X_1615_ _1613_/A _1672_/S _1674_/S _1674_/X _1714_/S vssd1 vssd1 vccd1 vccd1 _1615_/X
+ sky130_fd_sc_hd__a32o_2
X_1546_ _1760_/Q _1551_/C _1545_/X vssd1 vssd1 vccd1 vccd1 _1547_/A sky130_fd_sc_hd__a21bo_2
X_1477_ _1681_/S _1598_/B _1576_/A vssd1 vssd1 vccd1 vccd1 _1591_/B sky130_fd_sc_hd__or3_2
XFILLER_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1400_ _1711_/X _1195_/X _1789_/Q _1397_/X vssd1 vssd1 vccd1 vccd1 _1789_/D sky130_fd_sc_hd__o22a_2
X_1331_ _1340_/A vssd1 vssd1 vccd1 vccd1 _1332_/A sky130_fd_sc_hd__buf_1
XFILLER_36_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1262_ _1592_/A _1683_/S vssd1 vssd1 vccd1 vccd1 _1270_/A sky130_fd_sc_hd__or2_2
X_1193_ _1548_/A _1395_/B _1793_/Q vssd1 vssd1 vccd1 vccd1 _1193_/X sky130_fd_sc_hd__or3_2
XANTENNA__1020__A _1784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0977_ _0977_/A vssd1 vssd1 vccd1 vccd1 _0977_/X sky130_fd_sc_hd__buf_1
X_1529_ _1529_/A vssd1 vssd1 vccd1 vccd1 _1529_/X sky130_fd_sc_hd__buf_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1880_ _1883_/CLK _1880_/D _1041_/X vssd1 vssd1 vccd1 vccd1 _1880_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0900_ _0906_/A vssd1 vssd1 vccd1 vccd1 _0901_/A sky130_fd_sc_hd__buf_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1314_ _1314_/A vssd1 vssd1 vccd1 vccd1 _1361_/A sky130_fd_sc_hd__buf_1
XFILLER_2_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1245_ _1522_/B vssd1 vssd1 vccd1 vccd1 _1249_/A sky130_fd_sc_hd__inv_2
X_1176_ _1176_/A _1756_/Q _1176_/C _1176_/D vssd1 vssd1 vccd1 vccd1 _1177_/B sky130_fd_sc_hd__or4_2
XFILLER_15_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1030_ _1800_/Q _1686_/X _1784_/Q _1029_/X vssd1 vssd1 vccd1 vccd1 _1030_/Y sky130_fd_sc_hd__a22oi_2
X_1863_ _1908_/CLK _1863_/D vssd1 vssd1 vccd1 vccd1 _1863_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1794_ _1904_/CLK _1794_/D _1394_/X vssd1 vssd1 vccd1 vccd1 _1794_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1228_ _1439_/A _1598_/B _1581_/A vssd1 vssd1 vccd1 vccd1 _1261_/A sky130_fd_sc_hd__or3_2
X_1159_ _1883_/Q _1208_/B vssd1 vssd1 vccd1 vccd1 _1159_/X sky130_fd_sc_hd__and2_2
XANTENNA__1295__B1 _1780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1013_ _1796_/Q _1797_/Q _1013_/C vssd1 vssd1 vccd1 vccd1 _1428_/B sky130_fd_sc_hd__or3_2
X_1777_ _1895_/CLK _1777_/D vssd1 vssd1 vccd1 vccd1 _1777_/Q sky130_fd_sc_hd__dfxtp_2
X_1846_ _1895_/CLK _1846_/D vssd1 vssd1 vccd1 vccd1 _1846_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1631_ vssd1 vssd1 vccd1 vccd1 data_be_o[1] _1631_/LO sky130_fd_sc_hd__conb_1
X_1700_ _1699_/X _1858_/Q _1798_/Q vssd1 vssd1 vccd1 vccd1 _1700_/X sky130_fd_sc_hd__mux2_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ rx_i _1493_/B vssd1 vssd1 vccd1 vccd1 _1494_/A sky130_fd_sc_hd__and2_2
X_1562_ _1563_/B vssd1 vssd1 vccd1 vccd1 _1562_/Y sky130_fd_sc_hd__inv_2
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1722__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1829_ _1830_/CLK _1829_/D vssd1 vssd1 vccd1 vccd1 _1829_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0993_ _0995_/B vssd1 vssd1 vccd1 vccd1 _0993_/Y sky130_fd_sc_hd__inv_2
X_1614_ _1644_/X _1714_/S _1837_/Q _1725_/S vssd1 vssd1 vccd1 vccd1 _1614_/X sky130_fd_sc_hd__a22o_2
XANTENNA__1717__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_14_0_clk_i clkbuf_3_7_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1904_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1545_ _1760_/Q _1551_/C vssd1 vssd1 vccd1 vccd1 _1545_/X sky130_fd_sc_hd__or2_2
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1476_ _1521_/A _1766_/Q vssd1 vssd1 vccd1 vccd1 _1476_/Y sky130_fd_sc_hd__nor2_2
XFILLER_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1330_ _1361_/A vssd1 vssd1 vccd1 vccd1 _1340_/A sky130_fd_sc_hd__buf_1
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1261_ _1261_/A vssd1 vssd1 vccd1 vccd1 _1592_/A sky130_fd_sc_hd__buf_1
X_1192_ _1804_/Q vssd1 vssd1 vccd1 vccd1 _1395_/B sky130_fd_sc_hd__inv_2
X_0976_ _0976_/A vssd1 vssd1 vccd1 vccd1 _0977_/A sky130_fd_sc_hd__buf_1
X_1528_ _1837_/Q _1528_/B vssd1 vssd1 vccd1 vccd1 _1529_/A sky130_fd_sc_hd__or2_2
XFILLER_19_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1459_ _1740_/Q _1458_/B _1460_/B vssd1 vssd1 vccd1 vccd1 _1459_/X sky130_fd_sc_hd__a21bo_2
XFILLER_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1313_ data_wdata_o[31] _1310_/X _1784_/Q _1312_/X vssd1 vssd1 vccd1 vccd1 _1820_/D
+ sky130_fd_sc_hd__a22o_2
X_1244_ _1776_/Q _1243_/Y _1776_/Q _1243_/Y vssd1 vssd1 vccd1 vccd1 _1522_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1175_ _1763_/Q _1764_/Q _1757_/Q _1758_/Q vssd1 vssd1 vccd1 vccd1 _1176_/C sky130_fd_sc_hd__or4_2
X_0959_ _0959_/A vssd1 vssd1 vccd1 vccd1 _0959_/X sky130_fd_sc_hd__buf_1
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1862_ _1908_/CLK _1862_/D vssd1 vssd1 vccd1 vccd1 _1862_/Q sky130_fd_sc_hd__dfxtp_2
X_1793_ _1840_/CLK _1793_/D vssd1 vssd1 vccd1 vccd1 _1793_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1725__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1158_ _1164_/A vssd1 vssd1 vccd1 vccd1 _1208_/B sky130_fd_sc_hd__buf_1
X_1227_ _1227_/A vssd1 vssd1 vccd1 vccd1 _1581_/A sky130_fd_sc_hd__buf_1
X_1089_ _1872_/Q _1086_/X data_rdata_i[31] _1088_/X _0881_/X vssd1 vssd1 vccd1 vccd1
+ _1872_/D sky130_fd_sc_hd__o221a_2
XFILLER_12_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1012_ _1800_/Q vssd1 vssd1 vccd1 vccd1 _1422_/A sky130_fd_sc_hd__inv_2
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1776_ _1851_/CLK _1776_/D vssd1 vssd1 vccd1 vccd1 _1776_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1845_ _1852_/CLK _1845_/D vssd1 vssd1 vccd1 vccd1 _1845_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__0960__B1 _1781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1630_ vssd1 vssd1 vccd1 vccd1 data_be_o[0] _1630_/LO sky130_fd_sc_hd__conb_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1492_/A vssd1 vssd1 vccd1 vccd1 _1493_/B sky130_fd_sc_hd__buf_1
X_1561_ _1763_/Q _1560_/B _1560_/Y vssd1 vssd1 vccd1 vccd1 _1563_/B sky130_fd_sc_hd__a21oi_2
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_10_0_clk_i clkbuf_3_5_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1881_/CLK sky130_fd_sc_hd__clkbuf_2
X_1759_ _1771_/CLK _1759_/D vssd1 vssd1 vccd1 vccd1 _1759_/Q sky130_fd_sc_hd__dfxtp_2
X_1828_ _1895_/CLK _1828_/D vssd1 vssd1 vccd1 vccd1 _1828_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1101__B1 data_rdata_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0992_ _1468_/A _0980_/X _1023_/C _0991_/X vssd1 vssd1 vccd1 vccd1 _0995_/B sky130_fd_sc_hd__a31o_2
X_1613_ _1613_/A _1613_/B vssd1 vssd1 vccd1 vccd1 _1666_/S sky130_fd_sc_hd__nor2_2
X_1544_ _1544_/A vssd1 vssd1 vccd1 vccd1 _1544_/X sky130_fd_sc_hd__buf_1
X_1475_ _1595_/A vssd1 vssd1 vccd1 vccd1 _1521_/A sky130_fd_sc_hd__buf_1
XANTENNA__1643__A1 _1006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1020__C_N _1782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1260_ _1216_/Y _1258_/X _1257_/A _1259_/X vssd1 vssd1 vccd1 vccd1 _1830_/D sky130_fd_sc_hd__o22ai_2
X_1191_ _1837_/Q vssd1 vssd1 vccd1 vccd1 _1548_/A sky130_fd_sc_hd__inv_2
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0975_ data_wdata_o[0] _0963_/X _1777_/Q _0964_/X vssd1 vssd1 vccd1 vccd1 _1885_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1527_ _1527_/A vssd1 vssd1 vccd1 vccd1 _1528_/B sky130_fd_sc_hd__buf_1
XANTENNA__1313__B1 _1784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1389_ _1391_/A vssd1 vssd1 vccd1 vccd1 _1390_/A sky130_fd_sc_hd__buf_1
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1458_ _1740_/Q _1458_/B vssd1 vssd1 vccd1 vccd1 _1460_/B sky130_fd_sc_hd__or2_2
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1312_ _1328_/A vssd1 vssd1 vccd1 vccd1 _1312_/X sky130_fd_sc_hd__buf_1
X_1243_ _1774_/Q _1775_/Q _1510_/B _1490_/A vssd1 vssd1 vccd1 vccd1 _1243_/Y sky130_fd_sc_hd__nor4_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1174_ _1755_/Q vssd1 vssd1 vccd1 vccd1 _1176_/A sky130_fd_sc_hd__inv_2
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0889_ _0889_/A vssd1 vssd1 vccd1 vccd1 _0889_/X sky130_fd_sc_hd__buf_1
X_0958_ _0961_/A vssd1 vssd1 vccd1 vccd1 _0959_/A sky130_fd_sc_hd__buf_1
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1792_ _1881_/CLK _1792_/D vssd1 vssd1 vccd1 vccd1 _1792_/Q sky130_fd_sc_hd__dfxtp_2
X_1861_ _1904_/CLK _1861_/D vssd1 vssd1 vccd1 vccd1 _1861_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1157_ _1160_/A _1672_/S vssd1 vssd1 vccd1 vccd1 _1164_/A sky130_fd_sc_hd__or2_2
X_1226_ rst_i _1226_/B vssd1 vssd1 vccd1 vccd1 _1227_/A sky130_fd_sc_hd__or2_2
XFILLER_16_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1088_ _1111_/A vssd1 vssd1 vccd1 vccd1 _1088_/X sky130_fd_sc_hd__buf_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1011_ _1275_/A _1017_/A vssd1 vssd1 vccd1 vccd1 _1343_/A sky130_fd_sc_hd__or2_2
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1775_ _1888_/CLK _1775_/D vssd1 vssd1 vccd1 vccd1 _1775_/Q sky130_fd_sc_hd__dfxtp_2
X_1844_ _1852_/CLK _1844_/D vssd1 vssd1 vccd1 vccd1 _1844_/Q sky130_fd_sc_hd__dfxtp_2
X_1209_ _1186_/A _1208_/Y _1833_/Q _1187_/X vssd1 vssd1 vccd1 vccd1 _1833_/D sky130_fd_sc_hd__o22a_2
XANTENNA__1826__CLK _1875_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1560_ _1763_/Q _1560_/B vssd1 vssd1 vccd1 vccd1 _1560_/Y sky130_fd_sc_hd__nor2_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ _1769_/Q _1242_/B _1510_/A vssd1 vssd1 vccd1 vccd1 _1492_/A sky130_fd_sc_hd__a21bo_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1827_ _1852_/CLK _1827_/D vssd1 vssd1 vccd1 vccd1 _1827_/Q sky130_fd_sc_hd__dfxtp_2
X_1758_ _1771_/CLK _1758_/D vssd1 vssd1 vccd1 vccd1 _1758_/Q sky130_fd_sc_hd__dfxtp_2
X_1689_ _1747_/Q _1442_/X _1692_/S vssd1 vssd1 vccd1 vccd1 _1689_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0991_ _0991_/A uart_error _1468_/B vssd1 vssd1 vccd1 vccd1 _0991_/X sky130_fd_sc_hd__or3_2
XFILLER_12_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1543_ _1543_/A _1543_/B vssd1 vssd1 vccd1 vccd1 _1544_/A sky130_fd_sc_hd__and2_2
X_1474_ rx_i vssd1 vssd1 vccd1 vccd1 _1595_/A sky130_fd_sc_hd__inv_2
X_1612_ _1650_/X _1584_/X _1688_/X _1592_/X vssd1 vssd1 vccd1 vccd1 _1612_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__1315__A _1361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk_i clkbuf_4_9_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1835_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1190_ _1190_/A vssd1 vssd1 vccd1 vccd1 _1714_/S sky130_fd_sc_hd__buf_1
X_0974_ _0974_/A vssd1 vssd1 vccd1 vccd1 _0974_/X sky130_fd_sc_hd__buf_1
X_1526_ _1652_/S _1526_/B vssd1 vssd1 vccd1 vccd1 _1527_/A sky130_fd_sc_hd__or2_2
X_1457_ _1738_/Q _1739_/Q _1458_/B vssd1 vssd1 vccd1 vccd1 _1457_/X sky130_fd_sc_hd__a21bo_2
X_1388_ _1388_/A vssd1 vssd1 vccd1 vccd1 _1388_/X sky130_fd_sc_hd__buf_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1311_ _1327_/A vssd1 vssd1 vccd1 vccd1 _1328_/A sky130_fd_sc_hd__inv_2
X_1242_ _1769_/Q _1242_/B vssd1 vssd1 vccd1 vccd1 _1490_/A sky130_fd_sc_hd__or2_2
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1173_ _1568_/B vssd1 vssd1 vccd1 vccd1 _1177_/A sky130_fd_sc_hd__inv_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0888_ _0891_/A vssd1 vssd1 vccd1 vccd1 _0889_/A sky130_fd_sc_hd__buf_1
X_0957_ data_wdata_o[5] _0947_/X _1782_/Q _0949_/X vssd1 vssd1 vccd1 vccd1 _1890_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1509_ _1773_/Q vssd1 vssd1 vccd1 vccd1 _1509_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1503__A rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
X_1860_ _1903_/CLK _1860_/D vssd1 vssd1 vccd1 vccd1 _1860_/Q sky130_fd_sc_hd__dfxtp_2
X_1791_ _1881_/CLK _1791_/D vssd1 vssd1 vccd1 vccd1 _1791_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1156_ _1613_/B vssd1 vssd1 vccd1 vccd1 _1672_/S sky130_fd_sc_hd__inv_2
X_1087_ _1119_/A vssd1 vssd1 vccd1 vccd1 _1111_/A sky130_fd_sc_hd__buf_1
X_1225_ _1587_/C vssd1 vssd1 vccd1 vccd1 _1598_/B sky130_fd_sc_hd__inv_2
XFILLER_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1233__A rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0982__A _1782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1010_ _1801_/Q vssd1 vssd1 vccd1 vccd1 _1275_/A sky130_fd_sc_hd__inv_2
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1843_ _1852_/CLK _1843_/D vssd1 vssd1 vccd1 vccd1 _1843_/Q sky130_fd_sc_hd__dfxtp_2
X_1774_ _1888_/CLK _1774_/D vssd1 vssd1 vccd1 vccd1 _1774_/Q sky130_fd_sc_hd__dfxtp_2
X_1208_ _1833_/Q _1208_/B vssd1 vssd1 vccd1 vccd1 _1208_/Y sky130_fd_sc_hd__nor2_2
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1139_ _1845_/Q _1133_/X data_rdata_i[4] _1134_/X _1138_/X vssd1 vssd1 vccd1 vccd1
+ _1845_/D sky130_fd_sc_hd__o221a_2
XFILLER_25_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1416__B1 _1780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1490_ _1490_/A vssd1 vssd1 vccd1 vccd1 _1510_/A sky130_fd_sc_hd__buf_1
XFILLER_3_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1826_ _1875_/CLK _1826_/D _1273_/X vssd1 vssd1 vccd1 vccd1 _1826_/Q sky130_fd_sc_hd__dfrtp_2
X_1688_ _1453_/Y _1454_/X _1692_/S vssd1 vssd1 vccd1 vccd1 _1688_/X sky130_fd_sc_hd__mux2_1
X_1757_ _1771_/CLK _1757_/D vssd1 vssd1 vccd1 vccd1 _1757_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_4_4_0_clk_i clkbuf_4_5_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1851_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_13_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0990_ _1006_/A vssd1 vssd1 vccd1 vccd1 _1468_/B sky130_fd_sc_hd__inv_2
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1611_ _1611_/A vssd1 vssd1 vccd1 vccd1 _1611_/X sky130_fd_sc_hd__buf_1
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1542_ _1542_/A vssd1 vssd1 vccd1 vccd1 _1543_/B sky130_fd_sc_hd__buf_1
X_1473_ _0945_/B _1423_/X _1436_/Y _1425_/X vssd1 vssd1 vccd1 vccd1 _1797_/D sky130_fd_sc_hd__o22ai_2
XFILLER_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1809_ _1892_/CLK _1809_/D _1354_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[4] sky130_fd_sc_hd__dfrtp_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0973_ _0976_/A vssd1 vssd1 vccd1 vccd1 _0974_/A sky130_fd_sc_hd__buf_1
X_1525_ _1176_/A _1756_/Q _1755_/Q _1524_/Y vssd1 vssd1 vccd1 vccd1 _1526_/B sky130_fd_sc_hd__o22a_2
XFILLER_19_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1456_ _1738_/Q _1739_/Q vssd1 vssd1 vccd1 vccd1 _1458_/B sky130_fd_sc_hd__or2_2
X_1387_ _1391_/A vssd1 vssd1 vccd1 vccd1 _1388_/A sky130_fd_sc_hd__buf_1
XFILLER_27_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1310_ _1327_/A vssd1 vssd1 vccd1 vccd1 _1310_/X sky130_fd_sc_hd__buf_1
X_1241_ _1768_/Q _1241_/B vssd1 vssd1 vccd1 vccd1 _1242_/B sky130_fd_sc_hd__or2_2
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1172_ _1765_/Q _1171_/X _1765_/Q _1171_/X vssd1 vssd1 vccd1 vccd1 _1568_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_32_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0956_ _0956_/A vssd1 vssd1 vccd1 vccd1 _0956_/X sky130_fd_sc_hd__buf_1
X_0887_ data_wdata_o[21] _0874_/X _1782_/Q _0876_/X vssd1 vssd1 vccd1 vccd1 _1906_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_46_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1508_ _1521_/A _1508_/B vssd1 vssd1 vccd1 vccd1 _1508_/Y sky130_fd_sc_hd__nor2_2
X_1439_ _1439_/A vssd1 vssd1 vccd1 vccd1 _1681_/S sky130_fd_sc_hd__buf_1
XFILLER_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1790_ _1881_/CLK _1790_/D vssd1 vssd1 vccd1 vccd1 _1790_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__0972__B1 _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1224_ _1224_/A vssd1 vssd1 vccd1 vccd1 _1587_/C sky130_fd_sc_hd__buf_1
X_1086_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1086_/X sky130_fd_sc_hd__buf_1
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1155_ _1155_/A _1745_/Q vssd1 vssd1 vccd1 vccd1 _1613_/B sky130_fd_sc_hd__nand2_2
X_0939_ _0942_/A vssd1 vssd1 vccd1 vccd1 _0940_/A sky130_fd_sc_hd__buf_1
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0954__B1 _1783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0982__B _1781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1773_ _1888_/CLK _1773_/D vssd1 vssd1 vccd1 vccd1 _1773_/Q sky130_fd_sc_hd__dfxtp_2
X_1842_ _1851_/CLK _1842_/D vssd1 vssd1 vccd1 vccd1 _1842_/Q sky130_fd_sc_hd__dfxtp_2
X_1207_ _1190_/A _1206_/X _1203_/X _1834_/Q _1186_/A vssd1 vssd1 vccd1 vccd1 _1834_/D
+ sky130_fd_sc_hd__a32o_2
XANTENNA__1122__B1 data_rdata_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1370__B1 _1777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1138_ _1145_/A vssd1 vssd1 vccd1 vccd1 _1138_/X sky130_fd_sc_hd__buf_1
X_1069_ _1069_/A vssd1 vssd1 vccd1 vccd1 _1150_/B sky130_fd_sc_hd__inv_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_clk_i clkbuf_4_1_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1771_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__1113__B1 data_rdata_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1416__A1 _1779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1104__B1 data_rdata_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1352__B1 _1782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1825_ _1875_/CLK _1825_/D _1284_/X vssd1 vssd1 vccd1 vccd1 _1825_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1756_ _1771_/CLK _1756_/D vssd1 vssd1 vccd1 vccd1 _1756_/Q sky130_fd_sc_hd__dfxtp_2
X_1687_ _1581_/B rx_i _1695_/S vssd1 vssd1 vccd1 vccd1 _1687_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1582__B1 rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1610_ _1610_/A _1688_/X vssd1 vssd1 vccd1 vccd1 _1611_/A sky130_fd_sc_hd__or2_2
XFILLER_8_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1573__B1 _1782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1472_ _0873_/B _1425_/X _1309_/A _1471_/X vssd1 vssd1 vccd1 vccd1 _1798_/D sky130_fd_sc_hd__o22ai_2
X_1541_ _1759_/Q _1540_/B _1551_/C vssd1 vssd1 vccd1 vccd1 _1542_/A sky130_fd_sc_hd__a21bo_2
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1808_ _1840_/CLK _1808_/D _1357_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[3] sky130_fd_sc_hd__dfrtp_2
X_1739_ _1840_/CLK _1739_/D vssd1 vssd1 vccd1 vccd1 _1739_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0972_ data_wdata_o[1] _0963_/X _1778_/Q _0964_/X vssd1 vssd1 vccd1 vccd1 _1886_/D
+ sky130_fd_sc_hd__a22o_2
X_1524_ _1756_/Q vssd1 vssd1 vccd1 vccd1 _1524_/Y sky130_fd_sc_hd__inv_2
X_1386_ _1386_/A vssd1 vssd1 vccd1 vccd1 _1386_/X sky130_fd_sc_hd__buf_1
X_1455_ _1455_/A vssd1 vssd1 vccd1 vccd1 _1725_/S sky130_fd_sc_hd__buf_1
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1517__A rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0985__B _1777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1240_ _1766_/Q _1767_/Q vssd1 vssd1 vccd1 vccd1 _1241_/B sky130_fd_sc_hd__or2_2
X_1171_ _1763_/Q _1764_/Q _1560_/B vssd1 vssd1 vccd1 vccd1 _1171_/X sky130_fd_sc_hd__or3_2
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0886_ _0886_/A vssd1 vssd1 vccd1 vccd1 _0886_/X sky130_fd_sc_hd__buf_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0955_ _0961_/A vssd1 vssd1 vccd1 vccd1 _0956_/A sky130_fd_sc_hd__buf_1
X_1507_ _1508_/B vssd1 vssd1 vccd1 vccd1 _1507_/Y sky130_fd_sc_hd__inv_2
X_1369_ _1369_/A vssd1 vssd1 vccd1 vccd1 _1369_/X sky130_fd_sc_hd__buf_1
X_1438_ _1436_/Y _1423_/X _1428_/A _1437_/X vssd1 vssd1 vccd1 vccd1 _1795_/D sky130_fd_sc_hd__o22ai_2
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1154_ _1154_/A _1744_/Q vssd1 vssd1 vccd1 vccd1 _1160_/A sky130_fd_sc_hd__nand2_2
X_1223_ rst_i _1605_/A vssd1 vssd1 vccd1 vccd1 _1224_/A sky130_fd_sc_hd__or2_2
X_1085_ _1117_/A vssd1 vssd1 vccd1 vccd1 _1110_/A sky130_fd_sc_hd__buf_1
X_0938_ data_wdata_o[9] _0929_/X _1778_/Q _0930_/X vssd1 vssd1 vccd1 vccd1 _1894_/D
+ sky130_fd_sc_hd__a22o_2
X_0869_ _1754_/Q vssd1 vssd1 vccd1 vccd1 _1002_/A sky130_fd_sc_hd__inv_2
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0890__B1 _1781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0982__C _1780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1772_ _1888_/CLK _1772_/D vssd1 vssd1 vccd1 vccd1 _1772_/Q sky130_fd_sc_hd__dfxtp_2
X_1841_ _1852_/CLK _1841_/D vssd1 vssd1 vccd1 vccd1 _1841_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1206_ _1834_/Q _1833_/Q _1201_/Y vssd1 vssd1 vccd1 vccd1 _1206_/X sky130_fd_sc_hd__a21o_2
XANTENNA_clkbuf_0_clk_i_A clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1137_ _1846_/Q _1133_/X data_rdata_i[5] _1134_/X _1131_/X vssd1 vssd1 vccd1 vccd1
+ _1846_/D sky130_fd_sc_hd__o221a_2
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1068_ _1831_/Q _1795_/Q _1884_/Q vssd1 vssd1 vccd1 vccd1 _1069_/A sky130_fd_sc_hd__o21ai_2
XANTENNA_clkbuf_3_2_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0985__C_N _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1686_ _1685_/X _1872_/Q _1794_/Q vssd1 vssd1 vccd1 vccd1 _1686_/X sky130_fd_sc_hd__mux2_1
X_1824_ _1875_/CLK _1824_/D _1290_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[11] sky130_fd_sc_hd__dfrtp_2
XFILLER_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1755_ _1840_/CLK _1755_/D vssd1 vssd1 vccd1 vccd1 _1755_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1098__B1 data_rdata_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1540_ _1759_/Q _1540_/B vssd1 vssd1 vccd1 vccd1 _1551_/C sky130_fd_sc_hd__or2_2
XFILLER_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1471_ _1471_/A _1471_/B vssd1 vssd1 vccd1 vccd1 _1471_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1089__B1 data_rdata_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1807_ _1888_/CLK _1807_/D _1363_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[2] sky130_fd_sc_hd__dfrtp_2
X_1738_ _1840_/CLK _1738_/D vssd1 vssd1 vccd1 vccd1 _1738_/Q sky130_fd_sc_hd__dfxtp_2
X_1669_ _1622_/X _1652_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1740_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0971_ _0971_/A vssd1 vssd1 vccd1 vccd1 _0971_/X sky130_fd_sc_hd__buf_1
X_1454_ _1450_/Y _1448_/Y _1751_/Q _1453_/Y _1451_/X vssd1 vssd1 vccd1 vccd1 _1454_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1523_ _1837_/Q _1755_/Q vssd1 vssd1 vccd1 vccd1 _1523_/Y sky130_fd_sc_hd__nor2_2
X_1385_ _1391_/A vssd1 vssd1 vccd1 vccd1 _1386_/A sky130_fd_sc_hd__buf_1
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1170_ _1540_/B _1176_/D vssd1 vssd1 vccd1 vccd1 _1560_/B sky130_fd_sc_hd__or2_2
X_0885_ _0891_/A vssd1 vssd1 vccd1 vccd1 _0886_/A sky130_fd_sc_hd__buf_1
X_0954_ data_wdata_o[6] _0947_/X _1783_/Q _0949_/X vssd1 vssd1 vccd1 vccd1 _1891_/D
+ sky130_fd_sc_hd__a22o_2
X_1437_ _1275_/X _1420_/B _1471_/A _0871_/A _1280_/X vssd1 vssd1 vccd1 vccd1 _1437_/X
+ sky130_fd_sc_hd__o2111a_2
X_1506_ _1772_/Q _1505_/B _1505_/Y vssd1 vssd1 vccd1 vccd1 _1508_/B sky130_fd_sc_hd__a21oi_2
X_1299_ data_addr_o[10] _1292_/X _1779_/Q _1294_/X vssd1 vssd1 vccd1 vccd1 _1823_/D
+ sky130_fd_sc_hd__a22o_2
X_1368_ _1373_/A vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__buf_1
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1084_ _1119_/A vssd1 vssd1 vccd1 vccd1 _1117_/A sky130_fd_sc_hd__inv_2
X_1222_ _1581_/B vssd1 vssd1 vccd1 vccd1 _1439_/A sky130_fd_sc_hd__inv_2
X_1153_ data_req_o _1152_/A _1737_/X _1152_/Y _1145_/X vssd1 vssd1 vccd1 vccd1 _1839_/D
+ sky130_fd_sc_hd__o221a_2
X_0937_ _0937_/A vssd1 vssd1 vccd1 vccd1 _0937_/X sky130_fd_sc_hd__buf_1
X_0868_ _1753_/Q vssd1 vssd1 vccd1 vccd1 _1226_/B sky130_fd_sc_hd__inv_2
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0982__D _1779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1840_ _1840_/CLK _1840_/D vssd1 vssd1 vccd1 vccd1 data_we_o sky130_fd_sc_hd__dfxtp_2
X_1771_ _1771_/CLK _1771_/D vssd1 vssd1 vccd1 vccd1 _1771_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1205_ _1205_/A vssd1 vssd1 vccd1 vccd1 _1835_/D sky130_fd_sc_hd__inv_2
X_1136_ _1847_/Q _1133_/X data_rdata_i[6] _1134_/X _1131_/X vssd1 vssd1 vccd1 vccd1
+ _1847_/D sky130_fd_sc_hd__o221a_2
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1067_ _1067_/A _1067_/B _1080_/A vssd1 vssd1 vccd1 vccd1 _1083_/A sky130_fd_sc_hd__or3b_2
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_6_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1823_ _1883_/CLK _1823_/D _1298_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[10] sky130_fd_sc_hd__dfrtp_2
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1685_ _1684_/X _1864_/Q _1798_/Q vssd1 vssd1 vccd1 vccd1 _1685_/X sky130_fd_sc_hd__mux2_1
X_1754_ _1851_/CLK _1754_/D vssd1 vssd1 vccd1 vccd1 _1754_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1361__A _1361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1119_ _1119_/A vssd1 vssd1 vccd1 vccd1 _1141_/A sky130_fd_sc_hd__buf_1
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1470_ _0980_/X _0993_/Y _1802_/Q _1469_/X vssd1 vssd1 vccd1 vccd1 _1802_/D sky130_fd_sc_hd__a22o_2
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1806_ _1888_/CLK _1806_/D _1366_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[1] sky130_fd_sc_hd__dfrtp_2
X_1599_ rx_i _1591_/B _1683_/X _1584_/A _1598_/X vssd1 vssd1 vccd1 vccd1 _1599_/Y
+ sky130_fd_sc_hd__o221ai_2
X_1668_ _1620_/X _1645_/X _1672_/S vssd1 vssd1 vccd1 vccd1 _1739_/D sky130_fd_sc_hd__mux2_1
X_1737_ _1065_/Y _1149_/Y _1737_/S vssd1 vssd1 vccd1 vccd1 _1737_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0970_ _0976_/A vssd1 vssd1 vccd1 vccd1 _0971_/A sky130_fd_sc_hd__buf_1
X_1453_ _1751_/Q vssd1 vssd1 vccd1 vccd1 _1453_/Y sky130_fd_sc_hd__inv_2
X_1522_ _1600_/A _1522_/B vssd1 vssd1 vccd1 vccd1 _1522_/Y sky130_fd_sc_hd__nor2_2
X_1384_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1391_/A sky130_fd_sc_hd__buf_1
XFILLER_50_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0884_ _1384_/A vssd1 vssd1 vccd1 vccd1 _0891_/A sky130_fd_sc_hd__buf_1
XANTENNA__0975__B1 _1777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0953_ _0953_/A vssd1 vssd1 vccd1 vccd1 _0953_/X sky130_fd_sc_hd__buf_1
X_1505_ _1772_/Q _1505_/B vssd1 vssd1 vccd1 vccd1 _1505_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__1634__A tx_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1367_ data_addr_o[1] _1358_/X _1778_/Q _1359_/X vssd1 vssd1 vccd1 vccd1 _1806_/D
+ sky130_fd_sc_hd__a22o_2
X_1436_ _1797_/Q vssd1 vssd1 vccd1 vccd1 _1436_/Y sky130_fd_sc_hd__inv_2
X_1298_ _1298_/A vssd1 vssd1 vccd1 vccd1 _1298_/X sky130_fd_sc_hd__buf_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1875__CLK _1875_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1694__A1 rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1143__B1 data_rdata_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0957__B1 _1782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1221_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1581_/B sky130_fd_sc_hd__buf_1
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1083_ _1083_/A _1150_/B vssd1 vssd1 vccd1 vccd1 _1119_/A sky130_fd_sc_hd__or2_2
X_1152_ _1152_/A vssd1 vssd1 vccd1 vccd1 _1152_/Y sky130_fd_sc_hd__inv_2
X_0936_ _0942_/A vssd1 vssd1 vccd1 vccd1 _0937_/A sky130_fd_sc_hd__buf_1
X_0867_ _1803_/Q vssd1 vssd1 vccd1 vccd1 _0871_/A sky130_fd_sc_hd__inv_2
X_1419_ _1419_/A vssd1 vssd1 vccd1 vccd1 _1420_/B sky130_fd_sc_hd__buf_1
XANTENNA__1125__B1 data_rdata_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1364__B1 _1779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1116__B1 data_rdata_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1770_ _1888_/CLK _1770_/D vssd1 vssd1 vccd1 vccd1 _1770_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1204_ _1208_/B _1202_/X _1195_/A _1200_/Y _1203_/X vssd1 vssd1 vccd1 vccd1 _1205_/A
+ sky130_fd_sc_hd__o32a_2
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1355__B1 _1781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1135_ _1848_/Q _1133_/X data_rdata_i[7] _1134_/X _1131_/X vssd1 vssd1 vccd1 vccd1
+ _1848_/D sky130_fd_sc_hd__o221a_2
X_1066_ _1873_/Q data_gnt_i _1065_/Y vssd1 vssd1 vccd1 vccd1 _1080_/A sky130_fd_sc_hd__a21oi_2
X_1899_ _1903_/CLK _1899_/D _0919_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[14] sky130_fd_sc_hd__dfrtp_2
X_0919_ _0919_/A vssd1 vssd1 vccd1 vccd1 _0919_/X sky130_fd_sc_hd__buf_1
XFILLER_17_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1822_ _1904_/CLK _1822_/D _1301_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[9] sky130_fd_sc_hd__dfrtp_2
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1753_ _1851_/CLK _1753_/D vssd1 vssd1 vccd1 vccd1 _1753_/Q sky130_fd_sc_hd__dfxtp_2
X_1684_ _1848_/Q _1856_/Q _1796_/Q vssd1 vssd1 vccd1 vccd1 _1684_/X sky130_fd_sc_hd__mux2_1
X_1049_ _1879_/Q _1047_/X _1047_/X _1048_/Y vssd1 vssd1 vccd1 vccd1 _1879_/D sky130_fd_sc_hd__o2bb2ai_2
X_1118_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1118_/X sky130_fd_sc_hd__buf_1
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1736_ _1247_/C _1476_/Y _1736_/S vssd1 vssd1 vccd1 vccd1 _1766_/D sky130_fd_sc_hd__mux2_1
X_1805_ _1888_/CLK _1805_/D _1369_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[0] sky130_fd_sc_hd__dfrtp_2
X_1598_ _1681_/S _1598_/B _1598_/C vssd1 vssd1 vccd1 vccd1 _1598_/X sky130_fd_sc_hd__or3_2
X_1667_ _1618_/X _1617_/B _1672_/S vssd1 vssd1 vccd1 vccd1 _1738_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1383_ _1383_/A vssd1 vssd1 vccd1 vccd1 _1383_/X sky130_fd_sc_hd__buf_1
X_1452_ _1450_/Y _1448_/Y _1451_/X vssd1 vssd1 vccd1 vccd1 _1452_/X sky130_fd_sc_hd__o21a_2
X_1521_ _1521_/A _1521_/B vssd1 vssd1 vccd1 vccd1 _1521_/Y sky130_fd_sc_hd__nor2_2
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1719_ _1554_/B _1555_/X _1725_/S vssd1 vssd1 vccd1 vccd1 _1761_/D sky130_fd_sc_hd__mux2_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0952_ _0961_/A vssd1 vssd1 vccd1 vccd1 _0953_/A sky130_fd_sc_hd__buf_1
X_0883_ _1154_/A vssd1 vssd1 vccd1 vccd1 _1384_/A sky130_fd_sc_hd__buf_1
X_1504_ _1504_/A vssd1 vssd1 vccd1 vccd1 _1504_/X sky130_fd_sc_hd__buf_1
XANTENNA__0975__A1 data_wdata_o[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1435_ _1435_/A vssd1 vssd1 vccd1 vccd1 _1794_/D sky130_fd_sc_hd__buf_1
X_1366_ _1366_/A vssd1 vssd1 vccd1 vccd1 _1366_/X sky130_fd_sc_hd__buf_1
X_1297_ _1306_/A vssd1 vssd1 vccd1 vccd1 _1298_/A sky130_fd_sc_hd__buf_1
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0957__A1 data_wdata_o[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1220_ rst_i _1220_/B vssd1 vssd1 vccd1 vccd1 _1221_/A sky130_fd_sc_hd__or2_2
X_1151_ _1149_/Y _1076_/A _1080_/Y _1150_/X vssd1 vssd1 vccd1 vccd1 _1152_/A sky130_fd_sc_hd__a211o_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1082_ rst_i _1082_/B vssd1 vssd1 vccd1 vccd1 _1873_/D sky130_fd_sc_hd__nor2_2
X_0866_ _1798_/Q vssd1 vssd1 vccd1 vccd1 _0873_/B sky130_fd_sc_hd__inv_2
X_0935_ data_wdata_o[10] _0929_/X _1779_/Q _0930_/X vssd1 vssd1 vccd1 vccd1 _1895_/D
+ sky130_fd_sc_hd__a22o_2
X_1349_ data_addr_o[6] _1342_/X _1783_/Q _1344_/X vssd1 vssd1 vccd1 vccd1 _1811_/D
+ sky130_fd_sc_hd__a22o_2
X_1418_ _1777_/Q _1413_/X _1778_/Q _1414_/X vssd1 vssd1 vccd1 vccd1 _1777_/D sky130_fd_sc_hd__a22o_2
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1052__B1 _1779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1203_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1203_/X sky130_fd_sc_hd__buf_1
X_1134_ _1141_/A vssd1 vssd1 vccd1 vccd1 _1134_/X sky130_fd_sc_hd__buf_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1065_ _1873_/Q _1065_/B vssd1 vssd1 vccd1 vccd1 _1065_/Y sky130_fd_sc_hd__nor2_2
XFILLER_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0918_ _0927_/A vssd1 vssd1 vccd1 vccd1 _0919_/A sky130_fd_sc_hd__buf_1
X_1898_ _1903_/CLK _1898_/D _0922_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[13] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1821_ _1883_/CLK _1821_/D _1304_/X vssd1 vssd1 vccd1 vccd1 data_addr_o[8] sky130_fd_sc_hd__dfrtp_2
XFILLER_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1683_ _1597_/X _1598_/C _1683_/S vssd1 vssd1 vccd1 vccd1 _1683_/X sky130_fd_sc_hd__mux2_1
X_1752_ _1851_/CLK _1752_/D vssd1 vssd1 vccd1 vccd1 _1752_/Q sky130_fd_sc_hd__dfxtp_2
X_1117_ _1117_/A vssd1 vssd1 vccd1 vccd1 _1140_/A sky130_fd_sc_hd__buf_1
X_1048_ _1800_/Q _1707_/X _1780_/Q _1029_/X vssd1 vssd1 vccd1 vccd1 _1048_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_0_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1007__B1 _1006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1666_ _1615_/X _1672_/S _1666_/S vssd1 vssd1 vccd1 vccd1 _1745_/D sky130_fd_sc_hd__mux2_1
X_1735_ _1484_/B _1485_/X _1736_/S vssd1 vssd1 vccd1 vccd1 _1767_/D sky130_fd_sc_hd__mux2_1
X_1804_ _1840_/CLK _1804_/D vssd1 vssd1 vccd1 vccd1 _1804_/Q sky130_fd_sc_hd__dfxtp_2
X_1597_ _1597_/A vssd1 vssd1 vccd1 vccd1 _1597_/X sky130_fd_sc_hd__buf_1
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1520_ _1521_/B vssd1 vssd1 vccd1 vccd1 _1520_/Y sky130_fd_sc_hd__inv_2
X_1382_ _1382_/A vssd1 vssd1 vccd1 vccd1 _1383_/A sky130_fd_sc_hd__buf_1
X_1451_ _1750_/Q _1451_/B vssd1 vssd1 vccd1 vccd1 _1451_/X sky130_fd_sc_hd__or2_2
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1649_ _1575_/X _1007_/X _1649_/S vssd1 vssd1 vccd1 vccd1 _1649_/X sky130_fd_sc_hd__mux2_1
X_1718_ _1558_/B _1559_/X _1725_/S vssd1 vssd1 vccd1 vccd1 _1762_/D sky130_fd_sc_hd__mux2_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0882_ data_wdata_o[22] _0874_/X _1783_/Q _0876_/X vssd1 vssd1 vccd1 vccd1 _1907_/D
+ sky130_fd_sc_hd__a22o_2
X_0951_ _0966_/A vssd1 vssd1 vccd1 vccd1 _0961_/A sky130_fd_sc_hd__buf_1
X_1503_ rx_i _1503_/B vssd1 vssd1 vccd1 vccd1 _1504_/A sky130_fd_sc_hd__and2_2
X_1296_ _1296_/A vssd1 vssd1 vccd1 vccd1 _1306_/A sky130_fd_sc_hd__buf_1
X_1434_ _1799_/Q _1434_/B _1434_/C vssd1 vssd1 vccd1 vccd1 _1435_/A sky130_fd_sc_hd__or3_2
X_1365_ _1373_/A vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__buf_1
XFILLER_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1150_ data_gnt_i _1150_/B vssd1 vssd1 vccd1 vccd1 _1150_/X sky130_fd_sc_hd__and2_2
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1081_ _1873_/Q _1065_/B _1076_/A _1079_/Y _1080_/Y vssd1 vssd1 vccd1 vccd1 _1082_/B
+ sky130_fd_sc_hd__o32a_2
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0934_ _0934_/A vssd1 vssd1 vccd1 vccd1 _0934_/X sky130_fd_sc_hd__buf_1
X_1417_ _1778_/Q _1413_/X _1779_/Q _1414_/X vssd1 vssd1 vccd1 vccd1 _1778_/D sky130_fd_sc_hd__a22o_2
X_1279_ _1873_/Q _1419_/A _1278_/X vssd1 vssd1 vccd1 vccd1 _1279_/X sky130_fd_sc_hd__o21a_2
X_1348_ _1348_/A vssd1 vssd1 vccd1 vccd1 _1348_/X sky130_fd_sc_hd__buf_1
XFILLER_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1202_ _1835_/Q _1201_/A _1200_/Y _1201_/Y vssd1 vssd1 vccd1 vccd1 _1202_/X sky130_fd_sc_hd__o22a_2
X_1064_ _1826_/Q vssd1 vssd1 vccd1 vccd1 _1065_/B sky130_fd_sc_hd__inv_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1133_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1133_/X sky130_fd_sc_hd__buf_1
X_1897_ _1903_/CLK _1897_/D _0925_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[12] sky130_fd_sc_hd__dfrtp_2
X_0917_ _0966_/A vssd1 vssd1 vccd1 vccd1 _0927_/A sky130_fd_sc_hd__buf_1
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1820_ _1908_/CLK _1820_/D _1307_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[31] sky130_fd_sc_hd__dfrtp_2
XFILLER_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1682_ _1589_/B _1590_/X _1695_/S vssd1 vssd1 vccd1 vccd1 _1682_/X sky130_fd_sc_hd__mux2_1
X_1751_ _1830_/CLK _1751_/D vssd1 vssd1 vccd1 vccd1 _1751_/Q sky130_fd_sc_hd__dfxtp_2
X_1047_ _1047_/A vssd1 vssd1 vccd1 vccd1 _1047_/X sky130_fd_sc_hd__buf_1
X_1116_ _1857_/Q _1110_/X data_rdata_i[16] _1111_/X _1115_/X vssd1 vssd1 vccd1 vccd1
+ _1857_/D sky130_fd_sc_hd__o221a_2
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1803_ _1892_/CLK _1803_/D _1374_/X vssd1 vssd1 vccd1 vccd1 _1803_/Q sky130_fd_sc_hd__dfrtp_2
X_1665_ _1614_/X _1181_/Y _1666_/S vssd1 vssd1 vccd1 vccd1 _1744_/D sky130_fd_sc_hd__mux2_1
X_1734_ _1488_/B _1489_/X _1736_/S vssd1 vssd1 vccd1 vccd1 _1768_/D sky130_fd_sc_hd__mux2_1
X_1596_ _1610_/A _1598_/C vssd1 vssd1 vccd1 vccd1 _1597_/A sky130_fd_sc_hd__or2_2
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0920__B1 _1783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1450_ _1750_/Q vssd1 vssd1 vccd1 vccd1 _1450_/Y sky130_fd_sc_hd__inv_4
X_1381_ _1381_/A vssd1 vssd1 vccd1 vccd1 _1381_/X sky130_fd_sc_hd__buf_1
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_clk_i clkbuf_3_6_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _1903_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1717_ _1562_/Y _1563_/Y _1725_/S vssd1 vssd1 vccd1 vccd1 _1763_/D sky130_fd_sc_hd__mux2_1
X_1579_ _1579_/A vssd1 vssd1 vccd1 vccd1 _1579_/X sky130_fd_sc_hd__buf_1
X_1648_ _1743_/Q _1466_/X _1652_/S vssd1 vssd1 vccd1 vccd1 _1648_/X sky130_fd_sc_hd__mux2_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0902__B1 _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0969__B1 _1779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1146__B1 data_rdata_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0881_ _1145_/A vssd1 vssd1 vccd1 vccd1 _0881_/X sky130_fd_sc_hd__buf_1
X_0950_ data_wdata_o[7] _0947_/X _1784_/Q _0949_/X vssd1 vssd1 vccd1 vccd1 _1892_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1433_ _1275_/A _1424_/X _1309_/A vssd1 vssd1 vccd1 vccd1 _1434_/C sky130_fd_sc_hd__a21oi_2
X_1502_ _1502_/A vssd1 vssd1 vccd1 vccd1 _1503_/B sky130_fd_sc_hd__buf_1
XANTENNA__1137__B1 data_rdata_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1295_ data_addr_o[11] _1292_/X _1780_/Q _1294_/X vssd1 vssd1 vccd1 vccd1 _1824_/D
+ sky130_fd_sc_hd__a22o_2
X_1364_ data_addr_o[2] _1358_/X _1779_/Q _1359_/X vssd1 vssd1 vccd1 vccd1 _1807_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_11_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1128__B1 data_rdata_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1367__B1 _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1080_ _1080_/A _1150_/B vssd1 vssd1 vccd1 vccd1 _1080_/Y sky130_fd_sc_hd__nor2_2
X_0933_ _0942_/A vssd1 vssd1 vccd1 vccd1 _0934_/A sky130_fd_sc_hd__buf_1
X_1416_ _1779_/Q _1413_/X _1780_/Q _1414_/X vssd1 vssd1 vccd1 vccd1 _1779_/D sky130_fd_sc_hd__a22o_2
X_1347_ _1356_/A vssd1 vssd1 vccd1 vccd1 _1348_/A sky130_fd_sc_hd__buf_1
X_1278_ _1278_/A _1469_/A vssd1 vssd1 vccd1 vccd1 _1278_/X sky130_fd_sc_hd__or2_2
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1349__B1 _1783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1201_ _1201_/A vssd1 vssd1 vccd1 vccd1 _1201_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1132_ _1849_/Q _1126_/X data_rdata_i[8] _1127_/X _1131_/X vssd1 vssd1 vccd1 vccd1
+ _1849_/D sky130_fd_sc_hd__o221a_2
X_1063_ data_rvalid_i vssd1 vssd1 vccd1 vccd1 _1067_/B sky130_fd_sc_hd__inv_2
X_0916_ _1314_/A vssd1 vssd1 vccd1 vccd1 _0966_/A sky130_fd_sc_hd__buf_1
X_1896_ _1903_/CLK _1896_/D _0928_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[11] sky130_fd_sc_hd__dfrtp_2
XFILLER_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1750_ _1830_/CLK _1750_/D vssd1 vssd1 vccd1 vccd1 _1750_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1681_ _1598_/B _1576_/A _1681_/S vssd1 vssd1 vccd1 vccd1 _1681_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1046_ _1046_/A vssd1 vssd1 vccd1 vccd1 _1046_/X sky130_fd_sc_hd__buf_1
X_1115_ _1131_/A vssd1 vssd1 vccd1 vccd1 _1115_/X sky130_fd_sc_hd__buf_1
X_1879_ _1883_/CLK _1879_/D _1046_/X vssd1 vssd1 vccd1 vccd1 _1879_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1802_ _1883_/CLK _1802_/D _1377_/X vssd1 vssd1 vccd1 vccd1 _1802_/Q sky130_fd_sc_hd__dfrtp_2
X_1733_ _1493_/B _1494_/X _1736_/S vssd1 vssd1 vccd1 vccd1 _1769_/D sky130_fd_sc_hd__mux2_1
X_1595_ _1595_/A vssd1 vssd1 vccd1 vccd1 _1610_/A sky130_fd_sc_hd__buf_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1664_ _1587_/C _1521_/A _1695_/S vssd1 vssd1 vccd1 vccd1 _1664_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1029_ _1570_/A vssd1 vssd1 vccd1 vccd1 _1029_/X sky130_fd_sc_hd__buf_1
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1380_ _1382_/A vssd1 vssd1 vccd1 vccd1 _1381_/A sky130_fd_sc_hd__buf_1
X_1716_ _1566_/B _1567_/X _1725_/S vssd1 vssd1 vccd1 vccd1 _1764_/D sky130_fd_sc_hd__mux2_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _1828_/Q _1578_/B _1830_/Q _1829_/Q vssd1 vssd1 vccd1 vccd1 _1579_/A sky130_fd_sc_hd__or4_2
X_1647_ _1742_/Q _1464_/X _1652_/S vssd1 vssd1 vccd1 vccd1 _1647_/X sky130_fd_sc_hd__mux2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1091__B1 data_rdata_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0969__A1 data_wdata_o[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0880_ _1154_/A vssd1 vssd1 vccd1 vccd1 _1145_/A sky130_fd_sc_hd__buf_1
X_1432_ _1432_/A vssd1 vssd1 vccd1 vccd1 _1799_/D sky130_fd_sc_hd__buf_1
X_1501_ _1771_/Q _1500_/B _1505_/B vssd1 vssd1 vccd1 vccd1 _1502_/A sky130_fd_sc_hd__a21bo_2
X_1363_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1363_/X sky130_fd_sc_hd__buf_1
X_1294_ _1294_/A vssd1 vssd1 vccd1 vccd1 _1294_/X sky130_fd_sc_hd__buf_1
XFILLER_11_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0887__B1 _1782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0932_ _0966_/A vssd1 vssd1 vccd1 vccd1 _0942_/A sky130_fd_sc_hd__buf_1
XFILLER_3_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1415_ _1780_/Q _1413_/X _1781_/Q _1414_/X vssd1 vssd1 vccd1 vccd1 _1780_/D sky130_fd_sc_hd__a22o_2
X_1346_ _1361_/A vssd1 vssd1 vccd1 vccd1 _1356_/A sky130_fd_sc_hd__buf_1
X_1277_ _1884_/Q vssd1 vssd1 vccd1 vccd1 _1278_/A sky130_fd_sc_hd__inv_2
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1200_ _1835_/Q vssd1 vssd1 vccd1 vccd1 _1200_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1131_ _1131_/A vssd1 vssd1 vccd1 vccd1 _1131_/X sky130_fd_sc_hd__buf_1
X_1062_ _1874_/Q vssd1 vssd1 vccd1 vccd1 _1067_/A sky130_fd_sc_hd__inv_2
X_0915_ _1154_/A vssd1 vssd1 vccd1 vccd1 _1314_/A sky130_fd_sc_hd__buf_1
X_1895_ _1895_/CLK _1895_/D _0934_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[10] sky130_fd_sc_hd__dfrtp_2
X_1329_ data_wdata_o[27] _1327_/X _1780_/Q _1328_/X vssd1 vssd1 vccd1 vccd1 _1816_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1680_ _1679_/X _1867_/Q _1794_/Q vssd1 vssd1 vccd1 vccd1 _1680_/X sky130_fd_sc_hd__mux2_1
X_1114_ _1858_/Q _1110_/X data_rdata_i[17] _1111_/X _1108_/X vssd1 vssd1 vccd1 vccd1
+ _1858_/D sky130_fd_sc_hd__o221a_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1045_ _1058_/A vssd1 vssd1 vccd1 vccd1 _1046_/A sky130_fd_sc_hd__buf_1
X_1878_ _1883_/CLK _1878_/D _1051_/X vssd1 vssd1 vccd1 vccd1 _1878_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1412__B1 _1782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1801_ _1875_/CLK _1801_/D _1379_/X vssd1 vssd1 vccd1 vccd1 _1801_/Q sky130_fd_sc_hd__dfrtp_2
X_1732_ _1498_/B _1499_/X _1736_/S vssd1 vssd1 vccd1 vccd1 _1770_/D sky130_fd_sc_hd__mux2_1
X_1663_ _1612_/Y _1238_/B _1681_/X vssd1 vssd1 vccd1 vccd1 _1751_/D sky130_fd_sc_hd__mux2_1
X_1594_ _1689_/X vssd1 vssd1 vccd1 vccd1 _1598_/C sky130_fd_sc_hd__inv_2
XFILLER_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1028_ _1047_/A vssd1 vssd1 vccd1 vccd1 _1028_/X sky130_fd_sc_hd__buf_1
XFILLER_14_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1498__A rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1646_ _1604_/X _1691_/X _1683_/S vssd1 vssd1 vccd1 vccd1 _1646_/X sky130_fd_sc_hd__mux2_1
X_1715_ _1177_/A _1568_/Y _1725_/S vssd1 vssd1 vccd1 vccd1 _1765_/D sky130_fd_sc_hd__mux2_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ _1577_/A vssd1 vssd1 vccd1 vccd1 _1656_/S sky130_fd_sc_hd__buf_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_7_0_clk_i clkbuf_4_7_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1895_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1500_ _1771_/Q _1500_/B vssd1 vssd1 vccd1 vccd1 _1505_/B sky130_fd_sc_hd__or2_2
X_1293_ _1293_/A vssd1 vssd1 vccd1 vccd1 _1294_/A sky130_fd_sc_hd__inv_2
X_1431_ _1431_/A _1431_/B vssd1 vssd1 vccd1 vccd1 _1432_/A sky130_fd_sc_hd__or2_2
X_1362_ _1373_/A vssd1 vssd1 vccd1 vccd1 _1363_/A sky130_fd_sc_hd__buf_1
XFILLER_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1720__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1629_ _1629_/A vssd1 vssd1 vccd1 vccd1 _1629_/X sky130_fd_sc_hd__buf_1
XFILLER_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0931_ data_wdata_o[11] _0929_/X _1780_/Q _0930_/X vssd1 vssd1 vccd1 vccd1 _1896_/D
+ sky130_fd_sc_hd__a22o_2
XANTENNA__1715__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1276_ _1276_/A vssd1 vssd1 vccd1 vccd1 _1419_/A sky130_fd_sc_hd__buf_1
XFILLER_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1345_ data_addr_o[7] _1342_/X _1784_/Q _1344_/X vssd1 vssd1 vccd1 vccd1 _1812_/D
+ sky130_fd_sc_hd__a22o_2
X_1414_ _1414_/A vssd1 vssd1 vccd1 vccd1 _1414_/X sky130_fd_sc_hd__buf_1
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_4_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_1130_ _1850_/Q _1126_/X data_rdata_i[9] _1127_/X _1124_/X vssd1 vssd1 vccd1 vccd1
+ _1850_/D sky130_fd_sc_hd__o221a_2
X_1061_ _1061_/A vssd1 vssd1 vccd1 vccd1 _1876_/D sky130_fd_sc_hd__buf_1
XFILLER_18_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0914_ data_wdata_o[15] _0911_/X _1784_/Q _0913_/X vssd1 vssd1 vccd1 vccd1 _1900_/D
+ sky130_fd_sc_hd__a22o_2
X_1894_ _1903_/CLK _1894_/D _0937_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[9] sky130_fd_sc_hd__dfrtp_2
X_1328_ _1328_/A vssd1 vssd1 vccd1 vccd1 _1328_/X sky130_fd_sc_hd__buf_1
X_1259_ _1829_/Q _1219_/A _1830_/Q _1229_/Y vssd1 vssd1 vccd1 vccd1 _1259_/X sky130_fd_sc_hd__o31a_2
XANTENNA__0950__B1 _1784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0941__B1 _1777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1044_ _1296_/A vssd1 vssd1 vccd1 vccd1 _1058_/A sky130_fd_sc_hd__buf_1
X_1113_ _1859_/Q _1110_/X data_rdata_i[18] _1111_/X _1108_/X vssd1 vssd1 vccd1 vccd1
+ _1859_/D sky130_fd_sc_hd__o221a_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1877_ _1881_/CLK _1877_/D _1055_/X vssd1 vssd1 vccd1 vccd1 _1877_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1412__A1 _1781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0923__B1 _1782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1800_ _1875_/CLK _1800_/D _1381_/X vssd1 vssd1 vccd1 vccd1 _1800_/Q sky130_fd_sc_hd__dfrtp_2
X_1662_ _1609_/Y _1238_/C _1681_/X vssd1 vssd1 vccd1 vccd1 _1750_/D sky130_fd_sc_hd__mux2_1
X_1731_ _1503_/B _1504_/X _1736_/S vssd1 vssd1 vccd1 vccd1 _1771_/D sky130_fd_sc_hd__mux2_1
XANTENNA__0914__B1 _1784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1593_ _1682_/X _1584_/X _1589_/B _1592_/X vssd1 vssd1 vccd1 vccd1 _1593_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__1723__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1027_ _1060_/S vssd1 vssd1 vccd1 vccd1 _1047_/A sky130_fd_sc_hd__buf_1
XANTENNA__0905__B1 _1777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_clk_i clkbuf_4_3_0_clk_i/A vssd1 vssd1 vccd1 vccd1 _1892_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_44_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1321__B1 _1782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1714_ _1876_/Q _1787_/Q _1714_/S vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1718__S _1725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1576_ _1576_/A _1681_/S _1754_/Q vssd1 vssd1 vccd1 vccd1 _1577_/A sky130_fd_sc_hd__and3_2
X_1645_ _1739_/Q _1457_/X _1652_/S vssd1 vssd1 vccd1 vccd1 _1645_/X sky130_fd_sc_hd__mux2_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1741__CLK _1875_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1430_ _0991_/A _1006_/X _1422_/A _1428_/X _0963_/A vssd1 vssd1 vccd1 vccd1 _1431_/B
+ sky130_fd_sc_hd__o221ai_2
X_1292_ _1293_/A vssd1 vssd1 vccd1 vccd1 _1292_/X sky130_fd_sc_hd__buf_1
X_1361_ _1361_/A vssd1 vssd1 vccd1 vccd1 _1373_/A sky130_fd_sc_hd__buf_1
XFILLER_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1021__B uart_error vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1628_ _1628_/A vssd1 vssd1 vccd1 vccd1 _1629_/A sky130_fd_sc_hd__buf_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1559_ _1559_/A vssd1 vssd1 vccd1 vccd1 _1559_/X sky130_fd_sc_hd__buf_1
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_0_0_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0930_ _0930_/A vssd1 vssd1 vccd1 vccd1 _0930_/X sky130_fd_sc_hd__buf_1
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1413_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1413_/X sky130_fd_sc_hd__buf_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1275_ _1275_/A vssd1 vssd1 vccd1 vccd1 _1275_/X sky130_fd_sc_hd__buf_1
X_1344_ _1434_/B vssd1 vssd1 vccd1 vccd1 _1344_/X sky130_fd_sc_hd__buf_1
XFILLER_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1060_ _1640_/X _1876_/Q _1060_/S vssd1 vssd1 vccd1 vccd1 _1061_/A sky130_fd_sc_hd__mux2_2
X_0913_ _0930_/A vssd1 vssd1 vccd1 vccd1 _0913_/X sky130_fd_sc_hd__buf_1
X_1893_ _1903_/CLK _1893_/D _0940_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[8] sky130_fd_sc_hd__dfrtp_2
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1327_ _1327_/A vssd1 vssd1 vccd1 vccd1 _1327_/X sky130_fd_sc_hd__buf_1
X_1189_ _1189_/A vssd1 vssd1 vccd1 vccd1 _1190_/A sky130_fd_sc_hd__buf_1
X_1258_ _1258_/A _1258_/B _1258_/C vssd1 vssd1 vccd1 vccd1 _1258_/X sky130_fd_sc_hd__and3_2
XFILLER_33_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0950__A1 data_wdata_o[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1825__CLK _1875_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1430__A2 _1006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0941__A1 data_wdata_o[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1043_ _1880_/Q _1028_/X _1028_/X _1042_/Y vssd1 vssd1 vccd1 vccd1 _1880_/D sky130_fd_sc_hd__o2bb2ai_2
X_1112_ _1860_/Q _1110_/X data_rdata_i[19] _1111_/X _1108_/X vssd1 vssd1 vccd1 vccd1
+ _1860_/D sky130_fd_sc_hd__o221a_2
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1876_ _1881_/CLK _1876_/D _1059_/X vssd1 vssd1 vccd1 vccd1 _1876_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1220__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0923__A1 data_wdata_o[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1661_ _1606_/Y _1253_/B _1681_/X vssd1 vssd1 vccd1 vccd1 _1749_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1730_ _1507_/Y _1508_/Y _1736_/S vssd1 vssd1 vccd1 vccd1 _1772_/D sky130_fd_sc_hd__mux2_1
X_1592_ _1592_/A _1592_/B vssd1 vssd1 vccd1 vccd1 _1592_/X sky130_fd_sc_hd__and2_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1026_ _0991_/A _1007_/X _1015_/X _1019_/Y _1025_/Y vssd1 vssd1 vccd1 vccd1 _1060_/S
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_14_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1859_ _1859_/CLK _1859_/D vssd1 vssd1 vccd1 vccd1 _1859_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0905__A1 data_wdata_o[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1215__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1094__B1 data_rdata_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1321__A1 data_wdata_o[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1713_ _1877_/Q _1788_/Q _1714_/S vssd1 vssd1 vccd1 vccd1 _1713_/X sky130_fd_sc_hd__mux2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0899__B1 _1779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1575_ _1471_/A _1016_/Y _1420_/B _1570_/X vssd1 vssd1 vccd1 vccd1 _1575_/X sky130_fd_sc_hd__a2bb2o_2
X_1644_ _1196_/A _1181_/Y _1674_/S vssd1 vssd1 vccd1 vccd1 _1644_/X sky130_fd_sc_hd__mux2_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1009_ _1800_/Q _1018_/A vssd1 vssd1 vccd1 vccd1 _1569_/A sky130_fd_sc_hd__or2_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1360_ data_addr_o[3] _1358_/X _1780_/Q _1359_/X vssd1 vssd1 vccd1 vccd1 _1808_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1291_ _1469_/A _1469_/B _1802_/Q vssd1 vssd1 vccd1 vccd1 _1293_/A sky130_fd_sc_hd__or3b_2
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _1489_/A vssd1 vssd1 vccd1 vccd1 _1489_/X sky130_fd_sc_hd__buf_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1558_ _1566_/A _1558_/B vssd1 vssd1 vccd1 vccd1 _1559_/A sky130_fd_sc_hd__and2_2
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1627_ _1627_/A vssd1 vssd1 vccd1 vccd1 _1627_/X sky130_fd_sc_hd__buf_1
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_1_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1343_ _1343_/A vssd1 vssd1 vccd1 vccd1 _1434_/B sky130_fd_sc_hd__inv_2
XFILLER_3_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1412_ _1781_/Q _1407_/X _1782_/Q _1408_/X vssd1 vssd1 vccd1 vccd1 _1781_/D sky130_fd_sc_hd__a22o_2
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1274_ _1343_/A vssd1 vssd1 vccd1 vccd1 _1358_/A sky130_fd_sc_hd__buf_1
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0989_ _1832_/Q _1276_/A vssd1 vssd1 vccd1 vccd1 _1006_/A sky130_fd_sc_hd__or2_2
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1223__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0912_ _0929_/A vssd1 vssd1 vccd1 vccd1 _0930_/A sky130_fd_sc_hd__inv_2
X_1892_ _1892_/CLK _1892_/D _0943_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[7] sky130_fd_sc_hd__dfrtp_2
X_1326_ _1326_/A vssd1 vssd1 vccd1 vccd1 _1326_/X sky130_fd_sc_hd__buf_1
X_1188_ _1159_/X _1186_/X _1838_/Q _1187_/X vssd1 vssd1 vccd1 vccd1 _1838_/D sky130_fd_sc_hd__o22a_2
X_1257_ _1257_/A vssd1 vssd1 vccd1 vccd1 _1258_/C sky130_fd_sc_hd__inv_2
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1415__B1 _1781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1042_ _1800_/Q _1704_/X _1781_/Q _1029_/X vssd1 vssd1 vccd1 vccd1 _1042_/Y sky130_fd_sc_hd__a22oi_2
X_1111_ _1111_/A vssd1 vssd1 vccd1 vccd1 _1111_/X sky130_fd_sc_hd__buf_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1406__B1 tx_o vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1875_ _1875_/CLK _1875_/D vssd1 vssd1 vccd1 vccd1 _1875_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1309_ _1309_/A _1471_/B vssd1 vssd1 vccd1 vccd1 _1327_/A sky130_fd_sc_hd__or2_2
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1591_ _1595_/A _1591_/B vssd1 vssd1 vccd1 vccd1 _1592_/B sky130_fd_sc_hd__or2_2
X_1660_ _1602_/Y _1600_/B _1681_/X vssd1 vssd1 vccd1 vccd1 _1748_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1025_ _1802_/Q _1276_/A _1469_/B _1431_/A vssd1 vssd1 vccd1 vccd1 _1025_/Y sky130_fd_sc_hd__a31oi_2
X_1858_ _1859_/CLK _1858_/D vssd1 vssd1 vccd1 vccd1 _1858_/Q sky130_fd_sc_hd__dfxtp_2
X_1789_ _1881_/CLK _1789_/D vssd1 vssd1 vccd1 vccd1 _1789_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1712_ _1878_/Q _1789_/Q _1714_/S vssd1 vssd1 vccd1 vccd1 _1712_/X sky130_fd_sc_hd__mux2_1
X_1643_ _1574_/X _1006_/X _1649_/S vssd1 vssd1 vccd1 vccd1 _1643_/X sky130_fd_sc_hd__mux2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ _1800_/Q _1698_/X _1783_/Q _1029_/X vssd1 vssd1 vccd1 vccd1 _1574_/X sky130_fd_sc_hd__a22o_2
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0899__A1 data_wdata_o[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1008_ _1801_/Q _1802_/Q _1803_/Q vssd1 vssd1 vccd1 vccd1 _1018_/A sky130_fd_sc_hd__or3_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1226__A rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1290_ _1290_/A vssd1 vssd1 vccd1 vccd1 _1290_/X sky130_fd_sc_hd__buf_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1626_ _1616_/X _1648_/X vssd1 vssd1 vccd1 vccd1 _1627_/A sky130_fd_sc_hd__and2b_2
XANTENNA__0885__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ rx_i _1488_/B vssd1 vssd1 vccd1 vccd1 _1489_/A sky130_fd_sc_hd__and2_2
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1557_ _1557_/A vssd1 vssd1 vccd1 vccd1 _1558_/B sky130_fd_sc_hd__buf_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_5_0_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1273_ _1273_/A vssd1 vssd1 vccd1 vccd1 _1273_/X sky130_fd_sc_hd__buf_1
X_1342_ _1358_/A vssd1 vssd1 vccd1 vccd1 _1342_/X sky130_fd_sc_hd__buf_1
X_1411_ _1782_/Q _1407_/X _1783_/Q _1408_/X vssd1 vssd1 vccd1 vccd1 _1782_/D sky130_fd_sc_hd__a22o_2
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0988_ _0988_/A vssd1 vssd1 vccd1 vccd1 uart_error sky130_fd_sc_hd__buf_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1609_ _1673_/X _1584_/X _1690_/X _1592_/X vssd1 vssd1 vccd1 vccd1 _1609_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1130__B1 data_rdata_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0911_ _0929_/A vssd1 vssd1 vccd1 vccd1 _0911_/X sky130_fd_sc_hd__buf_1
X_1891_ _1892_/CLK _1891_/D _0953_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[6] sky130_fd_sc_hd__dfrtp_2
X_1325_ _1325_/A vssd1 vssd1 vccd1 vccd1 _1326_/A sky130_fd_sc_hd__buf_1
X_1256_ _1229_/Y _1233_/Y _1695_/S vssd1 vssd1 vccd1 vccd1 _1257_/A sky130_fd_sc_hd__o21ai_2
X_1187_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1187_/X sky130_fd_sc_hd__buf_1
XFILLER_33_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1121__B1 data_rdata_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0935__B1 _1779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1112__B1 data_rdata_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1360__B1 _1780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1415__A1 _1780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0926__B1 _1781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1110_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1110_/X sky130_fd_sc_hd__buf_1
XFILLER_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1041_ _1041_/A vssd1 vssd1 vccd1 vccd1 _1041_/X sky130_fd_sc_hd__buf_1
XANTENNA__0983__A _1784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1874_ _1875_/CLK _1874_/D vssd1 vssd1 vccd1 vccd1 _1874_/Q sky130_fd_sc_hd__dfxtp_2
X_1308_ _1794_/Q vssd1 vssd1 vccd1 vccd1 _1309_/A sky130_fd_sc_hd__inv_2
X_1239_ _1770_/Q _1771_/Q _1772_/Q _1773_/Q vssd1 vssd1 vccd1 vccd1 _1510_/B sky130_fd_sc_hd__or4_2
XANTENNA__1333__B1 _1779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1572__B1 _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1590_ _1590_/A vssd1 vssd1 vccd1 vccd1 _1590_/X sky130_fd_sc_hd__buf_1
XANTENNA__1324__B1 _1781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1024_ _1799_/Q _1006_/X _1021_/X _1022_/Y _1023_/X vssd1 vssd1 vccd1 vccd1 _1431_/A
+ sky130_fd_sc_hd__a32o_2
XANTENNA__0888__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1788_ _1881_/CLK _1788_/D vssd1 vssd1 vccd1 vccd1 _1788_/Q sky130_fd_sc_hd__dfxtp_2
X_1857_ _1859_/CLK _1857_/D vssd1 vssd1 vccd1 vccd1 _1857_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1512__A rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1711_ _1879_/Q _1790_/Q _1714_/S vssd1 vssd1 vccd1 vccd1 _1711_/X sky130_fd_sc_hd__mux2_1
X_1642_ _1573_/X _1468_/B _1649_/S vssd1 vssd1 vccd1 vccd1 _1642_/X sky130_fd_sc_hd__mux2_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _1800_/Q _1677_/X _1782_/Q _1570_/X vssd1 vssd1 vccd1 vccd1 _1573_/X sky130_fd_sc_hd__a22o_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1007_ _1220_/B _1226_/B _1605_/A _1016_/B _1006_/X vssd1 vssd1 vccd1 vccd1 _1007_/X
+ sky130_fd_sc_hd__a41o_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1556_ _1762_/Q _1551_/X _1560_/B vssd1 vssd1 vccd1 vccd1 _1557_/A sky130_fd_sc_hd__a21bo_2
X_1625_ _1625_/A vssd1 vssd1 vccd1 vccd1 _1625_/X sky130_fd_sc_hd__buf_1
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _1487_/A vssd1 vssd1 vccd1 vccd1 _1488_/B sky130_fd_sc_hd__buf_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1410_ _1783_/Q _1407_/X _1784_/Q _1408_/X vssd1 vssd1 vccd1 vccd1 _1783_/D sky130_fd_sc_hd__a22o_2
X_1272_ _1289_/A vssd1 vssd1 vccd1 vccd1 _1273_/A sky130_fd_sc_hd__buf_1
X_1341_ _1341_/A vssd1 vssd1 vccd1 vccd1 _1341_/X sky130_fd_sc_hd__buf_1
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0987_ _1752_/Q _1226_/B _1754_/Q vssd1 vssd1 vccd1 vccd1 _0988_/A sky130_fd_sc_hd__and3_2
X_1608_ _1608_/A vssd1 vssd1 vccd1 vccd1 _1608_/X sky130_fd_sc_hd__buf_1
X_1539_ _1539_/A vssd1 vssd1 vccd1 vccd1 _1539_/X sky130_fd_sc_hd__buf_1
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0910_ _0945_/B _1013_/C _0910_/C vssd1 vssd1 vccd1 vccd1 _0929_/A sky130_fd_sc_hd__or3_2
X_1890_ _1892_/CLK _1890_/D _0956_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[5] sky130_fd_sc_hd__dfrtp_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1324_ data_wdata_o[28] _1310_/X _1781_/Q _1312_/X vssd1 vssd1 vccd1 vccd1 _1817_/D
+ sky130_fd_sc_hd__a22o_2
X_1186_ _1186_/A vssd1 vssd1 vccd1 vccd1 _1186_/X sky130_fd_sc_hd__buf_1
X_1255_ _1683_/S vssd1 vssd1 vccd1 vccd1 _1695_/S sky130_fd_sc_hd__inv_2
XFILLER_3_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0926__A1 data_wdata_o[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1040_ _1040_/A vssd1 vssd1 vccd1 vccd1 _1041_/A sky130_fd_sc_hd__buf_1
X_1873_ _1875_/CLK _1873_/D vssd1 vssd1 vccd1 vccd1 _1873_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__0984__C_N _1777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1307_ _1307_/A vssd1 vssd1 vccd1 vccd1 _1307_/X sky130_fd_sc_hd__buf_1
X_1169_ _1760_/Q _1761_/Q _1759_/Q _1762_/Q vssd1 vssd1 vccd1 vccd1 _1176_/D sky130_fd_sc_hd__or4_2
X_1238_ _1600_/B _1238_/B _1238_/C vssd1 vssd1 vccd1 vccd1 _1253_/C sky130_fd_sc_hd__or3_2
XANTENNA__1030__B1 _1784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1333__A1 data_wdata_o[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1097__B1 data_rdata_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1023_ _1021_/X _1799_/Q _1023_/C vssd1 vssd1 vccd1 vccd1 _1023_/X sky130_fd_sc_hd__and3b_2
X_1787_ _1881_/CLK _1787_/D vssd1 vssd1 vccd1 vccd1 _1787_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1856_ _1903_/CLK _1856_/D vssd1 vssd1 vccd1 vccd1 _1856_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_4_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1710_ _1880_/Q _1791_/Q _1714_/S vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__mux2_1
X_1572_ _1800_/Q _1701_/X _1778_/Q _1570_/X vssd1 vssd1 vccd1 vccd1 _1572_/X sky130_fd_sc_hd__a22o_2
X_1641_ _1572_/X _1022_/Y _1649_/S vssd1 vssd1 vccd1 vccd1 _1641_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1006_ _1006_/A vssd1 vssd1 vccd1 vccd1 _1006_/X sky130_fd_sc_hd__buf_1
XFILLER_34_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1908_ _1908_/CLK _1908_/D _1629_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[23] sky130_fd_sc_hd__dfrtp_2
X_1839_ _1840_/CLK _1839_/D vssd1 vssd1 vccd1 vccd1 data_req_o sky130_fd_sc_hd__dfxtp_2
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0991__B uart_error vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1555_ _1555_/A vssd1 vssd1 vccd1 vccd1 _1555_/X sky130_fd_sc_hd__buf_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1624_ _1616_/X _1647_/X vssd1 vssd1 vccd1 vccd1 _1625_/A sky130_fd_sc_hd__and2b_2
XFILLER_39_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1486_ _1768_/Q _1241_/B _1242_/B vssd1 vssd1 vccd1 vccd1 _1487_/A sky130_fd_sc_hd__a21bo_2
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1340_ _1340_/A vssd1 vssd1 vccd1 vccd1 _1341_/A sky130_fd_sc_hd__buf_1
X_1271_ _1827_/Q _1414_/A _1578_/B _1257_/A vssd1 vssd1 vccd1 vccd1 _1827_/D sky130_fd_sc_hd__o22a_2
X_0986_ _1799_/Q vssd1 vssd1 vccd1 vccd1 _0991_/A sky130_fd_sc_hd__inv_2
X_1469_ _1469_/A _1469_/B vssd1 vssd1 vccd1 vccd1 _1469_/X sky130_fd_sc_hd__or2_2
X_1538_ _1543_/A _1538_/B vssd1 vssd1 vccd1 vccd1 _1539_/A sky130_fd_sc_hd__and2_2
X_1607_ _1610_/A _1690_/X vssd1 vssd1 vccd1 vccd1 _1608_/A sky130_fd_sc_hd__or2_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1418__B1 _1778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1323_ _1323_/A vssd1 vssd1 vccd1 vccd1 _1323_/X sky130_fd_sc_hd__buf_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1185_ _1195_/A vssd1 vssd1 vccd1 vccd1 _1186_/A sky130_fd_sc_hd__buf_1
X_1254_ _1254_/A vssd1 vssd1 vccd1 vccd1 _1683_/S sky130_fd_sc_hd__buf_1
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1409__B1 rx_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0969_ data_wdata_o[2] _0963_/X _1779_/Q _0964_/X vssd1 vssd1 vccd1 vccd1 _1887_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1872_ _1904_/CLK _1872_/D vssd1 vssd1 vccd1 vccd1 _1872_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1306_ _1306_/A vssd1 vssd1 vccd1 vccd1 _1307_/A sky130_fd_sc_hd__buf_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1099_ _1866_/Q _1095_/X data_rdata_i[25] _1096_/X _1093_/X vssd1 vssd1 vccd1 vccd1
+ _1866_/D sky130_fd_sc_hd__o221a_2
X_1237_ _1690_/X vssd1 vssd1 vccd1 vccd1 _1238_/C sky130_fd_sc_hd__inv_2
X_1168_ _1757_/Q _1758_/Q _1530_/B vssd1 vssd1 vccd1 vccd1 _1540_/B sky130_fd_sc_hd__or3_2
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1022_ _1022_/A _1468_/B vssd1 vssd1 vccd1 vccd1 _1022_/Y sky130_fd_sc_hd__nor2_2
X_1855_ _1859_/CLK _1855_/D vssd1 vssd1 vccd1 vccd1 _1855_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1786_ _1835_/CLK _1786_/D vssd1 vssd1 vccd1 vccd1 _1786_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1346__A _1361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1571_ _1800_/Q _1637_/X _1777_/Q _1570_/X vssd1 vssd1 vccd1 vccd1 _1571_/X sky130_fd_sc_hd__a22o_2
X_1640_ _1571_/X _1468_/Y _1649_/S vssd1 vssd1 vccd1 vccd1 _1640_/X sky130_fd_sc_hd__mux2_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1005_ _1428_/C vssd1 vssd1 vccd1 vccd1 _1016_/B sky130_fd_sc_hd__inv_2
X_1838_ _1881_/CLK _1838_/D vssd1 vssd1 vccd1 vccd1 _1838_/Q sky130_fd_sc_hd__dfxtp_2
X_1907_ _1908_/CLK _1907_/D _0881_/X vssd1 vssd1 vccd1 vccd1 data_wdata_o[22] sky130_fd_sc_hd__dfrtp_2
X_1769_ _1888_/CLK _1769_/D vssd1 vssd1 vccd1 vccd1 _1769_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1623_ _1543_/A _1725_/S _1651_/X _1653_/X _1190_/A vssd1 vssd1 vccd1 vccd1 _1623_/X
+ sky130_fd_sc_hd__a32o_2
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1485_ _1485_/A vssd1 vssd1 vccd1 vccd1 _1485_/X sky130_fd_sc_hd__buf_1
X_1554_ _1566_/A _1554_/B vssd1 vssd1 vccd1 vccd1 _1555_/A sky130_fd_sc_hd__and2_2
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

