magic
tech sky130A
magscale 1 2
timestamp 1640351255
<< obsli1 >>
rect 1104 2159 29595 30481
<< obsm1 >>
rect 14 1300 29886 30592
<< metal2 >>
rect 662 31889 718 32689
rect 1950 31889 2006 32689
rect 3238 31889 3294 32689
rect 4618 31889 4674 32689
rect 5906 31889 5962 32689
rect 7286 31889 7342 32689
rect 8574 31889 8630 32689
rect 9954 31889 10010 32689
rect 11242 31889 11298 32689
rect 12530 31889 12586 32689
rect 13910 31889 13966 32689
rect 15198 31889 15254 32689
rect 16578 31889 16634 32689
rect 17866 31889 17922 32689
rect 19246 31889 19302 32689
rect 20534 31889 20590 32689
rect 21822 31889 21878 32689
rect 23202 31889 23258 32689
rect 24490 31889 24546 32689
rect 25870 31889 25926 32689
rect 27158 31889 27214 32689
rect 28538 31889 28594 32689
rect 29826 31889 29882 32689
rect 570 0 626 800
rect 1766 0 1822 800
rect 2962 0 3018 800
rect 4158 0 4214 800
rect 5446 0 5502 800
rect 6642 0 6698 800
rect 7838 0 7894 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 11518 0 11574 800
rect 12714 0 12770 800
rect 14002 0 14058 800
rect 15198 0 15254 800
rect 16394 0 16450 800
rect 17590 0 17646 800
rect 18878 0 18934 800
rect 20074 0 20130 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 23754 0 23810 800
rect 24950 0 25006 800
rect 26146 0 26202 800
rect 27434 0 27490 800
rect 28630 0 28686 800
rect 29826 0 29882 800
<< obsm2 >>
rect 20 31833 606 32065
rect 774 31833 1894 32065
rect 2062 31833 3182 32065
rect 3350 31833 4562 32065
rect 4730 31833 5850 32065
rect 6018 31833 7230 32065
rect 7398 31833 8518 32065
rect 8686 31833 9898 32065
rect 10066 31833 11186 32065
rect 11354 31833 12474 32065
rect 12642 31833 13854 32065
rect 14022 31833 15142 32065
rect 15310 31833 16522 32065
rect 16690 31833 17810 32065
rect 17978 31833 19190 32065
rect 19358 31833 20478 32065
rect 20646 31833 21766 32065
rect 21934 31833 23146 32065
rect 23314 31833 24434 32065
rect 24602 31833 25814 32065
rect 25982 31833 27102 32065
rect 27270 31833 28482 32065
rect 28650 31833 29770 32065
rect 20 856 29880 31833
rect 20 711 514 856
rect 682 711 1710 856
rect 1878 711 2906 856
rect 3074 711 4102 856
rect 4270 711 5390 856
rect 5558 711 6586 856
rect 6754 711 7782 856
rect 7950 711 8978 856
rect 9146 711 10266 856
rect 10434 711 11462 856
rect 11630 711 12658 856
rect 12826 711 13946 856
rect 14114 711 15142 856
rect 15310 711 16338 856
rect 16506 711 17534 856
rect 17702 711 18822 856
rect 18990 711 20018 856
rect 20186 711 21214 856
rect 21382 711 22502 856
rect 22670 711 23698 856
rect 23866 711 24894 856
rect 25062 711 26090 856
rect 26258 711 27378 856
rect 27546 711 28574 856
rect 28742 711 29770 856
<< metal3 >>
rect 0 31968 800 32088
rect 29745 31560 30545 31680
rect 0 30608 800 30728
rect 29745 29656 30545 29776
rect 0 29248 800 29368
rect 0 27888 800 28008
rect 29745 27752 30545 27872
rect 0 26528 800 26648
rect 29745 25848 30545 25968
rect 0 25168 800 25288
rect 0 23808 800 23928
rect 29745 23944 30545 24064
rect 0 22448 800 22568
rect 29745 22040 30545 22160
rect 0 21088 800 21208
rect 29745 20136 30545 20256
rect 0 19728 800 19848
rect 0 18368 800 18488
rect 29745 18232 30545 18352
rect 0 17008 800 17128
rect 29745 16192 30545 16312
rect 0 15648 800 15768
rect 0 14288 800 14408
rect 29745 14288 30545 14408
rect 0 12928 800 13048
rect 29745 12384 30545 12504
rect 0 11568 800 11688
rect 29745 10480 30545 10600
rect 0 10208 800 10328
rect 0 8848 800 8968
rect 29745 8576 30545 8696
rect 0 7488 800 7608
rect 29745 6672 30545 6792
rect 0 6128 800 6248
rect 0 4768 800 4888
rect 29745 4768 30545 4888
rect 0 3408 800 3528
rect 29745 2864 30545 2984
rect 0 2048 800 2168
rect 29745 960 30545 1080
rect 0 688 800 808
<< obsm3 >>
rect 880 31888 29745 32061
rect 800 31760 29745 31888
rect 800 31480 29665 31760
rect 800 30808 29745 31480
rect 880 30528 29745 30808
rect 800 29856 29745 30528
rect 800 29576 29665 29856
rect 800 29448 29745 29576
rect 880 29168 29745 29448
rect 800 28088 29745 29168
rect 880 27952 29745 28088
rect 880 27808 29665 27952
rect 800 27672 29665 27808
rect 800 26728 29745 27672
rect 880 26448 29745 26728
rect 800 26048 29745 26448
rect 800 25768 29665 26048
rect 800 25368 29745 25768
rect 880 25088 29745 25368
rect 800 24144 29745 25088
rect 800 24008 29665 24144
rect 880 23864 29665 24008
rect 880 23728 29745 23864
rect 800 22648 29745 23728
rect 880 22368 29745 22648
rect 800 22240 29745 22368
rect 800 21960 29665 22240
rect 800 21288 29745 21960
rect 880 21008 29745 21288
rect 800 20336 29745 21008
rect 800 20056 29665 20336
rect 800 19928 29745 20056
rect 880 19648 29745 19928
rect 800 18568 29745 19648
rect 880 18432 29745 18568
rect 880 18288 29665 18432
rect 800 18152 29665 18288
rect 800 17208 29745 18152
rect 880 16928 29745 17208
rect 800 16392 29745 16928
rect 800 16112 29665 16392
rect 800 15848 29745 16112
rect 880 15568 29745 15848
rect 800 14488 29745 15568
rect 880 14208 29665 14488
rect 800 13128 29745 14208
rect 880 12848 29745 13128
rect 800 12584 29745 12848
rect 800 12304 29665 12584
rect 800 11768 29745 12304
rect 880 11488 29745 11768
rect 800 10680 29745 11488
rect 800 10408 29665 10680
rect 880 10400 29665 10408
rect 880 10128 29745 10400
rect 800 9048 29745 10128
rect 880 8776 29745 9048
rect 880 8768 29665 8776
rect 800 8496 29665 8768
rect 800 7688 29745 8496
rect 880 7408 29745 7688
rect 800 6872 29745 7408
rect 800 6592 29665 6872
rect 800 6328 29745 6592
rect 880 6048 29745 6328
rect 800 4968 29745 6048
rect 880 4688 29665 4968
rect 800 3608 29745 4688
rect 880 3328 29745 3608
rect 800 3064 29745 3328
rect 800 2784 29665 3064
rect 800 2248 29745 2784
rect 880 1968 29745 2248
rect 800 1160 29745 1968
rect 800 888 29665 1160
rect 880 880 29665 888
rect 880 715 29745 880
<< metal4 >>
rect 5667 2128 5987 30512
rect 10389 2128 10709 30512
rect 15112 2128 15432 30512
rect 19834 2128 20154 30512
rect 24557 2128 24877 30512
<< obsm4 >>
rect 6067 2128 10309 30512
rect 10789 2128 15032 30512
rect 15512 2128 19754 30512
rect 20234 2128 20365 30512
<< labels >>
rlabel metal2 s 570 0 626 800 6 clk_i
port 1 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 data_addr_o[0]
port 2 nsew signal output
rlabel metal2 s 13910 31889 13966 32689 6 data_addr_o[10]
port 3 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 data_addr_o[11]
port 4 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 data_addr_o[1]
port 5 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 data_addr_o[2]
port 6 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 data_addr_o[3]
port 7 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 data_addr_o[4]
port 8 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 data_addr_o[5]
port 9 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 data_addr_o[6]
port 10 nsew signal output
rlabel metal3 s 29745 10480 30545 10600 6 data_addr_o[7]
port 11 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 data_addr_o[8]
port 12 nsew signal output
rlabel metal2 s 12530 31889 12586 32689 6 data_addr_o[9]
port 13 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 data_be_o[0]
port 14 nsew signal output
rlabel metal2 s 3238 31889 3294 32689 6 data_be_o[1]
port 15 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 data_be_o[2]
port 16 nsew signal output
rlabel metal2 s 4618 31889 4674 32689 6 data_be_o[3]
port 17 nsew signal output
rlabel metal2 s 662 31889 718 32689 6 data_gnt_i
port 18 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 data_rdata_i[0]
port 19 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 data_rdata_i[10]
port 20 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 data_rdata_i[11]
port 21 nsew signal input
rlabel metal3 s 29745 16192 30545 16312 6 data_rdata_i[12]
port 22 nsew signal input
rlabel metal3 s 29745 18232 30545 18352 6 data_rdata_i[13]
port 23 nsew signal input
rlabel metal2 s 16578 31889 16634 32689 6 data_rdata_i[14]
port 24 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 data_rdata_i[15]
port 25 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 data_rdata_i[16]
port 26 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 data_rdata_i[17]
port 27 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 data_rdata_i[18]
port 28 nsew signal input
rlabel metal2 s 20534 31889 20590 32689 6 data_rdata_i[19]
port 29 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 data_rdata_i[1]
port 30 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 data_rdata_i[20]
port 31 nsew signal input
rlabel metal3 s 29745 22040 30545 22160 6 data_rdata_i[21]
port 32 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 data_rdata_i[22]
port 33 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 data_rdata_i[23]
port 34 nsew signal input
rlabel metal2 s 25870 31889 25926 32689 6 data_rdata_i[24]
port 35 nsew signal input
rlabel metal3 s 29745 25848 30545 25968 6 data_rdata_i[25]
port 36 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 data_rdata_i[26]
port 37 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 data_rdata_i[27]
port 38 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 data_rdata_i[28]
port 39 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 data_rdata_i[29]
port 40 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 data_rdata_i[2]
port 41 nsew signal input
rlabel metal3 s 29745 29656 30545 29776 6 data_rdata_i[30]
port 42 nsew signal input
rlabel metal3 s 29745 31560 30545 31680 6 data_rdata_i[31]
port 43 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 data_rdata_i[3]
port 44 nsew signal input
rlabel metal2 s 5906 31889 5962 32689 6 data_rdata_i[4]
port 45 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 data_rdata_i[5]
port 46 nsew signal input
rlabel metal3 s 29745 8576 30545 8696 6 data_rdata_i[6]
port 47 nsew signal input
rlabel metal2 s 7286 31889 7342 32689 6 data_rdata_i[7]
port 48 nsew signal input
rlabel metal2 s 9954 31889 10010 32689 6 data_rdata_i[8]
port 49 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 data_rdata_i[9]
port 50 nsew signal input
rlabel metal3 s 0 688 800 808 6 data_req_o
port 51 nsew signal output
rlabel metal3 s 29745 960 30545 1080 6 data_rvalid_i
port 52 nsew signal input
rlabel metal3 s 29745 2864 30545 2984 6 data_wdata_o[0]
port 53 nsew signal output
rlabel metal3 s 29745 12384 30545 12504 6 data_wdata_o[10]
port 54 nsew signal output
rlabel metal3 s 29745 14288 30545 14408 6 data_wdata_o[11]
port 55 nsew signal output
rlabel metal2 s 15198 31889 15254 32689 6 data_wdata_o[12]
port 56 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 data_wdata_o[13]
port 57 nsew signal output
rlabel metal3 s 29745 20136 30545 20256 6 data_wdata_o[14]
port 58 nsew signal output
rlabel metal2 s 17866 31889 17922 32689 6 data_wdata_o[15]
port 59 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 data_wdata_o[16]
port 60 nsew signal output
rlabel metal2 s 19246 31889 19302 32689 6 data_wdata_o[17]
port 61 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 data_wdata_o[18]
port 62 nsew signal output
rlabel metal2 s 21822 31889 21878 32689 6 data_wdata_o[19]
port 63 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 data_wdata_o[1]
port 64 nsew signal output
rlabel metal2 s 23202 31889 23258 32689 6 data_wdata_o[20]
port 65 nsew signal output
rlabel metal2 s 24490 31889 24546 32689 6 data_wdata_o[21]
port 66 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 data_wdata_o[22]
port 67 nsew signal output
rlabel metal3 s 29745 23944 30545 24064 6 data_wdata_o[23]
port 68 nsew signal output
rlabel metal2 s 27158 31889 27214 32689 6 data_wdata_o[24]
port 69 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 data_wdata_o[25]
port 70 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 data_wdata_o[26]
port 71 nsew signal output
rlabel metal3 s 29745 27752 30545 27872 6 data_wdata_o[27]
port 72 nsew signal output
rlabel metal2 s 28538 31889 28594 32689 6 data_wdata_o[28]
port 73 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 data_wdata_o[29]
port 74 nsew signal output
rlabel metal3 s 29745 4768 30545 4888 6 data_wdata_o[2]
port 75 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 data_wdata_o[30]
port 76 nsew signal output
rlabel metal2 s 29826 31889 29882 32689 6 data_wdata_o[31]
port 77 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 data_wdata_o[3]
port 78 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 data_wdata_o[4]
port 79 nsew signal output
rlabel metal3 s 29745 6672 30545 6792 6 data_wdata_o[5]
port 80 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 data_wdata_o[6]
port 81 nsew signal output
rlabel metal2 s 8574 31889 8630 32689 6 data_wdata_o[7]
port 82 nsew signal output
rlabel metal2 s 11242 31889 11298 32689 6 data_wdata_o[8]
port 83 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 data_wdata_o[9]
port 84 nsew signal output
rlabel metal2 s 1950 31889 2006 32689 6 data_we_o
port 85 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 rst_i
port 86 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 rx_i
port 87 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 tx_o
port 88 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 uart_error
port 89 nsew signal output
rlabel metal4 s 5667 2128 5987 30512 6 vccd1
port 90 nsew power input
rlabel metal4 s 15112 2128 15432 30512 6 vccd1
port 90 nsew power input
rlabel metal4 s 24557 2128 24877 30512 6 vccd1
port 90 nsew power input
rlabel metal4 s 10389 2128 10709 30512 6 vssd1
port 91 nsew ground input
rlabel metal4 s 19834 2128 20154 30512 6 vssd1
port 91 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 30545 32689
string LEFview TRUE
string GDS_FILE /project/openlane/uart_to_mem/runs/uart_to_mem/results/magic/uart_to_mem.gds
string GDS_END 2948858
string GDS_START 388486
<< end >>

