magic
tech sky130A
magscale 1 2
timestamp 1640350731
<< obsli1 >>
rect 1104 2159 26283 28475
<< obsm1 >>
rect 566 1300 26298 28484
<< metal2 >>
rect 570 28642 626 29442
rect 1674 28642 1730 29442
rect 2870 28642 2926 29442
rect 4066 28642 4122 29442
rect 5262 28642 5318 29442
rect 6458 28642 6514 29442
rect 7654 28642 7710 29442
rect 8850 28642 8906 29442
rect 10046 28642 10102 29442
rect 11242 28642 11298 29442
rect 12438 28642 12494 29442
rect 13634 28642 13690 29442
rect 14738 28642 14794 29442
rect 15934 28642 15990 29442
rect 17130 28642 17186 29442
rect 18326 28642 18382 29442
rect 19522 28642 19578 29442
rect 20718 28642 20774 29442
rect 21914 28642 21970 29442
rect 23110 28642 23166 29442
rect 24306 28642 24362 29442
rect 25502 28642 25558 29442
rect 26698 28642 26754 29442
rect 570 0 626 800
rect 1674 0 1730 800
rect 2870 0 2926 800
rect 4066 0 4122 800
rect 5262 0 5318 800
rect 6458 0 6514 800
rect 7654 0 7710 800
rect 8850 0 8906 800
rect 10046 0 10102 800
rect 11242 0 11298 800
rect 12438 0 12494 800
rect 13634 0 13690 800
rect 14738 0 14794 800
rect 15934 0 15990 800
rect 17130 0 17186 800
rect 18326 0 18382 800
rect 19522 0 19578 800
rect 20718 0 20774 800
rect 21914 0 21970 800
rect 23110 0 23166 800
rect 24306 0 24362 800
rect 25502 0 25558 800
rect 26698 0 26754 800
<< obsm2 >>
rect 682 28586 1618 28778
rect 1786 28586 2814 28778
rect 2982 28586 4010 28778
rect 4178 28586 5206 28778
rect 5374 28586 6402 28778
rect 6570 28586 7598 28778
rect 7766 28586 8794 28778
rect 8962 28586 9990 28778
rect 10158 28586 11186 28778
rect 11354 28586 12382 28778
rect 12550 28586 13578 28778
rect 13746 28586 14682 28778
rect 14850 28586 15878 28778
rect 16046 28586 17074 28778
rect 17242 28586 18270 28778
rect 18438 28586 19466 28778
rect 19634 28586 20662 28778
rect 20830 28586 21858 28778
rect 22026 28586 23054 28778
rect 23222 28586 24250 28778
rect 24418 28586 25446 28778
rect 25614 28586 26294 28778
rect 572 856 26294 28586
rect 682 711 1618 856
rect 1786 711 2814 856
rect 2982 711 4010 856
rect 4178 711 5206 856
rect 5374 711 6402 856
rect 6570 711 7598 856
rect 7766 711 8794 856
rect 8962 711 9990 856
rect 10158 711 11186 856
rect 11354 711 12382 856
rect 12550 711 13578 856
rect 13746 711 14682 856
rect 14850 711 15878 856
rect 16046 711 17074 856
rect 17242 711 18270 856
rect 18438 711 19466 856
rect 19634 711 20662 856
rect 20830 711 21858 856
rect 22026 711 23054 856
rect 23222 711 24250 856
rect 24418 711 25446 856
rect 25614 711 26294 856
<< metal3 >>
rect 0 28568 800 28688
rect 26498 28432 27298 28552
rect 0 27208 800 27328
rect 26498 26936 27298 27056
rect 0 25848 800 25968
rect 26498 25304 27298 25424
rect 0 24352 800 24472
rect 26498 23808 27298 23928
rect 0 22992 800 23112
rect 26498 22312 27298 22432
rect 0 21632 800 21752
rect 26498 20680 27298 20800
rect 0 20272 800 20392
rect 26498 19184 27298 19304
rect 0 18776 800 18896
rect 26498 17688 27298 17808
rect 0 17416 800 17536
rect 0 16056 800 16176
rect 26498 16056 27298 16176
rect 0 14560 800 14680
rect 26498 14560 27298 14680
rect 0 13200 800 13320
rect 26498 12928 27298 13048
rect 0 11840 800 11960
rect 26498 11432 27298 11552
rect 0 10480 800 10600
rect 26498 9936 27298 10056
rect 0 8984 800 9104
rect 26498 8304 27298 8424
rect 0 7624 800 7744
rect 26498 6808 27298 6928
rect 0 6264 800 6384
rect 26498 5312 27298 5432
rect 0 4768 800 4888
rect 26498 3680 27298 3800
rect 0 3408 800 3528
rect 0 2048 800 2168
rect 26498 2184 27298 2304
rect 0 688 800 808
rect 26498 688 27298 808
<< obsm3 >>
rect 880 28488 26418 28525
rect 800 28352 26418 28488
rect 800 27408 26498 28352
rect 880 27136 26498 27408
rect 880 27128 26418 27136
rect 800 26856 26418 27128
rect 800 26048 26498 26856
rect 880 25768 26498 26048
rect 800 25504 26498 25768
rect 800 25224 26418 25504
rect 800 24552 26498 25224
rect 880 24272 26498 24552
rect 800 24008 26498 24272
rect 800 23728 26418 24008
rect 800 23192 26498 23728
rect 880 22912 26498 23192
rect 800 22512 26498 22912
rect 800 22232 26418 22512
rect 800 21832 26498 22232
rect 880 21552 26498 21832
rect 800 20880 26498 21552
rect 800 20600 26418 20880
rect 800 20472 26498 20600
rect 880 20192 26498 20472
rect 800 19384 26498 20192
rect 800 19104 26418 19384
rect 800 18976 26498 19104
rect 880 18696 26498 18976
rect 800 17888 26498 18696
rect 800 17616 26418 17888
rect 880 17608 26418 17616
rect 880 17336 26498 17608
rect 800 16256 26498 17336
rect 880 15976 26418 16256
rect 800 14760 26498 15976
rect 880 14480 26418 14760
rect 800 13400 26498 14480
rect 880 13128 26498 13400
rect 880 13120 26418 13128
rect 800 12848 26418 13120
rect 800 12040 26498 12848
rect 880 11760 26498 12040
rect 800 11632 26498 11760
rect 800 11352 26418 11632
rect 800 10680 26498 11352
rect 880 10400 26498 10680
rect 800 10136 26498 10400
rect 800 9856 26418 10136
rect 800 9184 26498 9856
rect 880 8904 26498 9184
rect 800 8504 26498 8904
rect 800 8224 26418 8504
rect 800 7824 26498 8224
rect 880 7544 26498 7824
rect 800 7008 26498 7544
rect 800 6728 26418 7008
rect 800 6464 26498 6728
rect 880 6184 26498 6464
rect 800 5512 26498 6184
rect 800 5232 26418 5512
rect 800 4968 26498 5232
rect 880 4688 26498 4968
rect 800 3880 26498 4688
rect 800 3608 26418 3880
rect 880 3600 26418 3608
rect 880 3328 26498 3600
rect 800 2384 26498 3328
rect 800 2248 26418 2384
rect 880 2104 26418 2248
rect 880 1968 26498 2104
rect 800 888 26498 1968
rect 880 715 26418 888
<< metal4 >>
rect 5115 2128 5435 27248
rect 9285 2128 9605 27248
rect 13456 2128 13776 27248
rect 17626 2128 17946 27248
rect 21797 2128 22117 27248
<< labels >>
rlabel metal3 s 0 688 800 808 6 clk
port 1 nsew signal input
rlabel metal2 s 570 28642 626 29442 6 data_req_i
port 2 nsew signal input
rlabel metal2 s 570 0 626 800 6 reset
port 3 nsew signal input
rlabel metal3 s 26498 688 27298 808 6 rxd_uart
port 4 nsew signal input
rlabel metal2 s 1674 28642 1730 29442 6 slave_data_addr_i[0]
port 5 nsew signal input
rlabel metal2 s 4066 28642 4122 29442 6 slave_data_addr_i[1]
port 6 nsew signal input
rlabel metal3 s 26498 8304 27298 8424 6 slave_data_addr_i[2]
port 7 nsew signal input
rlabel metal2 s 8850 28642 8906 29442 6 slave_data_addr_i[3]
port 8 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 slave_data_addr_i[4]
port 9 nsew signal input
rlabel metal3 s 26498 11432 27298 11552 6 slave_data_addr_i[5]
port 10 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 slave_data_addr_i[6]
port 11 nsew signal input
rlabel metal3 s 26498 12928 27298 13048 6 slave_data_addr_i[7]
port 12 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 slave_data_addr_i[8]
port 13 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 slave_data_addr_i[9]
port 14 nsew signal input
rlabel metal3 s 26498 5312 27298 5432 6 slave_data_be_i[0]
port 15 nsew signal input
rlabel metal3 s 26498 6808 27298 6928 6 slave_data_be_i[1]
port 16 nsew signal input
rlabel metal2 s 5262 28642 5318 29442 6 slave_data_be_i[2]
port 17 nsew signal input
rlabel metal2 s 10046 28642 10102 29442 6 slave_data_be_i[3]
port 18 nsew signal input
rlabel metal3 s 26498 2184 27298 2304 6 slave_data_gnt_o
port 19 nsew signal output
rlabel metal2 s 2870 28642 2926 29442 6 slave_data_rdata_o[0]
port 20 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 slave_data_rdata_o[10]
port 21 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 slave_data_rdata_o[11]
port 22 nsew signal output
rlabel metal3 s 26498 16056 27298 16176 6 slave_data_rdata_o[12]
port 23 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 slave_data_rdata_o[13]
port 24 nsew signal output
rlabel metal3 s 26498 17688 27298 17808 6 slave_data_rdata_o[14]
port 25 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 slave_data_rdata_o[15]
port 26 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 slave_data_rdata_o[16]
port 27 nsew signal output
rlabel metal2 s 17130 28642 17186 29442 6 slave_data_rdata_o[17]
port 28 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 slave_data_rdata_o[18]
port 29 nsew signal output
rlabel metal3 s 0 21632 800 21752 6 slave_data_rdata_o[19]
port 30 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 slave_data_rdata_o[1]
port 31 nsew signal output
rlabel metal2 s 18326 28642 18382 29442 6 slave_data_rdata_o[20]
port 32 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 slave_data_rdata_o[21]
port 33 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 slave_data_rdata_o[22]
port 34 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 slave_data_rdata_o[23]
port 35 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 slave_data_rdata_o[24]
port 36 nsew signal output
rlabel metal3 s 26498 25304 27298 25424 6 slave_data_rdata_o[25]
port 37 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 slave_data_rdata_o[26]
port 38 nsew signal output
rlabel metal2 s 21914 28642 21970 29442 6 slave_data_rdata_o[27]
port 39 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 slave_data_rdata_o[28]
port 40 nsew signal output
rlabel metal2 s 23110 28642 23166 29442 6 slave_data_rdata_o[29]
port 41 nsew signal output
rlabel metal2 s 6458 28642 6514 29442 6 slave_data_rdata_o[2]
port 42 nsew signal output
rlabel metal2 s 25502 28642 25558 29442 6 slave_data_rdata_o[30]
port 43 nsew signal output
rlabel metal3 s 26498 28432 27298 28552 6 slave_data_rdata_o[31]
port 44 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 slave_data_rdata_o[3]
port 45 nsew signal output
rlabel metal2 s 11242 28642 11298 29442 6 slave_data_rdata_o[4]
port 46 nsew signal output
rlabel metal2 s 12438 28642 12494 29442 6 slave_data_rdata_o[5]
port 47 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 slave_data_rdata_o[6]
port 48 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 slave_data_rdata_o[7]
port 49 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 slave_data_rdata_o[8]
port 50 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 slave_data_rdata_o[9]
port 51 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 slave_data_rvalid_o
port 52 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 slave_data_wdata_i[0]
port 53 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 slave_data_wdata_i[10]
port 54 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 slave_data_wdata_i[11]
port 55 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 slave_data_wdata_i[12]
port 56 nsew signal input
rlabel metal2 s 14738 28642 14794 29442 6 slave_data_wdata_i[13]
port 57 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 slave_data_wdata_i[14]
port 58 nsew signal input
rlabel metal2 s 15934 28642 15990 29442 6 slave_data_wdata_i[15]
port 59 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 slave_data_wdata_i[16]
port 60 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 slave_data_wdata_i[17]
port 61 nsew signal input
rlabel metal3 s 26498 19184 27298 19304 6 slave_data_wdata_i[18]
port 62 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 slave_data_wdata_i[19]
port 63 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 slave_data_wdata_i[1]
port 64 nsew signal input
rlabel metal2 s 19522 28642 19578 29442 6 slave_data_wdata_i[20]
port 65 nsew signal input
rlabel metal2 s 20718 28642 20774 29442 6 slave_data_wdata_i[21]
port 66 nsew signal input
rlabel metal3 s 26498 20680 27298 20800 6 slave_data_wdata_i[22]
port 67 nsew signal input
rlabel metal3 s 26498 22312 27298 22432 6 slave_data_wdata_i[23]
port 68 nsew signal input
rlabel metal3 s 26498 23808 27298 23928 6 slave_data_wdata_i[24]
port 69 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 slave_data_wdata_i[25]
port 70 nsew signal input
rlabel metal3 s 26498 26936 27298 27056 6 slave_data_wdata_i[26]
port 71 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 slave_data_wdata_i[27]
port 72 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 slave_data_wdata_i[28]
port 73 nsew signal input
rlabel metal2 s 24306 28642 24362 29442 6 slave_data_wdata_i[29]
port 74 nsew signal input
rlabel metal2 s 7654 28642 7710 29442 6 slave_data_wdata_i[2]
port 75 nsew signal input
rlabel metal2 s 26698 28642 26754 29442 6 slave_data_wdata_i[30]
port 76 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 slave_data_wdata_i[31]
port 77 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 slave_data_wdata_i[3]
port 78 nsew signal input
rlabel metal3 s 26498 9936 27298 10056 6 slave_data_wdata_i[4]
port 79 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 slave_data_wdata_i[5]
port 80 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 slave_data_wdata_i[6]
port 81 nsew signal input
rlabel metal2 s 13634 28642 13690 29442 6 slave_data_wdata_i[7]
port 82 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 slave_data_wdata_i[8]
port 83 nsew signal input
rlabel metal3 s 26498 14560 27298 14680 6 slave_data_wdata_i[9]
port 84 nsew signal input
rlabel metal3 s 26498 3680 27298 3800 6 slave_data_we_i
port 85 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 txd_uart
port 86 nsew signal output
rlabel metal4 s 5115 2128 5435 27248 6 vccd1
port 87 nsew power input
rlabel metal4 s 13456 2128 13776 27248 6 vccd1
port 87 nsew power input
rlabel metal4 s 21797 2128 22117 27248 6 vccd1
port 87 nsew power input
rlabel metal4 s 9285 2128 9605 27248 6 vssd1
port 88 nsew ground input
rlabel metal4 s 17626 2128 17946 27248 6 vssd1
port 88 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 27298 29442
string LEFview TRUE
string GDS_FILE /project/openlane/peripheral/runs/peripheral/results/magic/peripheral.gds
string GDS_END 2284808
string GDS_START 241546
<< end >>

