magic
tech sky130A
magscale 1 2
timestamp 1640734602
<< obsli1 >>
rect 1104 2159 29687 30481
<< obsm1 >>
rect 566 1300 30070 30728
<< metal2 >>
rect 570 32056 626 32856
rect 1766 32056 1822 32856
rect 2962 32056 3018 32856
rect 4250 32056 4306 32856
rect 5446 32056 5502 32856
rect 6642 32056 6698 32856
rect 7930 32056 7986 32856
rect 9126 32056 9182 32856
rect 10322 32056 10378 32856
rect 11610 32056 11666 32856
rect 12806 32056 12862 32856
rect 14002 32056 14058 32856
rect 15290 32056 15346 32856
rect 16486 32056 16542 32856
rect 17774 32056 17830 32856
rect 18970 32056 19026 32856
rect 20166 32056 20222 32856
rect 21454 32056 21510 32856
rect 22650 32056 22706 32856
rect 23846 32056 23902 32856
rect 25134 32056 25190 32856
rect 26330 32056 26386 32856
rect 27526 32056 27582 32856
rect 28814 32056 28870 32856
rect 30010 32056 30066 32856
rect 846 0 902 800
rect 2502 0 2558 800
rect 4250 0 4306 800
rect 5906 0 5962 800
rect 7654 0 7710 800
rect 9310 0 9366 800
rect 11058 0 11114 800
rect 12714 0 12770 800
rect 14462 0 14518 800
rect 16210 0 16266 800
rect 17866 0 17922 800
rect 19614 0 19670 800
rect 21270 0 21326 800
rect 23018 0 23074 800
rect 24674 0 24730 800
rect 26422 0 26478 800
rect 28078 0 28134 800
rect 29826 0 29882 800
<< obsm2 >>
rect 682 32000 1710 32201
rect 1878 32000 2906 32201
rect 3074 32000 4194 32201
rect 4362 32000 5390 32201
rect 5558 32000 6586 32201
rect 6754 32000 7874 32201
rect 8042 32000 9070 32201
rect 9238 32000 10266 32201
rect 10434 32000 11554 32201
rect 11722 32000 12750 32201
rect 12918 32000 13946 32201
rect 14114 32000 15234 32201
rect 15402 32000 16430 32201
rect 16598 32000 17718 32201
rect 17886 32000 18914 32201
rect 19082 32000 20110 32201
rect 20278 32000 21398 32201
rect 21566 32000 22594 32201
rect 22762 32000 23790 32201
rect 23958 32000 25078 32201
rect 25246 32000 26274 32201
rect 26442 32000 27470 32201
rect 27638 32000 28758 32201
rect 28926 32000 29954 32201
rect 572 856 30064 32000
rect 572 711 790 856
rect 958 711 2446 856
rect 2614 711 4194 856
rect 4362 711 5850 856
rect 6018 711 7598 856
rect 7766 711 9254 856
rect 9422 711 11002 856
rect 11170 711 12658 856
rect 12826 711 14406 856
rect 14574 711 16154 856
rect 16322 711 17810 856
rect 17978 711 19558 856
rect 19726 711 21214 856
rect 21382 711 22962 856
rect 23130 711 24618 856
rect 24786 711 26366 856
rect 26534 711 28022 856
rect 28190 711 29770 856
rect 29938 711 30064 856
<< metal3 >>
rect 0 32104 800 32224
rect 29912 32104 30712 32224
rect 0 30744 800 30864
rect 29912 30608 30712 30728
rect 0 29384 800 29504
rect 29912 29112 30712 29232
rect 0 28024 800 28144
rect 29912 27616 30712 27736
rect 0 26664 800 26784
rect 29912 26120 30712 26240
rect 0 25304 800 25424
rect 29912 24624 30712 24744
rect 0 23944 800 24064
rect 29912 23128 30712 23248
rect 0 22584 800 22704
rect 29912 21632 30712 21752
rect 0 21224 800 21344
rect 29912 20136 30712 20256
rect 0 19864 800 19984
rect 0 18504 800 18624
rect 29912 18640 30712 18760
rect 0 17144 800 17264
rect 29912 17144 30712 17264
rect 0 15648 800 15768
rect 29912 15648 30712 15768
rect 0 14288 800 14408
rect 29912 14152 30712 14272
rect 0 12928 800 13048
rect 29912 12656 30712 12776
rect 0 11568 800 11688
rect 29912 11160 30712 11280
rect 0 10208 800 10328
rect 29912 9664 30712 9784
rect 0 8848 800 8968
rect 29912 8168 30712 8288
rect 0 7488 800 7608
rect 29912 6672 30712 6792
rect 0 6128 800 6248
rect 29912 5176 30712 5296
rect 0 4768 800 4888
rect 29912 3680 30712 3800
rect 0 3408 800 3528
rect 0 2048 800 2168
rect 29912 2184 30712 2304
rect 0 688 800 808
rect 29912 688 30712 808
<< obsm3 >>
rect 880 32024 29832 32197
rect 800 30944 29912 32024
rect 880 30808 29912 30944
rect 880 30664 29832 30808
rect 800 30528 29832 30664
rect 800 29584 29912 30528
rect 880 29312 29912 29584
rect 880 29304 29832 29312
rect 800 29032 29832 29304
rect 800 28224 29912 29032
rect 880 27944 29912 28224
rect 800 27816 29912 27944
rect 800 27536 29832 27816
rect 800 26864 29912 27536
rect 880 26584 29912 26864
rect 800 26320 29912 26584
rect 800 26040 29832 26320
rect 800 25504 29912 26040
rect 880 25224 29912 25504
rect 800 24824 29912 25224
rect 800 24544 29832 24824
rect 800 24144 29912 24544
rect 880 23864 29912 24144
rect 800 23328 29912 23864
rect 800 23048 29832 23328
rect 800 22784 29912 23048
rect 880 22504 29912 22784
rect 800 21832 29912 22504
rect 800 21552 29832 21832
rect 800 21424 29912 21552
rect 880 21144 29912 21424
rect 800 20336 29912 21144
rect 800 20064 29832 20336
rect 880 20056 29832 20064
rect 880 19784 29912 20056
rect 800 18840 29912 19784
rect 800 18704 29832 18840
rect 880 18560 29832 18704
rect 880 18424 29912 18560
rect 800 17344 29912 18424
rect 880 17064 29832 17344
rect 800 15848 29912 17064
rect 880 15568 29832 15848
rect 800 14488 29912 15568
rect 880 14352 29912 14488
rect 880 14208 29832 14352
rect 800 14072 29832 14208
rect 800 13128 29912 14072
rect 880 12856 29912 13128
rect 880 12848 29832 12856
rect 800 12576 29832 12848
rect 800 11768 29912 12576
rect 880 11488 29912 11768
rect 800 11360 29912 11488
rect 800 11080 29832 11360
rect 800 10408 29912 11080
rect 880 10128 29912 10408
rect 800 9864 29912 10128
rect 800 9584 29832 9864
rect 800 9048 29912 9584
rect 880 8768 29912 9048
rect 800 8368 29912 8768
rect 800 8088 29832 8368
rect 800 7688 29912 8088
rect 880 7408 29912 7688
rect 800 6872 29912 7408
rect 800 6592 29832 6872
rect 800 6328 29912 6592
rect 880 6048 29912 6328
rect 800 5376 29912 6048
rect 800 5096 29832 5376
rect 800 4968 29912 5096
rect 880 4688 29912 4968
rect 800 3880 29912 4688
rect 800 3608 29832 3880
rect 880 3600 29832 3608
rect 880 3328 29912 3600
rect 800 2384 29912 3328
rect 800 2248 29832 2384
rect 880 2104 29832 2248
rect 880 1968 29912 2104
rect 800 888 29912 1968
rect 880 715 29832 888
<< metal4 >>
rect 5681 2128 6001 30512
rect 10419 2128 10739 30512
rect 15157 2128 15477 30512
rect 19895 2128 20215 30512
rect 24633 2128 24953 30512
<< obsm4 >>
rect 6081 2128 10339 30512
rect 10819 2128 15077 30512
rect 15557 2128 19815 30512
rect 20295 2128 20549 30512
<< labels >>
rlabel metal3 s 29912 688 30712 808 6 clk_i
port 1 nsew signal input
rlabel metal2 s 1766 32056 1822 32856 6 data_addr_o[0]
port 2 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 data_addr_o[10]
port 3 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 data_addr_o[11]
port 4 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 data_addr_o[1]
port 5 nsew signal output
rlabel metal3 s 29912 5176 30712 5296 6 data_addr_o[2]
port 6 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 data_addr_o[3]
port 7 nsew signal output
rlabel metal2 s 7930 32056 7986 32856 6 data_addr_o[4]
port 8 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 data_addr_o[5]
port 9 nsew signal output
rlabel metal2 s 9126 32056 9182 32856 6 data_addr_o[6]
port 10 nsew signal output
rlabel metal2 s 10322 32056 10378 32856 6 data_addr_o[7]
port 11 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 data_addr_o[8]
port 12 nsew signal output
rlabel metal3 s 29912 17144 30712 17264 6 data_addr_o[9]
port 13 nsew signal output
rlabel metal2 s 2962 32056 3018 32856 6 data_be_o[0]
port 14 nsew signal output
rlabel metal2 s 4250 32056 4306 32856 6 data_be_o[1]
port 15 nsew signal output
rlabel metal2 s 6642 32056 6698 32856 6 data_be_o[2]
port 16 nsew signal output
rlabel metal3 s 29912 8168 30712 8288 6 data_be_o[3]
port 17 nsew signal output
rlabel metal2 s 846 0 902 800 6 data_gnt_i
port 18 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 data_rdata_i[0]
port 19 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 data_rdata_i[10]
port 20 nsew signal input
rlabel metal2 s 14002 32056 14058 32856 6 data_rdata_i[11]
port 21 nsew signal input
rlabel metal2 s 15290 32056 15346 32856 6 data_rdata_i[12]
port 22 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 data_rdata_i[13]
port 23 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 data_rdata_i[14]
port 24 nsew signal input
rlabel metal3 s 29912 23128 30712 23248 6 data_rdata_i[15]
port 25 nsew signal input
rlabel metal2 s 16486 32056 16542 32856 6 data_rdata_i[16]
port 26 nsew signal input
rlabel metal2 s 17774 32056 17830 32856 6 data_rdata_i[17]
port 27 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 data_rdata_i[18]
port 28 nsew signal input
rlabel metal3 s 29912 27616 30712 27736 6 data_rdata_i[19]
port 29 nsew signal input
rlabel metal2 s 5446 32056 5502 32856 6 data_rdata_i[1]
port 30 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 data_rdata_i[20]
port 31 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 data_rdata_i[21]
port 32 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 data_rdata_i[22]
port 33 nsew signal input
rlabel metal2 s 21454 32056 21510 32856 6 data_rdata_i[23]
port 34 nsew signal input
rlabel metal3 s 29912 29112 30712 29232 6 data_rdata_i[24]
port 35 nsew signal input
rlabel metal2 s 23846 32056 23902 32856 6 data_rdata_i[25]
port 36 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 data_rdata_i[26]
port 37 nsew signal input
rlabel metal2 s 26330 32056 26386 32856 6 data_rdata_i[27]
port 38 nsew signal input
rlabel metal2 s 27526 32056 27582 32856 6 data_rdata_i[28]
port 39 nsew signal input
rlabel metal2 s 28814 32056 28870 32856 6 data_rdata_i[29]
port 40 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 data_rdata_i[2]
port 41 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 data_rdata_i[30]
port 42 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 data_rdata_i[31]
port 43 nsew signal input
rlabel metal3 s 29912 9664 30712 9784 6 data_rdata_i[3]
port 44 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 data_rdata_i[4]
port 45 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 data_rdata_i[5]
port 46 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 data_rdata_i[6]
port 47 nsew signal input
rlabel metal3 s 29912 15648 30712 15768 6 data_rdata_i[7]
port 48 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 data_rdata_i[8]
port 49 nsew signal input
rlabel metal3 s 29912 18640 30712 18760 6 data_rdata_i[9]
port 50 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 data_req_o
port 51 nsew signal output
rlabel metal3 s 0 688 800 808 6 data_rvalid_i
port 52 nsew signal input
rlabel metal3 s 29912 3680 30712 3800 6 data_wdata_o[0]
port 53 nsew signal output
rlabel metal2 s 12806 32056 12862 32856 6 data_wdata_o[10]
port 54 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 data_wdata_o[11]
port 55 nsew signal output
rlabel metal3 s 29912 21632 30712 21752 6 data_wdata_o[12]
port 56 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 data_wdata_o[13]
port 57 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 data_wdata_o[14]
port 58 nsew signal output
rlabel metal3 s 29912 24624 30712 24744 6 data_wdata_o[15]
port 59 nsew signal output
rlabel metal3 s 29912 26120 30712 26240 6 data_wdata_o[16]
port 60 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 data_wdata_o[17]
port 61 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 data_wdata_o[18]
port 62 nsew signal output
rlabel metal2 s 18970 32056 19026 32856 6 data_wdata_o[19]
port 63 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 data_wdata_o[1]
port 64 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 data_wdata_o[20]
port 65 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 data_wdata_o[21]
port 66 nsew signal output
rlabel metal2 s 20166 32056 20222 32856 6 data_wdata_o[22]
port 67 nsew signal output
rlabel metal2 s 22650 32056 22706 32856 6 data_wdata_o[23]
port 68 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 data_wdata_o[24]
port 69 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 data_wdata_o[25]
port 70 nsew signal output
rlabel metal2 s 25134 32056 25190 32856 6 data_wdata_o[26]
port 71 nsew signal output
rlabel metal3 s 29912 30608 30712 30728 6 data_wdata_o[27]
port 72 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 data_wdata_o[28]
port 73 nsew signal output
rlabel metal2 s 30010 32056 30066 32856 6 data_wdata_o[29]
port 74 nsew signal output
rlabel metal3 s 29912 6672 30712 6792 6 data_wdata_o[2]
port 75 nsew signal output
rlabel metal3 s 29912 32104 30712 32224 6 data_wdata_o[30]
port 76 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 data_wdata_o[31]
port 77 nsew signal output
rlabel metal3 s 29912 11160 30712 11280 6 data_wdata_o[3]
port 78 nsew signal output
rlabel metal3 s 29912 12656 30712 12776 6 data_wdata_o[4]
port 79 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 data_wdata_o[5]
port 80 nsew signal output
rlabel metal3 s 29912 14152 30712 14272 6 data_wdata_o[6]
port 81 nsew signal output
rlabel metal2 s 11610 32056 11666 32856 6 data_wdata_o[7]
port 82 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 data_wdata_o[8]
port 83 nsew signal output
rlabel metal3 s 29912 20136 30712 20256 6 data_wdata_o[9]
port 84 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 data_we_o
port 85 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 rst_i
port 86 nsew signal input
rlabel metal3 s 29912 2184 30712 2304 6 rx_i
port 87 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 tx_o
port 88 nsew signal output
rlabel metal2 s 570 32056 626 32856 6 uart_error
port 89 nsew signal output
rlabel metal4 s 5681 2128 6001 30512 6 vccd1
port 90 nsew power input
rlabel metal4 s 15157 2128 15477 30512 6 vccd1
port 90 nsew power input
rlabel metal4 s 24633 2128 24953 30512 6 vccd1
port 90 nsew power input
rlabel metal4 s 10419 2128 10739 30512 6 vssd1
port 91 nsew ground input
rlabel metal4 s 19895 2128 20215 30512 6 vssd1
port 91 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 30712 32856
string LEFview TRUE
string GDS_FILE /project/openlane/uart_to_mem/runs/uart_to_mem/results/magic/uart_to_mem.gds
string GDS_END 2941210
string GDS_START 389658
<< end >>

