VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO soric_soc
  CLASS BLOCK ;
  FOREIGN soric_soc ;
  ORIGIN 0.000 0.000 ;
  SIZE 1700.000 BY 300.000 ;
  PIN error_uart_to_mem
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 24.520 1700.000 25.120 ;
    END
  END error_uart_to_mem
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 0.000 1058.830 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.470 0.000 1197.750 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.110 296.000 1627.390 300.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 96.600 1700.000 97.200 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 0.000 1227.650 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 0.000 1257.550 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.050 0.000 1277.330 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.830 0.000 1297.110 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.330 0.000 1078.610 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 129.920 1700.000 130.520 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.630 0.000 1356.910 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 136.040 1700.000 136.640 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.410 0.000 1376.690 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.130 296.000 1644.410 300.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.970 296.000 1646.250 300.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.430 0.000 1416.710 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.110 296.000 1650.390 300.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 0.000 1436.490 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.410 296.000 1652.690 300.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 157.800 1700.000 158.400 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 169.360 1700.000 169.960 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 52.400 1700.000 53.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 57.840 1700.000 58.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 63.280 1700.000 63.880 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 69.400 1700.000 70.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.790 0.000 1148.070 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 80.280 1700.000 80.880 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1624.810 296.000 1625.090 300.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 29.960 1700.000 30.560 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 0.000 1188.090 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.490 0.000 1237.770 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 108.160 1700.000 108.760 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.170 0.000 1287.450 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 119.040 1700.000 119.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 36.080 1700.000 36.680 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 124.480 1700.000 125.080 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.550 296.000 1633.830 300.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.390 296.000 1635.670 300.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.530 296.000 1639.810 300.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.750 0.000 1367.030 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 141.480 1700.000 142.080 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.530 0.000 1386.810 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.190 0.000 1396.470 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 46.960 1700.000 47.560 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.090 0.000 1426.370 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 152.360 1700.000 152.960 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.250 296.000 1654.530 300.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.550 296.000 1656.830 300.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 0.000 1456.270 4.000 ;
    END
  END io_out[35]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.230 0.000 1108.510 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 0.000 1128.290 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 296.000 1623.250 300.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 85.720 1700.000 86.320 ;
    END
  END io_out[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.210 0.000 1068.490 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.050 0.000 1645.330 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 263.200 1700.000 263.800 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.990 296.000 1686.270 300.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.290 296.000 1688.570 300.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.590 296.000 1690.870 300.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.710 0.000 1654.990 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.830 0.000 1665.110 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 269.320 1700.000 269.920 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.950 0.000 1675.230 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 274.760 1700.000 275.360 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 280.200 1700.000 280.800 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.430 296.000 1692.710 300.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.610 0.000 1684.890 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.730 0.000 1695.010 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 91.160 1700.000 91.760 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 285.640 1700.000 286.240 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.730 296.000 1695.010 300.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 291.080 1700.000 291.680 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 296.520 1700.000 297.120 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.570 296.000 1696.850 300.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.870 296.000 1699.150 300.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 0.000 1217.530 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 102.720 1700.000 103.320 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.950 296.000 1629.230 300.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1631.250 296.000 1631.530 300.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.150 0.000 1247.430 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 0.000 1267.210 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 113.600 1700.000 114.200 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.950 0.000 1307.230 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 41.520 1700.000 42.120 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.850 0.000 1337.130 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.510 0.000 1346.790 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1637.690 296.000 1637.970 300.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.830 296.000 1642.110 300.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 146.920 1700.000 147.520 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.310 0.000 1406.590 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.270 296.000 1648.550 300.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 0.000 1446.610 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 296.000 1659.130 300.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 163.240 1700.000 163.840 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 174.800 1700.000 175.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.110 0.000 1466.390 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.770 0.000 1476.050 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.690 296.000 1660.970 300.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.890 0.000 1486.170 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 180.240 1700.000 180.840 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.010 0.000 1496.290 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.890 0.000 1118.170 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 185.680 1700.000 186.280 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.990 296.000 1663.270 300.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.830 296.000 1665.110 300.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 191.120 1700.000 191.720 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.130 296.000 1667.410 300.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1505.670 0.000 1505.950 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.790 0.000 1516.070 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.430 296.000 1669.710 300.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 0.000 1138.410 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.450 0.000 1525.730 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 296.000 1671.550 300.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 196.560 1700.000 197.160 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.570 0.000 1535.850 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 0.000 1545.970 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1673.570 296.000 1673.850 300.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.410 296.000 1675.690 300.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 74.840 1700.000 75.440 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.710 296.000 1677.990 300.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 202.680 1700.000 203.280 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.010 296.000 1680.290 300.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 208.120 1700.000 208.720 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 0.000 1555.630 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 213.560 1700.000 214.160 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 219.000 1700.000 219.600 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.910 0.000 1158.190 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 224.440 1700.000 225.040 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.470 0.000 1565.750 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.590 0.000 1575.870 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.250 0.000 1585.530 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.850 296.000 1682.130 300.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 229.880 1700.000 230.480 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.370 0.000 1595.650 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.030 0.000 1605.310 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 4.000 247.480 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.570 0.000 1167.850 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1615.150 0.000 1615.430 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 236.000 1700.000 236.600 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.270 0.000 1625.550 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.930 0.000 1635.210 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 241.440 1700.000 242.040 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.150 296.000 1684.430 300.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 246.880 1700.000 247.480 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 252.320 1700.000 252.920 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 257.760 1700.000 258.360 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.690 0.000 1177.970 4.000 ;
    END
  END la_data_out[9]
  PIN master_data_addr_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 296.000 1.290 300.000 ;
    END
  END master_data_addr_to_inter_i[0]
  PIN master_data_addr_to_inter_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 296.000 153.090 300.000 ;
    END
  END master_data_addr_to_inter_i[10]
  PIN master_data_addr_to_inter_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 296.000 163.670 300.000 ;
    END
  END master_data_addr_to_inter_i[11]
  PIN master_data_addr_to_inter_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 296.000 174.250 300.000 ;
    END
  END master_data_addr_to_inter_i[12]
  PIN master_data_addr_to_inter_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 296.000 184.830 300.000 ;
    END
  END master_data_addr_to_inter_i[13]
  PIN master_data_addr_to_inter_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 296.000 195.410 300.000 ;
    END
  END master_data_addr_to_inter_i[14]
  PIN master_data_addr_to_inter_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 296.000 205.990 300.000 ;
    END
  END master_data_addr_to_inter_i[15]
  PIN master_data_addr_to_inter_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 296.000 216.570 300.000 ;
    END
  END master_data_addr_to_inter_i[16]
  PIN master_data_addr_to_inter_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 296.000 227.150 300.000 ;
    END
  END master_data_addr_to_inter_i[17]
  PIN master_data_addr_to_inter_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 296.000 237.730 300.000 ;
    END
  END master_data_addr_to_inter_i[18]
  PIN master_data_addr_to_inter_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 296.000 248.310 300.000 ;
    END
  END master_data_addr_to_inter_i[19]
  PIN master_data_addr_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 296.000 28.430 300.000 ;
    END
  END master_data_addr_to_inter_i[1]
  PIN master_data_addr_to_inter_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 296.000 258.890 300.000 ;
    END
  END master_data_addr_to_inter_i[20]
  PIN master_data_addr_to_inter_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 296.000 269.470 300.000 ;
    END
  END master_data_addr_to_inter_i[21]
  PIN master_data_addr_to_inter_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 296.000 280.050 300.000 ;
    END
  END master_data_addr_to_inter_i[22]
  PIN master_data_addr_to_inter_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 296.000 290.630 300.000 ;
    END
  END master_data_addr_to_inter_i[23]
  PIN master_data_addr_to_inter_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 296.000 300.750 300.000 ;
    END
  END master_data_addr_to_inter_i[24]
  PIN master_data_addr_to_inter_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 296.000 311.330 300.000 ;
    END
  END master_data_addr_to_inter_i[25]
  PIN master_data_addr_to_inter_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 296.000 321.910 300.000 ;
    END
  END master_data_addr_to_inter_i[26]
  PIN master_data_addr_to_inter_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 296.000 330.650 300.000 ;
    END
  END master_data_addr_to_inter_i[27]
  PIN master_data_addr_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 296.000 56.030 300.000 ;
    END
  END master_data_addr_to_inter_i[2]
  PIN master_data_addr_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 296.000 68.450 300.000 ;
    END
  END master_data_addr_to_inter_i[3]
  PIN master_data_addr_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 296.000 81.330 300.000 ;
    END
  END master_data_addr_to_inter_i[4]
  PIN master_data_addr_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 296.000 94.210 300.000 ;
    END
  END master_data_addr_to_inter_i[5]
  PIN master_data_addr_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 296.000 106.630 300.000 ;
    END
  END master_data_addr_to_inter_i[6]
  PIN master_data_addr_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 296.000 119.510 300.000 ;
    END
  END master_data_addr_to_inter_i[7]
  PIN master_data_addr_to_inter_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 296.000 131.930 300.000 ;
    END
  END master_data_addr_to_inter_i[8]
  PIN master_data_addr_to_inter_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 296.000 142.510 300.000 ;
    END
  END master_data_addr_to_inter_i[9]
  PIN master_data_addr_to_inter_ro_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 296.000 3.130 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[0]
  PIN master_data_addr_to_inter_ro_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 296.000 155.390 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[10]
  PIN master_data_addr_to_inter_ro_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 296.000 165.970 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[11]
  PIN master_data_addr_to_inter_ro_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 296.000 176.550 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[12]
  PIN master_data_addr_to_inter_ro_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 296.000 187.130 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[13]
  PIN master_data_addr_to_inter_ro_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 296.000 197.250 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[14]
  PIN master_data_addr_to_inter_ro_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 296.000 207.830 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[15]
  PIN master_data_addr_to_inter_ro_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 296.000 218.410 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[16]
  PIN master_data_addr_to_inter_ro_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 296.000 228.990 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[17]
  PIN master_data_addr_to_inter_ro_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 296.000 239.570 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[18]
  PIN master_data_addr_to_inter_ro_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 296.000 250.150 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[19]
  PIN master_data_addr_to_inter_ro_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 296.000 30.730 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[1]
  PIN master_data_addr_to_inter_ro_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 296.000 260.730 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[20]
  PIN master_data_addr_to_inter_ro_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 296.000 271.310 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[21]
  PIN master_data_addr_to_inter_ro_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 296.000 281.890 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[22]
  PIN master_data_addr_to_inter_ro_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 296.000 292.470 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[23]
  PIN master_data_addr_to_inter_ro_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 296.000 303.050 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[24]
  PIN master_data_addr_to_inter_ro_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 296.000 313.630 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[25]
  PIN master_data_addr_to_inter_ro_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 296.000 57.870 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[2]
  PIN master_data_addr_to_inter_ro_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 296.000 70.750 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[3]
  PIN master_data_addr_to_inter_ro_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 296.000 83.630 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[4]
  PIN master_data_addr_to_inter_ro_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 296.000 96.050 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[5]
  PIN master_data_addr_to_inter_ro_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 296.000 108.930 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[6]
  PIN master_data_addr_to_inter_ro_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 296.000 121.350 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[7]
  PIN master_data_addr_to_inter_ro_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 296.000 134.230 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[8]
  PIN master_data_addr_to_inter_ro_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 296.000 144.810 300.000 ;
    END
  END master_data_addr_to_inter_ro_i[9]
  PIN master_data_be_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 296.000 5.430 300.000 ;
    END
  END master_data_be_to_inter_i[0]
  PIN master_data_be_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 296.000 32.570 300.000 ;
    END
  END master_data_be_to_inter_i[1]
  PIN master_data_be_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 296.000 60.170 300.000 ;
    END
  END master_data_be_to_inter_i[2]
  PIN master_data_be_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 296.000 73.050 300.000 ;
    END
  END master_data_be_to_inter_i[3]
  PIN master_data_be_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 296.000 85.470 300.000 ;
    END
  END master_data_be_to_inter_i[4]
  PIN master_data_be_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 296.000 98.350 300.000 ;
    END
  END master_data_be_to_inter_i[5]
  PIN master_data_be_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 296.000 110.770 300.000 ;
    END
  END master_data_be_to_inter_i[6]
  PIN master_data_be_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 296.000 123.650 300.000 ;
    END
  END master_data_be_to_inter_i[7]
  PIN master_data_gnt_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 296.000 7.270 300.000 ;
    END
  END master_data_gnt_to_inter_o[0]
  PIN master_data_gnt_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 296.000 34.870 300.000 ;
    END
  END master_data_gnt_to_inter_o[1]
  PIN master_data_gnt_to_inter_ro_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 296.000 9.570 300.000 ;
    END
  END master_data_gnt_to_inter_ro_o[0]
  PIN master_data_gnt_to_inter_ro_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 296.000 37.170 300.000 ;
    END
  END master_data_gnt_to_inter_ro_o[1]
  PIN master_data_rdata_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 296.000 11.410 300.000 ;
    END
  END master_data_rdata_to_inter_o[0]
  PIN master_data_rdata_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 296.000 157.230 300.000 ;
    END
  END master_data_rdata_to_inter_o[10]
  PIN master_data_rdata_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 296.000 167.810 300.000 ;
    END
  END master_data_rdata_to_inter_o[11]
  PIN master_data_rdata_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 296.000 178.390 300.000 ;
    END
  END master_data_rdata_to_inter_o[12]
  PIN master_data_rdata_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 296.000 188.970 300.000 ;
    END
  END master_data_rdata_to_inter_o[13]
  PIN master_data_rdata_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 296.000 199.550 300.000 ;
    END
  END master_data_rdata_to_inter_o[14]
  PIN master_data_rdata_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 296.000 210.130 300.000 ;
    END
  END master_data_rdata_to_inter_o[15]
  PIN master_data_rdata_to_inter_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 296.000 220.710 300.000 ;
    END
  END master_data_rdata_to_inter_o[16]
  PIN master_data_rdata_to_inter_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 296.000 231.290 300.000 ;
    END
  END master_data_rdata_to_inter_o[17]
  PIN master_data_rdata_to_inter_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 296.000 241.870 300.000 ;
    END
  END master_data_rdata_to_inter_o[18]
  PIN master_data_rdata_to_inter_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 296.000 252.450 300.000 ;
    END
  END master_data_rdata_to_inter_o[19]
  PIN master_data_rdata_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 296.000 39.010 300.000 ;
    END
  END master_data_rdata_to_inter_o[1]
  PIN master_data_rdata_to_inter_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 296.000 263.030 300.000 ;
    END
  END master_data_rdata_to_inter_o[20]
  PIN master_data_rdata_to_inter_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 296.000 273.610 300.000 ;
    END
  END master_data_rdata_to_inter_o[21]
  PIN master_data_rdata_to_inter_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 296.000 284.190 300.000 ;
    END
  END master_data_rdata_to_inter_o[22]
  PIN master_data_rdata_to_inter_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 296.000 294.770 300.000 ;
    END
  END master_data_rdata_to_inter_o[23]
  PIN master_data_rdata_to_inter_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 296.000 305.350 300.000 ;
    END
  END master_data_rdata_to_inter_o[24]
  PIN master_data_rdata_to_inter_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 296.000 315.930 300.000 ;
    END
  END master_data_rdata_to_inter_o[25]
  PIN master_data_rdata_to_inter_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 296.000 324.210 300.000 ;
    END
  END master_data_rdata_to_inter_o[26]
  PIN master_data_rdata_to_inter_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 296.000 332.490 300.000 ;
    END
  END master_data_rdata_to_inter_o[27]
  PIN master_data_rdata_to_inter_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 296.000 338.930 300.000 ;
    END
  END master_data_rdata_to_inter_o[28]
  PIN master_data_rdata_to_inter_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 296.000 345.370 300.000 ;
    END
  END master_data_rdata_to_inter_o[29]
  PIN master_data_rdata_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 296.000 62.470 300.000 ;
    END
  END master_data_rdata_to_inter_o[2]
  PIN master_data_rdata_to_inter_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 296.000 351.810 300.000 ;
    END
  END master_data_rdata_to_inter_o[30]
  PIN master_data_rdata_to_inter_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 296.000 357.790 300.000 ;
    END
  END master_data_rdata_to_inter_o[31]
  PIN master_data_rdata_to_inter_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 296.000 364.230 300.000 ;
    END
  END master_data_rdata_to_inter_o[32]
  PIN master_data_rdata_to_inter_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 296.000 370.670 300.000 ;
    END
  END master_data_rdata_to_inter_o[33]
  PIN master_data_rdata_to_inter_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 296.000 377.110 300.000 ;
    END
  END master_data_rdata_to_inter_o[34]
  PIN master_data_rdata_to_inter_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 296.000 383.550 300.000 ;
    END
  END master_data_rdata_to_inter_o[35]
  PIN master_data_rdata_to_inter_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 296.000 389.530 300.000 ;
    END
  END master_data_rdata_to_inter_o[36]
  PIN master_data_rdata_to_inter_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 296.000 395.970 300.000 ;
    END
  END master_data_rdata_to_inter_o[37]
  PIN master_data_rdata_to_inter_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 296.000 402.410 300.000 ;
    END
  END master_data_rdata_to_inter_o[38]
  PIN master_data_rdata_to_inter_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 296.000 408.850 300.000 ;
    END
  END master_data_rdata_to_inter_o[39]
  PIN master_data_rdata_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 296.000 74.890 300.000 ;
    END
  END master_data_rdata_to_inter_o[3]
  PIN master_data_rdata_to_inter_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 296.000 414.830 300.000 ;
    END
  END master_data_rdata_to_inter_o[40]
  PIN master_data_rdata_to_inter_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 296.000 421.270 300.000 ;
    END
  END master_data_rdata_to_inter_o[41]
  PIN master_data_rdata_to_inter_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 296.000 427.710 300.000 ;
    END
  END master_data_rdata_to_inter_o[42]
  PIN master_data_rdata_to_inter_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 296.000 434.150 300.000 ;
    END
  END master_data_rdata_to_inter_o[43]
  PIN master_data_rdata_to_inter_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 296.000 440.130 300.000 ;
    END
  END master_data_rdata_to_inter_o[44]
  PIN master_data_rdata_to_inter_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 296.000 446.570 300.000 ;
    END
  END master_data_rdata_to_inter_o[45]
  PIN master_data_rdata_to_inter_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 296.000 453.010 300.000 ;
    END
  END master_data_rdata_to_inter_o[46]
  PIN master_data_rdata_to_inter_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 296.000 459.450 300.000 ;
    END
  END master_data_rdata_to_inter_o[47]
  PIN master_data_rdata_to_inter_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 296.000 465.890 300.000 ;
    END
  END master_data_rdata_to_inter_o[48]
  PIN master_data_rdata_to_inter_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 296.000 471.870 300.000 ;
    END
  END master_data_rdata_to_inter_o[49]
  PIN master_data_rdata_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 296.000 87.770 300.000 ;
    END
  END master_data_rdata_to_inter_o[4]
  PIN master_data_rdata_to_inter_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 296.000 478.310 300.000 ;
    END
  END master_data_rdata_to_inter_o[50]
  PIN master_data_rdata_to_inter_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 296.000 484.750 300.000 ;
    END
  END master_data_rdata_to_inter_o[51]
  PIN master_data_rdata_to_inter_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 296.000 491.190 300.000 ;
    END
  END master_data_rdata_to_inter_o[52]
  PIN master_data_rdata_to_inter_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 296.000 497.170 300.000 ;
    END
  END master_data_rdata_to_inter_o[53]
  PIN master_data_rdata_to_inter_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 296.000 503.610 300.000 ;
    END
  END master_data_rdata_to_inter_o[54]
  PIN master_data_rdata_to_inter_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 296.000 510.050 300.000 ;
    END
  END master_data_rdata_to_inter_o[55]
  PIN master_data_rdata_to_inter_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 296.000 516.490 300.000 ;
    END
  END master_data_rdata_to_inter_o[56]
  PIN master_data_rdata_to_inter_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 296.000 522.930 300.000 ;
    END
  END master_data_rdata_to_inter_o[57]
  PIN master_data_rdata_to_inter_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 296.000 528.910 300.000 ;
    END
  END master_data_rdata_to_inter_o[58]
  PIN master_data_rdata_to_inter_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 296.000 535.350 300.000 ;
    END
  END master_data_rdata_to_inter_o[59]
  PIN master_data_rdata_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 296.000 100.190 300.000 ;
    END
  END master_data_rdata_to_inter_o[5]
  PIN master_data_rdata_to_inter_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 296.000 541.790 300.000 ;
    END
  END master_data_rdata_to_inter_o[60]
  PIN master_data_rdata_to_inter_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 296.000 548.230 300.000 ;
    END
  END master_data_rdata_to_inter_o[61]
  PIN master_data_rdata_to_inter_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 296.000 554.210 300.000 ;
    END
  END master_data_rdata_to_inter_o[62]
  PIN master_data_rdata_to_inter_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 296.000 560.650 300.000 ;
    END
  END master_data_rdata_to_inter_o[63]
  PIN master_data_rdata_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 296.000 113.070 300.000 ;
    END
  END master_data_rdata_to_inter_o[6]
  PIN master_data_rdata_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 296.000 125.490 300.000 ;
    END
  END master_data_rdata_to_inter_o[7]
  PIN master_data_rdata_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 296.000 136.070 300.000 ;
    END
  END master_data_rdata_to_inter_o[8]
  PIN master_data_rdata_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 296.000 146.650 300.000 ;
    END
  END master_data_rdata_to_inter_o[9]
  PIN master_data_rdata_to_inter_ro_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 296.000 13.710 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[0]
  PIN master_data_rdata_to_inter_ro_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 296.000 159.530 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[10]
  PIN master_data_rdata_to_inter_ro_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 296.000 170.110 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[11]
  PIN master_data_rdata_to_inter_ro_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 296.000 180.690 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[12]
  PIN master_data_rdata_to_inter_ro_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 296.000 191.270 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[13]
  PIN master_data_rdata_to_inter_ro_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 296.000 201.850 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[14]
  PIN master_data_rdata_to_inter_ro_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 296.000 212.430 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[15]
  PIN master_data_rdata_to_inter_ro_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 296.000 223.010 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[16]
  PIN master_data_rdata_to_inter_ro_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 296.000 233.590 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[17]
  PIN master_data_rdata_to_inter_ro_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 296.000 244.170 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[18]
  PIN master_data_rdata_to_inter_ro_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 296.000 254.290 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[19]
  PIN master_data_rdata_to_inter_ro_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 296.000 41.310 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[1]
  PIN master_data_rdata_to_inter_ro_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 296.000 264.870 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[20]
  PIN master_data_rdata_to_inter_ro_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 296.000 275.450 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[21]
  PIN master_data_rdata_to_inter_ro_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 296.000 286.030 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[22]
  PIN master_data_rdata_to_inter_ro_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 296.000 296.610 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[23]
  PIN master_data_rdata_to_inter_ro_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 296.000 307.190 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[24]
  PIN master_data_rdata_to_inter_ro_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 296.000 317.770 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[25]
  PIN master_data_rdata_to_inter_ro_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 296.000 326.510 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[26]
  PIN master_data_rdata_to_inter_ro_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 296.000 334.790 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[27]
  PIN master_data_rdata_to_inter_ro_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 296.000 341.230 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[28]
  PIN master_data_rdata_to_inter_ro_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 296.000 347.210 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[29]
  PIN master_data_rdata_to_inter_ro_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 296.000 64.310 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[2]
  PIN master_data_rdata_to_inter_ro_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 296.000 353.650 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[30]
  PIN master_data_rdata_to_inter_ro_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 296.000 360.090 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[31]
  PIN master_data_rdata_to_inter_ro_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 296.000 366.530 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[32]
  PIN master_data_rdata_to_inter_ro_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 296.000 372.970 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[33]
  PIN master_data_rdata_to_inter_ro_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 296.000 378.950 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[34]
  PIN master_data_rdata_to_inter_ro_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 296.000 385.390 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[35]
  PIN master_data_rdata_to_inter_ro_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 296.000 391.830 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[36]
  PIN master_data_rdata_to_inter_ro_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 296.000 398.270 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[37]
  PIN master_data_rdata_to_inter_ro_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 296.000 404.250 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[38]
  PIN master_data_rdata_to_inter_ro_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 296.000 410.690 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[39]
  PIN master_data_rdata_to_inter_ro_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 296.000 77.190 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[3]
  PIN master_data_rdata_to_inter_ro_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 296.000 417.130 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[40]
  PIN master_data_rdata_to_inter_ro_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 296.000 423.570 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[41]
  PIN master_data_rdata_to_inter_ro_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 296.000 430.010 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[42]
  PIN master_data_rdata_to_inter_ro_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 296.000 435.990 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[43]
  PIN master_data_rdata_to_inter_ro_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 296.000 442.430 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[44]
  PIN master_data_rdata_to_inter_ro_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 296.000 448.870 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[45]
  PIN master_data_rdata_to_inter_ro_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 296.000 455.310 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[46]
  PIN master_data_rdata_to_inter_ro_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 296.000 461.290 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[47]
  PIN master_data_rdata_to_inter_ro_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 296.000 467.730 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[48]
  PIN master_data_rdata_to_inter_ro_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 296.000 474.170 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[49]
  PIN master_data_rdata_to_inter_ro_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 296.000 89.610 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[4]
  PIN master_data_rdata_to_inter_ro_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 296.000 480.610 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[50]
  PIN master_data_rdata_to_inter_ro_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 296.000 487.050 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[51]
  PIN master_data_rdata_to_inter_ro_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 296.000 493.030 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[52]
  PIN master_data_rdata_to_inter_ro_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 296.000 499.470 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[53]
  PIN master_data_rdata_to_inter_ro_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 296.000 505.910 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[54]
  PIN master_data_rdata_to_inter_ro_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 296.000 512.350 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[55]
  PIN master_data_rdata_to_inter_ro_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 296.000 518.330 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[56]
  PIN master_data_rdata_to_inter_ro_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 296.000 524.770 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[57]
  PIN master_data_rdata_to_inter_ro_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 296.000 531.210 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[58]
  PIN master_data_rdata_to_inter_ro_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 296.000 537.650 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[59]
  PIN master_data_rdata_to_inter_ro_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 296.000 102.490 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[5]
  PIN master_data_rdata_to_inter_ro_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 296.000 543.630 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[60]
  PIN master_data_rdata_to_inter_ro_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 296.000 550.070 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[61]
  PIN master_data_rdata_to_inter_ro_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 296.000 556.510 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[62]
  PIN master_data_rdata_to_inter_ro_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 296.000 562.950 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[63]
  PIN master_data_rdata_to_inter_ro_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 296.000 114.910 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[6]
  PIN master_data_rdata_to_inter_ro_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 296.000 127.790 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[7]
  PIN master_data_rdata_to_inter_ro_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 296.000 138.370 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[8]
  PIN master_data_rdata_to_inter_ro_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 296.000 148.950 300.000 ;
    END
  END master_data_rdata_to_inter_ro_o[9]
  PIN master_data_req_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 296.000 16.010 300.000 ;
    END
  END master_data_req_to_inter_i[0]
  PIN master_data_req_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 296.000 43.150 300.000 ;
    END
  END master_data_req_to_inter_i[1]
  PIN master_data_req_to_inter_ro_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 296.000 17.850 300.000 ;
    END
  END master_data_req_to_inter_ro_i[0]
  PIN master_data_req_to_inter_ro_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 296.000 45.450 300.000 ;
    END
  END master_data_req_to_inter_ro_i[1]
  PIN master_data_rvalid_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 296.000 20.150 300.000 ;
    END
  END master_data_rvalid_to_inter_o[0]
  PIN master_data_rvalid_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 296.000 47.750 300.000 ;
    END
  END master_data_rvalid_to_inter_o[1]
  PIN master_data_rvalid_to_inter_ro_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 296.000 21.990 300.000 ;
    END
  END master_data_rvalid_to_inter_ro_o[0]
  PIN master_data_rvalid_to_inter_ro_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 296.000 49.590 300.000 ;
    END
  END master_data_rvalid_to_inter_ro_o[1]
  PIN master_data_wdata_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 296.000 24.290 300.000 ;
    END
  END master_data_wdata_to_inter_i[0]
  PIN master_data_wdata_to_inter_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 296.000 161.370 300.000 ;
    END
  END master_data_wdata_to_inter_i[10]
  PIN master_data_wdata_to_inter_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 296.000 171.950 300.000 ;
    END
  END master_data_wdata_to_inter_i[11]
  PIN master_data_wdata_to_inter_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 296.000 182.530 300.000 ;
    END
  END master_data_wdata_to_inter_i[12]
  PIN master_data_wdata_to_inter_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 296.000 193.110 300.000 ;
    END
  END master_data_wdata_to_inter_i[13]
  PIN master_data_wdata_to_inter_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 296.000 203.690 300.000 ;
    END
  END master_data_wdata_to_inter_i[14]
  PIN master_data_wdata_to_inter_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 296.000 214.270 300.000 ;
    END
  END master_data_wdata_to_inter_i[15]
  PIN master_data_wdata_to_inter_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 296.000 224.850 300.000 ;
    END
  END master_data_wdata_to_inter_i[16]
  PIN master_data_wdata_to_inter_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 296.000 235.430 300.000 ;
    END
  END master_data_wdata_to_inter_i[17]
  PIN master_data_wdata_to_inter_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 296.000 246.010 300.000 ;
    END
  END master_data_wdata_to_inter_i[18]
  PIN master_data_wdata_to_inter_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 296.000 256.590 300.000 ;
    END
  END master_data_wdata_to_inter_i[19]
  PIN master_data_wdata_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 296.000 51.890 300.000 ;
    END
  END master_data_wdata_to_inter_i[1]
  PIN master_data_wdata_to_inter_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 296.000 267.170 300.000 ;
    END
  END master_data_wdata_to_inter_i[20]
  PIN master_data_wdata_to_inter_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 296.000 277.750 300.000 ;
    END
  END master_data_wdata_to_inter_i[21]
  PIN master_data_wdata_to_inter_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 296.000 288.330 300.000 ;
    END
  END master_data_wdata_to_inter_i[22]
  PIN master_data_wdata_to_inter_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 296.000 298.910 300.000 ;
    END
  END master_data_wdata_to_inter_i[23]
  PIN master_data_wdata_to_inter_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 296.000 309.490 300.000 ;
    END
  END master_data_wdata_to_inter_i[24]
  PIN master_data_wdata_to_inter_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 296.000 320.070 300.000 ;
    END
  END master_data_wdata_to_inter_i[25]
  PIN master_data_wdata_to_inter_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 296.000 328.350 300.000 ;
    END
  END master_data_wdata_to_inter_i[26]
  PIN master_data_wdata_to_inter_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 296.000 337.090 300.000 ;
    END
  END master_data_wdata_to_inter_i[27]
  PIN master_data_wdata_to_inter_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 296.000 343.070 300.000 ;
    END
  END master_data_wdata_to_inter_i[28]
  PIN master_data_wdata_to_inter_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 296.000 349.510 300.000 ;
    END
  END master_data_wdata_to_inter_i[29]
  PIN master_data_wdata_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 296.000 66.610 300.000 ;
    END
  END master_data_wdata_to_inter_i[2]
  PIN master_data_wdata_to_inter_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 296.000 355.950 300.000 ;
    END
  END master_data_wdata_to_inter_i[30]
  PIN master_data_wdata_to_inter_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 296.000 362.390 300.000 ;
    END
  END master_data_wdata_to_inter_i[31]
  PIN master_data_wdata_to_inter_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 296.000 368.370 300.000 ;
    END
  END master_data_wdata_to_inter_i[32]
  PIN master_data_wdata_to_inter_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 296.000 374.810 300.000 ;
    END
  END master_data_wdata_to_inter_i[33]
  PIN master_data_wdata_to_inter_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 296.000 381.250 300.000 ;
    END
  END master_data_wdata_to_inter_i[34]
  PIN master_data_wdata_to_inter_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 296.000 387.690 300.000 ;
    END
  END master_data_wdata_to_inter_i[35]
  PIN master_data_wdata_to_inter_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 296.000 393.670 300.000 ;
    END
  END master_data_wdata_to_inter_i[36]
  PIN master_data_wdata_to_inter_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 296.000 400.110 300.000 ;
    END
  END master_data_wdata_to_inter_i[37]
  PIN master_data_wdata_to_inter_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 296.000 406.550 300.000 ;
    END
  END master_data_wdata_to_inter_i[38]
  PIN master_data_wdata_to_inter_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 296.000 412.990 300.000 ;
    END
  END master_data_wdata_to_inter_i[39]
  PIN master_data_wdata_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 296.000 79.030 300.000 ;
    END
  END master_data_wdata_to_inter_i[3]
  PIN master_data_wdata_to_inter_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 296.000 419.430 300.000 ;
    END
  END master_data_wdata_to_inter_i[40]
  PIN master_data_wdata_to_inter_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 296.000 425.410 300.000 ;
    END
  END master_data_wdata_to_inter_i[41]
  PIN master_data_wdata_to_inter_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 296.000 431.850 300.000 ;
    END
  END master_data_wdata_to_inter_i[42]
  PIN master_data_wdata_to_inter_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 296.000 438.290 300.000 ;
    END
  END master_data_wdata_to_inter_i[43]
  PIN master_data_wdata_to_inter_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 296.000 444.730 300.000 ;
    END
  END master_data_wdata_to_inter_i[44]
  PIN master_data_wdata_to_inter_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 296.000 450.710 300.000 ;
    END
  END master_data_wdata_to_inter_i[45]
  PIN master_data_wdata_to_inter_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 296.000 457.150 300.000 ;
    END
  END master_data_wdata_to_inter_i[46]
  PIN master_data_wdata_to_inter_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 296.000 463.590 300.000 ;
    END
  END master_data_wdata_to_inter_i[47]
  PIN master_data_wdata_to_inter_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 296.000 470.030 300.000 ;
    END
  END master_data_wdata_to_inter_i[48]
  PIN master_data_wdata_to_inter_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 296.000 476.470 300.000 ;
    END
  END master_data_wdata_to_inter_i[49]
  PIN master_data_wdata_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 296.000 91.910 300.000 ;
    END
  END master_data_wdata_to_inter_i[4]
  PIN master_data_wdata_to_inter_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 296.000 482.450 300.000 ;
    END
  END master_data_wdata_to_inter_i[50]
  PIN master_data_wdata_to_inter_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 296.000 488.890 300.000 ;
    END
  END master_data_wdata_to_inter_i[51]
  PIN master_data_wdata_to_inter_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 296.000 495.330 300.000 ;
    END
  END master_data_wdata_to_inter_i[52]
  PIN master_data_wdata_to_inter_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 296.000 501.770 300.000 ;
    END
  END master_data_wdata_to_inter_i[53]
  PIN master_data_wdata_to_inter_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 296.000 507.750 300.000 ;
    END
  END master_data_wdata_to_inter_i[54]
  PIN master_data_wdata_to_inter_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 296.000 514.190 300.000 ;
    END
  END master_data_wdata_to_inter_i[55]
  PIN master_data_wdata_to_inter_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 296.000 520.630 300.000 ;
    END
  END master_data_wdata_to_inter_i[56]
  PIN master_data_wdata_to_inter_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 296.000 527.070 300.000 ;
    END
  END master_data_wdata_to_inter_i[57]
  PIN master_data_wdata_to_inter_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 296.000 533.510 300.000 ;
    END
  END master_data_wdata_to_inter_i[58]
  PIN master_data_wdata_to_inter_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 296.000 539.490 300.000 ;
    END
  END master_data_wdata_to_inter_i[59]
  PIN master_data_wdata_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 296.000 104.330 300.000 ;
    END
  END master_data_wdata_to_inter_i[5]
  PIN master_data_wdata_to_inter_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 296.000 545.930 300.000 ;
    END
  END master_data_wdata_to_inter_i[60]
  PIN master_data_wdata_to_inter_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 296.000 552.370 300.000 ;
    END
  END master_data_wdata_to_inter_i[61]
  PIN master_data_wdata_to_inter_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 296.000 558.810 300.000 ;
    END
  END master_data_wdata_to_inter_i[62]
  PIN master_data_wdata_to_inter_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 296.000 564.790 300.000 ;
    END
  END master_data_wdata_to_inter_i[63]
  PIN master_data_wdata_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 296.000 117.210 300.000 ;
    END
  END master_data_wdata_to_inter_i[6]
  PIN master_data_wdata_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 296.000 130.090 300.000 ;
    END
  END master_data_wdata_to_inter_i[7]
  PIN master_data_wdata_to_inter_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 296.000 140.670 300.000 ;
    END
  END master_data_wdata_to_inter_i[8]
  PIN master_data_wdata_to_inter_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 296.000 150.790 300.000 ;
    END
  END master_data_wdata_to_inter_i[9]
  PIN master_data_we_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 296.000 26.590 300.000 ;
    END
  END master_data_we_to_inter_i[0]
  PIN master_data_we_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 296.000 53.730 300.000 ;
    END
  END master_data_we_to_inter_i[1]
  PIN rxd_uart
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 2.760 1700.000 3.360 ;
    END
  END rxd_uart
  PIN rxd_uart_to_mem
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 8.200 1700.000 8.800 ;
    END
  END rxd_uart_to_mem
  PIN slave_data_addr_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 296.000 567.090 300.000 ;
    END
  END slave_data_addr_to_inter_o[0]
  PIN slave_data_addr_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 296.000 719.350 300.000 ;
    END
  END slave_data_addr_to_inter_o[10]
  PIN slave_data_addr_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 296.000 731.770 300.000 ;
    END
  END slave_data_addr_to_inter_o[11]
  PIN slave_data_addr_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 296.000 744.650 300.000 ;
    END
  END slave_data_addr_to_inter_o[12]
  PIN slave_data_addr_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 296.000 757.070 300.000 ;
    END
  END slave_data_addr_to_inter_o[13]
  PIN slave_data_addr_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 296.000 769.950 300.000 ;
    END
  END slave_data_addr_to_inter_o[14]
  PIN slave_data_addr_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 296.000 782.370 300.000 ;
    END
  END slave_data_addr_to_inter_o[15]
  PIN slave_data_addr_to_inter_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 296.000 795.250 300.000 ;
    END
  END slave_data_addr_to_inter_o[16]
  PIN slave_data_addr_to_inter_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 296.000 805.830 300.000 ;
    END
  END slave_data_addr_to_inter_o[17]
  PIN slave_data_addr_to_inter_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 296.000 816.410 300.000 ;
    END
  END slave_data_addr_to_inter_o[18]
  PIN slave_data_addr_to_inter_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 296.000 826.990 300.000 ;
    END
  END slave_data_addr_to_inter_o[19]
  PIN slave_data_addr_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 296.000 585.950 300.000 ;
    END
  END slave_data_addr_to_inter_o[1]
  PIN slave_data_addr_to_inter_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 296.000 837.570 300.000 ;
    END
  END slave_data_addr_to_inter_o[20]
  PIN slave_data_addr_to_inter_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.870 296.000 848.150 300.000 ;
    END
  END slave_data_addr_to_inter_o[21]
  PIN slave_data_addr_to_inter_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 296.000 858.730 300.000 ;
    END
  END slave_data_addr_to_inter_o[22]
  PIN slave_data_addr_to_inter_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.030 296.000 869.310 300.000 ;
    END
  END slave_data_addr_to_inter_o[23]
  PIN slave_data_addr_to_inter_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 296.000 879.430 300.000 ;
    END
  END slave_data_addr_to_inter_o[24]
  PIN slave_data_addr_to_inter_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 296.000 890.010 300.000 ;
    END
  END slave_data_addr_to_inter_o[25]
  PIN slave_data_addr_to_inter_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 296.000 900.590 300.000 ;
    END
  END slave_data_addr_to_inter_o[26]
  PIN slave_data_addr_to_inter_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 296.000 911.170 300.000 ;
    END
  END slave_data_addr_to_inter_o[27]
  PIN slave_data_addr_to_inter_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 296.000 921.750 300.000 ;
    END
  END slave_data_addr_to_inter_o[28]
  PIN slave_data_addr_to_inter_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 296.000 932.330 300.000 ;
    END
  END slave_data_addr_to_inter_o[29]
  PIN slave_data_addr_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 296.000 605.270 300.000 ;
    END
  END slave_data_addr_to_inter_o[2]
  PIN slave_data_addr_to_inter_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 296.000 942.910 300.000 ;
    END
  END slave_data_addr_to_inter_o[30]
  PIN slave_data_addr_to_inter_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 296.000 953.490 300.000 ;
    END
  END slave_data_addr_to_inter_o[31]
  PIN slave_data_addr_to_inter_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 296.000 964.070 300.000 ;
    END
  END slave_data_addr_to_inter_o[32]
  PIN slave_data_addr_to_inter_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.370 296.000 974.650 300.000 ;
    END
  END slave_data_addr_to_inter_o[33]
  PIN slave_data_addr_to_inter_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 296.000 985.230 300.000 ;
    END
  END slave_data_addr_to_inter_o[34]
  PIN slave_data_addr_to_inter_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.530 296.000 995.810 300.000 ;
    END
  END slave_data_addr_to_inter_o[35]
  PIN slave_data_addr_to_inter_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.110 296.000 1006.390 300.000 ;
    END
  END slave_data_addr_to_inter_o[36]
  PIN slave_data_addr_to_inter_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 296.000 1016.970 300.000 ;
    END
  END slave_data_addr_to_inter_o[37]
  PIN slave_data_addr_to_inter_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 296.000 1027.550 300.000 ;
    END
  END slave_data_addr_to_inter_o[38]
  PIN slave_data_addr_to_inter_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 296.000 1038.130 300.000 ;
    END
  END slave_data_addr_to_inter_o[39]
  PIN slave_data_addr_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 296.000 624.130 300.000 ;
    END
  END slave_data_addr_to_inter_o[3]
  PIN slave_data_addr_to_inter_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.430 296.000 1048.710 300.000 ;
    END
  END slave_data_addr_to_inter_o[40]
  PIN slave_data_addr_to_inter_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 296.000 1059.290 300.000 ;
    END
  END slave_data_addr_to_inter_o[41]
  PIN slave_data_addr_to_inter_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 296.000 1069.870 300.000 ;
    END
  END slave_data_addr_to_inter_o[42]
  PIN slave_data_addr_to_inter_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.170 296.000 1080.450 300.000 ;
    END
  END slave_data_addr_to_inter_o[43]
  PIN slave_data_addr_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 296.000 642.990 300.000 ;
    END
  END slave_data_addr_to_inter_o[4]
  PIN slave_data_addr_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 296.000 655.870 300.000 ;
    END
  END slave_data_addr_to_inter_o[5]
  PIN slave_data_addr_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 296.000 668.290 300.000 ;
    END
  END slave_data_addr_to_inter_o[6]
  PIN slave_data_addr_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 296.000 681.170 300.000 ;
    END
  END slave_data_addr_to_inter_o[7]
  PIN slave_data_addr_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 296.000 693.590 300.000 ;
    END
  END slave_data_addr_to_inter_o[8]
  PIN slave_data_addr_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 296.000 706.470 300.000 ;
    END
  END slave_data_addr_to_inter_o[9]
  PIN slave_data_addr_to_inter_ro_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 296.000 569.390 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[0]
  PIN slave_data_addr_to_inter_ro_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 296.000 721.190 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[10]
  PIN slave_data_addr_to_inter_ro_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 296.000 734.070 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[11]
  PIN slave_data_addr_to_inter_ro_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 296.000 746.490 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[12]
  PIN slave_data_addr_to_inter_ro_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 296.000 759.370 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[13]
  PIN slave_data_addr_to_inter_ro_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 296.000 771.790 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[14]
  PIN slave_data_addr_to_inter_ro_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 296.000 784.670 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[15]
  PIN slave_data_addr_to_inter_ro_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 296.000 797.090 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[16]
  PIN slave_data_addr_to_inter_ro_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 296.000 807.670 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[17]
  PIN slave_data_addr_to_inter_ro_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 296.000 818.250 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[18]
  PIN slave_data_addr_to_inter_ro_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 296.000 828.830 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[19]
  PIN slave_data_addr_to_inter_ro_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 296.000 588.250 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[1]
  PIN slave_data_addr_to_inter_ro_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 296.000 839.410 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[20]
  PIN slave_data_addr_to_inter_ro_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 296.000 849.990 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[21]
  PIN slave_data_addr_to_inter_ro_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 296.000 860.570 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[22]
  PIN slave_data_addr_to_inter_ro_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 296.000 871.150 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[23]
  PIN slave_data_addr_to_inter_ro_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 296.000 881.730 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[24]
  PIN slave_data_addr_to_inter_ro_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 296.000 892.310 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[25]
  PIN slave_data_addr_to_inter_ro_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 296.000 902.890 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[26]
  PIN slave_data_addr_to_inter_ro_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.190 296.000 913.470 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[27]
  PIN slave_data_addr_to_inter_ro_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 296.000 924.050 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[28]
  PIN slave_data_addr_to_inter_ro_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 296.000 934.630 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[29]
  PIN slave_data_addr_to_inter_ro_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 296.000 607.110 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[2]
  PIN slave_data_addr_to_inter_ro_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 296.000 945.210 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[30]
  PIN slave_data_addr_to_inter_ro_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.510 296.000 955.790 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[31]
  PIN slave_data_addr_to_inter_ro_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 296.000 966.370 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[32]
  PIN slave_data_addr_to_inter_ro_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 296.000 976.950 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[33]
  PIN slave_data_addr_to_inter_ro_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 296.000 987.530 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[34]
  PIN slave_data_addr_to_inter_ro_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.830 296.000 998.110 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[35]
  PIN slave_data_addr_to_inter_ro_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.410 296.000 1008.690 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[36]
  PIN slave_data_addr_to_inter_ro_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 296.000 1019.270 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[37]
  PIN slave_data_addr_to_inter_ro_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 296.000 1029.390 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[38]
  PIN slave_data_addr_to_inter_ro_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.690 296.000 1039.970 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[39]
  PIN slave_data_addr_to_inter_ro_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 296.000 626.430 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[3]
  PIN slave_data_addr_to_inter_ro_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 296.000 1050.550 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[40]
  PIN slave_data_addr_to_inter_ro_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.850 296.000 1061.130 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[41]
  PIN slave_data_addr_to_inter_ro_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 296.000 1071.710 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[42]
  PIN slave_data_addr_to_inter_ro_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 296.000 1082.290 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[43]
  PIN slave_data_addr_to_inter_ro_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 296.000 645.290 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[4]
  PIN slave_data_addr_to_inter_ro_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 296.000 657.710 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[5]
  PIN slave_data_addr_to_inter_ro_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 296.000 670.590 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[6]
  PIN slave_data_addr_to_inter_ro_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 296.000 683.010 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[7]
  PIN slave_data_addr_to_inter_ro_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 296.000 695.890 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[8]
  PIN slave_data_addr_to_inter_ro_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 296.000 708.770 300.000 ;
    END
  END slave_data_addr_to_inter_ro_o[9]
  PIN slave_data_be_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 296.000 571.230 300.000 ;
    END
  END slave_data_be_to_inter_o[0]
  PIN slave_data_be_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 296.000 723.490 300.000 ;
    END
  END slave_data_be_to_inter_o[10]
  PIN slave_data_be_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 296.000 735.910 300.000 ;
    END
  END slave_data_be_to_inter_o[11]
  PIN slave_data_be_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 296.000 748.790 300.000 ;
    END
  END slave_data_be_to_inter_o[12]
  PIN slave_data_be_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 296.000 761.210 300.000 ;
    END
  END slave_data_be_to_inter_o[13]
  PIN slave_data_be_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 296.000 774.090 300.000 ;
    END
  END slave_data_be_to_inter_o[14]
  PIN slave_data_be_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 296.000 786.510 300.000 ;
    END
  END slave_data_be_to_inter_o[15]
  PIN slave_data_be_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 296.000 590.090 300.000 ;
    END
  END slave_data_be_to_inter_o[1]
  PIN slave_data_be_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 296.000 609.410 300.000 ;
    END
  END slave_data_be_to_inter_o[2]
  PIN slave_data_be_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 296.000 628.270 300.000 ;
    END
  END slave_data_be_to_inter_o[3]
  PIN slave_data_be_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 296.000 647.130 300.000 ;
    END
  END slave_data_be_to_inter_o[4]
  PIN slave_data_be_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 296.000 660.010 300.000 ;
    END
  END slave_data_be_to_inter_o[5]
  PIN slave_data_be_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 296.000 672.890 300.000 ;
    END
  END slave_data_be_to_inter_o[6]
  PIN slave_data_be_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 296.000 685.310 300.000 ;
    END
  END slave_data_be_to_inter_o[7]
  PIN slave_data_be_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 296.000 698.190 300.000 ;
    END
  END slave_data_be_to_inter_o[8]
  PIN slave_data_be_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 296.000 710.610 300.000 ;
    END
  END slave_data_be_to_inter_o[9]
  PIN slave_data_rdata_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 296.000 573.530 300.000 ;
    END
  END slave_data_rdata_to_inter_i[0]
  PIN slave_data_rdata_to_inter_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.410 296.000 1445.690 300.000 ;
    END
  END slave_data_rdata_to_inter_i[100]
  PIN slave_data_rdata_to_inter_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.850 296.000 1452.130 300.000 ;
    END
  END slave_data_rdata_to_inter_i[101]
  PIN slave_data_rdata_to_inter_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.290 296.000 1458.570 300.000 ;
    END
  END slave_data_rdata_to_inter_i[102]
  PIN slave_data_rdata_to_inter_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.270 296.000 1464.550 300.000 ;
    END
  END slave_data_rdata_to_inter_i[103]
  PIN slave_data_rdata_to_inter_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.710 296.000 1470.990 300.000 ;
    END
  END slave_data_rdata_to_inter_i[104]
  PIN slave_data_rdata_to_inter_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.150 296.000 1477.430 300.000 ;
    END
  END slave_data_rdata_to_inter_i[105]
  PIN slave_data_rdata_to_inter_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.590 296.000 1483.870 300.000 ;
    END
  END slave_data_rdata_to_inter_i[106]
  PIN slave_data_rdata_to_inter_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.570 296.000 1489.850 300.000 ;
    END
  END slave_data_rdata_to_inter_i[107]
  PIN slave_data_rdata_to_inter_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.010 296.000 1496.290 300.000 ;
    END
  END slave_data_rdata_to_inter_i[108]
  PIN slave_data_rdata_to_inter_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1502.450 296.000 1502.730 300.000 ;
    END
  END slave_data_rdata_to_inter_i[109]
  PIN slave_data_rdata_to_inter_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 296.000 725.330 300.000 ;
    END
  END slave_data_rdata_to_inter_i[10]
  PIN slave_data_rdata_to_inter_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.890 296.000 1509.170 300.000 ;
    END
  END slave_data_rdata_to_inter_i[110]
  PIN slave_data_rdata_to_inter_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.870 296.000 1515.150 300.000 ;
    END
  END slave_data_rdata_to_inter_i[111]
  PIN slave_data_rdata_to_inter_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.310 296.000 1521.590 300.000 ;
    END
  END slave_data_rdata_to_inter_i[112]
  PIN slave_data_rdata_to_inter_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.750 296.000 1528.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[113]
  PIN slave_data_rdata_to_inter_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.190 296.000 1534.470 300.000 ;
    END
  END slave_data_rdata_to_inter_i[114]
  PIN slave_data_rdata_to_inter_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.630 296.000 1540.910 300.000 ;
    END
  END slave_data_rdata_to_inter_i[115]
  PIN slave_data_rdata_to_inter_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.610 296.000 1546.890 300.000 ;
    END
  END slave_data_rdata_to_inter_i[116]
  PIN slave_data_rdata_to_inter_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.050 296.000 1553.330 300.000 ;
    END
  END slave_data_rdata_to_inter_i[117]
  PIN slave_data_rdata_to_inter_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.490 296.000 1559.770 300.000 ;
    END
  END slave_data_rdata_to_inter_i[118]
  PIN slave_data_rdata_to_inter_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.930 296.000 1566.210 300.000 ;
    END
  END slave_data_rdata_to_inter_i[119]
  PIN slave_data_rdata_to_inter_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 296.000 738.210 300.000 ;
    END
  END slave_data_rdata_to_inter_i[11]
  PIN slave_data_rdata_to_inter_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.910 296.000 1572.190 300.000 ;
    END
  END slave_data_rdata_to_inter_i[120]
  PIN slave_data_rdata_to_inter_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.350 296.000 1578.630 300.000 ;
    END
  END slave_data_rdata_to_inter_i[121]
  PIN slave_data_rdata_to_inter_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.790 296.000 1585.070 300.000 ;
    END
  END slave_data_rdata_to_inter_i[122]
  PIN slave_data_rdata_to_inter_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.230 296.000 1591.510 300.000 ;
    END
  END slave_data_rdata_to_inter_i[123]
  PIN slave_data_rdata_to_inter_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.670 296.000 1597.950 300.000 ;
    END
  END slave_data_rdata_to_inter_i[124]
  PIN slave_data_rdata_to_inter_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 296.000 1603.930 300.000 ;
    END
  END slave_data_rdata_to_inter_i[125]
  PIN slave_data_rdata_to_inter_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 296.000 1610.370 300.000 ;
    END
  END slave_data_rdata_to_inter_i[126]
  PIN slave_data_rdata_to_inter_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 296.000 1616.810 300.000 ;
    END
  END slave_data_rdata_to_inter_i[127]
  PIN slave_data_rdata_to_inter_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 296.000 750.630 300.000 ;
    END
  END slave_data_rdata_to_inter_i[12]
  PIN slave_data_rdata_to_inter_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 296.000 763.510 300.000 ;
    END
  END slave_data_rdata_to_inter_i[13]
  PIN slave_data_rdata_to_inter_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 296.000 776.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[14]
  PIN slave_data_rdata_to_inter_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 296.000 788.810 300.000 ;
    END
  END slave_data_rdata_to_inter_i[15]
  PIN slave_data_rdata_to_inter_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 296.000 799.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[16]
  PIN slave_data_rdata_to_inter_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 296.000 809.970 300.000 ;
    END
  END slave_data_rdata_to_inter_i[17]
  PIN slave_data_rdata_to_inter_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 296.000 820.550 300.000 ;
    END
  END slave_data_rdata_to_inter_i[18]
  PIN slave_data_rdata_to_inter_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 296.000 831.130 300.000 ;
    END
  END slave_data_rdata_to_inter_i[19]
  PIN slave_data_rdata_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 296.000 592.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[1]
  PIN slave_data_rdata_to_inter_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.430 296.000 841.710 300.000 ;
    END
  END slave_data_rdata_to_inter_i[20]
  PIN slave_data_rdata_to_inter_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 296.000 852.290 300.000 ;
    END
  END slave_data_rdata_to_inter_i[21]
  PIN slave_data_rdata_to_inter_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 296.000 862.870 300.000 ;
    END
  END slave_data_rdata_to_inter_i[22]
  PIN slave_data_rdata_to_inter_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 296.000 873.450 300.000 ;
    END
  END slave_data_rdata_to_inter_i[23]
  PIN slave_data_rdata_to_inter_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.750 296.000 884.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[24]
  PIN slave_data_rdata_to_inter_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 296.000 894.610 300.000 ;
    END
  END slave_data_rdata_to_inter_i[25]
  PIN slave_data_rdata_to_inter_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 296.000 905.190 300.000 ;
    END
  END slave_data_rdata_to_inter_i[26]
  PIN slave_data_rdata_to_inter_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.490 296.000 915.770 300.000 ;
    END
  END slave_data_rdata_to_inter_i[27]
  PIN slave_data_rdata_to_inter_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 296.000 925.890 300.000 ;
    END
  END slave_data_rdata_to_inter_i[28]
  PIN slave_data_rdata_to_inter_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.190 296.000 936.470 300.000 ;
    END
  END slave_data_rdata_to_inter_i[29]
  PIN slave_data_rdata_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 296.000 611.250 300.000 ;
    END
  END slave_data_rdata_to_inter_i[2]
  PIN slave_data_rdata_to_inter_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 296.000 947.050 300.000 ;
    END
  END slave_data_rdata_to_inter_i[30]
  PIN slave_data_rdata_to_inter_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 296.000 957.630 300.000 ;
    END
  END slave_data_rdata_to_inter_i[31]
  PIN slave_data_rdata_to_inter_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 296.000 968.210 300.000 ;
    END
  END slave_data_rdata_to_inter_i[32]
  PIN slave_data_rdata_to_inter_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.510 296.000 978.790 300.000 ;
    END
  END slave_data_rdata_to_inter_i[33]
  PIN slave_data_rdata_to_inter_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.090 296.000 989.370 300.000 ;
    END
  END slave_data_rdata_to_inter_i[34]
  PIN slave_data_rdata_to_inter_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 296.000 999.950 300.000 ;
    END
  END slave_data_rdata_to_inter_i[35]
  PIN slave_data_rdata_to_inter_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 296.000 1010.530 300.000 ;
    END
  END slave_data_rdata_to_inter_i[36]
  PIN slave_data_rdata_to_inter_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 296.000 1021.110 300.000 ;
    END
  END slave_data_rdata_to_inter_i[37]
  PIN slave_data_rdata_to_inter_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.410 296.000 1031.690 300.000 ;
    END
  END slave_data_rdata_to_inter_i[38]
  PIN slave_data_rdata_to_inter_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.990 296.000 1042.270 300.000 ;
    END
  END slave_data_rdata_to_inter_i[39]
  PIN slave_data_rdata_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 296.000 630.570 300.000 ;
    END
  END slave_data_rdata_to_inter_i[3]
  PIN slave_data_rdata_to_inter_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.570 296.000 1052.850 300.000 ;
    END
  END slave_data_rdata_to_inter_i[40]
  PIN slave_data_rdata_to_inter_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.150 296.000 1063.430 300.000 ;
    END
  END slave_data_rdata_to_inter_i[41]
  PIN slave_data_rdata_to_inter_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 296.000 1074.010 300.000 ;
    END
  END slave_data_rdata_to_inter_i[42]
  PIN slave_data_rdata_to_inter_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 296.000 1084.590 300.000 ;
    END
  END slave_data_rdata_to_inter_i[43]
  PIN slave_data_rdata_to_inter_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.750 296.000 1091.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[44]
  PIN slave_data_rdata_to_inter_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.730 296.000 1097.010 300.000 ;
    END
  END slave_data_rdata_to_inter_i[45]
  PIN slave_data_rdata_to_inter_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.170 296.000 1103.450 300.000 ;
    END
  END slave_data_rdata_to_inter_i[46]
  PIN slave_data_rdata_to_inter_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 296.000 1109.890 300.000 ;
    END
  END slave_data_rdata_to_inter_i[47]
  PIN slave_data_rdata_to_inter_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.050 296.000 1116.330 300.000 ;
    END
  END slave_data_rdata_to_inter_i[48]
  PIN slave_data_rdata_to_inter_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.030 296.000 1122.310 300.000 ;
    END
  END slave_data_rdata_to_inter_i[49]
  PIN slave_data_rdata_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 296.000 649.430 300.000 ;
    END
  END slave_data_rdata_to_inter_i[4]
  PIN slave_data_rdata_to_inter_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 296.000 1128.750 300.000 ;
    END
  END slave_data_rdata_to_inter_i[50]
  PIN slave_data_rdata_to_inter_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 296.000 1135.190 300.000 ;
    END
  END slave_data_rdata_to_inter_i[51]
  PIN slave_data_rdata_to_inter_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 296.000 1141.630 300.000 ;
    END
  END slave_data_rdata_to_inter_i[52]
  PIN slave_data_rdata_to_inter_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.790 296.000 1148.070 300.000 ;
    END
  END slave_data_rdata_to_inter_i[53]
  PIN slave_data_rdata_to_inter_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.770 296.000 1154.050 300.000 ;
    END
  END slave_data_rdata_to_inter_i[54]
  PIN slave_data_rdata_to_inter_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.210 296.000 1160.490 300.000 ;
    END
  END slave_data_rdata_to_inter_i[55]
  PIN slave_data_rdata_to_inter_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.650 296.000 1166.930 300.000 ;
    END
  END slave_data_rdata_to_inter_i[56]
  PIN slave_data_rdata_to_inter_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.090 296.000 1173.370 300.000 ;
    END
  END slave_data_rdata_to_inter_i[57]
  PIN slave_data_rdata_to_inter_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.070 296.000 1179.350 300.000 ;
    END
  END slave_data_rdata_to_inter_i[58]
  PIN slave_data_rdata_to_inter_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.510 296.000 1185.790 300.000 ;
    END
  END slave_data_rdata_to_inter_i[59]
  PIN slave_data_rdata_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 296.000 662.310 300.000 ;
    END
  END slave_data_rdata_to_inter_i[5]
  PIN slave_data_rdata_to_inter_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 296.000 1192.230 300.000 ;
    END
  END slave_data_rdata_to_inter_i[60]
  PIN slave_data_rdata_to_inter_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.390 296.000 1198.670 300.000 ;
    END
  END slave_data_rdata_to_inter_i[61]
  PIN slave_data_rdata_to_inter_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.830 296.000 1205.110 300.000 ;
    END
  END slave_data_rdata_to_inter_i[62]
  PIN slave_data_rdata_to_inter_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 296.000 1211.090 300.000 ;
    END
  END slave_data_rdata_to_inter_i[63]
  PIN slave_data_rdata_to_inter_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 296.000 1217.530 300.000 ;
    END
  END slave_data_rdata_to_inter_i[64]
  PIN slave_data_rdata_to_inter_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 296.000 1223.970 300.000 ;
    END
  END slave_data_rdata_to_inter_i[65]
  PIN slave_data_rdata_to_inter_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 296.000 1230.410 300.000 ;
    END
  END slave_data_rdata_to_inter_i[66]
  PIN slave_data_rdata_to_inter_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.110 296.000 1236.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[67]
  PIN slave_data_rdata_to_inter_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 296.000 1242.830 300.000 ;
    END
  END slave_data_rdata_to_inter_i[68]
  PIN slave_data_rdata_to_inter_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.990 296.000 1249.270 300.000 ;
    END
  END slave_data_rdata_to_inter_i[69]
  PIN slave_data_rdata_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 296.000 674.730 300.000 ;
    END
  END slave_data_rdata_to_inter_i[6]
  PIN slave_data_rdata_to_inter_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.430 296.000 1255.710 300.000 ;
    END
  END slave_data_rdata_to_inter_i[70]
  PIN slave_data_rdata_to_inter_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.870 296.000 1262.150 300.000 ;
    END
  END slave_data_rdata_to_inter_i[71]
  PIN slave_data_rdata_to_inter_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.850 296.000 1268.130 300.000 ;
    END
  END slave_data_rdata_to_inter_i[72]
  PIN slave_data_rdata_to_inter_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.290 296.000 1274.570 300.000 ;
    END
  END slave_data_rdata_to_inter_i[73]
  PIN slave_data_rdata_to_inter_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.730 296.000 1281.010 300.000 ;
    END
  END slave_data_rdata_to_inter_i[74]
  PIN slave_data_rdata_to_inter_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.170 296.000 1287.450 300.000 ;
    END
  END slave_data_rdata_to_inter_i[75]
  PIN slave_data_rdata_to_inter_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.150 296.000 1293.430 300.000 ;
    END
  END slave_data_rdata_to_inter_i[76]
  PIN slave_data_rdata_to_inter_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.590 296.000 1299.870 300.000 ;
    END
  END slave_data_rdata_to_inter_i[77]
  PIN slave_data_rdata_to_inter_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.030 296.000 1306.310 300.000 ;
    END
  END slave_data_rdata_to_inter_i[78]
  PIN slave_data_rdata_to_inter_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.470 296.000 1312.750 300.000 ;
    END
  END slave_data_rdata_to_inter_i[79]
  PIN slave_data_rdata_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 296.000 687.610 300.000 ;
    END
  END slave_data_rdata_to_inter_i[7]
  PIN slave_data_rdata_to_inter_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.450 296.000 1318.730 300.000 ;
    END
  END slave_data_rdata_to_inter_i[80]
  PIN slave_data_rdata_to_inter_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.890 296.000 1325.170 300.000 ;
    END
  END slave_data_rdata_to_inter_i[81]
  PIN slave_data_rdata_to_inter_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.330 296.000 1331.610 300.000 ;
    END
  END slave_data_rdata_to_inter_i[82]
  PIN slave_data_rdata_to_inter_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.770 296.000 1338.050 300.000 ;
    END
  END slave_data_rdata_to_inter_i[83]
  PIN slave_data_rdata_to_inter_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 296.000 1344.490 300.000 ;
    END
  END slave_data_rdata_to_inter_i[84]
  PIN slave_data_rdata_to_inter_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.190 296.000 1350.470 300.000 ;
    END
  END slave_data_rdata_to_inter_i[85]
  PIN slave_data_rdata_to_inter_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.630 296.000 1356.910 300.000 ;
    END
  END slave_data_rdata_to_inter_i[86]
  PIN slave_data_rdata_to_inter_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.070 296.000 1363.350 300.000 ;
    END
  END slave_data_rdata_to_inter_i[87]
  PIN slave_data_rdata_to_inter_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.510 296.000 1369.790 300.000 ;
    END
  END slave_data_rdata_to_inter_i[88]
  PIN slave_data_rdata_to_inter_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.490 296.000 1375.770 300.000 ;
    END
  END slave_data_rdata_to_inter_i[89]
  PIN slave_data_rdata_to_inter_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 296.000 700.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[8]
  PIN slave_data_rdata_to_inter_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.930 296.000 1382.210 300.000 ;
    END
  END slave_data_rdata_to_inter_i[90]
  PIN slave_data_rdata_to_inter_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.370 296.000 1388.650 300.000 ;
    END
  END slave_data_rdata_to_inter_i[91]
  PIN slave_data_rdata_to_inter_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.810 296.000 1395.090 300.000 ;
    END
  END slave_data_rdata_to_inter_i[92]
  PIN slave_data_rdata_to_inter_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.250 296.000 1401.530 300.000 ;
    END
  END slave_data_rdata_to_inter_i[93]
  PIN slave_data_rdata_to_inter_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 296.000 1407.510 300.000 ;
    END
  END slave_data_rdata_to_inter_i[94]
  PIN slave_data_rdata_to_inter_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 296.000 1413.950 300.000 ;
    END
  END slave_data_rdata_to_inter_i[95]
  PIN slave_data_rdata_to_inter_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 296.000 1420.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[96]
  PIN slave_data_rdata_to_inter_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 296.000 1426.830 300.000 ;
    END
  END slave_data_rdata_to_inter_i[97]
  PIN slave_data_rdata_to_inter_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.530 296.000 1432.810 300.000 ;
    END
  END slave_data_rdata_to_inter_i[98]
  PIN slave_data_rdata_to_inter_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.970 296.000 1439.250 300.000 ;
    END
  END slave_data_rdata_to_inter_i[99]
  PIN slave_data_rdata_to_inter_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 296.000 712.910 300.000 ;
    END
  END slave_data_rdata_to_inter_i[9]
  PIN slave_data_rdata_to_inter_ro_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 296.000 575.370 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[0]
  PIN slave_data_rdata_to_inter_ro_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.710 296.000 1447.990 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[100]
  PIN slave_data_rdata_to_inter_ro_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.690 296.000 1453.970 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[101]
  PIN slave_data_rdata_to_inter_ro_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.130 296.000 1460.410 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[102]
  PIN slave_data_rdata_to_inter_ro_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.570 296.000 1466.850 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[103]
  PIN slave_data_rdata_to_inter_ro_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.010 296.000 1473.290 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[104]
  PIN slave_data_rdata_to_inter_ro_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.990 296.000 1479.270 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[105]
  PIN slave_data_rdata_to_inter_ro_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.430 296.000 1485.710 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[106]
  PIN slave_data_rdata_to_inter_ro_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.870 296.000 1492.150 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[107]
  PIN slave_data_rdata_to_inter_ro_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.310 296.000 1498.590 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[108]
  PIN slave_data_rdata_to_inter_ro_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.750 296.000 1505.030 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[109]
  PIN slave_data_rdata_to_inter_ro_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 296.000 727.630 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[10]
  PIN slave_data_rdata_to_inter_ro_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.730 296.000 1511.010 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[110]
  PIN slave_data_rdata_to_inter_ro_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.170 296.000 1517.450 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[111]
  PIN slave_data_rdata_to_inter_ro_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.610 296.000 1523.890 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[112]
  PIN slave_data_rdata_to_inter_ro_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.050 296.000 1530.330 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[113]
  PIN slave_data_rdata_to_inter_ro_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.030 296.000 1536.310 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[114]
  PIN slave_data_rdata_to_inter_ro_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 296.000 1542.750 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[115]
  PIN slave_data_rdata_to_inter_ro_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 296.000 1549.190 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[116]
  PIN slave_data_rdata_to_inter_ro_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 296.000 1555.630 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[117]
  PIN slave_data_rdata_to_inter_ro_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.330 296.000 1561.610 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[118]
  PIN slave_data_rdata_to_inter_ro_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.770 296.000 1568.050 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[119]
  PIN slave_data_rdata_to_inter_ro_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 296.000 740.050 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[11]
  PIN slave_data_rdata_to_inter_ro_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.210 296.000 1574.490 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[120]
  PIN slave_data_rdata_to_inter_ro_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.650 296.000 1580.930 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[121]
  PIN slave_data_rdata_to_inter_ro_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.090 296.000 1587.370 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[122]
  PIN slave_data_rdata_to_inter_ro_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.070 296.000 1593.350 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[123]
  PIN slave_data_rdata_to_inter_ro_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.510 296.000 1599.790 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[124]
  PIN slave_data_rdata_to_inter_ro_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.950 296.000 1606.230 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[125]
  PIN slave_data_rdata_to_inter_ro_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.390 296.000 1612.670 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[126]
  PIN slave_data_rdata_to_inter_ro_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.370 296.000 1618.650 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[127]
  PIN slave_data_rdata_to_inter_ro_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 296.000 752.930 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[12]
  PIN slave_data_rdata_to_inter_ro_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 296.000 765.810 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[13]
  PIN slave_data_rdata_to_inter_ro_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 296.000 778.230 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[14]
  PIN slave_data_rdata_to_inter_ro_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 296.000 791.110 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[15]
  PIN slave_data_rdata_to_inter_ro_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 296.000 801.690 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[16]
  PIN slave_data_rdata_to_inter_ro_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 296.000 812.270 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[17]
  PIN slave_data_rdata_to_inter_ro_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 296.000 822.850 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[18]
  PIN slave_data_rdata_to_inter_ro_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 296.000 832.970 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[19]
  PIN slave_data_rdata_to_inter_ro_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 296.000 594.690 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[1]
  PIN slave_data_rdata_to_inter_ro_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 296.000 843.550 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[20]
  PIN slave_data_rdata_to_inter_ro_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 296.000 854.130 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[21]
  PIN slave_data_rdata_to_inter_ro_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 296.000 864.710 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[22]
  PIN slave_data_rdata_to_inter_ro_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 296.000 875.290 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[23]
  PIN slave_data_rdata_to_inter_ro_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 296.000 885.870 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[24]
  PIN slave_data_rdata_to_inter_ro_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 296.000 896.450 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[25]
  PIN slave_data_rdata_to_inter_ro_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 296.000 907.030 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[26]
  PIN slave_data_rdata_to_inter_ro_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.330 296.000 917.610 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[27]
  PIN slave_data_rdata_to_inter_ro_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 296.000 928.190 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[28]
  PIN slave_data_rdata_to_inter_ro_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 296.000 938.770 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[29]
  PIN slave_data_rdata_to_inter_ro_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 296.000 613.550 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[2]
  PIN slave_data_rdata_to_inter_ro_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 296.000 949.350 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[30]
  PIN slave_data_rdata_to_inter_ro_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 296.000 959.930 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[31]
  PIN slave_data_rdata_to_inter_ro_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 296.000 970.510 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[32]
  PIN slave_data_rdata_to_inter_ro_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 296.000 981.090 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[33]
  PIN slave_data_rdata_to_inter_ro_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 296.000 991.670 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[34]
  PIN slave_data_rdata_to_inter_ro_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.970 296.000 1002.250 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[35]
  PIN slave_data_rdata_to_inter_ro_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 296.000 1012.830 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[36]
  PIN slave_data_rdata_to_inter_ro_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.130 296.000 1023.410 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[37]
  PIN slave_data_rdata_to_inter_ro_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 296.000 1033.990 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[38]
  PIN slave_data_rdata_to_inter_ro_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 296.000 1044.570 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[39]
  PIN slave_data_rdata_to_inter_ro_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 296.000 632.410 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[3]
  PIN slave_data_rdata_to_inter_ro_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.870 296.000 1055.150 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[40]
  PIN slave_data_rdata_to_inter_ro_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 296.000 1065.730 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[41]
  PIN slave_data_rdata_to_inter_ro_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 296.000 1075.850 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[42]
  PIN slave_data_rdata_to_inter_ro_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 296.000 1086.430 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[43]
  PIN slave_data_rdata_to_inter_ro_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 296.000 1092.870 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[44]
  PIN slave_data_rdata_to_inter_ro_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 296.000 1099.310 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[45]
  PIN slave_data_rdata_to_inter_ro_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.470 296.000 1105.750 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[46]
  PIN slave_data_rdata_to_inter_ro_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 296.000 1112.190 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[47]
  PIN slave_data_rdata_to_inter_ro_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.890 296.000 1118.170 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[48]
  PIN slave_data_rdata_to_inter_ro_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 296.000 1124.610 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[49]
  PIN slave_data_rdata_to_inter_ro_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 296.000 651.730 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[4]
  PIN slave_data_rdata_to_inter_ro_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.770 296.000 1131.050 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[50]
  PIN slave_data_rdata_to_inter_ro_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 296.000 1137.490 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[51]
  PIN slave_data_rdata_to_inter_ro_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 296.000 1143.470 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[52]
  PIN slave_data_rdata_to_inter_ro_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 296.000 1149.910 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[53]
  PIN slave_data_rdata_to_inter_ro_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 296.000 1156.350 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[54]
  PIN slave_data_rdata_to_inter_ro_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 296.000 1162.790 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[55]
  PIN slave_data_rdata_to_inter_ro_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.490 296.000 1168.770 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[56]
  PIN slave_data_rdata_to_inter_ro_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.930 296.000 1175.210 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[57]
  PIN slave_data_rdata_to_inter_ro_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.370 296.000 1181.650 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[58]
  PIN slave_data_rdata_to_inter_ro_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 296.000 1188.090 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[59]
  PIN slave_data_rdata_to_inter_ro_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 296.000 664.150 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[5]
  PIN slave_data_rdata_to_inter_ro_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 296.000 1194.530 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[60]
  PIN slave_data_rdata_to_inter_ro_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.230 296.000 1200.510 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[61]
  PIN slave_data_rdata_to_inter_ro_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.670 296.000 1206.950 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[62]
  PIN slave_data_rdata_to_inter_ro_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.110 296.000 1213.390 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[63]
  PIN slave_data_rdata_to_inter_ro_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 296.000 1219.830 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[64]
  PIN slave_data_rdata_to_inter_ro_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.530 296.000 1225.810 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[65]
  PIN slave_data_rdata_to_inter_ro_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.970 296.000 1232.250 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[66]
  PIN slave_data_rdata_to_inter_ro_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.410 296.000 1238.690 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[67]
  PIN slave_data_rdata_to_inter_ro_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.850 296.000 1245.130 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[68]
  PIN slave_data_rdata_to_inter_ro_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.290 296.000 1251.570 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[69]
  PIN slave_data_rdata_to_inter_ro_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 296.000 677.030 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[6]
  PIN slave_data_rdata_to_inter_ro_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 296.000 1257.550 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[70]
  PIN slave_data_rdata_to_inter_ro_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.710 296.000 1263.990 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[71]
  PIN slave_data_rdata_to_inter_ro_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1270.150 296.000 1270.430 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[72]
  PIN slave_data_rdata_to_inter_ro_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.590 296.000 1276.870 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[73]
  PIN slave_data_rdata_to_inter_ro_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.570 296.000 1282.850 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[74]
  PIN slave_data_rdata_to_inter_ro_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 296.000 1289.290 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[75]
  PIN slave_data_rdata_to_inter_ro_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.450 296.000 1295.730 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[76]
  PIN slave_data_rdata_to_inter_ro_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.890 296.000 1302.170 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[77]
  PIN slave_data_rdata_to_inter_ro_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.330 296.000 1308.610 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[78]
  PIN slave_data_rdata_to_inter_ro_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 296.000 1314.590 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[79]
  PIN slave_data_rdata_to_inter_ro_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 296.000 689.450 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[7]
  PIN slave_data_rdata_to_inter_ro_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.750 296.000 1321.030 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[80]
  PIN slave_data_rdata_to_inter_ro_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.190 296.000 1327.470 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[81]
  PIN slave_data_rdata_to_inter_ro_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 296.000 1333.910 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[82]
  PIN slave_data_rdata_to_inter_ro_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.610 296.000 1339.890 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[83]
  PIN slave_data_rdata_to_inter_ro_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 296.000 1346.330 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[84]
  PIN slave_data_rdata_to_inter_ro_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 296.000 1352.770 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[85]
  PIN slave_data_rdata_to_inter_ro_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 296.000 1359.210 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[86]
  PIN slave_data_rdata_to_inter_ro_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.910 296.000 1365.190 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[87]
  PIN slave_data_rdata_to_inter_ro_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.350 296.000 1371.630 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[88]
  PIN slave_data_rdata_to_inter_ro_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.790 296.000 1378.070 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[89]
  PIN slave_data_rdata_to_inter_ro_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 296.000 702.330 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[8]
  PIN slave_data_rdata_to_inter_ro_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.230 296.000 1384.510 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[90]
  PIN slave_data_rdata_to_inter_ro_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.670 296.000 1390.950 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[91]
  PIN slave_data_rdata_to_inter_ro_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.650 296.000 1396.930 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[92]
  PIN slave_data_rdata_to_inter_ro_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.090 296.000 1403.370 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[93]
  PIN slave_data_rdata_to_inter_ro_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.530 296.000 1409.810 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[94]
  PIN slave_data_rdata_to_inter_ro_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.970 296.000 1416.250 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[95]
  PIN slave_data_rdata_to_inter_ro_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.950 296.000 1422.230 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[96]
  PIN slave_data_rdata_to_inter_ro_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.390 296.000 1428.670 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[97]
  PIN slave_data_rdata_to_inter_ro_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.830 296.000 1435.110 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[98]
  PIN slave_data_rdata_to_inter_ro_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.270 296.000 1441.550 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[99]
  PIN slave_data_rdata_to_inter_ro_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 296.000 714.750 300.000 ;
    END
  END slave_data_rdata_to_inter_ro_i[9]
  PIN slave_data_req_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 296.000 577.670 300.000 ;
    END
  END slave_data_req_to_inter_o[0]
  PIN slave_data_req_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 296.000 596.530 300.000 ;
    END
  END slave_data_req_to_inter_o[1]
  PIN slave_data_req_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 296.000 615.850 300.000 ;
    END
  END slave_data_req_to_inter_o[2]
  PIN slave_data_req_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 296.000 634.710 300.000 ;
    END
  END slave_data_req_to_inter_o[3]
  PIN slave_data_req_to_inter_ro_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 296.000 579.970 300.000 ;
    END
  END slave_data_req_to_inter_ro_o[0]
  PIN slave_data_req_to_inter_ro_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 296.000 598.830 300.000 ;
    END
  END slave_data_req_to_inter_ro_o[1]
  PIN slave_data_req_to_inter_ro_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 296.000 617.690 300.000 ;
    END
  END slave_data_req_to_inter_ro_o[2]
  PIN slave_data_req_to_inter_ro_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 296.000 636.550 300.000 ;
    END
  END slave_data_req_to_inter_ro_o[3]
  PIN slave_data_wdata_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 296.000 581.810 300.000 ;
    END
  END slave_data_wdata_to_inter_o[0]
  PIN slave_data_wdata_to_inter_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.550 296.000 1449.830 300.000 ;
    END
  END slave_data_wdata_to_inter_o[100]
  PIN slave_data_wdata_to_inter_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 296.000 1456.270 300.000 ;
    END
  END slave_data_wdata_to_inter_o[101]
  PIN slave_data_wdata_to_inter_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.430 296.000 1462.710 300.000 ;
    END
  END slave_data_wdata_to_inter_o[102]
  PIN slave_data_wdata_to_inter_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 296.000 1468.690 300.000 ;
    END
  END slave_data_wdata_to_inter_o[103]
  PIN slave_data_wdata_to_inter_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 296.000 1475.130 300.000 ;
    END
  END slave_data_wdata_to_inter_o[104]
  PIN slave_data_wdata_to_inter_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 296.000 1481.570 300.000 ;
    END
  END slave_data_wdata_to_inter_o[105]
  PIN slave_data_wdata_to_inter_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 296.000 1488.010 300.000 ;
    END
  END slave_data_wdata_to_inter_o[106]
  PIN slave_data_wdata_to_inter_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 296.000 1494.450 300.000 ;
    END
  END slave_data_wdata_to_inter_o[107]
  PIN slave_data_wdata_to_inter_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.150 296.000 1500.430 300.000 ;
    END
  END slave_data_wdata_to_inter_o[108]
  PIN slave_data_wdata_to_inter_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.590 296.000 1506.870 300.000 ;
    END
  END slave_data_wdata_to_inter_o[109]
  PIN slave_data_wdata_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 296.000 729.930 300.000 ;
    END
  END slave_data_wdata_to_inter_o[10]
  PIN slave_data_wdata_to_inter_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.030 296.000 1513.310 300.000 ;
    END
  END slave_data_wdata_to_inter_o[110]
  PIN slave_data_wdata_to_inter_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.470 296.000 1519.750 300.000 ;
    END
  END slave_data_wdata_to_inter_o[111]
  PIN slave_data_wdata_to_inter_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.450 296.000 1525.730 300.000 ;
    END
  END slave_data_wdata_to_inter_o[112]
  PIN slave_data_wdata_to_inter_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.890 296.000 1532.170 300.000 ;
    END
  END slave_data_wdata_to_inter_o[113]
  PIN slave_data_wdata_to_inter_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.330 296.000 1538.610 300.000 ;
    END
  END slave_data_wdata_to_inter_o[114]
  PIN slave_data_wdata_to_inter_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.770 296.000 1545.050 300.000 ;
    END
  END slave_data_wdata_to_inter_o[115]
  PIN slave_data_wdata_to_inter_o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.210 296.000 1551.490 300.000 ;
    END
  END slave_data_wdata_to_inter_o[116]
  PIN slave_data_wdata_to_inter_o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 296.000 1557.470 300.000 ;
    END
  END slave_data_wdata_to_inter_o[117]
  PIN slave_data_wdata_to_inter_o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.630 296.000 1563.910 300.000 ;
    END
  END slave_data_wdata_to_inter_o[118]
  PIN slave_data_wdata_to_inter_o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.070 296.000 1570.350 300.000 ;
    END
  END slave_data_wdata_to_inter_o[119]
  PIN slave_data_wdata_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 296.000 742.350 300.000 ;
    END
  END slave_data_wdata_to_inter_o[11]
  PIN slave_data_wdata_to_inter_o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.510 296.000 1576.790 300.000 ;
    END
  END slave_data_wdata_to_inter_o[120]
  PIN slave_data_wdata_to_inter_o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.490 296.000 1582.770 300.000 ;
    END
  END slave_data_wdata_to_inter_o[121]
  PIN slave_data_wdata_to_inter_o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.930 296.000 1589.210 300.000 ;
    END
  END slave_data_wdata_to_inter_o[122]
  PIN slave_data_wdata_to_inter_o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.370 296.000 1595.650 300.000 ;
    END
  END slave_data_wdata_to_inter_o[123]
  PIN slave_data_wdata_to_inter_o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1601.810 296.000 1602.090 300.000 ;
    END
  END slave_data_wdata_to_inter_o[124]
  PIN slave_data_wdata_to_inter_o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.790 296.000 1608.070 300.000 ;
    END
  END slave_data_wdata_to_inter_o[125]
  PIN slave_data_wdata_to_inter_o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.230 296.000 1614.510 300.000 ;
    END
  END slave_data_wdata_to_inter_o[126]
  PIN slave_data_wdata_to_inter_o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.670 296.000 1620.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[127]
  PIN slave_data_wdata_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 296.000 755.230 300.000 ;
    END
  END slave_data_wdata_to_inter_o[12]
  PIN slave_data_wdata_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 296.000 767.650 300.000 ;
    END
  END slave_data_wdata_to_inter_o[13]
  PIN slave_data_wdata_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 296.000 780.530 300.000 ;
    END
  END slave_data_wdata_to_inter_o[14]
  PIN slave_data_wdata_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 296.000 792.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[15]
  PIN slave_data_wdata_to_inter_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 296.000 803.530 300.000 ;
    END
  END slave_data_wdata_to_inter_o[16]
  PIN slave_data_wdata_to_inter_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 296.000 814.110 300.000 ;
    END
  END slave_data_wdata_to_inter_o[17]
  PIN slave_data_wdata_to_inter_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 296.000 824.690 300.000 ;
    END
  END slave_data_wdata_to_inter_o[18]
  PIN slave_data_wdata_to_inter_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 296.000 835.270 300.000 ;
    END
  END slave_data_wdata_to_inter_o[19]
  PIN slave_data_wdata_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 296.000 600.670 300.000 ;
    END
  END slave_data_wdata_to_inter_o[1]
  PIN slave_data_wdata_to_inter_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 296.000 845.850 300.000 ;
    END
  END slave_data_wdata_to_inter_o[20]
  PIN slave_data_wdata_to_inter_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 296.000 856.430 300.000 ;
    END
  END slave_data_wdata_to_inter_o[21]
  PIN slave_data_wdata_to_inter_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 296.000 867.010 300.000 ;
    END
  END slave_data_wdata_to_inter_o[22]
  PIN slave_data_wdata_to_inter_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 296.000 877.590 300.000 ;
    END
  END slave_data_wdata_to_inter_o[23]
  PIN slave_data_wdata_to_inter_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 296.000 888.170 300.000 ;
    END
  END slave_data_wdata_to_inter_o[24]
  PIN slave_data_wdata_to_inter_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 296.000 898.750 300.000 ;
    END
  END slave_data_wdata_to_inter_o[25]
  PIN slave_data_wdata_to_inter_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050 296.000 909.330 300.000 ;
    END
  END slave_data_wdata_to_inter_o[26]
  PIN slave_data_wdata_to_inter_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.630 296.000 919.910 300.000 ;
    END
  END slave_data_wdata_to_inter_o[27]
  PIN slave_data_wdata_to_inter_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 296.000 930.490 300.000 ;
    END
  END slave_data_wdata_to_inter_o[28]
  PIN slave_data_wdata_to_inter_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.790 296.000 941.070 300.000 ;
    END
  END slave_data_wdata_to_inter_o[29]
  PIN slave_data_wdata_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 296.000 619.990 300.000 ;
    END
  END slave_data_wdata_to_inter_o[2]
  PIN slave_data_wdata_to_inter_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 296.000 951.650 300.000 ;
    END
  END slave_data_wdata_to_inter_o[30]
  PIN slave_data_wdata_to_inter_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.950 296.000 962.230 300.000 ;
    END
  END slave_data_wdata_to_inter_o[31]
  PIN slave_data_wdata_to_inter_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 296.000 972.810 300.000 ;
    END
  END slave_data_wdata_to_inter_o[32]
  PIN slave_data_wdata_to_inter_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 296.000 982.930 300.000 ;
    END
  END slave_data_wdata_to_inter_o[33]
  PIN slave_data_wdata_to_inter_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230 296.000 993.510 300.000 ;
    END
  END slave_data_wdata_to_inter_o[34]
  PIN slave_data_wdata_to_inter_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.810 296.000 1004.090 300.000 ;
    END
  END slave_data_wdata_to_inter_o[35]
  PIN slave_data_wdata_to_inter_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 296.000 1014.670 300.000 ;
    END
  END slave_data_wdata_to_inter_o[36]
  PIN slave_data_wdata_to_inter_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 296.000 1025.250 300.000 ;
    END
  END slave_data_wdata_to_inter_o[37]
  PIN slave_data_wdata_to_inter_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.550 296.000 1035.830 300.000 ;
    END
  END slave_data_wdata_to_inter_o[38]
  PIN slave_data_wdata_to_inter_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 296.000 1046.410 300.000 ;
    END
  END slave_data_wdata_to_inter_o[39]
  PIN slave_data_wdata_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 296.000 638.850 300.000 ;
    END
  END slave_data_wdata_to_inter_o[3]
  PIN slave_data_wdata_to_inter_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 296.000 1056.990 300.000 ;
    END
  END slave_data_wdata_to_inter_o[40]
  PIN slave_data_wdata_to_inter_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.290 296.000 1067.570 300.000 ;
    END
  END slave_data_wdata_to_inter_o[41]
  PIN slave_data_wdata_to_inter_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.870 296.000 1078.150 300.000 ;
    END
  END slave_data_wdata_to_inter_o[42]
  PIN slave_data_wdata_to_inter_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 296.000 1088.730 300.000 ;
    END
  END slave_data_wdata_to_inter_o[43]
  PIN slave_data_wdata_to_inter_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 296.000 1095.170 300.000 ;
    END
  END slave_data_wdata_to_inter_o[44]
  PIN slave_data_wdata_to_inter_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 296.000 1101.610 300.000 ;
    END
  END slave_data_wdata_to_inter_o[45]
  PIN slave_data_wdata_to_inter_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.310 296.000 1107.590 300.000 ;
    END
  END slave_data_wdata_to_inter_o[46]
  PIN slave_data_wdata_to_inter_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.750 296.000 1114.030 300.000 ;
    END
  END slave_data_wdata_to_inter_o[47]
  PIN slave_data_wdata_to_inter_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 296.000 1120.470 300.000 ;
    END
  END slave_data_wdata_to_inter_o[48]
  PIN slave_data_wdata_to_inter_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.630 296.000 1126.910 300.000 ;
    END
  END slave_data_wdata_to_inter_o[49]
  PIN slave_data_wdata_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 296.000 653.570 300.000 ;
    END
  END slave_data_wdata_to_inter_o[4]
  PIN slave_data_wdata_to_inter_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.610 296.000 1132.890 300.000 ;
    END
  END slave_data_wdata_to_inter_o[50]
  PIN slave_data_wdata_to_inter_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.050 296.000 1139.330 300.000 ;
    END
  END slave_data_wdata_to_inter_o[51]
  PIN slave_data_wdata_to_inter_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.490 296.000 1145.770 300.000 ;
    END
  END slave_data_wdata_to_inter_o[52]
  PIN slave_data_wdata_to_inter_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.930 296.000 1152.210 300.000 ;
    END
  END slave_data_wdata_to_inter_o[53]
  PIN slave_data_wdata_to_inter_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.370 296.000 1158.650 300.000 ;
    END
  END slave_data_wdata_to_inter_o[54]
  PIN slave_data_wdata_to_inter_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 296.000 1164.630 300.000 ;
    END
  END slave_data_wdata_to_inter_o[55]
  PIN slave_data_wdata_to_inter_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.790 296.000 1171.070 300.000 ;
    END
  END slave_data_wdata_to_inter_o[56]
  PIN slave_data_wdata_to_inter_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 296.000 1177.510 300.000 ;
    END
  END slave_data_wdata_to_inter_o[57]
  PIN slave_data_wdata_to_inter_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 296.000 1183.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[58]
  PIN slave_data_wdata_to_inter_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.650 296.000 1189.930 300.000 ;
    END
  END slave_data_wdata_to_inter_o[59]
  PIN slave_data_wdata_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 296.000 666.450 300.000 ;
    END
  END slave_data_wdata_to_inter_o[5]
  PIN slave_data_wdata_to_inter_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.090 296.000 1196.370 300.000 ;
    END
  END slave_data_wdata_to_inter_o[60]
  PIN slave_data_wdata_to_inter_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.530 296.000 1202.810 300.000 ;
    END
  END slave_data_wdata_to_inter_o[61]
  PIN slave_data_wdata_to_inter_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.970 296.000 1209.250 300.000 ;
    END
  END slave_data_wdata_to_inter_o[62]
  PIN slave_data_wdata_to_inter_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.410 296.000 1215.690 300.000 ;
    END
  END slave_data_wdata_to_inter_o[63]
  PIN slave_data_wdata_to_inter_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.390 296.000 1221.670 300.000 ;
    END
  END slave_data_wdata_to_inter_o[64]
  PIN slave_data_wdata_to_inter_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.830 296.000 1228.110 300.000 ;
    END
  END slave_data_wdata_to_inter_o[65]
  PIN slave_data_wdata_to_inter_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.270 296.000 1234.550 300.000 ;
    END
  END slave_data_wdata_to_inter_o[66]
  PIN slave_data_wdata_to_inter_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.710 296.000 1240.990 300.000 ;
    END
  END slave_data_wdata_to_inter_o[67]
  PIN slave_data_wdata_to_inter_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.690 296.000 1246.970 300.000 ;
    END
  END slave_data_wdata_to_inter_o[68]
  PIN slave_data_wdata_to_inter_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 296.000 1253.410 300.000 ;
    END
  END slave_data_wdata_to_inter_o[69]
  PIN slave_data_wdata_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 296.000 678.870 300.000 ;
    END
  END slave_data_wdata_to_inter_o[6]
  PIN slave_data_wdata_to_inter_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.570 296.000 1259.850 300.000 ;
    END
  END slave_data_wdata_to_inter_o[70]
  PIN slave_data_wdata_to_inter_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 296.000 1266.290 300.000 ;
    END
  END slave_data_wdata_to_inter_o[71]
  PIN slave_data_wdata_to_inter_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 296.000 1272.270 300.000 ;
    END
  END slave_data_wdata_to_inter_o[72]
  PIN slave_data_wdata_to_inter_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 296.000 1278.710 300.000 ;
    END
  END slave_data_wdata_to_inter_o[73]
  PIN slave_data_wdata_to_inter_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 296.000 1285.150 300.000 ;
    END
  END slave_data_wdata_to_inter_o[74]
  PIN slave_data_wdata_to_inter_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 296.000 1291.590 300.000 ;
    END
  END slave_data_wdata_to_inter_o[75]
  PIN slave_data_wdata_to_inter_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 296.000 1298.030 300.000 ;
    END
  END slave_data_wdata_to_inter_o[76]
  PIN slave_data_wdata_to_inter_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.730 296.000 1304.010 300.000 ;
    END
  END slave_data_wdata_to_inter_o[77]
  PIN slave_data_wdata_to_inter_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.170 296.000 1310.450 300.000 ;
    END
  END slave_data_wdata_to_inter_o[78]
  PIN slave_data_wdata_to_inter_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.610 296.000 1316.890 300.000 ;
    END
  END slave_data_wdata_to_inter_o[79]
  PIN slave_data_wdata_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 296.000 691.750 300.000 ;
    END
  END slave_data_wdata_to_inter_o[7]
  PIN slave_data_wdata_to_inter_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 296.000 1323.330 300.000 ;
    END
  END slave_data_wdata_to_inter_o[80]
  PIN slave_data_wdata_to_inter_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.030 296.000 1329.310 300.000 ;
    END
  END slave_data_wdata_to_inter_o[81]
  PIN slave_data_wdata_to_inter_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 296.000 1335.750 300.000 ;
    END
  END slave_data_wdata_to_inter_o[82]
  PIN slave_data_wdata_to_inter_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.910 296.000 1342.190 300.000 ;
    END
  END slave_data_wdata_to_inter_o[83]
  PIN slave_data_wdata_to_inter_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.350 296.000 1348.630 300.000 ;
    END
  END slave_data_wdata_to_inter_o[84]
  PIN slave_data_wdata_to_inter_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.790 296.000 1355.070 300.000 ;
    END
  END slave_data_wdata_to_inter_o[85]
  PIN slave_data_wdata_to_inter_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 296.000 1361.050 300.000 ;
    END
  END slave_data_wdata_to_inter_o[86]
  PIN slave_data_wdata_to_inter_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.210 296.000 1367.490 300.000 ;
    END
  END slave_data_wdata_to_inter_o[87]
  PIN slave_data_wdata_to_inter_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.650 296.000 1373.930 300.000 ;
    END
  END slave_data_wdata_to_inter_o[88]
  PIN slave_data_wdata_to_inter_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 296.000 1380.370 300.000 ;
    END
  END slave_data_wdata_to_inter_o[89]
  PIN slave_data_wdata_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 296.000 704.170 300.000 ;
    END
  END slave_data_wdata_to_inter_o[8]
  PIN slave_data_wdata_to_inter_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.070 296.000 1386.350 300.000 ;
    END
  END slave_data_wdata_to_inter_o[90]
  PIN slave_data_wdata_to_inter_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.510 296.000 1392.790 300.000 ;
    END
  END slave_data_wdata_to_inter_o[91]
  PIN slave_data_wdata_to_inter_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.950 296.000 1399.230 300.000 ;
    END
  END slave_data_wdata_to_inter_o[92]
  PIN slave_data_wdata_to_inter_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.390 296.000 1405.670 300.000 ;
    END
  END slave_data_wdata_to_inter_o[93]
  PIN slave_data_wdata_to_inter_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.370 296.000 1411.650 300.000 ;
    END
  END slave_data_wdata_to_inter_o[94]
  PIN slave_data_wdata_to_inter_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.810 296.000 1418.090 300.000 ;
    END
  END slave_data_wdata_to_inter_o[95]
  PIN slave_data_wdata_to_inter_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.250 296.000 1424.530 300.000 ;
    END
  END slave_data_wdata_to_inter_o[96]
  PIN slave_data_wdata_to_inter_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1430.690 296.000 1430.970 300.000 ;
    END
  END slave_data_wdata_to_inter_o[97]
  PIN slave_data_wdata_to_inter_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.130 296.000 1437.410 300.000 ;
    END
  END slave_data_wdata_to_inter_o[98]
  PIN slave_data_wdata_to_inter_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.110 296.000 1443.390 300.000 ;
    END
  END slave_data_wdata_to_inter_o[99]
  PIN slave_data_wdata_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 296.000 717.050 300.000 ;
    END
  END slave_data_wdata_to_inter_o[9]
  PIN slave_data_we_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 296.000 584.110 300.000 ;
    END
  END slave_data_we_to_inter_o[0]
  PIN slave_data_we_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 296.000 602.970 300.000 ;
    END
  END slave_data_we_to_inter_o[1]
  PIN slave_data_we_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 296.000 621.830 300.000 ;
    END
  END slave_data_we_to_inter_o[2]
  PIN slave_data_we_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 296.000 641.150 300.000 ;
    END
  END slave_data_we_to_inter_o[3]
  PIN txd_uart
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 13.640 1700.000 14.240 ;
    END
  END txd_uart
  PIN txd_uart_to_mem
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 19.080 1700.000 19.680 ;
    END
  END txd_uart_to_mem
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.990 0.000 1088.270 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.310 0.000 1038.590 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 0.000 621.370 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 0.000 740.510 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 0.000 770.410 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 0.000 859.650 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 0.000 889.550 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.170 0.000 919.450 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 0.000 949.350 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.870 0.000 1009.150 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 0.000 839.870 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 0.000 959.010 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.530 0.000 1018.810 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 0.000 611.250 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 0.000 849.990 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050 0.000 909.330 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.950 0.000 939.230 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 0.000 969.130 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 0.000 1028.930 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1694.180 288.405 ;
      LAYER met1 ;
        RECT 0.990 9.220 1699.170 299.840 ;
      LAYER met2 ;
        RECT 1.570 295.720 2.570 299.870 ;
        RECT 3.410 295.720 4.870 299.870 ;
        RECT 5.710 295.720 6.710 299.870 ;
        RECT 7.550 295.720 9.010 299.870 ;
        RECT 9.850 295.720 10.850 299.870 ;
        RECT 11.690 295.720 13.150 299.870 ;
        RECT 13.990 295.720 15.450 299.870 ;
        RECT 16.290 295.720 17.290 299.870 ;
        RECT 18.130 295.720 19.590 299.870 ;
        RECT 20.430 295.720 21.430 299.870 ;
        RECT 22.270 295.720 23.730 299.870 ;
        RECT 24.570 295.720 26.030 299.870 ;
        RECT 26.870 295.720 27.870 299.870 ;
        RECT 28.710 295.720 30.170 299.870 ;
        RECT 31.010 295.720 32.010 299.870 ;
        RECT 32.850 295.720 34.310 299.870 ;
        RECT 35.150 295.720 36.610 299.870 ;
        RECT 37.450 295.720 38.450 299.870 ;
        RECT 39.290 295.720 40.750 299.870 ;
        RECT 41.590 295.720 42.590 299.870 ;
        RECT 43.430 295.720 44.890 299.870 ;
        RECT 45.730 295.720 47.190 299.870 ;
        RECT 48.030 295.720 49.030 299.870 ;
        RECT 49.870 295.720 51.330 299.870 ;
        RECT 52.170 295.720 53.170 299.870 ;
        RECT 54.010 295.720 55.470 299.870 ;
        RECT 56.310 295.720 57.310 299.870 ;
        RECT 58.150 295.720 59.610 299.870 ;
        RECT 60.450 295.720 61.910 299.870 ;
        RECT 62.750 295.720 63.750 299.870 ;
        RECT 64.590 295.720 66.050 299.870 ;
        RECT 66.890 295.720 67.890 299.870 ;
        RECT 68.730 295.720 70.190 299.870 ;
        RECT 71.030 295.720 72.490 299.870 ;
        RECT 73.330 295.720 74.330 299.870 ;
        RECT 75.170 295.720 76.630 299.870 ;
        RECT 77.470 295.720 78.470 299.870 ;
        RECT 79.310 295.720 80.770 299.870 ;
        RECT 81.610 295.720 83.070 299.870 ;
        RECT 83.910 295.720 84.910 299.870 ;
        RECT 85.750 295.720 87.210 299.870 ;
        RECT 88.050 295.720 89.050 299.870 ;
        RECT 89.890 295.720 91.350 299.870 ;
        RECT 92.190 295.720 93.650 299.870 ;
        RECT 94.490 295.720 95.490 299.870 ;
        RECT 96.330 295.720 97.790 299.870 ;
        RECT 98.630 295.720 99.630 299.870 ;
        RECT 100.470 295.720 101.930 299.870 ;
        RECT 102.770 295.720 103.770 299.870 ;
        RECT 104.610 295.720 106.070 299.870 ;
        RECT 106.910 295.720 108.370 299.870 ;
        RECT 109.210 295.720 110.210 299.870 ;
        RECT 111.050 295.720 112.510 299.870 ;
        RECT 113.350 295.720 114.350 299.870 ;
        RECT 115.190 295.720 116.650 299.870 ;
        RECT 117.490 295.720 118.950 299.870 ;
        RECT 119.790 295.720 120.790 299.870 ;
        RECT 121.630 295.720 123.090 299.870 ;
        RECT 123.930 295.720 124.930 299.870 ;
        RECT 125.770 295.720 127.230 299.870 ;
        RECT 128.070 295.720 129.530 299.870 ;
        RECT 130.370 295.720 131.370 299.870 ;
        RECT 132.210 295.720 133.670 299.870 ;
        RECT 134.510 295.720 135.510 299.870 ;
        RECT 136.350 295.720 137.810 299.870 ;
        RECT 138.650 295.720 140.110 299.870 ;
        RECT 140.950 295.720 141.950 299.870 ;
        RECT 142.790 295.720 144.250 299.870 ;
        RECT 145.090 295.720 146.090 299.870 ;
        RECT 146.930 295.720 148.390 299.870 ;
        RECT 149.230 295.720 150.230 299.870 ;
        RECT 151.070 295.720 152.530 299.870 ;
        RECT 153.370 295.720 154.830 299.870 ;
        RECT 155.670 295.720 156.670 299.870 ;
        RECT 157.510 295.720 158.970 299.870 ;
        RECT 159.810 295.720 160.810 299.870 ;
        RECT 161.650 295.720 163.110 299.870 ;
        RECT 163.950 295.720 165.410 299.870 ;
        RECT 166.250 295.720 167.250 299.870 ;
        RECT 168.090 295.720 169.550 299.870 ;
        RECT 170.390 295.720 171.390 299.870 ;
        RECT 172.230 295.720 173.690 299.870 ;
        RECT 174.530 295.720 175.990 299.870 ;
        RECT 176.830 295.720 177.830 299.870 ;
        RECT 178.670 295.720 180.130 299.870 ;
        RECT 180.970 295.720 181.970 299.870 ;
        RECT 182.810 295.720 184.270 299.870 ;
        RECT 185.110 295.720 186.570 299.870 ;
        RECT 187.410 295.720 188.410 299.870 ;
        RECT 189.250 295.720 190.710 299.870 ;
        RECT 191.550 295.720 192.550 299.870 ;
        RECT 193.390 295.720 194.850 299.870 ;
        RECT 195.690 295.720 196.690 299.870 ;
        RECT 197.530 295.720 198.990 299.870 ;
        RECT 199.830 295.720 201.290 299.870 ;
        RECT 202.130 295.720 203.130 299.870 ;
        RECT 203.970 295.720 205.430 299.870 ;
        RECT 206.270 295.720 207.270 299.870 ;
        RECT 208.110 295.720 209.570 299.870 ;
        RECT 210.410 295.720 211.870 299.870 ;
        RECT 212.710 295.720 213.710 299.870 ;
        RECT 214.550 295.720 216.010 299.870 ;
        RECT 216.850 295.720 217.850 299.870 ;
        RECT 218.690 295.720 220.150 299.870 ;
        RECT 220.990 295.720 222.450 299.870 ;
        RECT 223.290 295.720 224.290 299.870 ;
        RECT 225.130 295.720 226.590 299.870 ;
        RECT 227.430 295.720 228.430 299.870 ;
        RECT 229.270 295.720 230.730 299.870 ;
        RECT 231.570 295.720 233.030 299.870 ;
        RECT 233.870 295.720 234.870 299.870 ;
        RECT 235.710 295.720 237.170 299.870 ;
        RECT 238.010 295.720 239.010 299.870 ;
        RECT 239.850 295.720 241.310 299.870 ;
        RECT 242.150 295.720 243.610 299.870 ;
        RECT 244.450 295.720 245.450 299.870 ;
        RECT 246.290 295.720 247.750 299.870 ;
        RECT 248.590 295.720 249.590 299.870 ;
        RECT 250.430 295.720 251.890 299.870 ;
        RECT 252.730 295.720 253.730 299.870 ;
        RECT 254.570 295.720 256.030 299.870 ;
        RECT 256.870 295.720 258.330 299.870 ;
        RECT 259.170 295.720 260.170 299.870 ;
        RECT 261.010 295.720 262.470 299.870 ;
        RECT 263.310 295.720 264.310 299.870 ;
        RECT 265.150 295.720 266.610 299.870 ;
        RECT 267.450 295.720 268.910 299.870 ;
        RECT 269.750 295.720 270.750 299.870 ;
        RECT 271.590 295.720 273.050 299.870 ;
        RECT 273.890 295.720 274.890 299.870 ;
        RECT 275.730 295.720 277.190 299.870 ;
        RECT 278.030 295.720 279.490 299.870 ;
        RECT 280.330 295.720 281.330 299.870 ;
        RECT 282.170 295.720 283.630 299.870 ;
        RECT 284.470 295.720 285.470 299.870 ;
        RECT 286.310 295.720 287.770 299.870 ;
        RECT 288.610 295.720 290.070 299.870 ;
        RECT 290.910 295.720 291.910 299.870 ;
        RECT 292.750 295.720 294.210 299.870 ;
        RECT 295.050 295.720 296.050 299.870 ;
        RECT 296.890 295.720 298.350 299.870 ;
        RECT 299.190 295.720 300.190 299.870 ;
        RECT 301.030 295.720 302.490 299.870 ;
        RECT 303.330 295.720 304.790 299.870 ;
        RECT 305.630 295.720 306.630 299.870 ;
        RECT 307.470 295.720 308.930 299.870 ;
        RECT 309.770 295.720 310.770 299.870 ;
        RECT 311.610 295.720 313.070 299.870 ;
        RECT 313.910 295.720 315.370 299.870 ;
        RECT 316.210 295.720 317.210 299.870 ;
        RECT 318.050 295.720 319.510 299.870 ;
        RECT 320.350 295.720 321.350 299.870 ;
        RECT 322.190 295.720 323.650 299.870 ;
        RECT 324.490 295.720 325.950 299.870 ;
        RECT 326.790 295.720 327.790 299.870 ;
        RECT 328.630 295.720 330.090 299.870 ;
        RECT 330.930 295.720 331.930 299.870 ;
        RECT 332.770 295.720 334.230 299.870 ;
        RECT 335.070 295.720 336.530 299.870 ;
        RECT 337.370 295.720 338.370 299.870 ;
        RECT 339.210 295.720 340.670 299.870 ;
        RECT 341.510 295.720 342.510 299.870 ;
        RECT 343.350 295.720 344.810 299.870 ;
        RECT 345.650 295.720 346.650 299.870 ;
        RECT 347.490 295.720 348.950 299.870 ;
        RECT 349.790 295.720 351.250 299.870 ;
        RECT 352.090 295.720 353.090 299.870 ;
        RECT 353.930 295.720 355.390 299.870 ;
        RECT 356.230 295.720 357.230 299.870 ;
        RECT 358.070 295.720 359.530 299.870 ;
        RECT 360.370 295.720 361.830 299.870 ;
        RECT 362.670 295.720 363.670 299.870 ;
        RECT 364.510 295.720 365.970 299.870 ;
        RECT 366.810 295.720 367.810 299.870 ;
        RECT 368.650 295.720 370.110 299.870 ;
        RECT 370.950 295.720 372.410 299.870 ;
        RECT 373.250 295.720 374.250 299.870 ;
        RECT 375.090 295.720 376.550 299.870 ;
        RECT 377.390 295.720 378.390 299.870 ;
        RECT 379.230 295.720 380.690 299.870 ;
        RECT 381.530 295.720 382.990 299.870 ;
        RECT 383.830 295.720 384.830 299.870 ;
        RECT 385.670 295.720 387.130 299.870 ;
        RECT 387.970 295.720 388.970 299.870 ;
        RECT 389.810 295.720 391.270 299.870 ;
        RECT 392.110 295.720 393.110 299.870 ;
        RECT 393.950 295.720 395.410 299.870 ;
        RECT 396.250 295.720 397.710 299.870 ;
        RECT 398.550 295.720 399.550 299.870 ;
        RECT 400.390 295.720 401.850 299.870 ;
        RECT 402.690 295.720 403.690 299.870 ;
        RECT 404.530 295.720 405.990 299.870 ;
        RECT 406.830 295.720 408.290 299.870 ;
        RECT 409.130 295.720 410.130 299.870 ;
        RECT 410.970 295.720 412.430 299.870 ;
        RECT 413.270 295.720 414.270 299.870 ;
        RECT 415.110 295.720 416.570 299.870 ;
        RECT 417.410 295.720 418.870 299.870 ;
        RECT 419.710 295.720 420.710 299.870 ;
        RECT 421.550 295.720 423.010 299.870 ;
        RECT 423.850 295.720 424.850 299.870 ;
        RECT 425.690 295.720 427.150 299.870 ;
        RECT 427.990 295.720 429.450 299.870 ;
        RECT 430.290 295.720 431.290 299.870 ;
        RECT 432.130 295.720 433.590 299.870 ;
        RECT 434.430 295.720 435.430 299.870 ;
        RECT 436.270 295.720 437.730 299.870 ;
        RECT 438.570 295.720 439.570 299.870 ;
        RECT 440.410 295.720 441.870 299.870 ;
        RECT 442.710 295.720 444.170 299.870 ;
        RECT 445.010 295.720 446.010 299.870 ;
        RECT 446.850 295.720 448.310 299.870 ;
        RECT 449.150 295.720 450.150 299.870 ;
        RECT 450.990 295.720 452.450 299.870 ;
        RECT 453.290 295.720 454.750 299.870 ;
        RECT 455.590 295.720 456.590 299.870 ;
        RECT 457.430 295.720 458.890 299.870 ;
        RECT 459.730 295.720 460.730 299.870 ;
        RECT 461.570 295.720 463.030 299.870 ;
        RECT 463.870 295.720 465.330 299.870 ;
        RECT 466.170 295.720 467.170 299.870 ;
        RECT 468.010 295.720 469.470 299.870 ;
        RECT 470.310 295.720 471.310 299.870 ;
        RECT 472.150 295.720 473.610 299.870 ;
        RECT 474.450 295.720 475.910 299.870 ;
        RECT 476.750 295.720 477.750 299.870 ;
        RECT 478.590 295.720 480.050 299.870 ;
        RECT 480.890 295.720 481.890 299.870 ;
        RECT 482.730 295.720 484.190 299.870 ;
        RECT 485.030 295.720 486.490 299.870 ;
        RECT 487.330 295.720 488.330 299.870 ;
        RECT 489.170 295.720 490.630 299.870 ;
        RECT 491.470 295.720 492.470 299.870 ;
        RECT 493.310 295.720 494.770 299.870 ;
        RECT 495.610 295.720 496.610 299.870 ;
        RECT 497.450 295.720 498.910 299.870 ;
        RECT 499.750 295.720 501.210 299.870 ;
        RECT 502.050 295.720 503.050 299.870 ;
        RECT 503.890 295.720 505.350 299.870 ;
        RECT 506.190 295.720 507.190 299.870 ;
        RECT 508.030 295.720 509.490 299.870 ;
        RECT 510.330 295.720 511.790 299.870 ;
        RECT 512.630 295.720 513.630 299.870 ;
        RECT 514.470 295.720 515.930 299.870 ;
        RECT 516.770 295.720 517.770 299.870 ;
        RECT 518.610 295.720 520.070 299.870 ;
        RECT 520.910 295.720 522.370 299.870 ;
        RECT 523.210 295.720 524.210 299.870 ;
        RECT 525.050 295.720 526.510 299.870 ;
        RECT 527.350 295.720 528.350 299.870 ;
        RECT 529.190 295.720 530.650 299.870 ;
        RECT 531.490 295.720 532.950 299.870 ;
        RECT 533.790 295.720 534.790 299.870 ;
        RECT 535.630 295.720 537.090 299.870 ;
        RECT 537.930 295.720 538.930 299.870 ;
        RECT 539.770 295.720 541.230 299.870 ;
        RECT 542.070 295.720 543.070 299.870 ;
        RECT 543.910 295.720 545.370 299.870 ;
        RECT 546.210 295.720 547.670 299.870 ;
        RECT 548.510 295.720 549.510 299.870 ;
        RECT 550.350 295.720 551.810 299.870 ;
        RECT 552.650 295.720 553.650 299.870 ;
        RECT 554.490 295.720 555.950 299.870 ;
        RECT 556.790 295.720 558.250 299.870 ;
        RECT 559.090 295.720 560.090 299.870 ;
        RECT 560.930 295.720 562.390 299.870 ;
        RECT 563.230 295.720 564.230 299.870 ;
        RECT 565.070 295.720 566.530 299.870 ;
        RECT 567.370 295.720 568.830 299.870 ;
        RECT 569.670 295.720 570.670 299.870 ;
        RECT 571.510 295.720 572.970 299.870 ;
        RECT 573.810 295.720 574.810 299.870 ;
        RECT 575.650 295.720 577.110 299.870 ;
        RECT 577.950 295.720 579.410 299.870 ;
        RECT 580.250 295.720 581.250 299.870 ;
        RECT 582.090 295.720 583.550 299.870 ;
        RECT 584.390 295.720 585.390 299.870 ;
        RECT 586.230 295.720 587.690 299.870 ;
        RECT 588.530 295.720 589.530 299.870 ;
        RECT 590.370 295.720 591.830 299.870 ;
        RECT 592.670 295.720 594.130 299.870 ;
        RECT 594.970 295.720 595.970 299.870 ;
        RECT 596.810 295.720 598.270 299.870 ;
        RECT 599.110 295.720 600.110 299.870 ;
        RECT 600.950 295.720 602.410 299.870 ;
        RECT 603.250 295.720 604.710 299.870 ;
        RECT 605.550 295.720 606.550 299.870 ;
        RECT 607.390 295.720 608.850 299.870 ;
        RECT 609.690 295.720 610.690 299.870 ;
        RECT 611.530 295.720 612.990 299.870 ;
        RECT 613.830 295.720 615.290 299.870 ;
        RECT 616.130 295.720 617.130 299.870 ;
        RECT 617.970 295.720 619.430 299.870 ;
        RECT 620.270 295.720 621.270 299.870 ;
        RECT 622.110 295.720 623.570 299.870 ;
        RECT 624.410 295.720 625.870 299.870 ;
        RECT 626.710 295.720 627.710 299.870 ;
        RECT 628.550 295.720 630.010 299.870 ;
        RECT 630.850 295.720 631.850 299.870 ;
        RECT 632.690 295.720 634.150 299.870 ;
        RECT 634.990 295.720 635.990 299.870 ;
        RECT 636.830 295.720 638.290 299.870 ;
        RECT 639.130 295.720 640.590 299.870 ;
        RECT 641.430 295.720 642.430 299.870 ;
        RECT 643.270 295.720 644.730 299.870 ;
        RECT 645.570 295.720 646.570 299.870 ;
        RECT 647.410 295.720 648.870 299.870 ;
        RECT 649.710 295.720 651.170 299.870 ;
        RECT 652.010 295.720 653.010 299.870 ;
        RECT 653.850 295.720 655.310 299.870 ;
        RECT 656.150 295.720 657.150 299.870 ;
        RECT 657.990 295.720 659.450 299.870 ;
        RECT 660.290 295.720 661.750 299.870 ;
        RECT 662.590 295.720 663.590 299.870 ;
        RECT 664.430 295.720 665.890 299.870 ;
        RECT 666.730 295.720 667.730 299.870 ;
        RECT 668.570 295.720 670.030 299.870 ;
        RECT 670.870 295.720 672.330 299.870 ;
        RECT 673.170 295.720 674.170 299.870 ;
        RECT 675.010 295.720 676.470 299.870 ;
        RECT 677.310 295.720 678.310 299.870 ;
        RECT 679.150 295.720 680.610 299.870 ;
        RECT 681.450 295.720 682.450 299.870 ;
        RECT 683.290 295.720 684.750 299.870 ;
        RECT 685.590 295.720 687.050 299.870 ;
        RECT 687.890 295.720 688.890 299.870 ;
        RECT 689.730 295.720 691.190 299.870 ;
        RECT 692.030 295.720 693.030 299.870 ;
        RECT 693.870 295.720 695.330 299.870 ;
        RECT 696.170 295.720 697.630 299.870 ;
        RECT 698.470 295.720 699.470 299.870 ;
        RECT 700.310 295.720 701.770 299.870 ;
        RECT 702.610 295.720 703.610 299.870 ;
        RECT 704.450 295.720 705.910 299.870 ;
        RECT 706.750 295.720 708.210 299.870 ;
        RECT 709.050 295.720 710.050 299.870 ;
        RECT 710.890 295.720 712.350 299.870 ;
        RECT 713.190 295.720 714.190 299.870 ;
        RECT 715.030 295.720 716.490 299.870 ;
        RECT 717.330 295.720 718.790 299.870 ;
        RECT 719.630 295.720 720.630 299.870 ;
        RECT 721.470 295.720 722.930 299.870 ;
        RECT 723.770 295.720 724.770 299.870 ;
        RECT 725.610 295.720 727.070 299.870 ;
        RECT 727.910 295.720 729.370 299.870 ;
        RECT 730.210 295.720 731.210 299.870 ;
        RECT 732.050 295.720 733.510 299.870 ;
        RECT 734.350 295.720 735.350 299.870 ;
        RECT 736.190 295.720 737.650 299.870 ;
        RECT 738.490 295.720 739.490 299.870 ;
        RECT 740.330 295.720 741.790 299.870 ;
        RECT 742.630 295.720 744.090 299.870 ;
        RECT 744.930 295.720 745.930 299.870 ;
        RECT 746.770 295.720 748.230 299.870 ;
        RECT 749.070 295.720 750.070 299.870 ;
        RECT 750.910 295.720 752.370 299.870 ;
        RECT 753.210 295.720 754.670 299.870 ;
        RECT 755.510 295.720 756.510 299.870 ;
        RECT 757.350 295.720 758.810 299.870 ;
        RECT 759.650 295.720 760.650 299.870 ;
        RECT 761.490 295.720 762.950 299.870 ;
        RECT 763.790 295.720 765.250 299.870 ;
        RECT 766.090 295.720 767.090 299.870 ;
        RECT 767.930 295.720 769.390 299.870 ;
        RECT 770.230 295.720 771.230 299.870 ;
        RECT 772.070 295.720 773.530 299.870 ;
        RECT 774.370 295.720 775.830 299.870 ;
        RECT 776.670 295.720 777.670 299.870 ;
        RECT 778.510 295.720 779.970 299.870 ;
        RECT 780.810 295.720 781.810 299.870 ;
        RECT 782.650 295.720 784.110 299.870 ;
        RECT 784.950 295.720 785.950 299.870 ;
        RECT 786.790 295.720 788.250 299.870 ;
        RECT 789.090 295.720 790.550 299.870 ;
        RECT 791.390 295.720 792.390 299.870 ;
        RECT 793.230 295.720 794.690 299.870 ;
        RECT 795.530 295.720 796.530 299.870 ;
        RECT 797.370 295.720 798.830 299.870 ;
        RECT 799.670 295.720 801.130 299.870 ;
        RECT 801.970 295.720 802.970 299.870 ;
        RECT 803.810 295.720 805.270 299.870 ;
        RECT 806.110 295.720 807.110 299.870 ;
        RECT 807.950 295.720 809.410 299.870 ;
        RECT 810.250 295.720 811.710 299.870 ;
        RECT 812.550 295.720 813.550 299.870 ;
        RECT 814.390 295.720 815.850 299.870 ;
        RECT 816.690 295.720 817.690 299.870 ;
        RECT 818.530 295.720 819.990 299.870 ;
        RECT 820.830 295.720 822.290 299.870 ;
        RECT 823.130 295.720 824.130 299.870 ;
        RECT 824.970 295.720 826.430 299.870 ;
        RECT 827.270 295.720 828.270 299.870 ;
        RECT 829.110 295.720 830.570 299.870 ;
        RECT 831.410 295.720 832.410 299.870 ;
        RECT 833.250 295.720 834.710 299.870 ;
        RECT 835.550 295.720 837.010 299.870 ;
        RECT 837.850 295.720 838.850 299.870 ;
        RECT 839.690 295.720 841.150 299.870 ;
        RECT 841.990 295.720 842.990 299.870 ;
        RECT 843.830 295.720 845.290 299.870 ;
        RECT 846.130 295.720 847.590 299.870 ;
        RECT 848.430 295.720 849.430 299.870 ;
        RECT 850.270 295.720 851.730 299.870 ;
        RECT 852.570 295.720 853.570 299.870 ;
        RECT 854.410 295.720 855.870 299.870 ;
        RECT 856.710 295.720 858.170 299.870 ;
        RECT 859.010 295.720 860.010 299.870 ;
        RECT 860.850 295.720 862.310 299.870 ;
        RECT 863.150 295.720 864.150 299.870 ;
        RECT 864.990 295.720 866.450 299.870 ;
        RECT 867.290 295.720 868.750 299.870 ;
        RECT 869.590 295.720 870.590 299.870 ;
        RECT 871.430 295.720 872.890 299.870 ;
        RECT 873.730 295.720 874.730 299.870 ;
        RECT 875.570 295.720 877.030 299.870 ;
        RECT 877.870 295.720 878.870 299.870 ;
        RECT 879.710 295.720 881.170 299.870 ;
        RECT 882.010 295.720 883.470 299.870 ;
        RECT 884.310 295.720 885.310 299.870 ;
        RECT 886.150 295.720 887.610 299.870 ;
        RECT 888.450 295.720 889.450 299.870 ;
        RECT 890.290 295.720 891.750 299.870 ;
        RECT 892.590 295.720 894.050 299.870 ;
        RECT 894.890 295.720 895.890 299.870 ;
        RECT 896.730 295.720 898.190 299.870 ;
        RECT 899.030 295.720 900.030 299.870 ;
        RECT 900.870 295.720 902.330 299.870 ;
        RECT 903.170 295.720 904.630 299.870 ;
        RECT 905.470 295.720 906.470 299.870 ;
        RECT 907.310 295.720 908.770 299.870 ;
        RECT 909.610 295.720 910.610 299.870 ;
        RECT 911.450 295.720 912.910 299.870 ;
        RECT 913.750 295.720 915.210 299.870 ;
        RECT 916.050 295.720 917.050 299.870 ;
        RECT 917.890 295.720 919.350 299.870 ;
        RECT 920.190 295.720 921.190 299.870 ;
        RECT 922.030 295.720 923.490 299.870 ;
        RECT 924.330 295.720 925.330 299.870 ;
        RECT 926.170 295.720 927.630 299.870 ;
        RECT 928.470 295.720 929.930 299.870 ;
        RECT 930.770 295.720 931.770 299.870 ;
        RECT 932.610 295.720 934.070 299.870 ;
        RECT 934.910 295.720 935.910 299.870 ;
        RECT 936.750 295.720 938.210 299.870 ;
        RECT 939.050 295.720 940.510 299.870 ;
        RECT 941.350 295.720 942.350 299.870 ;
        RECT 943.190 295.720 944.650 299.870 ;
        RECT 945.490 295.720 946.490 299.870 ;
        RECT 947.330 295.720 948.790 299.870 ;
        RECT 949.630 295.720 951.090 299.870 ;
        RECT 951.930 295.720 952.930 299.870 ;
        RECT 953.770 295.720 955.230 299.870 ;
        RECT 956.070 295.720 957.070 299.870 ;
        RECT 957.910 295.720 959.370 299.870 ;
        RECT 960.210 295.720 961.670 299.870 ;
        RECT 962.510 295.720 963.510 299.870 ;
        RECT 964.350 295.720 965.810 299.870 ;
        RECT 966.650 295.720 967.650 299.870 ;
        RECT 968.490 295.720 969.950 299.870 ;
        RECT 970.790 295.720 972.250 299.870 ;
        RECT 973.090 295.720 974.090 299.870 ;
        RECT 974.930 295.720 976.390 299.870 ;
        RECT 977.230 295.720 978.230 299.870 ;
        RECT 979.070 295.720 980.530 299.870 ;
        RECT 981.370 295.720 982.370 299.870 ;
        RECT 983.210 295.720 984.670 299.870 ;
        RECT 985.510 295.720 986.970 299.870 ;
        RECT 987.810 295.720 988.810 299.870 ;
        RECT 989.650 295.720 991.110 299.870 ;
        RECT 991.950 295.720 992.950 299.870 ;
        RECT 993.790 295.720 995.250 299.870 ;
        RECT 996.090 295.720 997.550 299.870 ;
        RECT 998.390 295.720 999.390 299.870 ;
        RECT 1000.230 295.720 1001.690 299.870 ;
        RECT 1002.530 295.720 1003.530 299.870 ;
        RECT 1004.370 295.720 1005.830 299.870 ;
        RECT 1006.670 295.720 1008.130 299.870 ;
        RECT 1008.970 295.720 1009.970 299.870 ;
        RECT 1010.810 295.720 1012.270 299.870 ;
        RECT 1013.110 295.720 1014.110 299.870 ;
        RECT 1014.950 295.720 1016.410 299.870 ;
        RECT 1017.250 295.720 1018.710 299.870 ;
        RECT 1019.550 295.720 1020.550 299.870 ;
        RECT 1021.390 295.720 1022.850 299.870 ;
        RECT 1023.690 295.720 1024.690 299.870 ;
        RECT 1025.530 295.720 1026.990 299.870 ;
        RECT 1027.830 295.720 1028.830 299.870 ;
        RECT 1029.670 295.720 1031.130 299.870 ;
        RECT 1031.970 295.720 1033.430 299.870 ;
        RECT 1034.270 295.720 1035.270 299.870 ;
        RECT 1036.110 295.720 1037.570 299.870 ;
        RECT 1038.410 295.720 1039.410 299.870 ;
        RECT 1040.250 295.720 1041.710 299.870 ;
        RECT 1042.550 295.720 1044.010 299.870 ;
        RECT 1044.850 295.720 1045.850 299.870 ;
        RECT 1046.690 295.720 1048.150 299.870 ;
        RECT 1048.990 295.720 1049.990 299.870 ;
        RECT 1050.830 295.720 1052.290 299.870 ;
        RECT 1053.130 295.720 1054.590 299.870 ;
        RECT 1055.430 295.720 1056.430 299.870 ;
        RECT 1057.270 295.720 1058.730 299.870 ;
        RECT 1059.570 295.720 1060.570 299.870 ;
        RECT 1061.410 295.720 1062.870 299.870 ;
        RECT 1063.710 295.720 1065.170 299.870 ;
        RECT 1066.010 295.720 1067.010 299.870 ;
        RECT 1067.850 295.720 1069.310 299.870 ;
        RECT 1070.150 295.720 1071.150 299.870 ;
        RECT 1071.990 295.720 1073.450 299.870 ;
        RECT 1074.290 295.720 1075.290 299.870 ;
        RECT 1076.130 295.720 1077.590 299.870 ;
        RECT 1078.430 295.720 1079.890 299.870 ;
        RECT 1080.730 295.720 1081.730 299.870 ;
        RECT 1082.570 295.720 1084.030 299.870 ;
        RECT 1084.870 295.720 1085.870 299.870 ;
        RECT 1086.710 295.720 1088.170 299.870 ;
        RECT 1089.010 295.720 1090.470 299.870 ;
        RECT 1091.310 295.720 1092.310 299.870 ;
        RECT 1093.150 295.720 1094.610 299.870 ;
        RECT 1095.450 295.720 1096.450 299.870 ;
        RECT 1097.290 295.720 1098.750 299.870 ;
        RECT 1099.590 295.720 1101.050 299.870 ;
        RECT 1101.890 295.720 1102.890 299.870 ;
        RECT 1103.730 295.720 1105.190 299.870 ;
        RECT 1106.030 295.720 1107.030 299.870 ;
        RECT 1107.870 295.720 1109.330 299.870 ;
        RECT 1110.170 295.720 1111.630 299.870 ;
        RECT 1112.470 295.720 1113.470 299.870 ;
        RECT 1114.310 295.720 1115.770 299.870 ;
        RECT 1116.610 295.720 1117.610 299.870 ;
        RECT 1118.450 295.720 1119.910 299.870 ;
        RECT 1120.750 295.720 1121.750 299.870 ;
        RECT 1122.590 295.720 1124.050 299.870 ;
        RECT 1124.890 295.720 1126.350 299.870 ;
        RECT 1127.190 295.720 1128.190 299.870 ;
        RECT 1129.030 295.720 1130.490 299.870 ;
        RECT 1131.330 295.720 1132.330 299.870 ;
        RECT 1133.170 295.720 1134.630 299.870 ;
        RECT 1135.470 295.720 1136.930 299.870 ;
        RECT 1137.770 295.720 1138.770 299.870 ;
        RECT 1139.610 295.720 1141.070 299.870 ;
        RECT 1141.910 295.720 1142.910 299.870 ;
        RECT 1143.750 295.720 1145.210 299.870 ;
        RECT 1146.050 295.720 1147.510 299.870 ;
        RECT 1148.350 295.720 1149.350 299.870 ;
        RECT 1150.190 295.720 1151.650 299.870 ;
        RECT 1152.490 295.720 1153.490 299.870 ;
        RECT 1154.330 295.720 1155.790 299.870 ;
        RECT 1156.630 295.720 1158.090 299.870 ;
        RECT 1158.930 295.720 1159.930 299.870 ;
        RECT 1160.770 295.720 1162.230 299.870 ;
        RECT 1163.070 295.720 1164.070 299.870 ;
        RECT 1164.910 295.720 1166.370 299.870 ;
        RECT 1167.210 295.720 1168.210 299.870 ;
        RECT 1169.050 295.720 1170.510 299.870 ;
        RECT 1171.350 295.720 1172.810 299.870 ;
        RECT 1173.650 295.720 1174.650 299.870 ;
        RECT 1175.490 295.720 1176.950 299.870 ;
        RECT 1177.790 295.720 1178.790 299.870 ;
        RECT 1179.630 295.720 1181.090 299.870 ;
        RECT 1181.930 295.720 1183.390 299.870 ;
        RECT 1184.230 295.720 1185.230 299.870 ;
        RECT 1186.070 295.720 1187.530 299.870 ;
        RECT 1188.370 295.720 1189.370 299.870 ;
        RECT 1190.210 295.720 1191.670 299.870 ;
        RECT 1192.510 295.720 1193.970 299.870 ;
        RECT 1194.810 295.720 1195.810 299.870 ;
        RECT 1196.650 295.720 1198.110 299.870 ;
        RECT 1198.950 295.720 1199.950 299.870 ;
        RECT 1200.790 295.720 1202.250 299.870 ;
        RECT 1203.090 295.720 1204.550 299.870 ;
        RECT 1205.390 295.720 1206.390 299.870 ;
        RECT 1207.230 295.720 1208.690 299.870 ;
        RECT 1209.530 295.720 1210.530 299.870 ;
        RECT 1211.370 295.720 1212.830 299.870 ;
        RECT 1213.670 295.720 1215.130 299.870 ;
        RECT 1215.970 295.720 1216.970 299.870 ;
        RECT 1217.810 295.720 1219.270 299.870 ;
        RECT 1220.110 295.720 1221.110 299.870 ;
        RECT 1221.950 295.720 1223.410 299.870 ;
        RECT 1224.250 295.720 1225.250 299.870 ;
        RECT 1226.090 295.720 1227.550 299.870 ;
        RECT 1228.390 295.720 1229.850 299.870 ;
        RECT 1230.690 295.720 1231.690 299.870 ;
        RECT 1232.530 295.720 1233.990 299.870 ;
        RECT 1234.830 295.720 1235.830 299.870 ;
        RECT 1236.670 295.720 1238.130 299.870 ;
        RECT 1238.970 295.720 1240.430 299.870 ;
        RECT 1241.270 295.720 1242.270 299.870 ;
        RECT 1243.110 295.720 1244.570 299.870 ;
        RECT 1245.410 295.720 1246.410 299.870 ;
        RECT 1247.250 295.720 1248.710 299.870 ;
        RECT 1249.550 295.720 1251.010 299.870 ;
        RECT 1251.850 295.720 1252.850 299.870 ;
        RECT 1253.690 295.720 1255.150 299.870 ;
        RECT 1255.990 295.720 1256.990 299.870 ;
        RECT 1257.830 295.720 1259.290 299.870 ;
        RECT 1260.130 295.720 1261.590 299.870 ;
        RECT 1262.430 295.720 1263.430 299.870 ;
        RECT 1264.270 295.720 1265.730 299.870 ;
        RECT 1266.570 295.720 1267.570 299.870 ;
        RECT 1268.410 295.720 1269.870 299.870 ;
        RECT 1270.710 295.720 1271.710 299.870 ;
        RECT 1272.550 295.720 1274.010 299.870 ;
        RECT 1274.850 295.720 1276.310 299.870 ;
        RECT 1277.150 295.720 1278.150 299.870 ;
        RECT 1278.990 295.720 1280.450 299.870 ;
        RECT 1281.290 295.720 1282.290 299.870 ;
        RECT 1283.130 295.720 1284.590 299.870 ;
        RECT 1285.430 295.720 1286.890 299.870 ;
        RECT 1287.730 295.720 1288.730 299.870 ;
        RECT 1289.570 295.720 1291.030 299.870 ;
        RECT 1291.870 295.720 1292.870 299.870 ;
        RECT 1293.710 295.720 1295.170 299.870 ;
        RECT 1296.010 295.720 1297.470 299.870 ;
        RECT 1298.310 295.720 1299.310 299.870 ;
        RECT 1300.150 295.720 1301.610 299.870 ;
        RECT 1302.450 295.720 1303.450 299.870 ;
        RECT 1304.290 295.720 1305.750 299.870 ;
        RECT 1306.590 295.720 1308.050 299.870 ;
        RECT 1308.890 295.720 1309.890 299.870 ;
        RECT 1310.730 295.720 1312.190 299.870 ;
        RECT 1313.030 295.720 1314.030 299.870 ;
        RECT 1314.870 295.720 1316.330 299.870 ;
        RECT 1317.170 295.720 1318.170 299.870 ;
        RECT 1319.010 295.720 1320.470 299.870 ;
        RECT 1321.310 295.720 1322.770 299.870 ;
        RECT 1323.610 295.720 1324.610 299.870 ;
        RECT 1325.450 295.720 1326.910 299.870 ;
        RECT 1327.750 295.720 1328.750 299.870 ;
        RECT 1329.590 295.720 1331.050 299.870 ;
        RECT 1331.890 295.720 1333.350 299.870 ;
        RECT 1334.190 295.720 1335.190 299.870 ;
        RECT 1336.030 295.720 1337.490 299.870 ;
        RECT 1338.330 295.720 1339.330 299.870 ;
        RECT 1340.170 295.720 1341.630 299.870 ;
        RECT 1342.470 295.720 1343.930 299.870 ;
        RECT 1344.770 295.720 1345.770 299.870 ;
        RECT 1346.610 295.720 1348.070 299.870 ;
        RECT 1348.910 295.720 1349.910 299.870 ;
        RECT 1350.750 295.720 1352.210 299.870 ;
        RECT 1353.050 295.720 1354.510 299.870 ;
        RECT 1355.350 295.720 1356.350 299.870 ;
        RECT 1357.190 295.720 1358.650 299.870 ;
        RECT 1359.490 295.720 1360.490 299.870 ;
        RECT 1361.330 295.720 1362.790 299.870 ;
        RECT 1363.630 295.720 1364.630 299.870 ;
        RECT 1365.470 295.720 1366.930 299.870 ;
        RECT 1367.770 295.720 1369.230 299.870 ;
        RECT 1370.070 295.720 1371.070 299.870 ;
        RECT 1371.910 295.720 1373.370 299.870 ;
        RECT 1374.210 295.720 1375.210 299.870 ;
        RECT 1376.050 295.720 1377.510 299.870 ;
        RECT 1378.350 295.720 1379.810 299.870 ;
        RECT 1380.650 295.720 1381.650 299.870 ;
        RECT 1382.490 295.720 1383.950 299.870 ;
        RECT 1384.790 295.720 1385.790 299.870 ;
        RECT 1386.630 295.720 1388.090 299.870 ;
        RECT 1388.930 295.720 1390.390 299.870 ;
        RECT 1391.230 295.720 1392.230 299.870 ;
        RECT 1393.070 295.720 1394.530 299.870 ;
        RECT 1395.370 295.720 1396.370 299.870 ;
        RECT 1397.210 295.720 1398.670 299.870 ;
        RECT 1399.510 295.720 1400.970 299.870 ;
        RECT 1401.810 295.720 1402.810 299.870 ;
        RECT 1403.650 295.720 1405.110 299.870 ;
        RECT 1405.950 295.720 1406.950 299.870 ;
        RECT 1407.790 295.720 1409.250 299.870 ;
        RECT 1410.090 295.720 1411.090 299.870 ;
        RECT 1411.930 295.720 1413.390 299.870 ;
        RECT 1414.230 295.720 1415.690 299.870 ;
        RECT 1416.530 295.720 1417.530 299.870 ;
        RECT 1418.370 295.720 1419.830 299.870 ;
        RECT 1420.670 295.720 1421.670 299.870 ;
        RECT 1422.510 295.720 1423.970 299.870 ;
        RECT 1424.810 295.720 1426.270 299.870 ;
        RECT 1427.110 295.720 1428.110 299.870 ;
        RECT 1428.950 295.720 1430.410 299.870 ;
        RECT 1431.250 295.720 1432.250 299.870 ;
        RECT 1433.090 295.720 1434.550 299.870 ;
        RECT 1435.390 295.720 1436.850 299.870 ;
        RECT 1437.690 295.720 1438.690 299.870 ;
        RECT 1439.530 295.720 1440.990 299.870 ;
        RECT 1441.830 295.720 1442.830 299.870 ;
        RECT 1443.670 295.720 1445.130 299.870 ;
        RECT 1445.970 295.720 1447.430 299.870 ;
        RECT 1448.270 295.720 1449.270 299.870 ;
        RECT 1450.110 295.720 1451.570 299.870 ;
        RECT 1452.410 295.720 1453.410 299.870 ;
        RECT 1454.250 295.720 1455.710 299.870 ;
        RECT 1456.550 295.720 1458.010 299.870 ;
        RECT 1458.850 295.720 1459.850 299.870 ;
        RECT 1460.690 295.720 1462.150 299.870 ;
        RECT 1462.990 295.720 1463.990 299.870 ;
        RECT 1464.830 295.720 1466.290 299.870 ;
        RECT 1467.130 295.720 1468.130 299.870 ;
        RECT 1468.970 295.720 1470.430 299.870 ;
        RECT 1471.270 295.720 1472.730 299.870 ;
        RECT 1473.570 295.720 1474.570 299.870 ;
        RECT 1475.410 295.720 1476.870 299.870 ;
        RECT 1477.710 295.720 1478.710 299.870 ;
        RECT 1479.550 295.720 1481.010 299.870 ;
        RECT 1481.850 295.720 1483.310 299.870 ;
        RECT 1484.150 295.720 1485.150 299.870 ;
        RECT 1485.990 295.720 1487.450 299.870 ;
        RECT 1488.290 295.720 1489.290 299.870 ;
        RECT 1490.130 295.720 1491.590 299.870 ;
        RECT 1492.430 295.720 1493.890 299.870 ;
        RECT 1494.730 295.720 1495.730 299.870 ;
        RECT 1496.570 295.720 1498.030 299.870 ;
        RECT 1498.870 295.720 1499.870 299.870 ;
        RECT 1500.710 295.720 1502.170 299.870 ;
        RECT 1503.010 295.720 1504.470 299.870 ;
        RECT 1505.310 295.720 1506.310 299.870 ;
        RECT 1507.150 295.720 1508.610 299.870 ;
        RECT 1509.450 295.720 1510.450 299.870 ;
        RECT 1511.290 295.720 1512.750 299.870 ;
        RECT 1513.590 295.720 1514.590 299.870 ;
        RECT 1515.430 295.720 1516.890 299.870 ;
        RECT 1517.730 295.720 1519.190 299.870 ;
        RECT 1520.030 295.720 1521.030 299.870 ;
        RECT 1521.870 295.720 1523.330 299.870 ;
        RECT 1524.170 295.720 1525.170 299.870 ;
        RECT 1526.010 295.720 1527.470 299.870 ;
        RECT 1528.310 295.720 1529.770 299.870 ;
        RECT 1530.610 295.720 1531.610 299.870 ;
        RECT 1532.450 295.720 1533.910 299.870 ;
        RECT 1534.750 295.720 1535.750 299.870 ;
        RECT 1536.590 295.720 1538.050 299.870 ;
        RECT 1538.890 295.720 1540.350 299.870 ;
        RECT 1541.190 295.720 1542.190 299.870 ;
        RECT 1543.030 295.720 1544.490 299.870 ;
        RECT 1545.330 295.720 1546.330 299.870 ;
        RECT 1547.170 295.720 1548.630 299.870 ;
        RECT 1549.470 295.720 1550.930 299.870 ;
        RECT 1551.770 295.720 1552.770 299.870 ;
        RECT 1553.610 295.720 1555.070 299.870 ;
        RECT 1555.910 295.720 1556.910 299.870 ;
        RECT 1557.750 295.720 1559.210 299.870 ;
        RECT 1560.050 295.720 1561.050 299.870 ;
        RECT 1561.890 295.720 1563.350 299.870 ;
        RECT 1564.190 295.720 1565.650 299.870 ;
        RECT 1566.490 295.720 1567.490 299.870 ;
        RECT 1568.330 295.720 1569.790 299.870 ;
        RECT 1570.630 295.720 1571.630 299.870 ;
        RECT 1572.470 295.720 1573.930 299.870 ;
        RECT 1574.770 295.720 1576.230 299.870 ;
        RECT 1577.070 295.720 1578.070 299.870 ;
        RECT 1578.910 295.720 1580.370 299.870 ;
        RECT 1581.210 295.720 1582.210 299.870 ;
        RECT 1583.050 295.720 1584.510 299.870 ;
        RECT 1585.350 295.720 1586.810 299.870 ;
        RECT 1587.650 295.720 1588.650 299.870 ;
        RECT 1589.490 295.720 1590.950 299.870 ;
        RECT 1591.790 295.720 1592.790 299.870 ;
        RECT 1593.630 295.720 1595.090 299.870 ;
        RECT 1595.930 295.720 1597.390 299.870 ;
        RECT 1598.230 295.720 1599.230 299.870 ;
        RECT 1600.070 295.720 1601.530 299.870 ;
        RECT 1602.370 295.720 1603.370 299.870 ;
        RECT 1604.210 295.720 1605.670 299.870 ;
        RECT 1606.510 295.720 1607.510 299.870 ;
        RECT 1608.350 295.720 1609.810 299.870 ;
        RECT 1610.650 295.720 1612.110 299.870 ;
        RECT 1612.950 295.720 1613.950 299.870 ;
        RECT 1614.790 295.720 1616.250 299.870 ;
        RECT 1617.090 295.720 1618.090 299.870 ;
        RECT 1618.930 295.720 1620.390 299.870 ;
        RECT 1621.230 295.720 1622.690 299.870 ;
        RECT 1623.530 295.720 1624.530 299.870 ;
        RECT 1625.370 295.720 1626.830 299.870 ;
        RECT 1627.670 295.720 1628.670 299.870 ;
        RECT 1629.510 295.720 1630.970 299.870 ;
        RECT 1631.810 295.720 1633.270 299.870 ;
        RECT 1634.110 295.720 1635.110 299.870 ;
        RECT 1635.950 295.720 1637.410 299.870 ;
        RECT 1638.250 295.720 1639.250 299.870 ;
        RECT 1640.090 295.720 1641.550 299.870 ;
        RECT 1642.390 295.720 1643.850 299.870 ;
        RECT 1644.690 295.720 1645.690 299.870 ;
        RECT 1646.530 295.720 1647.990 299.870 ;
        RECT 1648.830 295.720 1649.830 299.870 ;
        RECT 1650.670 295.720 1652.130 299.870 ;
        RECT 1652.970 295.720 1653.970 299.870 ;
        RECT 1654.810 295.720 1656.270 299.870 ;
        RECT 1657.110 295.720 1658.570 299.870 ;
        RECT 1659.410 295.720 1660.410 299.870 ;
        RECT 1661.250 295.720 1662.710 299.870 ;
        RECT 1663.550 295.720 1664.550 299.870 ;
        RECT 1665.390 295.720 1666.850 299.870 ;
        RECT 1667.690 295.720 1669.150 299.870 ;
        RECT 1669.990 295.720 1670.990 299.870 ;
        RECT 1671.830 295.720 1673.290 299.870 ;
        RECT 1674.130 295.720 1675.130 299.870 ;
        RECT 1675.970 295.720 1677.430 299.870 ;
        RECT 1678.270 295.720 1679.730 299.870 ;
        RECT 1680.570 295.720 1681.570 299.870 ;
        RECT 1682.410 295.720 1683.870 299.870 ;
        RECT 1684.710 295.720 1685.710 299.870 ;
        RECT 1686.550 295.720 1688.010 299.870 ;
        RECT 1688.850 295.720 1690.310 299.870 ;
        RECT 1691.150 295.720 1692.150 299.870 ;
        RECT 1692.990 295.720 1694.450 299.870 ;
        RECT 1695.290 295.720 1696.290 299.870 ;
        RECT 1697.130 295.720 1698.590 299.870 ;
        RECT 1.020 4.280 1699.140 295.720 ;
        RECT 1.020 2.875 4.410 4.280 ;
        RECT 5.250 2.875 14.070 4.280 ;
        RECT 14.910 2.875 24.190 4.280 ;
        RECT 25.030 2.875 33.850 4.280 ;
        RECT 34.690 2.875 43.970 4.280 ;
        RECT 44.810 2.875 54.090 4.280 ;
        RECT 54.930 2.875 63.750 4.280 ;
        RECT 64.590 2.875 73.870 4.280 ;
        RECT 74.710 2.875 83.530 4.280 ;
        RECT 84.370 2.875 93.650 4.280 ;
        RECT 94.490 2.875 103.770 4.280 ;
        RECT 104.610 2.875 113.430 4.280 ;
        RECT 114.270 2.875 123.550 4.280 ;
        RECT 124.390 2.875 133.210 4.280 ;
        RECT 134.050 2.875 143.330 4.280 ;
        RECT 144.170 2.875 153.450 4.280 ;
        RECT 154.290 2.875 163.110 4.280 ;
        RECT 163.950 2.875 173.230 4.280 ;
        RECT 174.070 2.875 183.350 4.280 ;
        RECT 184.190 2.875 193.010 4.280 ;
        RECT 193.850 2.875 203.130 4.280 ;
        RECT 203.970 2.875 212.790 4.280 ;
        RECT 213.630 2.875 222.910 4.280 ;
        RECT 223.750 2.875 233.030 4.280 ;
        RECT 233.870 2.875 242.690 4.280 ;
        RECT 243.530 2.875 252.810 4.280 ;
        RECT 253.650 2.875 262.470 4.280 ;
        RECT 263.310 2.875 272.590 4.280 ;
        RECT 273.430 2.875 282.710 4.280 ;
        RECT 283.550 2.875 292.370 4.280 ;
        RECT 293.210 2.875 302.490 4.280 ;
        RECT 303.330 2.875 312.610 4.280 ;
        RECT 313.450 2.875 322.270 4.280 ;
        RECT 323.110 2.875 332.390 4.280 ;
        RECT 333.230 2.875 342.050 4.280 ;
        RECT 342.890 2.875 352.170 4.280 ;
        RECT 353.010 2.875 362.290 4.280 ;
        RECT 363.130 2.875 371.950 4.280 ;
        RECT 372.790 2.875 382.070 4.280 ;
        RECT 382.910 2.875 391.730 4.280 ;
        RECT 392.570 2.875 401.850 4.280 ;
        RECT 402.690 2.875 411.970 4.280 ;
        RECT 412.810 2.875 421.630 4.280 ;
        RECT 422.470 2.875 431.750 4.280 ;
        RECT 432.590 2.875 441.870 4.280 ;
        RECT 442.710 2.875 451.530 4.280 ;
        RECT 452.370 2.875 461.650 4.280 ;
        RECT 462.490 2.875 471.310 4.280 ;
        RECT 472.150 2.875 481.430 4.280 ;
        RECT 482.270 2.875 491.550 4.280 ;
        RECT 492.390 2.875 501.210 4.280 ;
        RECT 502.050 2.875 511.330 4.280 ;
        RECT 512.170 2.875 520.990 4.280 ;
        RECT 521.830 2.875 531.110 4.280 ;
        RECT 531.950 2.875 541.230 4.280 ;
        RECT 542.070 2.875 550.890 4.280 ;
        RECT 551.730 2.875 561.010 4.280 ;
        RECT 561.850 2.875 571.130 4.280 ;
        RECT 571.970 2.875 580.790 4.280 ;
        RECT 581.630 2.875 590.910 4.280 ;
        RECT 591.750 2.875 600.570 4.280 ;
        RECT 601.410 2.875 610.690 4.280 ;
        RECT 611.530 2.875 620.810 4.280 ;
        RECT 621.650 2.875 630.470 4.280 ;
        RECT 631.310 2.875 640.590 4.280 ;
        RECT 641.430 2.875 650.250 4.280 ;
        RECT 651.090 2.875 660.370 4.280 ;
        RECT 661.210 2.875 670.490 4.280 ;
        RECT 671.330 2.875 680.150 4.280 ;
        RECT 680.990 2.875 690.270 4.280 ;
        RECT 691.110 2.875 699.930 4.280 ;
        RECT 700.770 2.875 710.050 4.280 ;
        RECT 710.890 2.875 720.170 4.280 ;
        RECT 721.010 2.875 729.830 4.280 ;
        RECT 730.670 2.875 739.950 4.280 ;
        RECT 740.790 2.875 750.070 4.280 ;
        RECT 750.910 2.875 759.730 4.280 ;
        RECT 760.570 2.875 769.850 4.280 ;
        RECT 770.690 2.875 779.510 4.280 ;
        RECT 780.350 2.875 789.630 4.280 ;
        RECT 790.470 2.875 799.750 4.280 ;
        RECT 800.590 2.875 809.410 4.280 ;
        RECT 810.250 2.875 819.530 4.280 ;
        RECT 820.370 2.875 829.190 4.280 ;
        RECT 830.030 2.875 839.310 4.280 ;
        RECT 840.150 2.875 849.430 4.280 ;
        RECT 850.270 2.875 859.090 4.280 ;
        RECT 859.930 2.875 869.210 4.280 ;
        RECT 870.050 2.875 879.330 4.280 ;
        RECT 880.170 2.875 888.990 4.280 ;
        RECT 889.830 2.875 899.110 4.280 ;
        RECT 899.950 2.875 908.770 4.280 ;
        RECT 909.610 2.875 918.890 4.280 ;
        RECT 919.730 2.875 929.010 4.280 ;
        RECT 929.850 2.875 938.670 4.280 ;
        RECT 939.510 2.875 948.790 4.280 ;
        RECT 949.630 2.875 958.450 4.280 ;
        RECT 959.290 2.875 968.570 4.280 ;
        RECT 969.410 2.875 978.690 4.280 ;
        RECT 979.530 2.875 988.350 4.280 ;
        RECT 989.190 2.875 998.470 4.280 ;
        RECT 999.310 2.875 1008.590 4.280 ;
        RECT 1009.430 2.875 1018.250 4.280 ;
        RECT 1019.090 2.875 1028.370 4.280 ;
        RECT 1029.210 2.875 1038.030 4.280 ;
        RECT 1038.870 2.875 1048.150 4.280 ;
        RECT 1048.990 2.875 1058.270 4.280 ;
        RECT 1059.110 2.875 1067.930 4.280 ;
        RECT 1068.770 2.875 1078.050 4.280 ;
        RECT 1078.890 2.875 1087.710 4.280 ;
        RECT 1088.550 2.875 1097.830 4.280 ;
        RECT 1098.670 2.875 1107.950 4.280 ;
        RECT 1108.790 2.875 1117.610 4.280 ;
        RECT 1118.450 2.875 1127.730 4.280 ;
        RECT 1128.570 2.875 1137.850 4.280 ;
        RECT 1138.690 2.875 1147.510 4.280 ;
        RECT 1148.350 2.875 1157.630 4.280 ;
        RECT 1158.470 2.875 1167.290 4.280 ;
        RECT 1168.130 2.875 1177.410 4.280 ;
        RECT 1178.250 2.875 1187.530 4.280 ;
        RECT 1188.370 2.875 1197.190 4.280 ;
        RECT 1198.030 2.875 1207.310 4.280 ;
        RECT 1208.150 2.875 1216.970 4.280 ;
        RECT 1217.810 2.875 1227.090 4.280 ;
        RECT 1227.930 2.875 1237.210 4.280 ;
        RECT 1238.050 2.875 1246.870 4.280 ;
        RECT 1247.710 2.875 1256.990 4.280 ;
        RECT 1257.830 2.875 1266.650 4.280 ;
        RECT 1267.490 2.875 1276.770 4.280 ;
        RECT 1277.610 2.875 1286.890 4.280 ;
        RECT 1287.730 2.875 1296.550 4.280 ;
        RECT 1297.390 2.875 1306.670 4.280 ;
        RECT 1307.510 2.875 1316.790 4.280 ;
        RECT 1317.630 2.875 1326.450 4.280 ;
        RECT 1327.290 2.875 1336.570 4.280 ;
        RECT 1337.410 2.875 1346.230 4.280 ;
        RECT 1347.070 2.875 1356.350 4.280 ;
        RECT 1357.190 2.875 1366.470 4.280 ;
        RECT 1367.310 2.875 1376.130 4.280 ;
        RECT 1376.970 2.875 1386.250 4.280 ;
        RECT 1387.090 2.875 1395.910 4.280 ;
        RECT 1396.750 2.875 1406.030 4.280 ;
        RECT 1406.870 2.875 1416.150 4.280 ;
        RECT 1416.990 2.875 1425.810 4.280 ;
        RECT 1426.650 2.875 1435.930 4.280 ;
        RECT 1436.770 2.875 1446.050 4.280 ;
        RECT 1446.890 2.875 1455.710 4.280 ;
        RECT 1456.550 2.875 1465.830 4.280 ;
        RECT 1466.670 2.875 1475.490 4.280 ;
        RECT 1476.330 2.875 1485.610 4.280 ;
        RECT 1486.450 2.875 1495.730 4.280 ;
        RECT 1496.570 2.875 1505.390 4.280 ;
        RECT 1506.230 2.875 1515.510 4.280 ;
        RECT 1516.350 2.875 1525.170 4.280 ;
        RECT 1526.010 2.875 1535.290 4.280 ;
        RECT 1536.130 2.875 1545.410 4.280 ;
        RECT 1546.250 2.875 1555.070 4.280 ;
        RECT 1555.910 2.875 1565.190 4.280 ;
        RECT 1566.030 2.875 1575.310 4.280 ;
        RECT 1576.150 2.875 1584.970 4.280 ;
        RECT 1585.810 2.875 1595.090 4.280 ;
        RECT 1595.930 2.875 1604.750 4.280 ;
        RECT 1605.590 2.875 1614.870 4.280 ;
        RECT 1615.710 2.875 1624.990 4.280 ;
        RECT 1625.830 2.875 1634.650 4.280 ;
        RECT 1635.490 2.875 1644.770 4.280 ;
        RECT 1645.610 2.875 1654.430 4.280 ;
        RECT 1655.270 2.875 1664.550 4.280 ;
        RECT 1665.390 2.875 1674.670 4.280 ;
        RECT 1675.510 2.875 1684.330 4.280 ;
        RECT 1685.170 2.875 1694.450 4.280 ;
        RECT 1695.290 2.875 1699.140 4.280 ;
      LAYER met3 ;
        RECT 4.400 296.120 1695.600 296.985 ;
        RECT 4.000 292.080 1696.000 296.120 ;
        RECT 4.400 290.680 1695.600 292.080 ;
        RECT 4.000 286.640 1696.000 290.680 ;
        RECT 4.400 285.240 1695.600 286.640 ;
        RECT 4.000 281.200 1696.000 285.240 ;
        RECT 4.400 279.800 1695.600 281.200 ;
        RECT 4.000 275.760 1696.000 279.800 ;
        RECT 4.400 274.360 1695.600 275.760 ;
        RECT 4.000 270.320 1696.000 274.360 ;
        RECT 4.400 268.920 1695.600 270.320 ;
        RECT 4.000 264.200 1696.000 268.920 ;
        RECT 4.400 262.800 1695.600 264.200 ;
        RECT 4.000 258.760 1696.000 262.800 ;
        RECT 4.400 257.360 1695.600 258.760 ;
        RECT 4.000 253.320 1696.000 257.360 ;
        RECT 4.400 251.920 1695.600 253.320 ;
        RECT 4.000 247.880 1696.000 251.920 ;
        RECT 4.400 246.480 1695.600 247.880 ;
        RECT 4.000 242.440 1696.000 246.480 ;
        RECT 4.400 241.040 1695.600 242.440 ;
        RECT 4.000 237.000 1696.000 241.040 ;
        RECT 4.400 235.600 1695.600 237.000 ;
        RECT 4.000 230.880 1696.000 235.600 ;
        RECT 4.400 229.480 1695.600 230.880 ;
        RECT 4.000 225.440 1696.000 229.480 ;
        RECT 4.400 224.040 1695.600 225.440 ;
        RECT 4.000 220.000 1696.000 224.040 ;
        RECT 4.400 218.600 1695.600 220.000 ;
        RECT 4.000 214.560 1696.000 218.600 ;
        RECT 4.400 213.160 1695.600 214.560 ;
        RECT 4.000 209.120 1696.000 213.160 ;
        RECT 4.400 207.720 1695.600 209.120 ;
        RECT 4.000 203.680 1696.000 207.720 ;
        RECT 4.400 202.280 1695.600 203.680 ;
        RECT 4.000 197.560 1696.000 202.280 ;
        RECT 4.400 196.160 1695.600 197.560 ;
        RECT 4.000 192.120 1696.000 196.160 ;
        RECT 4.400 190.720 1695.600 192.120 ;
        RECT 4.000 186.680 1696.000 190.720 ;
        RECT 4.400 185.280 1695.600 186.680 ;
        RECT 4.000 181.240 1696.000 185.280 ;
        RECT 4.400 179.840 1695.600 181.240 ;
        RECT 4.000 175.800 1696.000 179.840 ;
        RECT 4.400 174.400 1695.600 175.800 ;
        RECT 4.000 170.360 1696.000 174.400 ;
        RECT 4.400 168.960 1695.600 170.360 ;
        RECT 4.000 164.240 1696.000 168.960 ;
        RECT 4.400 162.840 1695.600 164.240 ;
        RECT 4.000 158.800 1696.000 162.840 ;
        RECT 4.400 157.400 1695.600 158.800 ;
        RECT 4.000 153.360 1696.000 157.400 ;
        RECT 4.400 151.960 1695.600 153.360 ;
        RECT 4.000 147.920 1696.000 151.960 ;
        RECT 4.400 146.520 1695.600 147.920 ;
        RECT 4.000 142.480 1696.000 146.520 ;
        RECT 4.400 141.080 1695.600 142.480 ;
        RECT 4.000 137.040 1696.000 141.080 ;
        RECT 4.400 135.640 1695.600 137.040 ;
        RECT 4.000 130.920 1696.000 135.640 ;
        RECT 4.400 129.520 1695.600 130.920 ;
        RECT 4.000 125.480 1696.000 129.520 ;
        RECT 4.400 124.080 1695.600 125.480 ;
        RECT 4.000 120.040 1696.000 124.080 ;
        RECT 4.400 118.640 1695.600 120.040 ;
        RECT 4.000 114.600 1696.000 118.640 ;
        RECT 4.400 113.200 1695.600 114.600 ;
        RECT 4.000 109.160 1696.000 113.200 ;
        RECT 4.400 107.760 1695.600 109.160 ;
        RECT 4.000 103.720 1696.000 107.760 ;
        RECT 4.400 102.320 1695.600 103.720 ;
        RECT 4.000 97.600 1696.000 102.320 ;
        RECT 4.400 96.200 1695.600 97.600 ;
        RECT 4.000 92.160 1696.000 96.200 ;
        RECT 4.400 90.760 1695.600 92.160 ;
        RECT 4.000 86.720 1696.000 90.760 ;
        RECT 4.400 85.320 1695.600 86.720 ;
        RECT 4.000 81.280 1696.000 85.320 ;
        RECT 4.400 79.880 1695.600 81.280 ;
        RECT 4.000 75.840 1696.000 79.880 ;
        RECT 4.400 74.440 1695.600 75.840 ;
        RECT 4.000 70.400 1696.000 74.440 ;
        RECT 4.400 69.000 1695.600 70.400 ;
        RECT 4.000 64.280 1696.000 69.000 ;
        RECT 4.400 62.880 1695.600 64.280 ;
        RECT 4.000 58.840 1696.000 62.880 ;
        RECT 4.400 57.440 1695.600 58.840 ;
        RECT 4.000 53.400 1696.000 57.440 ;
        RECT 4.400 52.000 1695.600 53.400 ;
        RECT 4.000 47.960 1696.000 52.000 ;
        RECT 4.400 46.560 1695.600 47.960 ;
        RECT 4.000 42.520 1696.000 46.560 ;
        RECT 4.400 41.120 1695.600 42.520 ;
        RECT 4.000 37.080 1696.000 41.120 ;
        RECT 4.400 35.680 1695.600 37.080 ;
        RECT 4.000 30.960 1696.000 35.680 ;
        RECT 4.400 29.560 1695.600 30.960 ;
        RECT 4.000 25.520 1696.000 29.560 ;
        RECT 4.400 24.120 1695.600 25.520 ;
        RECT 4.000 20.080 1696.000 24.120 ;
        RECT 4.400 18.680 1695.600 20.080 ;
        RECT 4.000 14.640 1696.000 18.680 ;
        RECT 4.400 13.240 1695.600 14.640 ;
        RECT 4.000 9.200 1696.000 13.240 ;
        RECT 4.400 7.800 1695.600 9.200 ;
        RECT 4.000 3.760 1696.000 7.800 ;
        RECT 4.400 2.895 1695.600 3.760 ;
      LAYER met4 ;
        RECT 164.975 288.960 1514.025 293.585 ;
        RECT 164.975 11.735 174.240 288.960 ;
        RECT 176.640 11.735 251.040 288.960 ;
        RECT 253.440 11.735 327.840 288.960 ;
        RECT 330.240 11.735 404.640 288.960 ;
        RECT 407.040 11.735 481.440 288.960 ;
        RECT 483.840 11.735 558.240 288.960 ;
        RECT 560.640 11.735 635.040 288.960 ;
        RECT 637.440 11.735 711.840 288.960 ;
        RECT 714.240 11.735 788.640 288.960 ;
        RECT 791.040 11.735 865.440 288.960 ;
        RECT 867.840 11.735 942.240 288.960 ;
        RECT 944.640 11.735 1019.040 288.960 ;
        RECT 1021.440 11.735 1095.840 288.960 ;
        RECT 1098.240 11.735 1172.640 288.960 ;
        RECT 1175.040 11.735 1249.440 288.960 ;
        RECT 1251.840 11.735 1326.240 288.960 ;
        RECT 1328.640 11.735 1403.040 288.960 ;
        RECT 1405.440 11.735 1479.840 288.960 ;
        RECT 1482.240 11.735 1514.025 288.960 ;
  END
END soric_soc
END LIBRARY

