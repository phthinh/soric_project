VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO uart_to_mem
  CLASS BLOCK ;
  FOREIGN uart_to_mem ;
  ORIGIN 0.000 0.000 ;
  SIZE 153.560 BY 164.280 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 3.440 153.560 4.040 ;
    END
  END clk_i
  PIN data_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 160.280 9.110 164.280 ;
    END
  END data_addr_o[0]
  PIN data_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 25.880 153.560 26.480 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 160.280 39.930 164.280 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 160.280 45.910 164.280 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 160.280 51.890 164.280 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 85.720 153.560 86.320 ;
    END
  END data_addr_o[9]
  PIN data_be_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 160.280 15.090 164.280 ;
    END
  END data_be_o[0]
  PIN data_be_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 160.280 21.530 164.280 ;
    END
  END data_be_o[1]
  PIN data_be_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 160.280 33.490 164.280 ;
    END
  END data_be_o[2]
  PIN data_be_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 40.840 153.560 41.440 ;
    END
  END data_be_o[3]
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END data_gnt_i
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END data_rdata_i[0]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 160.280 70.290 164.280 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 160.280 76.730 164.280 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 115.640 153.560 116.240 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 160.280 82.710 164.280 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 160.280 89.150 164.280 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 138.080 153.560 138.680 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 160.280 27.510 164.280 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 160.280 107.550 164.280 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 145.560 153.560 146.160 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 160.280 119.510 164.280 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 160.280 131.930 164.280 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 160.280 137.910 164.280 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 160.280 144.350 164.280 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 48.320 153.560 48.920 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 78.240 153.560 78.840 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 93.200 153.560 93.800 ;
    END
  END data_rdata_i[9]
  PIN data_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END data_req_o
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END data_rvalid_i
  PIN data_wdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 18.400 153.560 19.000 ;
    END
  END data_wdata_o[0]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 160.280 64.310 164.280 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 108.160 153.560 108.760 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 123.120 153.560 123.720 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 130.600 153.560 131.200 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 160.280 95.130 164.280 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 160.280 101.110 164.280 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 160.280 113.530 164.280 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 160.280 125.950 164.280 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 153.040 153.560 153.640 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 160.280 150.330 164.280 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 33.360 153.560 33.960 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 160.520 153.560 161.120 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 55.800 153.560 56.400 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 63.280 153.560 63.880 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 70.760 153.560 71.360 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 160.280 58.330 164.280 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 100.680 153.560 101.280 ;
    END
  END data_wdata_o[9]
  PIN data_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END data_we_o
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END rst_i
  PIN rx_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.560 10.920 153.560 11.520 ;
    END
  END rx_i
  PIN tx_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END tx_o
  PIN uart_error
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 160.280 3.130 164.280 ;
    END
  END uart_error
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.405 10.640 30.005 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.785 10.640 77.385 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.165 10.640 124.765 152.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 52.095 10.640 53.695 152.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.475 10.640 101.075 152.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 148.435 152.405 ;
      LAYER met1 ;
        RECT 2.830 6.500 150.350 153.640 ;
      LAYER met2 ;
        RECT 3.410 160.000 8.550 161.005 ;
        RECT 9.390 160.000 14.530 161.005 ;
        RECT 15.370 160.000 20.970 161.005 ;
        RECT 21.810 160.000 26.950 161.005 ;
        RECT 27.790 160.000 32.930 161.005 ;
        RECT 33.770 160.000 39.370 161.005 ;
        RECT 40.210 160.000 45.350 161.005 ;
        RECT 46.190 160.000 51.330 161.005 ;
        RECT 52.170 160.000 57.770 161.005 ;
        RECT 58.610 160.000 63.750 161.005 ;
        RECT 64.590 160.000 69.730 161.005 ;
        RECT 70.570 160.000 76.170 161.005 ;
        RECT 77.010 160.000 82.150 161.005 ;
        RECT 82.990 160.000 88.590 161.005 ;
        RECT 89.430 160.000 94.570 161.005 ;
        RECT 95.410 160.000 100.550 161.005 ;
        RECT 101.390 160.000 106.990 161.005 ;
        RECT 107.830 160.000 112.970 161.005 ;
        RECT 113.810 160.000 118.950 161.005 ;
        RECT 119.790 160.000 125.390 161.005 ;
        RECT 126.230 160.000 131.370 161.005 ;
        RECT 132.210 160.000 137.350 161.005 ;
        RECT 138.190 160.000 143.790 161.005 ;
        RECT 144.630 160.000 149.770 161.005 ;
        RECT 2.860 4.280 150.320 160.000 ;
        RECT 2.860 3.555 3.950 4.280 ;
        RECT 4.790 3.555 12.230 4.280 ;
        RECT 13.070 3.555 20.970 4.280 ;
        RECT 21.810 3.555 29.250 4.280 ;
        RECT 30.090 3.555 37.990 4.280 ;
        RECT 38.830 3.555 46.270 4.280 ;
        RECT 47.110 3.555 55.010 4.280 ;
        RECT 55.850 3.555 63.290 4.280 ;
        RECT 64.130 3.555 72.030 4.280 ;
        RECT 72.870 3.555 80.770 4.280 ;
        RECT 81.610 3.555 89.050 4.280 ;
        RECT 89.890 3.555 97.790 4.280 ;
        RECT 98.630 3.555 106.070 4.280 ;
        RECT 106.910 3.555 114.810 4.280 ;
        RECT 115.650 3.555 123.090 4.280 ;
        RECT 123.930 3.555 131.830 4.280 ;
        RECT 132.670 3.555 140.110 4.280 ;
        RECT 140.950 3.555 148.850 4.280 ;
        RECT 149.690 3.555 150.320 4.280 ;
      LAYER met3 ;
        RECT 4.400 160.120 149.160 160.985 ;
        RECT 4.000 154.720 149.560 160.120 ;
        RECT 4.400 154.040 149.560 154.720 ;
        RECT 4.400 153.320 149.160 154.040 ;
        RECT 4.000 152.640 149.160 153.320 ;
        RECT 4.000 147.920 149.560 152.640 ;
        RECT 4.400 146.560 149.560 147.920 ;
        RECT 4.400 146.520 149.160 146.560 ;
        RECT 4.000 145.160 149.160 146.520 ;
        RECT 4.000 141.120 149.560 145.160 ;
        RECT 4.400 139.720 149.560 141.120 ;
        RECT 4.000 139.080 149.560 139.720 ;
        RECT 4.000 137.680 149.160 139.080 ;
        RECT 4.000 134.320 149.560 137.680 ;
        RECT 4.400 132.920 149.560 134.320 ;
        RECT 4.000 131.600 149.560 132.920 ;
        RECT 4.000 130.200 149.160 131.600 ;
        RECT 4.000 127.520 149.560 130.200 ;
        RECT 4.400 126.120 149.560 127.520 ;
        RECT 4.000 124.120 149.560 126.120 ;
        RECT 4.000 122.720 149.160 124.120 ;
        RECT 4.000 120.720 149.560 122.720 ;
        RECT 4.400 119.320 149.560 120.720 ;
        RECT 4.000 116.640 149.560 119.320 ;
        RECT 4.000 115.240 149.160 116.640 ;
        RECT 4.000 113.920 149.560 115.240 ;
        RECT 4.400 112.520 149.560 113.920 ;
        RECT 4.000 109.160 149.560 112.520 ;
        RECT 4.000 107.760 149.160 109.160 ;
        RECT 4.000 107.120 149.560 107.760 ;
        RECT 4.400 105.720 149.560 107.120 ;
        RECT 4.000 101.680 149.560 105.720 ;
        RECT 4.000 100.320 149.160 101.680 ;
        RECT 4.400 100.280 149.160 100.320 ;
        RECT 4.400 98.920 149.560 100.280 ;
        RECT 4.000 94.200 149.560 98.920 ;
        RECT 4.000 93.520 149.160 94.200 ;
        RECT 4.400 92.800 149.160 93.520 ;
        RECT 4.400 92.120 149.560 92.800 ;
        RECT 4.000 86.720 149.560 92.120 ;
        RECT 4.400 85.320 149.160 86.720 ;
        RECT 4.000 79.240 149.560 85.320 ;
        RECT 4.400 77.840 149.160 79.240 ;
        RECT 4.000 72.440 149.560 77.840 ;
        RECT 4.400 71.760 149.560 72.440 ;
        RECT 4.400 71.040 149.160 71.760 ;
        RECT 4.000 70.360 149.160 71.040 ;
        RECT 4.000 65.640 149.560 70.360 ;
        RECT 4.400 64.280 149.560 65.640 ;
        RECT 4.400 64.240 149.160 64.280 ;
        RECT 4.000 62.880 149.160 64.240 ;
        RECT 4.000 58.840 149.560 62.880 ;
        RECT 4.400 57.440 149.560 58.840 ;
        RECT 4.000 56.800 149.560 57.440 ;
        RECT 4.000 55.400 149.160 56.800 ;
        RECT 4.000 52.040 149.560 55.400 ;
        RECT 4.400 50.640 149.560 52.040 ;
        RECT 4.000 49.320 149.560 50.640 ;
        RECT 4.000 47.920 149.160 49.320 ;
        RECT 4.000 45.240 149.560 47.920 ;
        RECT 4.400 43.840 149.560 45.240 ;
        RECT 4.000 41.840 149.560 43.840 ;
        RECT 4.000 40.440 149.160 41.840 ;
        RECT 4.000 38.440 149.560 40.440 ;
        RECT 4.400 37.040 149.560 38.440 ;
        RECT 4.000 34.360 149.560 37.040 ;
        RECT 4.000 32.960 149.160 34.360 ;
        RECT 4.000 31.640 149.560 32.960 ;
        RECT 4.400 30.240 149.560 31.640 ;
        RECT 4.000 26.880 149.560 30.240 ;
        RECT 4.000 25.480 149.160 26.880 ;
        RECT 4.000 24.840 149.560 25.480 ;
        RECT 4.400 23.440 149.560 24.840 ;
        RECT 4.000 19.400 149.560 23.440 ;
        RECT 4.000 18.040 149.160 19.400 ;
        RECT 4.400 18.000 149.160 18.040 ;
        RECT 4.400 16.640 149.560 18.000 ;
        RECT 4.000 11.920 149.560 16.640 ;
        RECT 4.000 11.240 149.160 11.920 ;
        RECT 4.400 10.520 149.160 11.240 ;
        RECT 4.400 9.840 149.560 10.520 ;
        RECT 4.000 4.440 149.560 9.840 ;
        RECT 4.400 3.575 149.160 4.440 ;
      LAYER met4 ;
        RECT 30.405 10.640 51.695 152.560 ;
        RECT 54.095 10.640 75.385 152.560 ;
        RECT 77.785 10.640 99.075 152.560 ;
        RECT 101.475 10.640 102.745 152.560 ;
  END
END uart_to_mem
END LIBRARY

