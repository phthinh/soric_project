VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO soric_soc
  CLASS BLOCK ;
  FOREIGN soric_soc ;
  ORIGIN 0.000 0.000 ;
  SIZE 1700.000 BY 300.000 ;
  PIN error_uart_to_mem
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 49.680 1700.000 50.280 ;
    END
  END error_uart_to_mem
  PIN master_data_addr_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 296.000 1.290 300.000 ;
    END
  END master_data_addr_to_inter_i[0]
  PIN master_data_addr_to_inter_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 296.000 160.450 300.000 ;
    END
  END master_data_addr_to_inter_i[10]
  PIN master_data_addr_to_inter_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 296.000 171.490 300.000 ;
    END
  END master_data_addr_to_inter_i[11]
  PIN master_data_addr_to_inter_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 296.000 182.530 300.000 ;
    END
  END master_data_addr_to_inter_i[12]
  PIN master_data_addr_to_inter_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 296.000 193.570 300.000 ;
    END
  END master_data_addr_to_inter_i[13]
  PIN master_data_addr_to_inter_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 296.000 204.610 300.000 ;
    END
  END master_data_addr_to_inter_i[14]
  PIN master_data_addr_to_inter_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 296.000 215.650 300.000 ;
    END
  END master_data_addr_to_inter_i[15]
  PIN master_data_addr_to_inter_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 296.000 226.690 300.000 ;
    END
  END master_data_addr_to_inter_i[16]
  PIN master_data_addr_to_inter_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 296.000 237.730 300.000 ;
    END
  END master_data_addr_to_inter_i[17]
  PIN master_data_addr_to_inter_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 296.000 248.770 300.000 ;
    END
  END master_data_addr_to_inter_i[18]
  PIN master_data_addr_to_inter_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 296.000 259.810 300.000 ;
    END
  END master_data_addr_to_inter_i[19]
  PIN master_data_addr_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 296.000 29.810 300.000 ;
    END
  END master_data_addr_to_inter_i[1]
  PIN master_data_addr_to_inter_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 296.000 270.850 300.000 ;
    END
  END master_data_addr_to_inter_i[20]
  PIN master_data_addr_to_inter_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 296.000 281.890 300.000 ;
    END
  END master_data_addr_to_inter_i[21]
  PIN master_data_addr_to_inter_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 296.000 292.930 300.000 ;
    END
  END master_data_addr_to_inter_i[22]
  PIN master_data_addr_to_inter_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 296.000 303.970 300.000 ;
    END
  END master_data_addr_to_inter_i[23]
  PIN master_data_addr_to_inter_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 296.000 315.010 300.000 ;
    END
  END master_data_addr_to_inter_i[24]
  PIN master_data_addr_to_inter_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 296.000 326.050 300.000 ;
    END
  END master_data_addr_to_inter_i[25]
  PIN master_data_addr_to_inter_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 296.000 337.090 300.000 ;
    END
  END master_data_addr_to_inter_i[26]
  PIN master_data_addr_to_inter_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 296.000 345.830 300.000 ;
    END
  END master_data_addr_to_inter_i[27]
  PIN master_data_addr_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 296.000 58.330 300.000 ;
    END
  END master_data_addr_to_inter_i[2]
  PIN master_data_addr_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 296.000 71.670 300.000 ;
    END
  END master_data_addr_to_inter_i[3]
  PIN master_data_addr_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 296.000 85.010 300.000 ;
    END
  END master_data_addr_to_inter_i[4]
  PIN master_data_addr_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 296.000 98.350 300.000 ;
    END
  END master_data_addr_to_inter_i[5]
  PIN master_data_addr_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 296.000 111.690 300.000 ;
    END
  END master_data_addr_to_inter_i[6]
  PIN master_data_addr_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 296.000 125.030 300.000 ;
    END
  END master_data_addr_to_inter_i[7]
  PIN master_data_addr_to_inter_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 296.000 137.910 300.000 ;
    END
  END master_data_addr_to_inter_i[8]
  PIN master_data_addr_to_inter_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 296.000 149.410 300.000 ;
    END
  END master_data_addr_to_inter_i[9]
  PIN master_data_addr_to_inter_ro[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 296.000 3.130 300.000 ;
    END
  END master_data_addr_to_inter_ro[0]
  PIN master_data_addr_to_inter_ro[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 296.000 162.290 300.000 ;
    END
  END master_data_addr_to_inter_ro[10]
  PIN master_data_addr_to_inter_ro[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 296.000 173.330 300.000 ;
    END
  END master_data_addr_to_inter_ro[11]
  PIN master_data_addr_to_inter_ro[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 296.000 184.370 300.000 ;
    END
  END master_data_addr_to_inter_ro[12]
  PIN master_data_addr_to_inter_ro[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 296.000 195.410 300.000 ;
    END
  END master_data_addr_to_inter_ro[13]
  PIN master_data_addr_to_inter_ro[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 296.000 206.450 300.000 ;
    END
  END master_data_addr_to_inter_ro[14]
  PIN master_data_addr_to_inter_ro[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 296.000 217.950 300.000 ;
    END
  END master_data_addr_to_inter_ro[15]
  PIN master_data_addr_to_inter_ro[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 296.000 228.990 300.000 ;
    END
  END master_data_addr_to_inter_ro[16]
  PIN master_data_addr_to_inter_ro[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 296.000 240.030 300.000 ;
    END
  END master_data_addr_to_inter_ro[17]
  PIN master_data_addr_to_inter_ro[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 296.000 251.070 300.000 ;
    END
  END master_data_addr_to_inter_ro[18]
  PIN master_data_addr_to_inter_ro[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 296.000 262.110 300.000 ;
    END
  END master_data_addr_to_inter_ro[19]
  PIN master_data_addr_to_inter_ro[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 296.000 32.110 300.000 ;
    END
  END master_data_addr_to_inter_ro[1]
  PIN master_data_addr_to_inter_ro[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 296.000 273.150 300.000 ;
    END
  END master_data_addr_to_inter_ro[20]
  PIN master_data_addr_to_inter_ro[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 296.000 284.190 300.000 ;
    END
  END master_data_addr_to_inter_ro[21]
  PIN master_data_addr_to_inter_ro[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 296.000 295.230 300.000 ;
    END
  END master_data_addr_to_inter_ro[22]
  PIN master_data_addr_to_inter_ro[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 296.000 306.270 300.000 ;
    END
  END master_data_addr_to_inter_ro[23]
  PIN master_data_addr_to_inter_ro[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 296.000 317.310 300.000 ;
    END
  END master_data_addr_to_inter_ro[24]
  PIN master_data_addr_to_inter_ro[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 296.000 328.350 300.000 ;
    END
  END master_data_addr_to_inter_ro[25]
  PIN master_data_addr_to_inter_ro[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 296.000 60.630 300.000 ;
    END
  END master_data_addr_to_inter_ro[2]
  PIN master_data_addr_to_inter_ro[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 296.000 73.970 300.000 ;
    END
  END master_data_addr_to_inter_ro[3]
  PIN master_data_addr_to_inter_ro[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 296.000 87.310 300.000 ;
    END
  END master_data_addr_to_inter_ro[4]
  PIN master_data_addr_to_inter_ro[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 296.000 100.650 300.000 ;
    END
  END master_data_addr_to_inter_ro[5]
  PIN master_data_addr_to_inter_ro[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 296.000 113.990 300.000 ;
    END
  END master_data_addr_to_inter_ro[6]
  PIN master_data_addr_to_inter_ro[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 296.000 126.870 300.000 ;
    END
  END master_data_addr_to_inter_ro[7]
  PIN master_data_addr_to_inter_ro[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 296.000 140.210 300.000 ;
    END
  END master_data_addr_to_inter_ro[8]
  PIN master_data_addr_to_inter_ro[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 296.000 151.250 300.000 ;
    END
  END master_data_addr_to_inter_ro[9]
  PIN master_data_be_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 296.000 5.430 300.000 ;
    END
  END master_data_be_to_inter_i[0]
  PIN master_data_be_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 296.000 34.410 300.000 ;
    END
  END master_data_be_to_inter_i[1]
  PIN master_data_be_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 296.000 62.930 300.000 ;
    END
  END master_data_be_to_inter_i[2]
  PIN master_data_be_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 296.000 76.270 300.000 ;
    END
  END master_data_be_to_inter_i[3]
  PIN master_data_be_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 296.000 89.610 300.000 ;
    END
  END master_data_be_to_inter_i[4]
  PIN master_data_be_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 296.000 102.950 300.000 ;
    END
  END master_data_be_to_inter_i[5]
  PIN master_data_be_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 296.000 115.830 300.000 ;
    END
  END master_data_be_to_inter_i[6]
  PIN master_data_be_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 296.000 129.170 300.000 ;
    END
  END master_data_be_to_inter_i[7]
  PIN master_data_gnt_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 296.000 7.730 300.000 ;
    END
  END master_data_gnt_to_inter_o[0]
  PIN master_data_gnt_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 296.000 36.250 300.000 ;
    END
  END master_data_gnt_to_inter_o[1]
  PIN master_data_gnt_to_inter_ro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 296.000 10.030 300.000 ;
    END
  END master_data_gnt_to_inter_ro[0]
  PIN master_data_gnt_to_inter_ro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 296.000 38.550 300.000 ;
    END
  END master_data_gnt_to_inter_ro[1]
  PIN master_data_rdata_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 296.000 12.330 300.000 ;
    END
  END master_data_rdata_to_inter_o[0]
  PIN master_data_rdata_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 296.000 164.590 300.000 ;
    END
  END master_data_rdata_to_inter_o[10]
  PIN master_data_rdata_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 296.000 175.630 300.000 ;
    END
  END master_data_rdata_to_inter_o[11]
  PIN master_data_rdata_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 296.000 186.670 300.000 ;
    END
  END master_data_rdata_to_inter_o[12]
  PIN master_data_rdata_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 296.000 197.710 300.000 ;
    END
  END master_data_rdata_to_inter_o[13]
  PIN master_data_rdata_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 296.000 208.750 300.000 ;
    END
  END master_data_rdata_to_inter_o[14]
  PIN master_data_rdata_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 296.000 219.790 300.000 ;
    END
  END master_data_rdata_to_inter_o[15]
  PIN master_data_rdata_to_inter_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 296.000 230.830 300.000 ;
    END
  END master_data_rdata_to_inter_o[16]
  PIN master_data_rdata_to_inter_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 296.000 241.870 300.000 ;
    END
  END master_data_rdata_to_inter_o[17]
  PIN master_data_rdata_to_inter_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 296.000 252.910 300.000 ;
    END
  END master_data_rdata_to_inter_o[18]
  PIN master_data_rdata_to_inter_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 296.000 263.950 300.000 ;
    END
  END master_data_rdata_to_inter_o[19]
  PIN master_data_rdata_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 296.000 40.850 300.000 ;
    END
  END master_data_rdata_to_inter_o[1]
  PIN master_data_rdata_to_inter_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 296.000 274.990 300.000 ;
    END
  END master_data_rdata_to_inter_o[20]
  PIN master_data_rdata_to_inter_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 296.000 286.490 300.000 ;
    END
  END master_data_rdata_to_inter_o[21]
  PIN master_data_rdata_to_inter_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 296.000 297.530 300.000 ;
    END
  END master_data_rdata_to_inter_o[22]
  PIN master_data_rdata_to_inter_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 296.000 308.570 300.000 ;
    END
  END master_data_rdata_to_inter_o[23]
  PIN master_data_rdata_to_inter_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 296.000 319.610 300.000 ;
    END
  END master_data_rdata_to_inter_o[24]
  PIN master_data_rdata_to_inter_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 296.000 330.650 300.000 ;
    END
  END master_data_rdata_to_inter_o[25]
  PIN master_data_rdata_to_inter_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 296.000 339.390 300.000 ;
    END
  END master_data_rdata_to_inter_o[26]
  PIN master_data_rdata_to_inter_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 296.000 348.130 300.000 ;
    END
  END master_data_rdata_to_inter_o[27]
  PIN master_data_rdata_to_inter_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 296.000 354.570 300.000 ;
    END
  END master_data_rdata_to_inter_o[28]
  PIN master_data_rdata_to_inter_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 296.000 361.470 300.000 ;
    END
  END master_data_rdata_to_inter_o[29]
  PIN master_data_rdata_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 296.000 65.230 300.000 ;
    END
  END master_data_rdata_to_inter_o[2]
  PIN master_data_rdata_to_inter_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 296.000 367.910 300.000 ;
    END
  END master_data_rdata_to_inter_o[30]
  PIN master_data_rdata_to_inter_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 296.000 374.810 300.000 ;
    END
  END master_data_rdata_to_inter_o[31]
  PIN master_data_rdata_to_inter_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 296.000 381.250 300.000 ;
    END
  END master_data_rdata_to_inter_o[32]
  PIN master_data_rdata_to_inter_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 296.000 388.150 300.000 ;
    END
  END master_data_rdata_to_inter_o[33]
  PIN master_data_rdata_to_inter_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 296.000 394.590 300.000 ;
    END
  END master_data_rdata_to_inter_o[34]
  PIN master_data_rdata_to_inter_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 296.000 401.030 300.000 ;
    END
  END master_data_rdata_to_inter_o[35]
  PIN master_data_rdata_to_inter_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 296.000 407.930 300.000 ;
    END
  END master_data_rdata_to_inter_o[36]
  PIN master_data_rdata_to_inter_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 296.000 414.370 300.000 ;
    END
  END master_data_rdata_to_inter_o[37]
  PIN master_data_rdata_to_inter_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 296.000 421.270 300.000 ;
    END
  END master_data_rdata_to_inter_o[38]
  PIN master_data_rdata_to_inter_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 296.000 427.710 300.000 ;
    END
  END master_data_rdata_to_inter_o[39]
  PIN master_data_rdata_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 296.000 78.570 300.000 ;
    END
  END master_data_rdata_to_inter_o[3]
  PIN master_data_rdata_to_inter_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 296.000 434.610 300.000 ;
    END
  END master_data_rdata_to_inter_o[40]
  PIN master_data_rdata_to_inter_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 296.000 441.050 300.000 ;
    END
  END master_data_rdata_to_inter_o[41]
  PIN master_data_rdata_to_inter_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 296.000 447.490 300.000 ;
    END
  END master_data_rdata_to_inter_o[42]
  PIN master_data_rdata_to_inter_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 296.000 454.390 300.000 ;
    END
  END master_data_rdata_to_inter_o[43]
  PIN master_data_rdata_to_inter_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 296.000 460.830 300.000 ;
    END
  END master_data_rdata_to_inter_o[44]
  PIN master_data_rdata_to_inter_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 296.000 467.730 300.000 ;
    END
  END master_data_rdata_to_inter_o[45]
  PIN master_data_rdata_to_inter_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 296.000 474.170 300.000 ;
    END
  END master_data_rdata_to_inter_o[46]
  PIN master_data_rdata_to_inter_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 296.000 480.610 300.000 ;
    END
  END master_data_rdata_to_inter_o[47]
  PIN master_data_rdata_to_inter_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 296.000 487.510 300.000 ;
    END
  END master_data_rdata_to_inter_o[48]
  PIN master_data_rdata_to_inter_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 296.000 493.950 300.000 ;
    END
  END master_data_rdata_to_inter_o[49]
  PIN master_data_rdata_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 296.000 91.910 300.000 ;
    END
  END master_data_rdata_to_inter_o[4]
  PIN master_data_rdata_to_inter_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 296.000 500.850 300.000 ;
    END
  END master_data_rdata_to_inter_o[50]
  PIN master_data_rdata_to_inter_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 296.000 507.290 300.000 ;
    END
  END master_data_rdata_to_inter_o[51]
  PIN master_data_rdata_to_inter_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 296.000 514.190 300.000 ;
    END
  END master_data_rdata_to_inter_o[52]
  PIN master_data_rdata_to_inter_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 296.000 520.630 300.000 ;
    END
  END master_data_rdata_to_inter_o[53]
  PIN master_data_rdata_to_inter_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 296.000 527.070 300.000 ;
    END
  END master_data_rdata_to_inter_o[54]
  PIN master_data_rdata_to_inter_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 296.000 533.970 300.000 ;
    END
  END master_data_rdata_to_inter_o[55]
  PIN master_data_rdata_to_inter_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 296.000 540.410 300.000 ;
    END
  END master_data_rdata_to_inter_o[56]
  PIN master_data_rdata_to_inter_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 296.000 547.310 300.000 ;
    END
  END master_data_rdata_to_inter_o[57]
  PIN master_data_rdata_to_inter_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 296.000 553.750 300.000 ;
    END
  END master_data_rdata_to_inter_o[58]
  PIN master_data_rdata_to_inter_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 296.000 560.190 300.000 ;
    END
  END master_data_rdata_to_inter_o[59]
  PIN master_data_rdata_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 296.000 104.790 300.000 ;
    END
  END master_data_rdata_to_inter_o[5]
  PIN master_data_rdata_to_inter_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 296.000 567.090 300.000 ;
    END
  END master_data_rdata_to_inter_o[60]
  PIN master_data_rdata_to_inter_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 296.000 573.530 300.000 ;
    END
  END master_data_rdata_to_inter_o[61]
  PIN master_data_rdata_to_inter_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 296.000 580.430 300.000 ;
    END
  END master_data_rdata_to_inter_o[62]
  PIN master_data_rdata_to_inter_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 296.000 586.870 300.000 ;
    END
  END master_data_rdata_to_inter_o[63]
  PIN master_data_rdata_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 296.000 118.130 300.000 ;
    END
  END master_data_rdata_to_inter_o[6]
  PIN master_data_rdata_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 296.000 131.470 300.000 ;
    END
  END master_data_rdata_to_inter_o[7]
  PIN master_data_rdata_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 296.000 142.510 300.000 ;
    END
  END master_data_rdata_to_inter_o[8]
  PIN master_data_rdata_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 296.000 153.550 300.000 ;
    END
  END master_data_rdata_to_inter_o[9]
  PIN master_data_rdata_to_inter_ro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 296.000 14.170 300.000 ;
    END
  END master_data_rdata_to_inter_ro[0]
  PIN master_data_rdata_to_inter_ro[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 296.000 166.890 300.000 ;
    END
  END master_data_rdata_to_inter_ro[10]
  PIN master_data_rdata_to_inter_ro[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 296.000 177.930 300.000 ;
    END
  END master_data_rdata_to_inter_ro[11]
  PIN master_data_rdata_to_inter_ro[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 296.000 188.970 300.000 ;
    END
  END master_data_rdata_to_inter_ro[12]
  PIN master_data_rdata_to_inter_ro[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 296.000 200.010 300.000 ;
    END
  END master_data_rdata_to_inter_ro[13]
  PIN master_data_rdata_to_inter_ro[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 296.000 211.050 300.000 ;
    END
  END master_data_rdata_to_inter_ro[14]
  PIN master_data_rdata_to_inter_ro[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 296.000 222.090 300.000 ;
    END
  END master_data_rdata_to_inter_ro[15]
  PIN master_data_rdata_to_inter_ro[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 296.000 233.130 300.000 ;
    END
  END master_data_rdata_to_inter_ro[16]
  PIN master_data_rdata_to_inter_ro[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 296.000 244.170 300.000 ;
    END
  END master_data_rdata_to_inter_ro[17]
  PIN master_data_rdata_to_inter_ro[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 296.000 255.210 300.000 ;
    END
  END master_data_rdata_to_inter_ro[18]
  PIN master_data_rdata_to_inter_ro[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 296.000 266.250 300.000 ;
    END
  END master_data_rdata_to_inter_ro[19]
  PIN master_data_rdata_to_inter_ro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 296.000 43.150 300.000 ;
    END
  END master_data_rdata_to_inter_ro[1]
  PIN master_data_rdata_to_inter_ro[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 296.000 277.290 300.000 ;
    END
  END master_data_rdata_to_inter_ro[20]
  PIN master_data_rdata_to_inter_ro[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 296.000 288.330 300.000 ;
    END
  END master_data_rdata_to_inter_ro[21]
  PIN master_data_rdata_to_inter_ro[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 296.000 299.370 300.000 ;
    END
  END master_data_rdata_to_inter_ro[22]
  PIN master_data_rdata_to_inter_ro[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 296.000 310.410 300.000 ;
    END
  END master_data_rdata_to_inter_ro[23]
  PIN master_data_rdata_to_inter_ro[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 296.000 321.450 300.000 ;
    END
  END master_data_rdata_to_inter_ro[24]
  PIN master_data_rdata_to_inter_ro[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 296.000 332.490 300.000 ;
    END
  END master_data_rdata_to_inter_ro[25]
  PIN master_data_rdata_to_inter_ro[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 296.000 341.690 300.000 ;
    END
  END master_data_rdata_to_inter_ro[26]
  PIN master_data_rdata_to_inter_ro[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 296.000 350.430 300.000 ;
    END
  END master_data_rdata_to_inter_ro[27]
  PIN master_data_rdata_to_inter_ro[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 296.000 356.870 300.000 ;
    END
  END master_data_rdata_to_inter_ro[28]
  PIN master_data_rdata_to_inter_ro[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 296.000 363.770 300.000 ;
    END
  END master_data_rdata_to_inter_ro[29]
  PIN master_data_rdata_to_inter_ro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 296.000 67.530 300.000 ;
    END
  END master_data_rdata_to_inter_ro[2]
  PIN master_data_rdata_to_inter_ro[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 296.000 370.210 300.000 ;
    END
  END master_data_rdata_to_inter_ro[30]
  PIN master_data_rdata_to_inter_ro[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 296.000 377.110 300.000 ;
    END
  END master_data_rdata_to_inter_ro[31]
  PIN master_data_rdata_to_inter_ro[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 296.000 383.550 300.000 ;
    END
  END master_data_rdata_to_inter_ro[32]
  PIN master_data_rdata_to_inter_ro[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 296.000 389.990 300.000 ;
    END
  END master_data_rdata_to_inter_ro[33]
  PIN master_data_rdata_to_inter_ro[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 296.000 396.890 300.000 ;
    END
  END master_data_rdata_to_inter_ro[34]
  PIN master_data_rdata_to_inter_ro[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 296.000 403.330 300.000 ;
    END
  END master_data_rdata_to_inter_ro[35]
  PIN master_data_rdata_to_inter_ro[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 296.000 410.230 300.000 ;
    END
  END master_data_rdata_to_inter_ro[36]
  PIN master_data_rdata_to_inter_ro[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 296.000 416.670 300.000 ;
    END
  END master_data_rdata_to_inter_ro[37]
  PIN master_data_rdata_to_inter_ro[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 296.000 423.110 300.000 ;
    END
  END master_data_rdata_to_inter_ro[38]
  PIN master_data_rdata_to_inter_ro[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 296.000 430.010 300.000 ;
    END
  END master_data_rdata_to_inter_ro[39]
  PIN master_data_rdata_to_inter_ro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 296.000 80.870 300.000 ;
    END
  END master_data_rdata_to_inter_ro[3]
  PIN master_data_rdata_to_inter_ro[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 296.000 436.450 300.000 ;
    END
  END master_data_rdata_to_inter_ro[40]
  PIN master_data_rdata_to_inter_ro[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 296.000 443.350 300.000 ;
    END
  END master_data_rdata_to_inter_ro[41]
  PIN master_data_rdata_to_inter_ro[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 296.000 449.790 300.000 ;
    END
  END master_data_rdata_to_inter_ro[42]
  PIN master_data_rdata_to_inter_ro[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 296.000 456.690 300.000 ;
    END
  END master_data_rdata_to_inter_ro[43]
  PIN master_data_rdata_to_inter_ro[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 296.000 463.130 300.000 ;
    END
  END master_data_rdata_to_inter_ro[44]
  PIN master_data_rdata_to_inter_ro[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 296.000 469.570 300.000 ;
    END
  END master_data_rdata_to_inter_ro[45]
  PIN master_data_rdata_to_inter_ro[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 296.000 476.470 300.000 ;
    END
  END master_data_rdata_to_inter_ro[46]
  PIN master_data_rdata_to_inter_ro[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 296.000 482.910 300.000 ;
    END
  END master_data_rdata_to_inter_ro[47]
  PIN master_data_rdata_to_inter_ro[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 296.000 489.810 300.000 ;
    END
  END master_data_rdata_to_inter_ro[48]
  PIN master_data_rdata_to_inter_ro[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 296.000 496.250 300.000 ;
    END
  END master_data_rdata_to_inter_ro[49]
  PIN master_data_rdata_to_inter_ro[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 296.000 93.750 300.000 ;
    END
  END master_data_rdata_to_inter_ro[4]
  PIN master_data_rdata_to_inter_ro[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 296.000 503.150 300.000 ;
    END
  END master_data_rdata_to_inter_ro[50]
  PIN master_data_rdata_to_inter_ro[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 296.000 509.590 300.000 ;
    END
  END master_data_rdata_to_inter_ro[51]
  PIN master_data_rdata_to_inter_ro[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 296.000 516.030 300.000 ;
    END
  END master_data_rdata_to_inter_ro[52]
  PIN master_data_rdata_to_inter_ro[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 296.000 522.930 300.000 ;
    END
  END master_data_rdata_to_inter_ro[53]
  PIN master_data_rdata_to_inter_ro[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 296.000 529.370 300.000 ;
    END
  END master_data_rdata_to_inter_ro[54]
  PIN master_data_rdata_to_inter_ro[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 296.000 536.270 300.000 ;
    END
  END master_data_rdata_to_inter_ro[55]
  PIN master_data_rdata_to_inter_ro[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 296.000 542.710 300.000 ;
    END
  END master_data_rdata_to_inter_ro[56]
  PIN master_data_rdata_to_inter_ro[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 296.000 549.150 300.000 ;
    END
  END master_data_rdata_to_inter_ro[57]
  PIN master_data_rdata_to_inter_ro[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 296.000 556.050 300.000 ;
    END
  END master_data_rdata_to_inter_ro[58]
  PIN master_data_rdata_to_inter_ro[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 296.000 562.490 300.000 ;
    END
  END master_data_rdata_to_inter_ro[59]
  PIN master_data_rdata_to_inter_ro[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 296.000 107.090 300.000 ;
    END
  END master_data_rdata_to_inter_ro[5]
  PIN master_data_rdata_to_inter_ro[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 296.000 569.390 300.000 ;
    END
  END master_data_rdata_to_inter_ro[60]
  PIN master_data_rdata_to_inter_ro[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 296.000 575.830 300.000 ;
    END
  END master_data_rdata_to_inter_ro[61]
  PIN master_data_rdata_to_inter_ro[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 296.000 582.730 300.000 ;
    END
  END master_data_rdata_to_inter_ro[62]
  PIN master_data_rdata_to_inter_ro[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 296.000 589.170 300.000 ;
    END
  END master_data_rdata_to_inter_ro[63]
  PIN master_data_rdata_to_inter_ro[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 296.000 120.430 300.000 ;
    END
  END master_data_rdata_to_inter_ro[6]
  PIN master_data_rdata_to_inter_ro[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 296.000 133.770 300.000 ;
    END
  END master_data_rdata_to_inter_ro[7]
  PIN master_data_rdata_to_inter_ro[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 296.000 144.810 300.000 ;
    END
  END master_data_rdata_to_inter_ro[8]
  PIN master_data_rdata_to_inter_ro[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 296.000 155.850 300.000 ;
    END
  END master_data_rdata_to_inter_ro[9]
  PIN master_data_req_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 296.000 16.470 300.000 ;
    END
  END master_data_req_to_inter_i[0]
  PIN master_data_req_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 296.000 45.450 300.000 ;
    END
  END master_data_req_to_inter_i[1]
  PIN master_data_req_to_inter_ro[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 296.000 18.770 300.000 ;
    END
  END master_data_req_to_inter_ro[0]
  PIN master_data_req_to_inter_ro[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 296.000 47.290 300.000 ;
    END
  END master_data_req_to_inter_ro[1]
  PIN master_data_rvalid_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 296.000 21.070 300.000 ;
    END
  END master_data_rvalid_to_inter_o[0]
  PIN master_data_rvalid_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 296.000 49.590 300.000 ;
    END
  END master_data_rvalid_to_inter_o[1]
  PIN master_data_rvalid_to_inter_ro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 296.000 23.370 300.000 ;
    END
  END master_data_rvalid_to_inter_ro[0]
  PIN master_data_rvalid_to_inter_ro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 296.000 51.890 300.000 ;
    END
  END master_data_rvalid_to_inter_ro[1]
  PIN master_data_wdata_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 296.000 25.210 300.000 ;
    END
  END master_data_wdata_to_inter_i[0]
  PIN master_data_wdata_to_inter_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 296.000 169.190 300.000 ;
    END
  END master_data_wdata_to_inter_i[10]
  PIN master_data_wdata_to_inter_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 296.000 180.230 300.000 ;
    END
  END master_data_wdata_to_inter_i[11]
  PIN master_data_wdata_to_inter_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 296.000 191.270 300.000 ;
    END
  END master_data_wdata_to_inter_i[12]
  PIN master_data_wdata_to_inter_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 296.000 202.310 300.000 ;
    END
  END master_data_wdata_to_inter_i[13]
  PIN master_data_wdata_to_inter_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 296.000 213.350 300.000 ;
    END
  END master_data_wdata_to_inter_i[14]
  PIN master_data_wdata_to_inter_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 296.000 224.390 300.000 ;
    END
  END master_data_wdata_to_inter_i[15]
  PIN master_data_wdata_to_inter_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 296.000 235.430 300.000 ;
    END
  END master_data_wdata_to_inter_i[16]
  PIN master_data_wdata_to_inter_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 296.000 246.470 300.000 ;
    END
  END master_data_wdata_to_inter_i[17]
  PIN master_data_wdata_to_inter_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 296.000 257.510 300.000 ;
    END
  END master_data_wdata_to_inter_i[18]
  PIN master_data_wdata_to_inter_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 296.000 268.550 300.000 ;
    END
  END master_data_wdata_to_inter_i[19]
  PIN master_data_wdata_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 296.000 54.190 300.000 ;
    END
  END master_data_wdata_to_inter_i[1]
  PIN master_data_wdata_to_inter_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 296.000 279.590 300.000 ;
    END
  END master_data_wdata_to_inter_i[20]
  PIN master_data_wdata_to_inter_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 296.000 290.630 300.000 ;
    END
  END master_data_wdata_to_inter_i[21]
  PIN master_data_wdata_to_inter_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 296.000 301.670 300.000 ;
    END
  END master_data_wdata_to_inter_i[22]
  PIN master_data_wdata_to_inter_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 296.000 312.710 300.000 ;
    END
  END master_data_wdata_to_inter_i[23]
  PIN master_data_wdata_to_inter_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 296.000 323.750 300.000 ;
    END
  END master_data_wdata_to_inter_i[24]
  PIN master_data_wdata_to_inter_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 296.000 334.790 300.000 ;
    END
  END master_data_wdata_to_inter_i[25]
  PIN master_data_wdata_to_inter_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 296.000 343.530 300.000 ;
    END
  END master_data_wdata_to_inter_i[26]
  PIN master_data_wdata_to_inter_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 296.000 352.730 300.000 ;
    END
  END master_data_wdata_to_inter_i[27]
  PIN master_data_wdata_to_inter_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 296.000 359.170 300.000 ;
    END
  END master_data_wdata_to_inter_i[28]
  PIN master_data_wdata_to_inter_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 296.000 366.070 300.000 ;
    END
  END master_data_wdata_to_inter_i[29]
  PIN master_data_wdata_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 296.000 69.370 300.000 ;
    END
  END master_data_wdata_to_inter_i[2]
  PIN master_data_wdata_to_inter_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 296.000 372.510 300.000 ;
    END
  END master_data_wdata_to_inter_i[30]
  PIN master_data_wdata_to_inter_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 296.000 378.950 300.000 ;
    END
  END master_data_wdata_to_inter_i[31]
  PIN master_data_wdata_to_inter_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 296.000 385.850 300.000 ;
    END
  END master_data_wdata_to_inter_i[32]
  PIN master_data_wdata_to_inter_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 296.000 392.290 300.000 ;
    END
  END master_data_wdata_to_inter_i[33]
  PIN master_data_wdata_to_inter_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 296.000 399.190 300.000 ;
    END
  END master_data_wdata_to_inter_i[34]
  PIN master_data_wdata_to_inter_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 296.000 405.630 300.000 ;
    END
  END master_data_wdata_to_inter_i[35]
  PIN master_data_wdata_to_inter_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 296.000 412.070 300.000 ;
    END
  END master_data_wdata_to_inter_i[36]
  PIN master_data_wdata_to_inter_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 296.000 418.970 300.000 ;
    END
  END master_data_wdata_to_inter_i[37]
  PIN master_data_wdata_to_inter_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 296.000 425.410 300.000 ;
    END
  END master_data_wdata_to_inter_i[38]
  PIN master_data_wdata_to_inter_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 296.000 432.310 300.000 ;
    END
  END master_data_wdata_to_inter_i[39]
  PIN master_data_wdata_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 296.000 82.710 300.000 ;
    END
  END master_data_wdata_to_inter_i[3]
  PIN master_data_wdata_to_inter_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 296.000 438.750 300.000 ;
    END
  END master_data_wdata_to_inter_i[40]
  PIN master_data_wdata_to_inter_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 296.000 445.650 300.000 ;
    END
  END master_data_wdata_to_inter_i[41]
  PIN master_data_wdata_to_inter_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 296.000 452.090 300.000 ;
    END
  END master_data_wdata_to_inter_i[42]
  PIN master_data_wdata_to_inter_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 296.000 458.530 300.000 ;
    END
  END master_data_wdata_to_inter_i[43]
  PIN master_data_wdata_to_inter_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 296.000 465.430 300.000 ;
    END
  END master_data_wdata_to_inter_i[44]
  PIN master_data_wdata_to_inter_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 296.000 471.870 300.000 ;
    END
  END master_data_wdata_to_inter_i[45]
  PIN master_data_wdata_to_inter_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 296.000 478.770 300.000 ;
    END
  END master_data_wdata_to_inter_i[46]
  PIN master_data_wdata_to_inter_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 296.000 485.210 300.000 ;
    END
  END master_data_wdata_to_inter_i[47]
  PIN master_data_wdata_to_inter_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 296.000 491.650 300.000 ;
    END
  END master_data_wdata_to_inter_i[48]
  PIN master_data_wdata_to_inter_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 296.000 498.550 300.000 ;
    END
  END master_data_wdata_to_inter_i[49]
  PIN master_data_wdata_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 296.000 96.050 300.000 ;
    END
  END master_data_wdata_to_inter_i[4]
  PIN master_data_wdata_to_inter_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 296.000 504.990 300.000 ;
    END
  END master_data_wdata_to_inter_i[50]
  PIN master_data_wdata_to_inter_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 296.000 511.890 300.000 ;
    END
  END master_data_wdata_to_inter_i[51]
  PIN master_data_wdata_to_inter_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 296.000 518.330 300.000 ;
    END
  END master_data_wdata_to_inter_i[52]
  PIN master_data_wdata_to_inter_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 296.000 525.230 300.000 ;
    END
  END master_data_wdata_to_inter_i[53]
  PIN master_data_wdata_to_inter_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 296.000 531.670 300.000 ;
    END
  END master_data_wdata_to_inter_i[54]
  PIN master_data_wdata_to_inter_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 296.000 538.110 300.000 ;
    END
  END master_data_wdata_to_inter_i[55]
  PIN master_data_wdata_to_inter_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 296.000 545.010 300.000 ;
    END
  END master_data_wdata_to_inter_i[56]
  PIN master_data_wdata_to_inter_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 296.000 551.450 300.000 ;
    END
  END master_data_wdata_to_inter_i[57]
  PIN master_data_wdata_to_inter_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 296.000 558.350 300.000 ;
    END
  END master_data_wdata_to_inter_i[58]
  PIN master_data_wdata_to_inter_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 296.000 564.790 300.000 ;
    END
  END master_data_wdata_to_inter_i[59]
  PIN master_data_wdata_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 296.000 109.390 300.000 ;
    END
  END master_data_wdata_to_inter_i[5]
  PIN master_data_wdata_to_inter_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 296.000 571.690 300.000 ;
    END
  END master_data_wdata_to_inter_i[60]
  PIN master_data_wdata_to_inter_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 296.000 578.130 300.000 ;
    END
  END master_data_wdata_to_inter_i[61]
  PIN master_data_wdata_to_inter_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 296.000 584.570 300.000 ;
    END
  END master_data_wdata_to_inter_i[62]
  PIN master_data_wdata_to_inter_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 296.000 591.470 300.000 ;
    END
  END master_data_wdata_to_inter_i[63]
  PIN master_data_wdata_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 296.000 122.730 300.000 ;
    END
  END master_data_wdata_to_inter_i[6]
  PIN master_data_wdata_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 296.000 136.070 300.000 ;
    END
  END master_data_wdata_to_inter_i[7]
  PIN master_data_wdata_to_inter_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 296.000 147.110 300.000 ;
    END
  END master_data_wdata_to_inter_i[8]
  PIN master_data_wdata_to_inter_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 296.000 158.150 300.000 ;
    END
  END master_data_wdata_to_inter_i[9]
  PIN master_data_we_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 296.000 27.510 300.000 ;
    END
  END master_data_we_to_inter_i[0]
  PIN master_data_we_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 296.000 56.490 300.000 ;
    END
  END master_data_we_to_inter_i[1]
  PIN rxd_uart
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 0.000 1692.250 4.000 ;
    END
  END rxd_uart
  PIN rxd_uart_to_mem
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.870 296.000 1699.150 300.000 ;
    END
  END rxd_uart_to_mem
  PIN slave_data_addr_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 296.000 593.770 300.000 ;
    END
  END slave_data_addr_to_inter_o[0]
  PIN slave_data_addr_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 296.000 752.930 300.000 ;
    END
  END slave_data_addr_to_inter_o[10]
  PIN slave_data_addr_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 296.000 765.810 300.000 ;
    END
  END slave_data_addr_to_inter_o[11]
  PIN slave_data_addr_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 296.000 779.150 300.000 ;
    END
  END slave_data_addr_to_inter_o[12]
  PIN slave_data_addr_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 296.000 792.490 300.000 ;
    END
  END slave_data_addr_to_inter_o[13]
  PIN slave_data_addr_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 296.000 805.830 300.000 ;
    END
  END slave_data_addr_to_inter_o[14]
  PIN slave_data_addr_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 296.000 819.170 300.000 ;
    END
  END slave_data_addr_to_inter_o[15]
  PIN slave_data_addr_to_inter_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.230 296.000 832.510 300.000 ;
    END
  END slave_data_addr_to_inter_o[16]
  PIN slave_data_addr_to_inter_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 296.000 843.550 300.000 ;
    END
  END slave_data_addr_to_inter_o[17]
  PIN slave_data_addr_to_inter_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 296.000 854.590 300.000 ;
    END
  END slave_data_addr_to_inter_o[18]
  PIN slave_data_addr_to_inter_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 296.000 865.630 300.000 ;
    END
  END slave_data_addr_to_inter_o[19]
  PIN slave_data_addr_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 296.000 613.550 300.000 ;
    END
  END slave_data_addr_to_inter_o[1]
  PIN slave_data_addr_to_inter_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 296.000 876.670 300.000 ;
    END
  END slave_data_addr_to_inter_o[20]
  PIN slave_data_addr_to_inter_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 296.000 887.710 300.000 ;
    END
  END slave_data_addr_to_inter_o[21]
  PIN slave_data_addr_to_inter_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 296.000 898.750 300.000 ;
    END
  END slave_data_addr_to_inter_o[22]
  PIN slave_data_addr_to_inter_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 296.000 909.790 300.000 ;
    END
  END slave_data_addr_to_inter_o[23]
  PIN slave_data_addr_to_inter_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 296.000 920.830 300.000 ;
    END
  END slave_data_addr_to_inter_o[24]
  PIN slave_data_addr_to_inter_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 296.000 931.870 300.000 ;
    END
  END slave_data_addr_to_inter_o[25]
  PIN slave_data_addr_to_inter_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 296.000 942.910 300.000 ;
    END
  END slave_data_addr_to_inter_o[26]
  PIN slave_data_addr_to_inter_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 296.000 953.950 300.000 ;
    END
  END slave_data_addr_to_inter_o[27]
  PIN slave_data_addr_to_inter_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 296.000 964.990 300.000 ;
    END
  END slave_data_addr_to_inter_o[28]
  PIN slave_data_addr_to_inter_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 296.000 976.030 300.000 ;
    END
  END slave_data_addr_to_inter_o[29]
  PIN slave_data_addr_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 296.000 633.330 300.000 ;
    END
  END slave_data_addr_to_inter_o[2]
  PIN slave_data_addr_to_inter_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 296.000 987.070 300.000 ;
    END
  END slave_data_addr_to_inter_o[30]
  PIN slave_data_addr_to_inter_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.830 296.000 998.110 300.000 ;
    END
  END slave_data_addr_to_inter_o[31]
  PIN slave_data_addr_to_inter_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.870 296.000 1009.150 300.000 ;
    END
  END slave_data_addr_to_inter_o[32]
  PIN slave_data_addr_to_inter_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.910 296.000 1020.190 300.000 ;
    END
  END slave_data_addr_to_inter_o[33]
  PIN slave_data_addr_to_inter_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 296.000 1031.230 300.000 ;
    END
  END slave_data_addr_to_inter_o[34]
  PIN slave_data_addr_to_inter_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.990 296.000 1042.270 300.000 ;
    END
  END slave_data_addr_to_inter_o[35]
  PIN slave_data_addr_to_inter_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 296.000 1053.310 300.000 ;
    END
  END slave_data_addr_to_inter_o[36]
  PIN slave_data_addr_to_inter_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.070 296.000 1064.350 300.000 ;
    END
  END slave_data_addr_to_inter_o[37]
  PIN slave_data_addr_to_inter_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.110 296.000 1075.390 300.000 ;
    END
  END slave_data_addr_to_inter_o[38]
  PIN slave_data_addr_to_inter_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 296.000 1086.430 300.000 ;
    END
  END slave_data_addr_to_inter_o[39]
  PIN slave_data_addr_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 296.000 653.110 300.000 ;
    END
  END slave_data_addr_to_inter_o[3]
  PIN slave_data_addr_to_inter_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.190 296.000 1097.470 300.000 ;
    END
  END slave_data_addr_to_inter_o[40]
  PIN slave_data_addr_to_inter_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.230 296.000 1108.510 300.000 ;
    END
  END slave_data_addr_to_inter_o[41]
  PIN slave_data_addr_to_inter_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.270 296.000 1119.550 300.000 ;
    END
  END slave_data_addr_to_inter_o[42]
  PIN slave_data_addr_to_inter_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 296.000 1130.590 300.000 ;
    END
  END slave_data_addr_to_inter_o[43]
  PIN slave_data_addr_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 296.000 673.350 300.000 ;
    END
  END slave_data_addr_to_inter_o[4]
  PIN slave_data_addr_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 296.000 686.230 300.000 ;
    END
  END slave_data_addr_to_inter_o[5]
  PIN slave_data_addr_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 296.000 699.570 300.000 ;
    END
  END slave_data_addr_to_inter_o[6]
  PIN slave_data_addr_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 296.000 712.910 300.000 ;
    END
  END slave_data_addr_to_inter_o[7]
  PIN slave_data_addr_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 296.000 726.250 300.000 ;
    END
  END slave_data_addr_to_inter_o[8]
  PIN slave_data_addr_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 296.000 739.590 300.000 ;
    END
  END slave_data_addr_to_inter_o[9]
  PIN slave_data_addr_to_inter_ro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 296.000 595.610 300.000 ;
    END
  END slave_data_addr_to_inter_ro[0]
  PIN slave_data_addr_to_inter_ro[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 296.000 754.770 300.000 ;
    END
  END slave_data_addr_to_inter_ro[10]
  PIN slave_data_addr_to_inter_ro[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 296.000 768.110 300.000 ;
    END
  END slave_data_addr_to_inter_ro[11]
  PIN slave_data_addr_to_inter_ro[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 296.000 781.450 300.000 ;
    END
  END slave_data_addr_to_inter_ro[12]
  PIN slave_data_addr_to_inter_ro[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 296.000 794.790 300.000 ;
    END
  END slave_data_addr_to_inter_ro[13]
  PIN slave_data_addr_to_inter_ro[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 296.000 808.130 300.000 ;
    END
  END slave_data_addr_to_inter_ro[14]
  PIN slave_data_addr_to_inter_ro[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 296.000 821.470 300.000 ;
    END
  END slave_data_addr_to_inter_ro[15]
  PIN slave_data_addr_to_inter_ro[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 296.000 834.350 300.000 ;
    END
  END slave_data_addr_to_inter_ro[16]
  PIN slave_data_addr_to_inter_ro[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 296.000 845.390 300.000 ;
    END
  END slave_data_addr_to_inter_ro[17]
  PIN slave_data_addr_to_inter_ro[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 296.000 856.890 300.000 ;
    END
  END slave_data_addr_to_inter_ro[18]
  PIN slave_data_addr_to_inter_ro[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.650 296.000 867.930 300.000 ;
    END
  END slave_data_addr_to_inter_ro[19]
  PIN slave_data_addr_to_inter_ro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 296.000 615.850 300.000 ;
    END
  END slave_data_addr_to_inter_ro[1]
  PIN slave_data_addr_to_inter_ro[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 296.000 878.970 300.000 ;
    END
  END slave_data_addr_to_inter_ro[20]
  PIN slave_data_addr_to_inter_ro[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 296.000 890.010 300.000 ;
    END
  END slave_data_addr_to_inter_ro[21]
  PIN slave_data_addr_to_inter_ro[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 296.000 901.050 300.000 ;
    END
  END slave_data_addr_to_inter_ro[22]
  PIN slave_data_addr_to_inter_ro[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 296.000 912.090 300.000 ;
    END
  END slave_data_addr_to_inter_ro[23]
  PIN slave_data_addr_to_inter_ro[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.850 296.000 923.130 300.000 ;
    END
  END slave_data_addr_to_inter_ro[24]
  PIN slave_data_addr_to_inter_ro[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 296.000 934.170 300.000 ;
    END
  END slave_data_addr_to_inter_ro[25]
  PIN slave_data_addr_to_inter_ro[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 296.000 945.210 300.000 ;
    END
  END slave_data_addr_to_inter_ro[26]
  PIN slave_data_addr_to_inter_ro[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 296.000 956.250 300.000 ;
    END
  END slave_data_addr_to_inter_ro[27]
  PIN slave_data_addr_to_inter_ro[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.010 296.000 967.290 300.000 ;
    END
  END slave_data_addr_to_inter_ro[28]
  PIN slave_data_addr_to_inter_ro[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.050 296.000 978.330 300.000 ;
    END
  END slave_data_addr_to_inter_ro[29]
  PIN slave_data_addr_to_inter_ro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 296.000 635.630 300.000 ;
    END
  END slave_data_addr_to_inter_ro[2]
  PIN slave_data_addr_to_inter_ro[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.090 296.000 989.370 300.000 ;
    END
  END slave_data_addr_to_inter_ro[30]
  PIN slave_data_addr_to_inter_ro[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.130 296.000 1000.410 300.000 ;
    END
  END slave_data_addr_to_inter_ro[31]
  PIN slave_data_addr_to_inter_ro[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 296.000 1011.450 300.000 ;
    END
  END slave_data_addr_to_inter_ro[32]
  PIN slave_data_addr_to_inter_ro[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 296.000 1022.490 300.000 ;
    END
  END slave_data_addr_to_inter_ro[33]
  PIN slave_data_addr_to_inter_ro[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 296.000 1033.530 300.000 ;
    END
  END slave_data_addr_to_inter_ro[34]
  PIN slave_data_addr_to_inter_ro[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 296.000 1044.570 300.000 ;
    END
  END slave_data_addr_to_inter_ro[35]
  PIN slave_data_addr_to_inter_ro[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.330 296.000 1055.610 300.000 ;
    END
  END slave_data_addr_to_inter_ro[36]
  PIN slave_data_addr_to_inter_ro[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.370 296.000 1066.650 300.000 ;
    END
  END slave_data_addr_to_inter_ro[37]
  PIN slave_data_addr_to_inter_ro[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.410 296.000 1077.690 300.000 ;
    END
  END slave_data_addr_to_inter_ro[38]
  PIN slave_data_addr_to_inter_ro[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 296.000 1088.730 300.000 ;
    END
  END slave_data_addr_to_inter_ro[39]
  PIN slave_data_addr_to_inter_ro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 296.000 655.410 300.000 ;
    END
  END slave_data_addr_to_inter_ro[3]
  PIN slave_data_addr_to_inter_ro[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.490 296.000 1099.770 300.000 ;
    END
  END slave_data_addr_to_inter_ro[40]
  PIN slave_data_addr_to_inter_ro[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.530 296.000 1110.810 300.000 ;
    END
  END slave_data_addr_to_inter_ro[41]
  PIN slave_data_addr_to_inter_ro[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.570 296.000 1121.850 300.000 ;
    END
  END slave_data_addr_to_inter_ro[42]
  PIN slave_data_addr_to_inter_ro[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.610 296.000 1132.890 300.000 ;
    END
  END slave_data_addr_to_inter_ro[43]
  PIN slave_data_addr_to_inter_ro[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 296.000 675.190 300.000 ;
    END
  END slave_data_addr_to_inter_ro[4]
  PIN slave_data_addr_to_inter_ro[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 296.000 688.530 300.000 ;
    END
  END slave_data_addr_to_inter_ro[5]
  PIN slave_data_addr_to_inter_ro[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 296.000 701.870 300.000 ;
    END
  END slave_data_addr_to_inter_ro[6]
  PIN slave_data_addr_to_inter_ro[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 296.000 715.210 300.000 ;
    END
  END slave_data_addr_to_inter_ro[7]
  PIN slave_data_addr_to_inter_ro[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 296.000 728.550 300.000 ;
    END
  END slave_data_addr_to_inter_ro[8]
  PIN slave_data_addr_to_inter_ro[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 296.000 741.890 300.000 ;
    END
  END slave_data_addr_to_inter_ro[9]
  PIN slave_data_be_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 296.000 597.910 300.000 ;
    END
  END slave_data_be_to_inter_o[0]
  PIN slave_data_be_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 296.000 757.070 300.000 ;
    END
  END slave_data_be_to_inter_o[10]
  PIN slave_data_be_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 296.000 770.410 300.000 ;
    END
  END slave_data_be_to_inter_o[11]
  PIN slave_data_be_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 296.000 783.750 300.000 ;
    END
  END slave_data_be_to_inter_o[12]
  PIN slave_data_be_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 296.000 797.090 300.000 ;
    END
  END slave_data_be_to_inter_o[13]
  PIN slave_data_be_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 296.000 810.430 300.000 ;
    END
  END slave_data_be_to_inter_o[14]
  PIN slave_data_be_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.030 296.000 823.310 300.000 ;
    END
  END slave_data_be_to_inter_o[15]
  PIN slave_data_be_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 296.000 617.690 300.000 ;
    END
  END slave_data_be_to_inter_o[1]
  PIN slave_data_be_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 296.000 637.930 300.000 ;
    END
  END slave_data_be_to_inter_o[2]
  PIN slave_data_be_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 296.000 657.710 300.000 ;
    END
  END slave_data_be_to_inter_o[3]
  PIN slave_data_be_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 296.000 677.490 300.000 ;
    END
  END slave_data_be_to_inter_o[4]
  PIN slave_data_be_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 296.000 690.830 300.000 ;
    END
  END slave_data_be_to_inter_o[5]
  PIN slave_data_be_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 296.000 704.170 300.000 ;
    END
  END slave_data_be_to_inter_o[6]
  PIN slave_data_be_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 296.000 717.510 300.000 ;
    END
  END slave_data_be_to_inter_o[7]
  PIN slave_data_be_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 296.000 730.850 300.000 ;
    END
  END slave_data_be_to_inter_o[8]
  PIN slave_data_be_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 296.000 743.730 300.000 ;
    END
  END slave_data_be_to_inter_o[9]
  PIN slave_data_rdata_to_inter_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 296.000 600.210 300.000 ;
    END
  END slave_data_rdata_to_inter_i[0]
  PIN slave_data_rdata_to_inter_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.030 296.000 1513.310 300.000 ;
    END
  END slave_data_rdata_to_inter_i[100]
  PIN slave_data_rdata_to_inter_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.470 296.000 1519.750 300.000 ;
    END
  END slave_data_rdata_to_inter_i[101]
  PIN slave_data_rdata_to_inter_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 296.000 1526.650 300.000 ;
    END
  END slave_data_rdata_to_inter_i[102]
  PIN slave_data_rdata_to_inter_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 296.000 1533.090 300.000 ;
    END
  END slave_data_rdata_to_inter_i[103]
  PIN slave_data_rdata_to_inter_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.710 296.000 1539.990 300.000 ;
    END
  END slave_data_rdata_to_inter_i[104]
  PIN slave_data_rdata_to_inter_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.150 296.000 1546.430 300.000 ;
    END
  END slave_data_rdata_to_inter_i[105]
  PIN slave_data_rdata_to_inter_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.590 296.000 1552.870 300.000 ;
    END
  END slave_data_rdata_to_inter_i[106]
  PIN slave_data_rdata_to_inter_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.490 296.000 1559.770 300.000 ;
    END
  END slave_data_rdata_to_inter_i[107]
  PIN slave_data_rdata_to_inter_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.930 296.000 1566.210 300.000 ;
    END
  END slave_data_rdata_to_inter_i[108]
  PIN slave_data_rdata_to_inter_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.830 296.000 1573.110 300.000 ;
    END
  END slave_data_rdata_to_inter_i[109]
  PIN slave_data_rdata_to_inter_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 296.000 759.370 300.000 ;
    END
  END slave_data_rdata_to_inter_i[10]
  PIN slave_data_rdata_to_inter_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.270 296.000 1579.550 300.000 ;
    END
  END slave_data_rdata_to_inter_i[110]
  PIN slave_data_rdata_to_inter_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.170 296.000 1586.450 300.000 ;
    END
  END slave_data_rdata_to_inter_i[111]
  PIN slave_data_rdata_to_inter_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.610 296.000 1592.890 300.000 ;
    END
  END slave_data_rdata_to_inter_i[112]
  PIN slave_data_rdata_to_inter_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.050 296.000 1599.330 300.000 ;
    END
  END slave_data_rdata_to_inter_i[113]
  PIN slave_data_rdata_to_inter_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.950 296.000 1606.230 300.000 ;
    END
  END slave_data_rdata_to_inter_i[114]
  PIN slave_data_rdata_to_inter_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.390 296.000 1612.670 300.000 ;
    END
  END slave_data_rdata_to_inter_i[115]
  PIN slave_data_rdata_to_inter_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.290 296.000 1619.570 300.000 ;
    END
  END slave_data_rdata_to_inter_i[116]
  PIN slave_data_rdata_to_inter_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 296.000 1626.010 300.000 ;
    END
  END slave_data_rdata_to_inter_i[117]
  PIN slave_data_rdata_to_inter_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 296.000 1632.910 300.000 ;
    END
  END slave_data_rdata_to_inter_i[118]
  PIN slave_data_rdata_to_inter_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 296.000 1639.350 300.000 ;
    END
  END slave_data_rdata_to_inter_i[119]
  PIN slave_data_rdata_to_inter_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.430 296.000 772.710 300.000 ;
    END
  END slave_data_rdata_to_inter_i[11]
  PIN slave_data_rdata_to_inter_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 296.000 1645.790 300.000 ;
    END
  END slave_data_rdata_to_inter_i[120]
  PIN slave_data_rdata_to_inter_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.410 296.000 1652.690 300.000 ;
    END
  END slave_data_rdata_to_inter_i[121]
  PIN slave_data_rdata_to_inter_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 296.000 1659.130 300.000 ;
    END
  END slave_data_rdata_to_inter_i[122]
  PIN slave_data_rdata_to_inter_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.750 296.000 1666.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[123]
  PIN slave_data_rdata_to_inter_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 296.000 1672.470 300.000 ;
    END
  END slave_data_rdata_to_inter_i[124]
  PIN slave_data_rdata_to_inter_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.630 296.000 1678.910 300.000 ;
    END
  END slave_data_rdata_to_inter_i[125]
  PIN slave_data_rdata_to_inter_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.530 296.000 1685.810 300.000 ;
    END
  END slave_data_rdata_to_inter_i[126]
  PIN slave_data_rdata_to_inter_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 296.000 1692.250 300.000 ;
    END
  END slave_data_rdata_to_inter_i[127]
  PIN slave_data_rdata_to_inter_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 296.000 786.050 300.000 ;
    END
  END slave_data_rdata_to_inter_i[12]
  PIN slave_data_rdata_to_inter_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 296.000 799.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[13]
  PIN slave_data_rdata_to_inter_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 296.000 812.270 300.000 ;
    END
  END slave_data_rdata_to_inter_i[14]
  PIN slave_data_rdata_to_inter_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 296.000 825.610 300.000 ;
    END
  END slave_data_rdata_to_inter_i[15]
  PIN slave_data_rdata_to_inter_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 296.000 836.650 300.000 ;
    END
  END slave_data_rdata_to_inter_i[16]
  PIN slave_data_rdata_to_inter_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 296.000 847.690 300.000 ;
    END
  END slave_data_rdata_to_inter_i[17]
  PIN slave_data_rdata_to_inter_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 296.000 858.730 300.000 ;
    END
  END slave_data_rdata_to_inter_i[18]
  PIN slave_data_rdata_to_inter_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 296.000 869.770 300.000 ;
    END
  END slave_data_rdata_to_inter_i[19]
  PIN slave_data_rdata_to_inter_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 296.000 619.990 300.000 ;
    END
  END slave_data_rdata_to_inter_i[1]
  PIN slave_data_rdata_to_inter_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.530 296.000 880.810 300.000 ;
    END
  END slave_data_rdata_to_inter_i[20]
  PIN slave_data_rdata_to_inter_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 296.000 891.850 300.000 ;
    END
  END slave_data_rdata_to_inter_i[21]
  PIN slave_data_rdata_to_inter_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 296.000 902.890 300.000 ;
    END
  END slave_data_rdata_to_inter_i[22]
  PIN slave_data_rdata_to_inter_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 296.000 913.930 300.000 ;
    END
  END slave_data_rdata_to_inter_i[23]
  PIN slave_data_rdata_to_inter_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.150 296.000 925.430 300.000 ;
    END
  END slave_data_rdata_to_inter_i[24]
  PIN slave_data_rdata_to_inter_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.190 296.000 936.470 300.000 ;
    END
  END slave_data_rdata_to_inter_i[25]
  PIN slave_data_rdata_to_inter_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 296.000 947.510 300.000 ;
    END
  END slave_data_rdata_to_inter_i[26]
  PIN slave_data_rdata_to_inter_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.270 296.000 958.550 300.000 ;
    END
  END slave_data_rdata_to_inter_i[27]
  PIN slave_data_rdata_to_inter_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 296.000 969.590 300.000 ;
    END
  END slave_data_rdata_to_inter_i[28]
  PIN slave_data_rdata_to_inter_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 296.000 980.630 300.000 ;
    END
  END slave_data_rdata_to_inter_i[29]
  PIN slave_data_rdata_to_inter_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 296.000 640.230 300.000 ;
    END
  END slave_data_rdata_to_inter_i[2]
  PIN slave_data_rdata_to_inter_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 296.000 991.670 300.000 ;
    END
  END slave_data_rdata_to_inter_i[30]
  PIN slave_data_rdata_to_inter_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 296.000 1002.710 300.000 ;
    END
  END slave_data_rdata_to_inter_i[31]
  PIN slave_data_rdata_to_inter_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.470 296.000 1013.750 300.000 ;
    END
  END slave_data_rdata_to_inter_i[32]
  PIN slave_data_rdata_to_inter_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.510 296.000 1024.790 300.000 ;
    END
  END slave_data_rdata_to_inter_i[33]
  PIN slave_data_rdata_to_inter_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.550 296.000 1035.830 300.000 ;
    END
  END slave_data_rdata_to_inter_i[34]
  PIN slave_data_rdata_to_inter_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 296.000 1046.870 300.000 ;
    END
  END slave_data_rdata_to_inter_i[35]
  PIN slave_data_rdata_to_inter_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.630 296.000 1057.910 300.000 ;
    END
  END slave_data_rdata_to_inter_i[36]
  PIN slave_data_rdata_to_inter_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.670 296.000 1068.950 300.000 ;
    END
  END slave_data_rdata_to_inter_i[37]
  PIN slave_data_rdata_to_inter_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 296.000 1079.990 300.000 ;
    END
  END slave_data_rdata_to_inter_i[38]
  PIN slave_data_rdata_to_inter_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.750 296.000 1091.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[39]
  PIN slave_data_rdata_to_inter_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 296.000 660.010 300.000 ;
    END
  END slave_data_rdata_to_inter_i[3]
  PIN slave_data_rdata_to_inter_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 296.000 1102.070 300.000 ;
    END
  END slave_data_rdata_to_inter_i[40]
  PIN slave_data_rdata_to_inter_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.830 296.000 1113.110 300.000 ;
    END
  END slave_data_rdata_to_inter_i[41]
  PIN slave_data_rdata_to_inter_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 296.000 1124.150 300.000 ;
    END
  END slave_data_rdata_to_inter_i[42]
  PIN slave_data_rdata_to_inter_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 296.000 1135.190 300.000 ;
    END
  END slave_data_rdata_to_inter_i[43]
  PIN slave_data_rdata_to_inter_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.810 296.000 1142.090 300.000 ;
    END
  END slave_data_rdata_to_inter_i[44]
  PIN slave_data_rdata_to_inter_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.250 296.000 1148.530 300.000 ;
    END
  END slave_data_rdata_to_inter_i[45]
  PIN slave_data_rdata_to_inter_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 296.000 1154.970 300.000 ;
    END
  END slave_data_rdata_to_inter_i[46]
  PIN slave_data_rdata_to_inter_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.590 296.000 1161.870 300.000 ;
    END
  END slave_data_rdata_to_inter_i[47]
  PIN slave_data_rdata_to_inter_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.030 296.000 1168.310 300.000 ;
    END
  END slave_data_rdata_to_inter_i[48]
  PIN slave_data_rdata_to_inter_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.930 296.000 1175.210 300.000 ;
    END
  END slave_data_rdata_to_inter_i[49]
  PIN slave_data_rdata_to_inter_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 296.000 679.790 300.000 ;
    END
  END slave_data_rdata_to_inter_i[4]
  PIN slave_data_rdata_to_inter_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.370 296.000 1181.650 300.000 ;
    END
  END slave_data_rdata_to_inter_i[50]
  PIN slave_data_rdata_to_inter_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 296.000 1188.090 300.000 ;
    END
  END slave_data_rdata_to_inter_i[51]
  PIN slave_data_rdata_to_inter_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 296.000 1194.990 300.000 ;
    END
  END slave_data_rdata_to_inter_i[52]
  PIN slave_data_rdata_to_inter_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 296.000 1201.430 300.000 ;
    END
  END slave_data_rdata_to_inter_i[53]
  PIN slave_data_rdata_to_inter_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.050 296.000 1208.330 300.000 ;
    END
  END slave_data_rdata_to_inter_i[54]
  PIN slave_data_rdata_to_inter_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.490 296.000 1214.770 300.000 ;
    END
  END slave_data_rdata_to_inter_i[55]
  PIN slave_data_rdata_to_inter_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.390 296.000 1221.670 300.000 ;
    END
  END slave_data_rdata_to_inter_i[56]
  PIN slave_data_rdata_to_inter_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.830 296.000 1228.110 300.000 ;
    END
  END slave_data_rdata_to_inter_i[57]
  PIN slave_data_rdata_to_inter_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.270 296.000 1234.550 300.000 ;
    END
  END slave_data_rdata_to_inter_i[58]
  PIN slave_data_rdata_to_inter_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.170 296.000 1241.450 300.000 ;
    END
  END slave_data_rdata_to_inter_i[59]
  PIN slave_data_rdata_to_inter_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 296.000 693.130 300.000 ;
    END
  END slave_data_rdata_to_inter_i[5]
  PIN slave_data_rdata_to_inter_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.610 296.000 1247.890 300.000 ;
    END
  END slave_data_rdata_to_inter_i[60]
  PIN slave_data_rdata_to_inter_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.510 296.000 1254.790 300.000 ;
    END
  END slave_data_rdata_to_inter_i[61]
  PIN slave_data_rdata_to_inter_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.950 296.000 1261.230 300.000 ;
    END
  END slave_data_rdata_to_inter_i[62]
  PIN slave_data_rdata_to_inter_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.390 296.000 1267.670 300.000 ;
    END
  END slave_data_rdata_to_inter_i[63]
  PIN slave_data_rdata_to_inter_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.290 296.000 1274.570 300.000 ;
    END
  END slave_data_rdata_to_inter_i[64]
  PIN slave_data_rdata_to_inter_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.730 296.000 1281.010 300.000 ;
    END
  END slave_data_rdata_to_inter_i[65]
  PIN slave_data_rdata_to_inter_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.630 296.000 1287.910 300.000 ;
    END
  END slave_data_rdata_to_inter_i[66]
  PIN slave_data_rdata_to_inter_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.070 296.000 1294.350 300.000 ;
    END
  END slave_data_rdata_to_inter_i[67]
  PIN slave_data_rdata_to_inter_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.970 296.000 1301.250 300.000 ;
    END
  END slave_data_rdata_to_inter_i[68]
  PIN slave_data_rdata_to_inter_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 296.000 1307.690 300.000 ;
    END
  END slave_data_rdata_to_inter_i[69]
  PIN slave_data_rdata_to_inter_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 296.000 706.470 300.000 ;
    END
  END slave_data_rdata_to_inter_i[6]
  PIN slave_data_rdata_to_inter_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 296.000 1314.130 300.000 ;
    END
  END slave_data_rdata_to_inter_i[70]
  PIN slave_data_rdata_to_inter_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.750 296.000 1321.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[71]
  PIN slave_data_rdata_to_inter_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.190 296.000 1327.470 300.000 ;
    END
  END slave_data_rdata_to_inter_i[72]
  PIN slave_data_rdata_to_inter_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.090 296.000 1334.370 300.000 ;
    END
  END slave_data_rdata_to_inter_i[73]
  PIN slave_data_rdata_to_inter_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.530 296.000 1340.810 300.000 ;
    END
  END slave_data_rdata_to_inter_i[74]
  PIN slave_data_rdata_to_inter_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.430 296.000 1347.710 300.000 ;
    END
  END slave_data_rdata_to_inter_i[75]
  PIN slave_data_rdata_to_inter_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.870 296.000 1354.150 300.000 ;
    END
  END slave_data_rdata_to_inter_i[76]
  PIN slave_data_rdata_to_inter_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.310 296.000 1360.590 300.000 ;
    END
  END slave_data_rdata_to_inter_i[77]
  PIN slave_data_rdata_to_inter_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.210 296.000 1367.490 300.000 ;
    END
  END slave_data_rdata_to_inter_i[78]
  PIN slave_data_rdata_to_inter_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.650 296.000 1373.930 300.000 ;
    END
  END slave_data_rdata_to_inter_i[79]
  PIN slave_data_rdata_to_inter_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 296.000 719.810 300.000 ;
    END
  END slave_data_rdata_to_inter_i[7]
  PIN slave_data_rdata_to_inter_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.550 296.000 1380.830 300.000 ;
    END
  END slave_data_rdata_to_inter_i[80]
  PIN slave_data_rdata_to_inter_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.990 296.000 1387.270 300.000 ;
    END
  END slave_data_rdata_to_inter_i[81]
  PIN slave_data_rdata_to_inter_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.430 296.000 1393.710 300.000 ;
    END
  END slave_data_rdata_to_inter_i[82]
  PIN slave_data_rdata_to_inter_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.330 296.000 1400.610 300.000 ;
    END
  END slave_data_rdata_to_inter_i[83]
  PIN slave_data_rdata_to_inter_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.770 296.000 1407.050 300.000 ;
    END
  END slave_data_rdata_to_inter_i[84]
  PIN slave_data_rdata_to_inter_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 296.000 1413.950 300.000 ;
    END
  END slave_data_rdata_to_inter_i[85]
  PIN slave_data_rdata_to_inter_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 296.000 1420.390 300.000 ;
    END
  END slave_data_rdata_to_inter_i[86]
  PIN slave_data_rdata_to_inter_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 296.000 1427.290 300.000 ;
    END
  END slave_data_rdata_to_inter_i[87]
  PIN slave_data_rdata_to_inter_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.450 296.000 1433.730 300.000 ;
    END
  END slave_data_rdata_to_inter_i[88]
  PIN slave_data_rdata_to_inter_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 296.000 1440.170 300.000 ;
    END
  END slave_data_rdata_to_inter_i[89]
  PIN slave_data_rdata_to_inter_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 296.000 732.690 300.000 ;
    END
  END slave_data_rdata_to_inter_i[8]
  PIN slave_data_rdata_to_inter_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.790 296.000 1447.070 300.000 ;
    END
  END slave_data_rdata_to_inter_i[90]
  PIN slave_data_rdata_to_inter_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.230 296.000 1453.510 300.000 ;
    END
  END slave_data_rdata_to_inter_i[91]
  PIN slave_data_rdata_to_inter_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.130 296.000 1460.410 300.000 ;
    END
  END slave_data_rdata_to_inter_i[92]
  PIN slave_data_rdata_to_inter_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.570 296.000 1466.850 300.000 ;
    END
  END slave_data_rdata_to_inter_i[93]
  PIN slave_data_rdata_to_inter_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.010 296.000 1473.290 300.000 ;
    END
  END slave_data_rdata_to_inter_i[94]
  PIN slave_data_rdata_to_inter_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.910 296.000 1480.190 300.000 ;
    END
  END slave_data_rdata_to_inter_i[95]
  PIN slave_data_rdata_to_inter_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.350 296.000 1486.630 300.000 ;
    END
  END slave_data_rdata_to_inter_i[96]
  PIN slave_data_rdata_to_inter_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.250 296.000 1493.530 300.000 ;
    END
  END slave_data_rdata_to_inter_i[97]
  PIN slave_data_rdata_to_inter_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 296.000 1499.970 300.000 ;
    END
  END slave_data_rdata_to_inter_i[98]
  PIN slave_data_rdata_to_inter_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.590 296.000 1506.870 300.000 ;
    END
  END slave_data_rdata_to_inter_i[99]
  PIN slave_data_rdata_to_inter_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 296.000 746.030 300.000 ;
    END
  END slave_data_rdata_to_inter_i[9]
  PIN slave_data_rdata_to_inter_ro[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 296.000 602.510 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[0]
  PIN slave_data_rdata_to_inter_ro[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.330 296.000 1515.610 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[100]
  PIN slave_data_rdata_to_inter_ro[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.770 296.000 1522.050 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[101]
  PIN slave_data_rdata_to_inter_ro[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.670 296.000 1528.950 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[102]
  PIN slave_data_rdata_to_inter_ro[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.110 296.000 1535.390 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[103]
  PIN slave_data_rdata_to_inter_ro[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.550 296.000 1541.830 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[104]
  PIN slave_data_rdata_to_inter_ro[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.450 296.000 1548.730 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[105]
  PIN slave_data_rdata_to_inter_ro[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.890 296.000 1555.170 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[106]
  PIN slave_data_rdata_to_inter_ro[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 296.000 1562.070 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[107]
  PIN slave_data_rdata_to_inter_ro[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 296.000 1568.510 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[108]
  PIN slave_data_rdata_to_inter_ro[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.130 296.000 1575.410 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[109]
  PIN slave_data_rdata_to_inter_ro[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 296.000 761.670 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[10]
  PIN slave_data_rdata_to_inter_ro[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.570 296.000 1581.850 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[110]
  PIN slave_data_rdata_to_inter_ro[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.010 296.000 1588.290 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[111]
  PIN slave_data_rdata_to_inter_ro[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.910 296.000 1595.190 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[112]
  PIN slave_data_rdata_to_inter_ro[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1601.350 296.000 1601.630 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[113]
  PIN slave_data_rdata_to_inter_ro[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1608.250 296.000 1608.530 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[114]
  PIN slave_data_rdata_to_inter_ro[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.690 296.000 1614.970 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[115]
  PIN slave_data_rdata_to_inter_ro[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.130 296.000 1621.410 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[116]
  PIN slave_data_rdata_to_inter_ro[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.030 296.000 1628.310 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[117]
  PIN slave_data_rdata_to_inter_ro[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.470 296.000 1634.750 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[118]
  PIN slave_data_rdata_to_inter_ro[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.370 296.000 1641.650 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[119]
  PIN slave_data_rdata_to_inter_ro[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 296.000 775.010 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[11]
  PIN slave_data_rdata_to_inter_ro[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.810 296.000 1648.090 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[120]
  PIN slave_data_rdata_to_inter_ro[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.710 296.000 1654.990 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[121]
  PIN slave_data_rdata_to_inter_ro[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.150 296.000 1661.430 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[122]
  PIN slave_data_rdata_to_inter_ro[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.590 296.000 1667.870 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[123]
  PIN slave_data_rdata_to_inter_ro[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 296.000 1674.770 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[124]
  PIN slave_data_rdata_to_inter_ro[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.930 296.000 1681.210 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[125]
  PIN slave_data_rdata_to_inter_ro[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.830 296.000 1688.110 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[126]
  PIN slave_data_rdata_to_inter_ro[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.270 296.000 1694.550 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[127]
  PIN slave_data_rdata_to_inter_ro[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 296.000 788.350 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[12]
  PIN slave_data_rdata_to_inter_ro[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 296.000 801.230 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[13]
  PIN slave_data_rdata_to_inter_ro[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 296.000 814.570 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[14]
  PIN slave_data_rdata_to_inter_ro[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 296.000 827.910 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[15]
  PIN slave_data_rdata_to_inter_ro[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 296.000 838.950 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[16]
  PIN slave_data_rdata_to_inter_ro[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 296.000 849.990 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[17]
  PIN slave_data_rdata_to_inter_ro[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 296.000 861.030 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[18]
  PIN slave_data_rdata_to_inter_ro[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 296.000 872.070 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[19]
  PIN slave_data_rdata_to_inter_ro[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 296.000 622.290 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[1]
  PIN slave_data_rdata_to_inter_ro[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 296.000 883.110 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[20]
  PIN slave_data_rdata_to_inter_ro[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 296.000 894.150 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[21]
  PIN slave_data_rdata_to_inter_ro[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 296.000 905.190 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[22]
  PIN slave_data_rdata_to_inter_ro[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 296.000 916.230 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[23]
  PIN slave_data_rdata_to_inter_ro[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 296.000 927.270 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[24]
  PIN slave_data_rdata_to_inter_ro[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 296.000 938.310 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[25]
  PIN slave_data_rdata_to_inter_ro[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 296.000 949.350 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[26]
  PIN slave_data_rdata_to_inter_ro[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 296.000 960.390 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[27]
  PIN slave_data_rdata_to_inter_ro[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.150 296.000 971.430 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[28]
  PIN slave_data_rdata_to_inter_ro[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 296.000 982.470 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[29]
  PIN slave_data_rdata_to_inter_ro[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 296.000 642.070 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[2]
  PIN slave_data_rdata_to_inter_ro[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 296.000 993.970 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[30]
  PIN slave_data_rdata_to_inter_ro[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 296.000 1005.010 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[31]
  PIN slave_data_rdata_to_inter_ro[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 296.000 1016.050 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[32]
  PIN slave_data_rdata_to_inter_ro[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.810 296.000 1027.090 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[33]
  PIN slave_data_rdata_to_inter_ro[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 296.000 1038.130 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[34]
  PIN slave_data_rdata_to_inter_ro[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.890 296.000 1049.170 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[35]
  PIN slave_data_rdata_to_inter_ro[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930 296.000 1060.210 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[36]
  PIN slave_data_rdata_to_inter_ro[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.970 296.000 1071.250 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[37]
  PIN slave_data_rdata_to_inter_ro[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 296.000 1082.290 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[38]
  PIN slave_data_rdata_to_inter_ro[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 296.000 1093.330 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[39]
  PIN slave_data_rdata_to_inter_ro[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 296.000 662.310 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[3]
  PIN slave_data_rdata_to_inter_ro[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 296.000 1104.370 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[40]
  PIN slave_data_rdata_to_inter_ro[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 296.000 1115.410 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[41]
  PIN slave_data_rdata_to_inter_ro[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.170 296.000 1126.450 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[42]
  PIN slave_data_rdata_to_inter_ro[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 296.000 1137.490 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[43]
  PIN slave_data_rdata_to_inter_ro[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.650 296.000 1143.930 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[44]
  PIN slave_data_rdata_to_inter_ro[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.550 296.000 1150.830 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[45]
  PIN slave_data_rdata_to_inter_ro[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.990 296.000 1157.270 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[46]
  PIN slave_data_rdata_to_inter_ro[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 296.000 1164.170 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[47]
  PIN slave_data_rdata_to_inter_ro[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.330 296.000 1170.610 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[48]
  PIN slave_data_rdata_to_inter_ro[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 296.000 1177.050 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[49]
  PIN slave_data_rdata_to_inter_ro[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 296.000 682.090 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[4]
  PIN slave_data_rdata_to_inter_ro[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 296.000 1183.950 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[50]
  PIN slave_data_rdata_to_inter_ro[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.110 296.000 1190.390 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[51]
  PIN slave_data_rdata_to_inter_ro[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.010 296.000 1197.290 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[52]
  PIN slave_data_rdata_to_inter_ro[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.450 296.000 1203.730 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[53]
  PIN slave_data_rdata_to_inter_ro[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.350 296.000 1210.630 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[54]
  PIN slave_data_rdata_to_inter_ro[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.790 296.000 1217.070 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[55]
  PIN slave_data_rdata_to_inter_ro[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.230 296.000 1223.510 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[56]
  PIN slave_data_rdata_to_inter_ro[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 296.000 1230.410 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[57]
  PIN slave_data_rdata_to_inter_ro[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 296.000 1236.850 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[58]
  PIN slave_data_rdata_to_inter_ro[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.470 296.000 1243.750 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[59]
  PIN slave_data_rdata_to_inter_ro[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 296.000 695.430 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[5]
  PIN slave_data_rdata_to_inter_ro[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 296.000 1250.190 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[60]
  PIN slave_data_rdata_to_inter_ro[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.350 296.000 1256.630 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[61]
  PIN slave_data_rdata_to_inter_ro[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.250 296.000 1263.530 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[62]
  PIN slave_data_rdata_to_inter_ro[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 296.000 1269.970 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[63]
  PIN slave_data_rdata_to_inter_ro[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.590 296.000 1276.870 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[64]
  PIN slave_data_rdata_to_inter_ro[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.030 296.000 1283.310 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[65]
  PIN slave_data_rdata_to_inter_ro[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.930 296.000 1290.210 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[66]
  PIN slave_data_rdata_to_inter_ro[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.370 296.000 1296.650 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[67]
  PIN slave_data_rdata_to_inter_ro[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.810 296.000 1303.090 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[68]
  PIN slave_data_rdata_to_inter_ro[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 296.000 1309.990 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[69]
  PIN slave_data_rdata_to_inter_ro[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 296.000 708.310 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[6]
  PIN slave_data_rdata_to_inter_ro[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 296.000 1316.430 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[70]
  PIN slave_data_rdata_to_inter_ro[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 296.000 1323.330 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[71]
  PIN slave_data_rdata_to_inter_ro[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.490 296.000 1329.770 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[72]
  PIN slave_data_rdata_to_inter_ro[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.930 296.000 1336.210 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[73]
  PIN slave_data_rdata_to_inter_ro[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 296.000 1343.110 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[74]
  PIN slave_data_rdata_to_inter_ro[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 296.000 1349.550 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[75]
  PIN slave_data_rdata_to_inter_ro[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.170 296.000 1356.450 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[76]
  PIN slave_data_rdata_to_inter_ro[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.610 296.000 1362.890 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[77]
  PIN slave_data_rdata_to_inter_ro[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.510 296.000 1369.790 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[78]
  PIN slave_data_rdata_to_inter_ro[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.950 296.000 1376.230 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[79]
  PIN slave_data_rdata_to_inter_ro[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 296.000 721.650 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[7]
  PIN slave_data_rdata_to_inter_ro[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.390 296.000 1382.670 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[80]
  PIN slave_data_rdata_to_inter_ro[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.290 296.000 1389.570 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[81]
  PIN slave_data_rdata_to_inter_ro[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.730 296.000 1396.010 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[82]
  PIN slave_data_rdata_to_inter_ro[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.630 296.000 1402.910 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[83]
  PIN slave_data_rdata_to_inter_ro[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.070 296.000 1409.350 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[84]
  PIN slave_data_rdata_to_inter_ro[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.510 296.000 1415.790 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[85]
  PIN slave_data_rdata_to_inter_ro[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.410 296.000 1422.690 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[86]
  PIN slave_data_rdata_to_inter_ro[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.850 296.000 1429.130 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[87]
  PIN slave_data_rdata_to_inter_ro[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.750 296.000 1436.030 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[88]
  PIN slave_data_rdata_to_inter_ro[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.190 296.000 1442.470 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[89]
  PIN slave_data_rdata_to_inter_ro[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 296.000 734.990 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[8]
  PIN slave_data_rdata_to_inter_ro[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 296.000 1449.370 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[90]
  PIN slave_data_rdata_to_inter_ro[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 296.000 1455.810 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[91]
  PIN slave_data_rdata_to_inter_ro[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 296.000 1462.250 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[92]
  PIN slave_data_rdata_to_inter_ro[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.870 296.000 1469.150 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[93]
  PIN slave_data_rdata_to_inter_ro[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 296.000 1475.590 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[94]
  PIN slave_data_rdata_to_inter_ro[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.210 296.000 1482.490 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[95]
  PIN slave_data_rdata_to_inter_ro[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.650 296.000 1488.930 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[96]
  PIN slave_data_rdata_to_inter_ro[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.550 296.000 1495.830 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[97]
  PIN slave_data_rdata_to_inter_ro[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.990 296.000 1502.270 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[98]
  PIN slave_data_rdata_to_inter_ro[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.430 296.000 1508.710 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[99]
  PIN slave_data_rdata_to_inter_ro[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 296.000 748.330 300.000 ;
    END
  END slave_data_rdata_to_inter_ro[9]
  PIN slave_data_req_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 296.000 604.810 300.000 ;
    END
  END slave_data_req_to_inter_o[0]
  PIN slave_data_req_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 296.000 624.590 300.000 ;
    END
  END slave_data_req_to_inter_o[1]
  PIN slave_data_req_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 296.000 644.370 300.000 ;
    END
  END slave_data_req_to_inter_o[2]
  PIN slave_data_req_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 296.000 664.150 300.000 ;
    END
  END slave_data_req_to_inter_o[3]
  PIN slave_data_req_to_inter_ro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 296.000 606.650 300.000 ;
    END
  END slave_data_req_to_inter_ro[0]
  PIN slave_data_req_to_inter_ro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 296.000 626.890 300.000 ;
    END
  END slave_data_req_to_inter_ro[1]
  PIN slave_data_req_to_inter_ro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 296.000 646.670 300.000 ;
    END
  END slave_data_req_to_inter_ro[2]
  PIN slave_data_req_to_inter_ro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 296.000 666.450 300.000 ;
    END
  END slave_data_req_to_inter_ro[3]
  PIN slave_data_wdata_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 296.000 608.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[0]
  PIN slave_data_wdata_to_inter_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.630 296.000 1517.910 300.000 ;
    END
  END slave_data_wdata_to_inter_o[100]
  PIN slave_data_wdata_to_inter_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.070 296.000 1524.350 300.000 ;
    END
  END slave_data_wdata_to_inter_o[101]
  PIN slave_data_wdata_to_inter_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.510 296.000 1530.790 300.000 ;
    END
  END slave_data_wdata_to_inter_o[102]
  PIN slave_data_wdata_to_inter_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1537.410 296.000 1537.690 300.000 ;
    END
  END slave_data_wdata_to_inter_o[103]
  PIN slave_data_wdata_to_inter_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1543.850 296.000 1544.130 300.000 ;
    END
  END slave_data_wdata_to_inter_o[104]
  PIN slave_data_wdata_to_inter_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.750 296.000 1551.030 300.000 ;
    END
  END slave_data_wdata_to_inter_o[105]
  PIN slave_data_wdata_to_inter_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 296.000 1557.470 300.000 ;
    END
  END slave_data_wdata_to_inter_o[106]
  PIN slave_data_wdata_to_inter_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.090 296.000 1564.370 300.000 ;
    END
  END slave_data_wdata_to_inter_o[107]
  PIN slave_data_wdata_to_inter_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.530 296.000 1570.810 300.000 ;
    END
  END slave_data_wdata_to_inter_o[108]
  PIN slave_data_wdata_to_inter_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.970 296.000 1577.250 300.000 ;
    END
  END slave_data_wdata_to_inter_o[109]
  PIN slave_data_wdata_to_inter_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 296.000 763.970 300.000 ;
    END
  END slave_data_wdata_to_inter_o[10]
  PIN slave_data_wdata_to_inter_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.870 296.000 1584.150 300.000 ;
    END
  END slave_data_wdata_to_inter_o[110]
  PIN slave_data_wdata_to_inter_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.310 296.000 1590.590 300.000 ;
    END
  END slave_data_wdata_to_inter_o[111]
  PIN slave_data_wdata_to_inter_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 296.000 1597.490 300.000 ;
    END
  END slave_data_wdata_to_inter_o[112]
  PIN slave_data_wdata_to_inter_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 296.000 1603.930 300.000 ;
    END
  END slave_data_wdata_to_inter_o[113]
  PIN slave_data_wdata_to_inter_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 296.000 1610.370 300.000 ;
    END
  END slave_data_wdata_to_inter_o[114]
  PIN slave_data_wdata_to_inter_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.990 296.000 1617.270 300.000 ;
    END
  END slave_data_wdata_to_inter_o[115]
  PIN slave_data_wdata_to_inter_o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.430 296.000 1623.710 300.000 ;
    END
  END slave_data_wdata_to_inter_o[116]
  PIN slave_data_wdata_to_inter_o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.330 296.000 1630.610 300.000 ;
    END
  END slave_data_wdata_to_inter_o[117]
  PIN slave_data_wdata_to_inter_o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.770 296.000 1637.050 300.000 ;
    END
  END slave_data_wdata_to_inter_o[118]
  PIN slave_data_wdata_to_inter_o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.670 296.000 1643.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[119]
  PIN slave_data_wdata_to_inter_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 296.000 776.850 300.000 ;
    END
  END slave_data_wdata_to_inter_o[11]
  PIN slave_data_wdata_to_inter_o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.110 296.000 1650.390 300.000 ;
    END
  END slave_data_wdata_to_inter_o[120]
  PIN slave_data_wdata_to_inter_o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.550 296.000 1656.830 300.000 ;
    END
  END slave_data_wdata_to_inter_o[121]
  PIN slave_data_wdata_to_inter_o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.450 296.000 1663.730 300.000 ;
    END
  END slave_data_wdata_to_inter_o[122]
  PIN slave_data_wdata_to_inter_o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.890 296.000 1670.170 300.000 ;
    END
  END slave_data_wdata_to_inter_o[123]
  PIN slave_data_wdata_to_inter_o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.790 296.000 1677.070 300.000 ;
    END
  END slave_data_wdata_to_inter_o[124]
  PIN slave_data_wdata_to_inter_o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.230 296.000 1683.510 300.000 ;
    END
  END slave_data_wdata_to_inter_o[125]
  PIN slave_data_wdata_to_inter_o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.670 296.000 1689.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[126]
  PIN slave_data_wdata_to_inter_o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.570 296.000 1696.850 300.000 ;
    END
  END slave_data_wdata_to_inter_o[127]
  PIN slave_data_wdata_to_inter_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 296.000 790.190 300.000 ;
    END
  END slave_data_wdata_to_inter_o[12]
  PIN slave_data_wdata_to_inter_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 296.000 803.530 300.000 ;
    END
  END slave_data_wdata_to_inter_o[13]
  PIN slave_data_wdata_to_inter_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 296.000 816.870 300.000 ;
    END
  END slave_data_wdata_to_inter_o[14]
  PIN slave_data_wdata_to_inter_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.930 296.000 830.210 300.000 ;
    END
  END slave_data_wdata_to_inter_o[15]
  PIN slave_data_wdata_to_inter_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.970 296.000 841.250 300.000 ;
    END
  END slave_data_wdata_to_inter_o[16]
  PIN slave_data_wdata_to_inter_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 296.000 852.290 300.000 ;
    END
  END slave_data_wdata_to_inter_o[17]
  PIN slave_data_wdata_to_inter_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 296.000 863.330 300.000 ;
    END
  END slave_data_wdata_to_inter_o[18]
  PIN slave_data_wdata_to_inter_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 296.000 874.370 300.000 ;
    END
  END slave_data_wdata_to_inter_o[19]
  PIN slave_data_wdata_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 296.000 628.730 300.000 ;
    END
  END slave_data_wdata_to_inter_o[1]
  PIN slave_data_wdata_to_inter_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 296.000 885.410 300.000 ;
    END
  END slave_data_wdata_to_inter_o[20]
  PIN slave_data_wdata_to_inter_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 296.000 896.450 300.000 ;
    END
  END slave_data_wdata_to_inter_o[21]
  PIN slave_data_wdata_to_inter_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 296.000 907.490 300.000 ;
    END
  END slave_data_wdata_to_inter_o[22]
  PIN slave_data_wdata_to_inter_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 296.000 918.530 300.000 ;
    END
  END slave_data_wdata_to_inter_o[23]
  PIN slave_data_wdata_to_inter_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 296.000 929.570 300.000 ;
    END
  END slave_data_wdata_to_inter_o[24]
  PIN slave_data_wdata_to_inter_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 296.000 940.610 300.000 ;
    END
  END slave_data_wdata_to_inter_o[25]
  PIN slave_data_wdata_to_inter_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 296.000 951.650 300.000 ;
    END
  END slave_data_wdata_to_inter_o[26]
  PIN slave_data_wdata_to_inter_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 296.000 962.690 300.000 ;
    END
  END slave_data_wdata_to_inter_o[27]
  PIN slave_data_wdata_to_inter_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.450 296.000 973.730 300.000 ;
    END
  END slave_data_wdata_to_inter_o[28]
  PIN slave_data_wdata_to_inter_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.490 296.000 984.770 300.000 ;
    END
  END slave_data_wdata_to_inter_o[29]
  PIN slave_data_wdata_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 296.000 648.970 300.000 ;
    END
  END slave_data_wdata_to_inter_o[2]
  PIN slave_data_wdata_to_inter_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.530 296.000 995.810 300.000 ;
    END
  END slave_data_wdata_to_inter_o[30]
  PIN slave_data_wdata_to_inter_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.570 296.000 1006.850 300.000 ;
    END
  END slave_data_wdata_to_inter_o[31]
  PIN slave_data_wdata_to_inter_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 296.000 1017.890 300.000 ;
    END
  END slave_data_wdata_to_inter_o[32]
  PIN slave_data_wdata_to_inter_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 296.000 1028.930 300.000 ;
    END
  END slave_data_wdata_to_inter_o[33]
  PIN slave_data_wdata_to_inter_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.690 296.000 1039.970 300.000 ;
    END
  END slave_data_wdata_to_inter_o[34]
  PIN slave_data_wdata_to_inter_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.730 296.000 1051.010 300.000 ;
    END
  END slave_data_wdata_to_inter_o[35]
  PIN slave_data_wdata_to_inter_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.770 296.000 1062.050 300.000 ;
    END
  END slave_data_wdata_to_inter_o[36]
  PIN slave_data_wdata_to_inter_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.270 296.000 1073.550 300.000 ;
    END
  END slave_data_wdata_to_inter_o[37]
  PIN slave_data_wdata_to_inter_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 296.000 1084.590 300.000 ;
    END
  END slave_data_wdata_to_inter_o[38]
  PIN slave_data_wdata_to_inter_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 296.000 1095.630 300.000 ;
    END
  END slave_data_wdata_to_inter_o[39]
  PIN slave_data_wdata_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 296.000 668.750 300.000 ;
    END
  END slave_data_wdata_to_inter_o[3]
  PIN slave_data_wdata_to_inter_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.390 296.000 1106.670 300.000 ;
    END
  END slave_data_wdata_to_inter_o[40]
  PIN slave_data_wdata_to_inter_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 296.000 1117.710 300.000 ;
    END
  END slave_data_wdata_to_inter_o[41]
  PIN slave_data_wdata_to_inter_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 296.000 1128.750 300.000 ;
    END
  END slave_data_wdata_to_inter_o[42]
  PIN slave_data_wdata_to_inter_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.510 296.000 1139.790 300.000 ;
    END
  END slave_data_wdata_to_inter_o[43]
  PIN slave_data_wdata_to_inter_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 296.000 1146.230 300.000 ;
    END
  END slave_data_wdata_to_inter_o[44]
  PIN slave_data_wdata_to_inter_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 296.000 1153.130 300.000 ;
    END
  END slave_data_wdata_to_inter_o[45]
  PIN slave_data_wdata_to_inter_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 296.000 1159.570 300.000 ;
    END
  END slave_data_wdata_to_inter_o[46]
  PIN slave_data_wdata_to_inter_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 296.000 1166.010 300.000 ;
    END
  END slave_data_wdata_to_inter_o[47]
  PIN slave_data_wdata_to_inter_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.630 296.000 1172.910 300.000 ;
    END
  END slave_data_wdata_to_inter_o[48]
  PIN slave_data_wdata_to_inter_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.070 296.000 1179.350 300.000 ;
    END
  END slave_data_wdata_to_inter_o[49]
  PIN slave_data_wdata_to_inter_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 296.000 684.390 300.000 ;
    END
  END slave_data_wdata_to_inter_o[4]
  PIN slave_data_wdata_to_inter_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.970 296.000 1186.250 300.000 ;
    END
  END slave_data_wdata_to_inter_o[50]
  PIN slave_data_wdata_to_inter_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.410 296.000 1192.690 300.000 ;
    END
  END slave_data_wdata_to_inter_o[51]
  PIN slave_data_wdata_to_inter_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.850 296.000 1199.130 300.000 ;
    END
  END slave_data_wdata_to_inter_o[52]
  PIN slave_data_wdata_to_inter_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.750 296.000 1206.030 300.000 ;
    END
  END slave_data_wdata_to_inter_o[53]
  PIN slave_data_wdata_to_inter_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.190 296.000 1212.470 300.000 ;
    END
  END slave_data_wdata_to_inter_o[54]
  PIN slave_data_wdata_to_inter_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.090 296.000 1219.370 300.000 ;
    END
  END slave_data_wdata_to_inter_o[55]
  PIN slave_data_wdata_to_inter_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.530 296.000 1225.810 300.000 ;
    END
  END slave_data_wdata_to_inter_o[56]
  PIN slave_data_wdata_to_inter_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.430 296.000 1232.710 300.000 ;
    END
  END slave_data_wdata_to_inter_o[57]
  PIN slave_data_wdata_to_inter_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.870 296.000 1239.150 300.000 ;
    END
  END slave_data_wdata_to_inter_o[58]
  PIN slave_data_wdata_to_inter_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.310 296.000 1245.590 300.000 ;
    END
  END slave_data_wdata_to_inter_o[59]
  PIN slave_data_wdata_to_inter_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 296.000 697.270 300.000 ;
    END
  END slave_data_wdata_to_inter_o[5]
  PIN slave_data_wdata_to_inter_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.210 296.000 1252.490 300.000 ;
    END
  END slave_data_wdata_to_inter_o[60]
  PIN slave_data_wdata_to_inter_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.650 296.000 1258.930 300.000 ;
    END
  END slave_data_wdata_to_inter_o[61]
  PIN slave_data_wdata_to_inter_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 296.000 1265.830 300.000 ;
    END
  END slave_data_wdata_to_inter_o[62]
  PIN slave_data_wdata_to_inter_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 296.000 1272.270 300.000 ;
    END
  END slave_data_wdata_to_inter_o[63]
  PIN slave_data_wdata_to_inter_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.890 296.000 1279.170 300.000 ;
    END
  END slave_data_wdata_to_inter_o[64]
  PIN slave_data_wdata_to_inter_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.330 296.000 1285.610 300.000 ;
    END
  END slave_data_wdata_to_inter_o[65]
  PIN slave_data_wdata_to_inter_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.770 296.000 1292.050 300.000 ;
    END
  END slave_data_wdata_to_inter_o[66]
  PIN slave_data_wdata_to_inter_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.670 296.000 1298.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[67]
  PIN slave_data_wdata_to_inter_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.110 296.000 1305.390 300.000 ;
    END
  END slave_data_wdata_to_inter_o[68]
  PIN slave_data_wdata_to_inter_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.010 296.000 1312.290 300.000 ;
    END
  END slave_data_wdata_to_inter_o[69]
  PIN slave_data_wdata_to_inter_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 296.000 710.610 300.000 ;
    END
  END slave_data_wdata_to_inter_o[6]
  PIN slave_data_wdata_to_inter_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.450 296.000 1318.730 300.000 ;
    END
  END slave_data_wdata_to_inter_o[70]
  PIN slave_data_wdata_to_inter_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.890 296.000 1325.170 300.000 ;
    END
  END slave_data_wdata_to_inter_o[71]
  PIN slave_data_wdata_to_inter_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.790 296.000 1332.070 300.000 ;
    END
  END slave_data_wdata_to_inter_o[72]
  PIN slave_data_wdata_to_inter_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.230 296.000 1338.510 300.000 ;
    END
  END slave_data_wdata_to_inter_o[73]
  PIN slave_data_wdata_to_inter_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.130 296.000 1345.410 300.000 ;
    END
  END slave_data_wdata_to_inter_o[74]
  PIN slave_data_wdata_to_inter_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.570 296.000 1351.850 300.000 ;
    END
  END slave_data_wdata_to_inter_o[75]
  PIN slave_data_wdata_to_inter_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.470 296.000 1358.750 300.000 ;
    END
  END slave_data_wdata_to_inter_o[76]
  PIN slave_data_wdata_to_inter_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.910 296.000 1365.190 300.000 ;
    END
  END slave_data_wdata_to_inter_o[77]
  PIN slave_data_wdata_to_inter_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.350 296.000 1371.630 300.000 ;
    END
  END slave_data_wdata_to_inter_o[78]
  PIN slave_data_wdata_to_inter_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 296.000 1378.530 300.000 ;
    END
  END slave_data_wdata_to_inter_o[79]
  PIN slave_data_wdata_to_inter_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 296.000 723.950 300.000 ;
    END
  END slave_data_wdata_to_inter_o[7]
  PIN slave_data_wdata_to_inter_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.690 296.000 1384.970 300.000 ;
    END
  END slave_data_wdata_to_inter_o[80]
  PIN slave_data_wdata_to_inter_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.590 296.000 1391.870 300.000 ;
    END
  END slave_data_wdata_to_inter_o[81]
  PIN slave_data_wdata_to_inter_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.030 296.000 1398.310 300.000 ;
    END
  END slave_data_wdata_to_inter_o[82]
  PIN slave_data_wdata_to_inter_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.470 296.000 1404.750 300.000 ;
    END
  END slave_data_wdata_to_inter_o[83]
  PIN slave_data_wdata_to_inter_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.370 296.000 1411.650 300.000 ;
    END
  END slave_data_wdata_to_inter_o[84]
  PIN slave_data_wdata_to_inter_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.810 296.000 1418.090 300.000 ;
    END
  END slave_data_wdata_to_inter_o[85]
  PIN slave_data_wdata_to_inter_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.710 296.000 1424.990 300.000 ;
    END
  END slave_data_wdata_to_inter_o[86]
  PIN slave_data_wdata_to_inter_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.150 296.000 1431.430 300.000 ;
    END
  END slave_data_wdata_to_inter_o[87]
  PIN slave_data_wdata_to_inter_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.050 296.000 1438.330 300.000 ;
    END
  END slave_data_wdata_to_inter_o[88]
  PIN slave_data_wdata_to_inter_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.490 296.000 1444.770 300.000 ;
    END
  END slave_data_wdata_to_inter_o[89]
  PIN slave_data_wdata_to_inter_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 296.000 737.290 300.000 ;
    END
  END slave_data_wdata_to_inter_o[8]
  PIN slave_data_wdata_to_inter_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.930 296.000 1451.210 300.000 ;
    END
  END slave_data_wdata_to_inter_o[90]
  PIN slave_data_wdata_to_inter_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.830 296.000 1458.110 300.000 ;
    END
  END slave_data_wdata_to_inter_o[91]
  PIN slave_data_wdata_to_inter_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.270 296.000 1464.550 300.000 ;
    END
  END slave_data_wdata_to_inter_o[92]
  PIN slave_data_wdata_to_inter_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.170 296.000 1471.450 300.000 ;
    END
  END slave_data_wdata_to_inter_o[93]
  PIN slave_data_wdata_to_inter_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.610 296.000 1477.890 300.000 ;
    END
  END slave_data_wdata_to_inter_o[94]
  PIN slave_data_wdata_to_inter_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.050 296.000 1484.330 300.000 ;
    END
  END slave_data_wdata_to_inter_o[95]
  PIN slave_data_wdata_to_inter_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 296.000 1491.230 300.000 ;
    END
  END slave_data_wdata_to_inter_o[96]
  PIN slave_data_wdata_to_inter_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 296.000 1497.670 300.000 ;
    END
  END slave_data_wdata_to_inter_o[97]
  PIN slave_data_wdata_to_inter_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.290 296.000 1504.570 300.000 ;
    END
  END slave_data_wdata_to_inter_o[98]
  PIN slave_data_wdata_to_inter_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.730 296.000 1511.010 300.000 ;
    END
  END slave_data_wdata_to_inter_o[99]
  PIN slave_data_wdata_to_inter_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 296.000 750.630 300.000 ;
    END
  END slave_data_wdata_to_inter_o[9]
  PIN slave_data_we_to_inter_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 296.000 611.250 300.000 ;
    END
  END slave_data_we_to_inter_o[0]
  PIN slave_data_we_to_inter_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 296.000 631.030 300.000 ;
    END
  END slave_data_we_to_inter_o[1]
  PIN slave_data_we_to_inter_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 296.000 651.270 300.000 ;
    END
  END slave_data_we_to_inter_o[2]
  PIN slave_data_we_to_inter_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 296.000 671.050 300.000 ;
    END
  END slave_data_we_to_inter_o[3]
  PIN txd_uart
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 149.640 1700.000 150.240 ;
    END
  END txd_uart
  PIN txd_uart_to_mem
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1696.000 249.600 1700.000 250.200 ;
    END
  END txd_uart_to_mem
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.230 0.000 1660.510 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.870 0.000 1676.150 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 0.000 611.710 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 0.000 659.550 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 0.000 849.990 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 0.000 945.210 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.770 0.000 993.050 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.610 0.000 1040.890 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.990 0.000 1088.270 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.830 0.000 1136.110 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 0.000 1183.950 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 0.000 1231.330 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.890 0.000 1279.170 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.270 0.000 1326.550 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.110 0.000 1374.390 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.950 0.000 1422.230 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1469.330 0.000 1469.610 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.170 0.000 1517.450 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 0.000 1565.290 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.390 0.000 1612.670 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 0.000 866.090 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.190 0.000 913.470 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 0.000 961.310 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.870 0.000 1009.150 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.310 0.000 1199.590 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.150 0.000 1247.430 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 0.000 1342.650 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.210 0.000 1390.490 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.590 0.000 1437.870 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.430 0.000 1485.710 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.270 0.000 1533.550 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.650 0.000 1580.930 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.490 0.000 1628.770 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 0.000 484.750 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 0.000 643.450 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 0.000 786.510 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.510 0.000 1024.790 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.730 0.000 1120.010 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.570 0.000 1167.850 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.410 0.000 1215.690 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.790 0.000 1263.070 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 0.000 1310.910 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.470 0.000 1358.750 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 0.000 1406.130 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.690 0.000 1453.970 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.070 0.000 1501.350 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 0.000 1549.190 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.750 0.000 1597.030 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.130 0.000 1644.410 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1695.875 299.795 ;
      LAYER met1 ;
        RECT 0.990 9.560 1699.170 299.840 ;
      LAYER met2 ;
        RECT 1.570 295.720 2.570 299.870 ;
        RECT 3.410 295.720 4.870 299.870 ;
        RECT 5.710 295.720 7.170 299.870 ;
        RECT 8.010 295.720 9.470 299.870 ;
        RECT 10.310 295.720 11.770 299.870 ;
        RECT 12.610 295.720 13.610 299.870 ;
        RECT 14.450 295.720 15.910 299.870 ;
        RECT 16.750 295.720 18.210 299.870 ;
        RECT 19.050 295.720 20.510 299.870 ;
        RECT 21.350 295.720 22.810 299.870 ;
        RECT 23.650 295.720 24.650 299.870 ;
        RECT 25.490 295.720 26.950 299.870 ;
        RECT 27.790 295.720 29.250 299.870 ;
        RECT 30.090 295.720 31.550 299.870 ;
        RECT 32.390 295.720 33.850 299.870 ;
        RECT 34.690 295.720 35.690 299.870 ;
        RECT 36.530 295.720 37.990 299.870 ;
        RECT 38.830 295.720 40.290 299.870 ;
        RECT 41.130 295.720 42.590 299.870 ;
        RECT 43.430 295.720 44.890 299.870 ;
        RECT 45.730 295.720 46.730 299.870 ;
        RECT 47.570 295.720 49.030 299.870 ;
        RECT 49.870 295.720 51.330 299.870 ;
        RECT 52.170 295.720 53.630 299.870 ;
        RECT 54.470 295.720 55.930 299.870 ;
        RECT 56.770 295.720 57.770 299.870 ;
        RECT 58.610 295.720 60.070 299.870 ;
        RECT 60.910 295.720 62.370 299.870 ;
        RECT 63.210 295.720 64.670 299.870 ;
        RECT 65.510 295.720 66.970 299.870 ;
        RECT 67.810 295.720 68.810 299.870 ;
        RECT 69.650 295.720 71.110 299.870 ;
        RECT 71.950 295.720 73.410 299.870 ;
        RECT 74.250 295.720 75.710 299.870 ;
        RECT 76.550 295.720 78.010 299.870 ;
        RECT 78.850 295.720 80.310 299.870 ;
        RECT 81.150 295.720 82.150 299.870 ;
        RECT 82.990 295.720 84.450 299.870 ;
        RECT 85.290 295.720 86.750 299.870 ;
        RECT 87.590 295.720 89.050 299.870 ;
        RECT 89.890 295.720 91.350 299.870 ;
        RECT 92.190 295.720 93.190 299.870 ;
        RECT 94.030 295.720 95.490 299.870 ;
        RECT 96.330 295.720 97.790 299.870 ;
        RECT 98.630 295.720 100.090 299.870 ;
        RECT 100.930 295.720 102.390 299.870 ;
        RECT 103.230 295.720 104.230 299.870 ;
        RECT 105.070 295.720 106.530 299.870 ;
        RECT 107.370 295.720 108.830 299.870 ;
        RECT 109.670 295.720 111.130 299.870 ;
        RECT 111.970 295.720 113.430 299.870 ;
        RECT 114.270 295.720 115.270 299.870 ;
        RECT 116.110 295.720 117.570 299.870 ;
        RECT 118.410 295.720 119.870 299.870 ;
        RECT 120.710 295.720 122.170 299.870 ;
        RECT 123.010 295.720 124.470 299.870 ;
        RECT 125.310 295.720 126.310 299.870 ;
        RECT 127.150 295.720 128.610 299.870 ;
        RECT 129.450 295.720 130.910 299.870 ;
        RECT 131.750 295.720 133.210 299.870 ;
        RECT 134.050 295.720 135.510 299.870 ;
        RECT 136.350 295.720 137.350 299.870 ;
        RECT 138.190 295.720 139.650 299.870 ;
        RECT 140.490 295.720 141.950 299.870 ;
        RECT 142.790 295.720 144.250 299.870 ;
        RECT 145.090 295.720 146.550 299.870 ;
        RECT 147.390 295.720 148.850 299.870 ;
        RECT 149.690 295.720 150.690 299.870 ;
        RECT 151.530 295.720 152.990 299.870 ;
        RECT 153.830 295.720 155.290 299.870 ;
        RECT 156.130 295.720 157.590 299.870 ;
        RECT 158.430 295.720 159.890 299.870 ;
        RECT 160.730 295.720 161.730 299.870 ;
        RECT 162.570 295.720 164.030 299.870 ;
        RECT 164.870 295.720 166.330 299.870 ;
        RECT 167.170 295.720 168.630 299.870 ;
        RECT 169.470 295.720 170.930 299.870 ;
        RECT 171.770 295.720 172.770 299.870 ;
        RECT 173.610 295.720 175.070 299.870 ;
        RECT 175.910 295.720 177.370 299.870 ;
        RECT 178.210 295.720 179.670 299.870 ;
        RECT 180.510 295.720 181.970 299.870 ;
        RECT 182.810 295.720 183.810 299.870 ;
        RECT 184.650 295.720 186.110 299.870 ;
        RECT 186.950 295.720 188.410 299.870 ;
        RECT 189.250 295.720 190.710 299.870 ;
        RECT 191.550 295.720 193.010 299.870 ;
        RECT 193.850 295.720 194.850 299.870 ;
        RECT 195.690 295.720 197.150 299.870 ;
        RECT 197.990 295.720 199.450 299.870 ;
        RECT 200.290 295.720 201.750 299.870 ;
        RECT 202.590 295.720 204.050 299.870 ;
        RECT 204.890 295.720 205.890 299.870 ;
        RECT 206.730 295.720 208.190 299.870 ;
        RECT 209.030 295.720 210.490 299.870 ;
        RECT 211.330 295.720 212.790 299.870 ;
        RECT 213.630 295.720 215.090 299.870 ;
        RECT 215.930 295.720 217.390 299.870 ;
        RECT 218.230 295.720 219.230 299.870 ;
        RECT 220.070 295.720 221.530 299.870 ;
        RECT 222.370 295.720 223.830 299.870 ;
        RECT 224.670 295.720 226.130 299.870 ;
        RECT 226.970 295.720 228.430 299.870 ;
        RECT 229.270 295.720 230.270 299.870 ;
        RECT 231.110 295.720 232.570 299.870 ;
        RECT 233.410 295.720 234.870 299.870 ;
        RECT 235.710 295.720 237.170 299.870 ;
        RECT 238.010 295.720 239.470 299.870 ;
        RECT 240.310 295.720 241.310 299.870 ;
        RECT 242.150 295.720 243.610 299.870 ;
        RECT 244.450 295.720 245.910 299.870 ;
        RECT 246.750 295.720 248.210 299.870 ;
        RECT 249.050 295.720 250.510 299.870 ;
        RECT 251.350 295.720 252.350 299.870 ;
        RECT 253.190 295.720 254.650 299.870 ;
        RECT 255.490 295.720 256.950 299.870 ;
        RECT 257.790 295.720 259.250 299.870 ;
        RECT 260.090 295.720 261.550 299.870 ;
        RECT 262.390 295.720 263.390 299.870 ;
        RECT 264.230 295.720 265.690 299.870 ;
        RECT 266.530 295.720 267.990 299.870 ;
        RECT 268.830 295.720 270.290 299.870 ;
        RECT 271.130 295.720 272.590 299.870 ;
        RECT 273.430 295.720 274.430 299.870 ;
        RECT 275.270 295.720 276.730 299.870 ;
        RECT 277.570 295.720 279.030 299.870 ;
        RECT 279.870 295.720 281.330 299.870 ;
        RECT 282.170 295.720 283.630 299.870 ;
        RECT 284.470 295.720 285.930 299.870 ;
        RECT 286.770 295.720 287.770 299.870 ;
        RECT 288.610 295.720 290.070 299.870 ;
        RECT 290.910 295.720 292.370 299.870 ;
        RECT 293.210 295.720 294.670 299.870 ;
        RECT 295.510 295.720 296.970 299.870 ;
        RECT 297.810 295.720 298.810 299.870 ;
        RECT 299.650 295.720 301.110 299.870 ;
        RECT 301.950 295.720 303.410 299.870 ;
        RECT 304.250 295.720 305.710 299.870 ;
        RECT 306.550 295.720 308.010 299.870 ;
        RECT 308.850 295.720 309.850 299.870 ;
        RECT 310.690 295.720 312.150 299.870 ;
        RECT 312.990 295.720 314.450 299.870 ;
        RECT 315.290 295.720 316.750 299.870 ;
        RECT 317.590 295.720 319.050 299.870 ;
        RECT 319.890 295.720 320.890 299.870 ;
        RECT 321.730 295.720 323.190 299.870 ;
        RECT 324.030 295.720 325.490 299.870 ;
        RECT 326.330 295.720 327.790 299.870 ;
        RECT 328.630 295.720 330.090 299.870 ;
        RECT 330.930 295.720 331.930 299.870 ;
        RECT 332.770 295.720 334.230 299.870 ;
        RECT 335.070 295.720 336.530 299.870 ;
        RECT 337.370 295.720 338.830 299.870 ;
        RECT 339.670 295.720 341.130 299.870 ;
        RECT 341.970 295.720 342.970 299.870 ;
        RECT 343.810 295.720 345.270 299.870 ;
        RECT 346.110 295.720 347.570 299.870 ;
        RECT 348.410 295.720 349.870 299.870 ;
        RECT 350.710 295.720 352.170 299.870 ;
        RECT 353.010 295.720 354.010 299.870 ;
        RECT 354.850 295.720 356.310 299.870 ;
        RECT 357.150 295.720 358.610 299.870 ;
        RECT 359.450 295.720 360.910 299.870 ;
        RECT 361.750 295.720 363.210 299.870 ;
        RECT 364.050 295.720 365.510 299.870 ;
        RECT 366.350 295.720 367.350 299.870 ;
        RECT 368.190 295.720 369.650 299.870 ;
        RECT 370.490 295.720 371.950 299.870 ;
        RECT 372.790 295.720 374.250 299.870 ;
        RECT 375.090 295.720 376.550 299.870 ;
        RECT 377.390 295.720 378.390 299.870 ;
        RECT 379.230 295.720 380.690 299.870 ;
        RECT 381.530 295.720 382.990 299.870 ;
        RECT 383.830 295.720 385.290 299.870 ;
        RECT 386.130 295.720 387.590 299.870 ;
        RECT 388.430 295.720 389.430 299.870 ;
        RECT 390.270 295.720 391.730 299.870 ;
        RECT 392.570 295.720 394.030 299.870 ;
        RECT 394.870 295.720 396.330 299.870 ;
        RECT 397.170 295.720 398.630 299.870 ;
        RECT 399.470 295.720 400.470 299.870 ;
        RECT 401.310 295.720 402.770 299.870 ;
        RECT 403.610 295.720 405.070 299.870 ;
        RECT 405.910 295.720 407.370 299.870 ;
        RECT 408.210 295.720 409.670 299.870 ;
        RECT 410.510 295.720 411.510 299.870 ;
        RECT 412.350 295.720 413.810 299.870 ;
        RECT 414.650 295.720 416.110 299.870 ;
        RECT 416.950 295.720 418.410 299.870 ;
        RECT 419.250 295.720 420.710 299.870 ;
        RECT 421.550 295.720 422.550 299.870 ;
        RECT 423.390 295.720 424.850 299.870 ;
        RECT 425.690 295.720 427.150 299.870 ;
        RECT 427.990 295.720 429.450 299.870 ;
        RECT 430.290 295.720 431.750 299.870 ;
        RECT 432.590 295.720 434.050 299.870 ;
        RECT 434.890 295.720 435.890 299.870 ;
        RECT 436.730 295.720 438.190 299.870 ;
        RECT 439.030 295.720 440.490 299.870 ;
        RECT 441.330 295.720 442.790 299.870 ;
        RECT 443.630 295.720 445.090 299.870 ;
        RECT 445.930 295.720 446.930 299.870 ;
        RECT 447.770 295.720 449.230 299.870 ;
        RECT 450.070 295.720 451.530 299.870 ;
        RECT 452.370 295.720 453.830 299.870 ;
        RECT 454.670 295.720 456.130 299.870 ;
        RECT 456.970 295.720 457.970 299.870 ;
        RECT 458.810 295.720 460.270 299.870 ;
        RECT 461.110 295.720 462.570 299.870 ;
        RECT 463.410 295.720 464.870 299.870 ;
        RECT 465.710 295.720 467.170 299.870 ;
        RECT 468.010 295.720 469.010 299.870 ;
        RECT 469.850 295.720 471.310 299.870 ;
        RECT 472.150 295.720 473.610 299.870 ;
        RECT 474.450 295.720 475.910 299.870 ;
        RECT 476.750 295.720 478.210 299.870 ;
        RECT 479.050 295.720 480.050 299.870 ;
        RECT 480.890 295.720 482.350 299.870 ;
        RECT 483.190 295.720 484.650 299.870 ;
        RECT 485.490 295.720 486.950 299.870 ;
        RECT 487.790 295.720 489.250 299.870 ;
        RECT 490.090 295.720 491.090 299.870 ;
        RECT 491.930 295.720 493.390 299.870 ;
        RECT 494.230 295.720 495.690 299.870 ;
        RECT 496.530 295.720 497.990 299.870 ;
        RECT 498.830 295.720 500.290 299.870 ;
        RECT 501.130 295.720 502.590 299.870 ;
        RECT 503.430 295.720 504.430 299.870 ;
        RECT 505.270 295.720 506.730 299.870 ;
        RECT 507.570 295.720 509.030 299.870 ;
        RECT 509.870 295.720 511.330 299.870 ;
        RECT 512.170 295.720 513.630 299.870 ;
        RECT 514.470 295.720 515.470 299.870 ;
        RECT 516.310 295.720 517.770 299.870 ;
        RECT 518.610 295.720 520.070 299.870 ;
        RECT 520.910 295.720 522.370 299.870 ;
        RECT 523.210 295.720 524.670 299.870 ;
        RECT 525.510 295.720 526.510 299.870 ;
        RECT 527.350 295.720 528.810 299.870 ;
        RECT 529.650 295.720 531.110 299.870 ;
        RECT 531.950 295.720 533.410 299.870 ;
        RECT 534.250 295.720 535.710 299.870 ;
        RECT 536.550 295.720 537.550 299.870 ;
        RECT 538.390 295.720 539.850 299.870 ;
        RECT 540.690 295.720 542.150 299.870 ;
        RECT 542.990 295.720 544.450 299.870 ;
        RECT 545.290 295.720 546.750 299.870 ;
        RECT 547.590 295.720 548.590 299.870 ;
        RECT 549.430 295.720 550.890 299.870 ;
        RECT 551.730 295.720 553.190 299.870 ;
        RECT 554.030 295.720 555.490 299.870 ;
        RECT 556.330 295.720 557.790 299.870 ;
        RECT 558.630 295.720 559.630 299.870 ;
        RECT 560.470 295.720 561.930 299.870 ;
        RECT 562.770 295.720 564.230 299.870 ;
        RECT 565.070 295.720 566.530 299.870 ;
        RECT 567.370 295.720 568.830 299.870 ;
        RECT 569.670 295.720 571.130 299.870 ;
        RECT 571.970 295.720 572.970 299.870 ;
        RECT 573.810 295.720 575.270 299.870 ;
        RECT 576.110 295.720 577.570 299.870 ;
        RECT 578.410 295.720 579.870 299.870 ;
        RECT 580.710 295.720 582.170 299.870 ;
        RECT 583.010 295.720 584.010 299.870 ;
        RECT 584.850 295.720 586.310 299.870 ;
        RECT 587.150 295.720 588.610 299.870 ;
        RECT 589.450 295.720 590.910 299.870 ;
        RECT 591.750 295.720 593.210 299.870 ;
        RECT 594.050 295.720 595.050 299.870 ;
        RECT 595.890 295.720 597.350 299.870 ;
        RECT 598.190 295.720 599.650 299.870 ;
        RECT 600.490 295.720 601.950 299.870 ;
        RECT 602.790 295.720 604.250 299.870 ;
        RECT 605.090 295.720 606.090 299.870 ;
        RECT 606.930 295.720 608.390 299.870 ;
        RECT 609.230 295.720 610.690 299.870 ;
        RECT 611.530 295.720 612.990 299.870 ;
        RECT 613.830 295.720 615.290 299.870 ;
        RECT 616.130 295.720 617.130 299.870 ;
        RECT 617.970 295.720 619.430 299.870 ;
        RECT 620.270 295.720 621.730 299.870 ;
        RECT 622.570 295.720 624.030 299.870 ;
        RECT 624.870 295.720 626.330 299.870 ;
        RECT 627.170 295.720 628.170 299.870 ;
        RECT 629.010 295.720 630.470 299.870 ;
        RECT 631.310 295.720 632.770 299.870 ;
        RECT 633.610 295.720 635.070 299.870 ;
        RECT 635.910 295.720 637.370 299.870 ;
        RECT 638.210 295.720 639.670 299.870 ;
        RECT 640.510 295.720 641.510 299.870 ;
        RECT 642.350 295.720 643.810 299.870 ;
        RECT 644.650 295.720 646.110 299.870 ;
        RECT 646.950 295.720 648.410 299.870 ;
        RECT 649.250 295.720 650.710 299.870 ;
        RECT 651.550 295.720 652.550 299.870 ;
        RECT 653.390 295.720 654.850 299.870 ;
        RECT 655.690 295.720 657.150 299.870 ;
        RECT 657.990 295.720 659.450 299.870 ;
        RECT 660.290 295.720 661.750 299.870 ;
        RECT 662.590 295.720 663.590 299.870 ;
        RECT 664.430 295.720 665.890 299.870 ;
        RECT 666.730 295.720 668.190 299.870 ;
        RECT 669.030 295.720 670.490 299.870 ;
        RECT 671.330 295.720 672.790 299.870 ;
        RECT 673.630 295.720 674.630 299.870 ;
        RECT 675.470 295.720 676.930 299.870 ;
        RECT 677.770 295.720 679.230 299.870 ;
        RECT 680.070 295.720 681.530 299.870 ;
        RECT 682.370 295.720 683.830 299.870 ;
        RECT 684.670 295.720 685.670 299.870 ;
        RECT 686.510 295.720 687.970 299.870 ;
        RECT 688.810 295.720 690.270 299.870 ;
        RECT 691.110 295.720 692.570 299.870 ;
        RECT 693.410 295.720 694.870 299.870 ;
        RECT 695.710 295.720 696.710 299.870 ;
        RECT 697.550 295.720 699.010 299.870 ;
        RECT 699.850 295.720 701.310 299.870 ;
        RECT 702.150 295.720 703.610 299.870 ;
        RECT 704.450 295.720 705.910 299.870 ;
        RECT 706.750 295.720 707.750 299.870 ;
        RECT 708.590 295.720 710.050 299.870 ;
        RECT 710.890 295.720 712.350 299.870 ;
        RECT 713.190 295.720 714.650 299.870 ;
        RECT 715.490 295.720 716.950 299.870 ;
        RECT 717.790 295.720 719.250 299.870 ;
        RECT 720.090 295.720 721.090 299.870 ;
        RECT 721.930 295.720 723.390 299.870 ;
        RECT 724.230 295.720 725.690 299.870 ;
        RECT 726.530 295.720 727.990 299.870 ;
        RECT 728.830 295.720 730.290 299.870 ;
        RECT 731.130 295.720 732.130 299.870 ;
        RECT 732.970 295.720 734.430 299.870 ;
        RECT 735.270 295.720 736.730 299.870 ;
        RECT 737.570 295.720 739.030 299.870 ;
        RECT 739.870 295.720 741.330 299.870 ;
        RECT 742.170 295.720 743.170 299.870 ;
        RECT 744.010 295.720 745.470 299.870 ;
        RECT 746.310 295.720 747.770 299.870 ;
        RECT 748.610 295.720 750.070 299.870 ;
        RECT 750.910 295.720 752.370 299.870 ;
        RECT 753.210 295.720 754.210 299.870 ;
        RECT 755.050 295.720 756.510 299.870 ;
        RECT 757.350 295.720 758.810 299.870 ;
        RECT 759.650 295.720 761.110 299.870 ;
        RECT 761.950 295.720 763.410 299.870 ;
        RECT 764.250 295.720 765.250 299.870 ;
        RECT 766.090 295.720 767.550 299.870 ;
        RECT 768.390 295.720 769.850 299.870 ;
        RECT 770.690 295.720 772.150 299.870 ;
        RECT 772.990 295.720 774.450 299.870 ;
        RECT 775.290 295.720 776.290 299.870 ;
        RECT 777.130 295.720 778.590 299.870 ;
        RECT 779.430 295.720 780.890 299.870 ;
        RECT 781.730 295.720 783.190 299.870 ;
        RECT 784.030 295.720 785.490 299.870 ;
        RECT 786.330 295.720 787.790 299.870 ;
        RECT 788.630 295.720 789.630 299.870 ;
        RECT 790.470 295.720 791.930 299.870 ;
        RECT 792.770 295.720 794.230 299.870 ;
        RECT 795.070 295.720 796.530 299.870 ;
        RECT 797.370 295.720 798.830 299.870 ;
        RECT 799.670 295.720 800.670 299.870 ;
        RECT 801.510 295.720 802.970 299.870 ;
        RECT 803.810 295.720 805.270 299.870 ;
        RECT 806.110 295.720 807.570 299.870 ;
        RECT 808.410 295.720 809.870 299.870 ;
        RECT 810.710 295.720 811.710 299.870 ;
        RECT 812.550 295.720 814.010 299.870 ;
        RECT 814.850 295.720 816.310 299.870 ;
        RECT 817.150 295.720 818.610 299.870 ;
        RECT 819.450 295.720 820.910 299.870 ;
        RECT 821.750 295.720 822.750 299.870 ;
        RECT 823.590 295.720 825.050 299.870 ;
        RECT 825.890 295.720 827.350 299.870 ;
        RECT 828.190 295.720 829.650 299.870 ;
        RECT 830.490 295.720 831.950 299.870 ;
        RECT 832.790 295.720 833.790 299.870 ;
        RECT 834.630 295.720 836.090 299.870 ;
        RECT 836.930 295.720 838.390 299.870 ;
        RECT 839.230 295.720 840.690 299.870 ;
        RECT 841.530 295.720 842.990 299.870 ;
        RECT 843.830 295.720 844.830 299.870 ;
        RECT 845.670 295.720 847.130 299.870 ;
        RECT 847.970 295.720 849.430 299.870 ;
        RECT 850.270 295.720 851.730 299.870 ;
        RECT 852.570 295.720 854.030 299.870 ;
        RECT 854.870 295.720 856.330 299.870 ;
        RECT 857.170 295.720 858.170 299.870 ;
        RECT 859.010 295.720 860.470 299.870 ;
        RECT 861.310 295.720 862.770 299.870 ;
        RECT 863.610 295.720 865.070 299.870 ;
        RECT 865.910 295.720 867.370 299.870 ;
        RECT 868.210 295.720 869.210 299.870 ;
        RECT 870.050 295.720 871.510 299.870 ;
        RECT 872.350 295.720 873.810 299.870 ;
        RECT 874.650 295.720 876.110 299.870 ;
        RECT 876.950 295.720 878.410 299.870 ;
        RECT 879.250 295.720 880.250 299.870 ;
        RECT 881.090 295.720 882.550 299.870 ;
        RECT 883.390 295.720 884.850 299.870 ;
        RECT 885.690 295.720 887.150 299.870 ;
        RECT 887.990 295.720 889.450 299.870 ;
        RECT 890.290 295.720 891.290 299.870 ;
        RECT 892.130 295.720 893.590 299.870 ;
        RECT 894.430 295.720 895.890 299.870 ;
        RECT 896.730 295.720 898.190 299.870 ;
        RECT 899.030 295.720 900.490 299.870 ;
        RECT 901.330 295.720 902.330 299.870 ;
        RECT 903.170 295.720 904.630 299.870 ;
        RECT 905.470 295.720 906.930 299.870 ;
        RECT 907.770 295.720 909.230 299.870 ;
        RECT 910.070 295.720 911.530 299.870 ;
        RECT 912.370 295.720 913.370 299.870 ;
        RECT 914.210 295.720 915.670 299.870 ;
        RECT 916.510 295.720 917.970 299.870 ;
        RECT 918.810 295.720 920.270 299.870 ;
        RECT 921.110 295.720 922.570 299.870 ;
        RECT 923.410 295.720 924.870 299.870 ;
        RECT 925.710 295.720 926.710 299.870 ;
        RECT 927.550 295.720 929.010 299.870 ;
        RECT 929.850 295.720 931.310 299.870 ;
        RECT 932.150 295.720 933.610 299.870 ;
        RECT 934.450 295.720 935.910 299.870 ;
        RECT 936.750 295.720 937.750 299.870 ;
        RECT 938.590 295.720 940.050 299.870 ;
        RECT 940.890 295.720 942.350 299.870 ;
        RECT 943.190 295.720 944.650 299.870 ;
        RECT 945.490 295.720 946.950 299.870 ;
        RECT 947.790 295.720 948.790 299.870 ;
        RECT 949.630 295.720 951.090 299.870 ;
        RECT 951.930 295.720 953.390 299.870 ;
        RECT 954.230 295.720 955.690 299.870 ;
        RECT 956.530 295.720 957.990 299.870 ;
        RECT 958.830 295.720 959.830 299.870 ;
        RECT 960.670 295.720 962.130 299.870 ;
        RECT 962.970 295.720 964.430 299.870 ;
        RECT 965.270 295.720 966.730 299.870 ;
        RECT 967.570 295.720 969.030 299.870 ;
        RECT 969.870 295.720 970.870 299.870 ;
        RECT 971.710 295.720 973.170 299.870 ;
        RECT 974.010 295.720 975.470 299.870 ;
        RECT 976.310 295.720 977.770 299.870 ;
        RECT 978.610 295.720 980.070 299.870 ;
        RECT 980.910 295.720 981.910 299.870 ;
        RECT 982.750 295.720 984.210 299.870 ;
        RECT 985.050 295.720 986.510 299.870 ;
        RECT 987.350 295.720 988.810 299.870 ;
        RECT 989.650 295.720 991.110 299.870 ;
        RECT 991.950 295.720 993.410 299.870 ;
        RECT 994.250 295.720 995.250 299.870 ;
        RECT 996.090 295.720 997.550 299.870 ;
        RECT 998.390 295.720 999.850 299.870 ;
        RECT 1000.690 295.720 1002.150 299.870 ;
        RECT 1002.990 295.720 1004.450 299.870 ;
        RECT 1005.290 295.720 1006.290 299.870 ;
        RECT 1007.130 295.720 1008.590 299.870 ;
        RECT 1009.430 295.720 1010.890 299.870 ;
        RECT 1011.730 295.720 1013.190 299.870 ;
        RECT 1014.030 295.720 1015.490 299.870 ;
        RECT 1016.330 295.720 1017.330 299.870 ;
        RECT 1018.170 295.720 1019.630 299.870 ;
        RECT 1020.470 295.720 1021.930 299.870 ;
        RECT 1022.770 295.720 1024.230 299.870 ;
        RECT 1025.070 295.720 1026.530 299.870 ;
        RECT 1027.370 295.720 1028.370 299.870 ;
        RECT 1029.210 295.720 1030.670 299.870 ;
        RECT 1031.510 295.720 1032.970 299.870 ;
        RECT 1033.810 295.720 1035.270 299.870 ;
        RECT 1036.110 295.720 1037.570 299.870 ;
        RECT 1038.410 295.720 1039.410 299.870 ;
        RECT 1040.250 295.720 1041.710 299.870 ;
        RECT 1042.550 295.720 1044.010 299.870 ;
        RECT 1044.850 295.720 1046.310 299.870 ;
        RECT 1047.150 295.720 1048.610 299.870 ;
        RECT 1049.450 295.720 1050.450 299.870 ;
        RECT 1051.290 295.720 1052.750 299.870 ;
        RECT 1053.590 295.720 1055.050 299.870 ;
        RECT 1055.890 295.720 1057.350 299.870 ;
        RECT 1058.190 295.720 1059.650 299.870 ;
        RECT 1060.490 295.720 1061.490 299.870 ;
        RECT 1062.330 295.720 1063.790 299.870 ;
        RECT 1064.630 295.720 1066.090 299.870 ;
        RECT 1066.930 295.720 1068.390 299.870 ;
        RECT 1069.230 295.720 1070.690 299.870 ;
        RECT 1071.530 295.720 1072.990 299.870 ;
        RECT 1073.830 295.720 1074.830 299.870 ;
        RECT 1075.670 295.720 1077.130 299.870 ;
        RECT 1077.970 295.720 1079.430 299.870 ;
        RECT 1080.270 295.720 1081.730 299.870 ;
        RECT 1082.570 295.720 1084.030 299.870 ;
        RECT 1084.870 295.720 1085.870 299.870 ;
        RECT 1086.710 295.720 1088.170 299.870 ;
        RECT 1089.010 295.720 1090.470 299.870 ;
        RECT 1091.310 295.720 1092.770 299.870 ;
        RECT 1093.610 295.720 1095.070 299.870 ;
        RECT 1095.910 295.720 1096.910 299.870 ;
        RECT 1097.750 295.720 1099.210 299.870 ;
        RECT 1100.050 295.720 1101.510 299.870 ;
        RECT 1102.350 295.720 1103.810 299.870 ;
        RECT 1104.650 295.720 1106.110 299.870 ;
        RECT 1106.950 295.720 1107.950 299.870 ;
        RECT 1108.790 295.720 1110.250 299.870 ;
        RECT 1111.090 295.720 1112.550 299.870 ;
        RECT 1113.390 295.720 1114.850 299.870 ;
        RECT 1115.690 295.720 1117.150 299.870 ;
        RECT 1117.990 295.720 1118.990 299.870 ;
        RECT 1119.830 295.720 1121.290 299.870 ;
        RECT 1122.130 295.720 1123.590 299.870 ;
        RECT 1124.430 295.720 1125.890 299.870 ;
        RECT 1126.730 295.720 1128.190 299.870 ;
        RECT 1129.030 295.720 1130.030 299.870 ;
        RECT 1130.870 295.720 1132.330 299.870 ;
        RECT 1133.170 295.720 1134.630 299.870 ;
        RECT 1135.470 295.720 1136.930 299.870 ;
        RECT 1137.770 295.720 1139.230 299.870 ;
        RECT 1140.070 295.720 1141.530 299.870 ;
        RECT 1142.370 295.720 1143.370 299.870 ;
        RECT 1144.210 295.720 1145.670 299.870 ;
        RECT 1146.510 295.720 1147.970 299.870 ;
        RECT 1148.810 295.720 1150.270 299.870 ;
        RECT 1151.110 295.720 1152.570 299.870 ;
        RECT 1153.410 295.720 1154.410 299.870 ;
        RECT 1155.250 295.720 1156.710 299.870 ;
        RECT 1157.550 295.720 1159.010 299.870 ;
        RECT 1159.850 295.720 1161.310 299.870 ;
        RECT 1162.150 295.720 1163.610 299.870 ;
        RECT 1164.450 295.720 1165.450 299.870 ;
        RECT 1166.290 295.720 1167.750 299.870 ;
        RECT 1168.590 295.720 1170.050 299.870 ;
        RECT 1170.890 295.720 1172.350 299.870 ;
        RECT 1173.190 295.720 1174.650 299.870 ;
        RECT 1175.490 295.720 1176.490 299.870 ;
        RECT 1177.330 295.720 1178.790 299.870 ;
        RECT 1179.630 295.720 1181.090 299.870 ;
        RECT 1181.930 295.720 1183.390 299.870 ;
        RECT 1184.230 295.720 1185.690 299.870 ;
        RECT 1186.530 295.720 1187.530 299.870 ;
        RECT 1188.370 295.720 1189.830 299.870 ;
        RECT 1190.670 295.720 1192.130 299.870 ;
        RECT 1192.970 295.720 1194.430 299.870 ;
        RECT 1195.270 295.720 1196.730 299.870 ;
        RECT 1197.570 295.720 1198.570 299.870 ;
        RECT 1199.410 295.720 1200.870 299.870 ;
        RECT 1201.710 295.720 1203.170 299.870 ;
        RECT 1204.010 295.720 1205.470 299.870 ;
        RECT 1206.310 295.720 1207.770 299.870 ;
        RECT 1208.610 295.720 1210.070 299.870 ;
        RECT 1210.910 295.720 1211.910 299.870 ;
        RECT 1212.750 295.720 1214.210 299.870 ;
        RECT 1215.050 295.720 1216.510 299.870 ;
        RECT 1217.350 295.720 1218.810 299.870 ;
        RECT 1219.650 295.720 1221.110 299.870 ;
        RECT 1221.950 295.720 1222.950 299.870 ;
        RECT 1223.790 295.720 1225.250 299.870 ;
        RECT 1226.090 295.720 1227.550 299.870 ;
        RECT 1228.390 295.720 1229.850 299.870 ;
        RECT 1230.690 295.720 1232.150 299.870 ;
        RECT 1232.990 295.720 1233.990 299.870 ;
        RECT 1234.830 295.720 1236.290 299.870 ;
        RECT 1237.130 295.720 1238.590 299.870 ;
        RECT 1239.430 295.720 1240.890 299.870 ;
        RECT 1241.730 295.720 1243.190 299.870 ;
        RECT 1244.030 295.720 1245.030 299.870 ;
        RECT 1245.870 295.720 1247.330 299.870 ;
        RECT 1248.170 295.720 1249.630 299.870 ;
        RECT 1250.470 295.720 1251.930 299.870 ;
        RECT 1252.770 295.720 1254.230 299.870 ;
        RECT 1255.070 295.720 1256.070 299.870 ;
        RECT 1256.910 295.720 1258.370 299.870 ;
        RECT 1259.210 295.720 1260.670 299.870 ;
        RECT 1261.510 295.720 1262.970 299.870 ;
        RECT 1263.810 295.720 1265.270 299.870 ;
        RECT 1266.110 295.720 1267.110 299.870 ;
        RECT 1267.950 295.720 1269.410 299.870 ;
        RECT 1270.250 295.720 1271.710 299.870 ;
        RECT 1272.550 295.720 1274.010 299.870 ;
        RECT 1274.850 295.720 1276.310 299.870 ;
        RECT 1277.150 295.720 1278.610 299.870 ;
        RECT 1279.450 295.720 1280.450 299.870 ;
        RECT 1281.290 295.720 1282.750 299.870 ;
        RECT 1283.590 295.720 1285.050 299.870 ;
        RECT 1285.890 295.720 1287.350 299.870 ;
        RECT 1288.190 295.720 1289.650 299.870 ;
        RECT 1290.490 295.720 1291.490 299.870 ;
        RECT 1292.330 295.720 1293.790 299.870 ;
        RECT 1294.630 295.720 1296.090 299.870 ;
        RECT 1296.930 295.720 1298.390 299.870 ;
        RECT 1299.230 295.720 1300.690 299.870 ;
        RECT 1301.530 295.720 1302.530 299.870 ;
        RECT 1303.370 295.720 1304.830 299.870 ;
        RECT 1305.670 295.720 1307.130 299.870 ;
        RECT 1307.970 295.720 1309.430 299.870 ;
        RECT 1310.270 295.720 1311.730 299.870 ;
        RECT 1312.570 295.720 1313.570 299.870 ;
        RECT 1314.410 295.720 1315.870 299.870 ;
        RECT 1316.710 295.720 1318.170 299.870 ;
        RECT 1319.010 295.720 1320.470 299.870 ;
        RECT 1321.310 295.720 1322.770 299.870 ;
        RECT 1323.610 295.720 1324.610 299.870 ;
        RECT 1325.450 295.720 1326.910 299.870 ;
        RECT 1327.750 295.720 1329.210 299.870 ;
        RECT 1330.050 295.720 1331.510 299.870 ;
        RECT 1332.350 295.720 1333.810 299.870 ;
        RECT 1334.650 295.720 1335.650 299.870 ;
        RECT 1336.490 295.720 1337.950 299.870 ;
        RECT 1338.790 295.720 1340.250 299.870 ;
        RECT 1341.090 295.720 1342.550 299.870 ;
        RECT 1343.390 295.720 1344.850 299.870 ;
        RECT 1345.690 295.720 1347.150 299.870 ;
        RECT 1347.990 295.720 1348.990 299.870 ;
        RECT 1349.830 295.720 1351.290 299.870 ;
        RECT 1352.130 295.720 1353.590 299.870 ;
        RECT 1354.430 295.720 1355.890 299.870 ;
        RECT 1356.730 295.720 1358.190 299.870 ;
        RECT 1359.030 295.720 1360.030 299.870 ;
        RECT 1360.870 295.720 1362.330 299.870 ;
        RECT 1363.170 295.720 1364.630 299.870 ;
        RECT 1365.470 295.720 1366.930 299.870 ;
        RECT 1367.770 295.720 1369.230 299.870 ;
        RECT 1370.070 295.720 1371.070 299.870 ;
        RECT 1371.910 295.720 1373.370 299.870 ;
        RECT 1374.210 295.720 1375.670 299.870 ;
        RECT 1376.510 295.720 1377.970 299.870 ;
        RECT 1378.810 295.720 1380.270 299.870 ;
        RECT 1381.110 295.720 1382.110 299.870 ;
        RECT 1382.950 295.720 1384.410 299.870 ;
        RECT 1385.250 295.720 1386.710 299.870 ;
        RECT 1387.550 295.720 1389.010 299.870 ;
        RECT 1389.850 295.720 1391.310 299.870 ;
        RECT 1392.150 295.720 1393.150 299.870 ;
        RECT 1393.990 295.720 1395.450 299.870 ;
        RECT 1396.290 295.720 1397.750 299.870 ;
        RECT 1398.590 295.720 1400.050 299.870 ;
        RECT 1400.890 295.720 1402.350 299.870 ;
        RECT 1403.190 295.720 1404.190 299.870 ;
        RECT 1405.030 295.720 1406.490 299.870 ;
        RECT 1407.330 295.720 1408.790 299.870 ;
        RECT 1409.630 295.720 1411.090 299.870 ;
        RECT 1411.930 295.720 1413.390 299.870 ;
        RECT 1414.230 295.720 1415.230 299.870 ;
        RECT 1416.070 295.720 1417.530 299.870 ;
        RECT 1418.370 295.720 1419.830 299.870 ;
        RECT 1420.670 295.720 1422.130 299.870 ;
        RECT 1422.970 295.720 1424.430 299.870 ;
        RECT 1425.270 295.720 1426.730 299.870 ;
        RECT 1427.570 295.720 1428.570 299.870 ;
        RECT 1429.410 295.720 1430.870 299.870 ;
        RECT 1431.710 295.720 1433.170 299.870 ;
        RECT 1434.010 295.720 1435.470 299.870 ;
        RECT 1436.310 295.720 1437.770 299.870 ;
        RECT 1438.610 295.720 1439.610 299.870 ;
        RECT 1440.450 295.720 1441.910 299.870 ;
        RECT 1442.750 295.720 1444.210 299.870 ;
        RECT 1445.050 295.720 1446.510 299.870 ;
        RECT 1447.350 295.720 1448.810 299.870 ;
        RECT 1449.650 295.720 1450.650 299.870 ;
        RECT 1451.490 295.720 1452.950 299.870 ;
        RECT 1453.790 295.720 1455.250 299.870 ;
        RECT 1456.090 295.720 1457.550 299.870 ;
        RECT 1458.390 295.720 1459.850 299.870 ;
        RECT 1460.690 295.720 1461.690 299.870 ;
        RECT 1462.530 295.720 1463.990 299.870 ;
        RECT 1464.830 295.720 1466.290 299.870 ;
        RECT 1467.130 295.720 1468.590 299.870 ;
        RECT 1469.430 295.720 1470.890 299.870 ;
        RECT 1471.730 295.720 1472.730 299.870 ;
        RECT 1473.570 295.720 1475.030 299.870 ;
        RECT 1475.870 295.720 1477.330 299.870 ;
        RECT 1478.170 295.720 1479.630 299.870 ;
        RECT 1480.470 295.720 1481.930 299.870 ;
        RECT 1482.770 295.720 1483.770 299.870 ;
        RECT 1484.610 295.720 1486.070 299.870 ;
        RECT 1486.910 295.720 1488.370 299.870 ;
        RECT 1489.210 295.720 1490.670 299.870 ;
        RECT 1491.510 295.720 1492.970 299.870 ;
        RECT 1493.810 295.720 1495.270 299.870 ;
        RECT 1496.110 295.720 1497.110 299.870 ;
        RECT 1497.950 295.720 1499.410 299.870 ;
        RECT 1500.250 295.720 1501.710 299.870 ;
        RECT 1502.550 295.720 1504.010 299.870 ;
        RECT 1504.850 295.720 1506.310 299.870 ;
        RECT 1507.150 295.720 1508.150 299.870 ;
        RECT 1508.990 295.720 1510.450 299.870 ;
        RECT 1511.290 295.720 1512.750 299.870 ;
        RECT 1513.590 295.720 1515.050 299.870 ;
        RECT 1515.890 295.720 1517.350 299.870 ;
        RECT 1518.190 295.720 1519.190 299.870 ;
        RECT 1520.030 295.720 1521.490 299.870 ;
        RECT 1522.330 295.720 1523.790 299.870 ;
        RECT 1524.630 295.720 1526.090 299.870 ;
        RECT 1526.930 295.720 1528.390 299.870 ;
        RECT 1529.230 295.720 1530.230 299.870 ;
        RECT 1531.070 295.720 1532.530 299.870 ;
        RECT 1533.370 295.720 1534.830 299.870 ;
        RECT 1535.670 295.720 1537.130 299.870 ;
        RECT 1537.970 295.720 1539.430 299.870 ;
        RECT 1540.270 295.720 1541.270 299.870 ;
        RECT 1542.110 295.720 1543.570 299.870 ;
        RECT 1544.410 295.720 1545.870 299.870 ;
        RECT 1546.710 295.720 1548.170 299.870 ;
        RECT 1549.010 295.720 1550.470 299.870 ;
        RECT 1551.310 295.720 1552.310 299.870 ;
        RECT 1553.150 295.720 1554.610 299.870 ;
        RECT 1555.450 295.720 1556.910 299.870 ;
        RECT 1557.750 295.720 1559.210 299.870 ;
        RECT 1560.050 295.720 1561.510 299.870 ;
        RECT 1562.350 295.720 1563.810 299.870 ;
        RECT 1564.650 295.720 1565.650 299.870 ;
        RECT 1566.490 295.720 1567.950 299.870 ;
        RECT 1568.790 295.720 1570.250 299.870 ;
        RECT 1571.090 295.720 1572.550 299.870 ;
        RECT 1573.390 295.720 1574.850 299.870 ;
        RECT 1575.690 295.720 1576.690 299.870 ;
        RECT 1577.530 295.720 1578.990 299.870 ;
        RECT 1579.830 295.720 1581.290 299.870 ;
        RECT 1582.130 295.720 1583.590 299.870 ;
        RECT 1584.430 295.720 1585.890 299.870 ;
        RECT 1586.730 295.720 1587.730 299.870 ;
        RECT 1588.570 295.720 1590.030 299.870 ;
        RECT 1590.870 295.720 1592.330 299.870 ;
        RECT 1593.170 295.720 1594.630 299.870 ;
        RECT 1595.470 295.720 1596.930 299.870 ;
        RECT 1597.770 295.720 1598.770 299.870 ;
        RECT 1599.610 295.720 1601.070 299.870 ;
        RECT 1601.910 295.720 1603.370 299.870 ;
        RECT 1604.210 295.720 1605.670 299.870 ;
        RECT 1606.510 295.720 1607.970 299.870 ;
        RECT 1608.810 295.720 1609.810 299.870 ;
        RECT 1610.650 295.720 1612.110 299.870 ;
        RECT 1612.950 295.720 1614.410 299.870 ;
        RECT 1615.250 295.720 1616.710 299.870 ;
        RECT 1617.550 295.720 1619.010 299.870 ;
        RECT 1619.850 295.720 1620.850 299.870 ;
        RECT 1621.690 295.720 1623.150 299.870 ;
        RECT 1623.990 295.720 1625.450 299.870 ;
        RECT 1626.290 295.720 1627.750 299.870 ;
        RECT 1628.590 295.720 1630.050 299.870 ;
        RECT 1630.890 295.720 1632.350 299.870 ;
        RECT 1633.190 295.720 1634.190 299.870 ;
        RECT 1635.030 295.720 1636.490 299.870 ;
        RECT 1637.330 295.720 1638.790 299.870 ;
        RECT 1639.630 295.720 1641.090 299.870 ;
        RECT 1641.930 295.720 1643.390 299.870 ;
        RECT 1644.230 295.720 1645.230 299.870 ;
        RECT 1646.070 295.720 1647.530 299.870 ;
        RECT 1648.370 295.720 1649.830 299.870 ;
        RECT 1650.670 295.720 1652.130 299.870 ;
        RECT 1652.970 295.720 1654.430 299.870 ;
        RECT 1655.270 295.720 1656.270 299.870 ;
        RECT 1657.110 295.720 1658.570 299.870 ;
        RECT 1659.410 295.720 1660.870 299.870 ;
        RECT 1661.710 295.720 1663.170 299.870 ;
        RECT 1664.010 295.720 1665.470 299.870 ;
        RECT 1666.310 295.720 1667.310 299.870 ;
        RECT 1668.150 295.720 1669.610 299.870 ;
        RECT 1670.450 295.720 1671.910 299.870 ;
        RECT 1672.750 295.720 1674.210 299.870 ;
        RECT 1675.050 295.720 1676.510 299.870 ;
        RECT 1677.350 295.720 1678.350 299.870 ;
        RECT 1679.190 295.720 1680.650 299.870 ;
        RECT 1681.490 295.720 1682.950 299.870 ;
        RECT 1683.790 295.720 1685.250 299.870 ;
        RECT 1686.090 295.720 1687.550 299.870 ;
        RECT 1688.390 295.720 1689.390 299.870 ;
        RECT 1690.230 295.720 1691.690 299.870 ;
        RECT 1692.530 295.720 1693.990 299.870 ;
        RECT 1694.830 295.720 1696.290 299.870 ;
        RECT 1697.130 295.720 1698.590 299.870 ;
        RECT 1.020 4.280 1699.140 295.720 ;
        RECT 1.020 3.670 7.630 4.280 ;
        RECT 8.470 3.670 23.270 4.280 ;
        RECT 24.110 3.670 39.370 4.280 ;
        RECT 40.210 3.670 55.010 4.280 ;
        RECT 55.850 3.670 71.110 4.280 ;
        RECT 71.950 3.670 86.750 4.280 ;
        RECT 87.590 3.670 102.850 4.280 ;
        RECT 103.690 3.670 118.490 4.280 ;
        RECT 119.330 3.670 134.590 4.280 ;
        RECT 135.430 3.670 150.230 4.280 ;
        RECT 151.070 3.670 166.330 4.280 ;
        RECT 167.170 3.670 181.970 4.280 ;
        RECT 182.810 3.670 198.070 4.280 ;
        RECT 198.910 3.670 214.170 4.280 ;
        RECT 215.010 3.670 229.810 4.280 ;
        RECT 230.650 3.670 245.910 4.280 ;
        RECT 246.750 3.670 261.550 4.280 ;
        RECT 262.390 3.670 277.650 4.280 ;
        RECT 278.490 3.670 293.290 4.280 ;
        RECT 294.130 3.670 309.390 4.280 ;
        RECT 310.230 3.670 325.030 4.280 ;
        RECT 325.870 3.670 341.130 4.280 ;
        RECT 341.970 3.670 356.770 4.280 ;
        RECT 357.610 3.670 372.870 4.280 ;
        RECT 373.710 3.670 388.970 4.280 ;
        RECT 389.810 3.670 404.610 4.280 ;
        RECT 405.450 3.670 420.710 4.280 ;
        RECT 421.550 3.670 436.350 4.280 ;
        RECT 437.190 3.670 452.450 4.280 ;
        RECT 453.290 3.670 468.090 4.280 ;
        RECT 468.930 3.670 484.190 4.280 ;
        RECT 485.030 3.670 499.830 4.280 ;
        RECT 500.670 3.670 515.930 4.280 ;
        RECT 516.770 3.670 531.570 4.280 ;
        RECT 532.410 3.670 547.670 4.280 ;
        RECT 548.510 3.670 563.310 4.280 ;
        RECT 564.150 3.670 579.410 4.280 ;
        RECT 580.250 3.670 595.510 4.280 ;
        RECT 596.350 3.670 611.150 4.280 ;
        RECT 611.990 3.670 627.250 4.280 ;
        RECT 628.090 3.670 642.890 4.280 ;
        RECT 643.730 3.670 658.990 4.280 ;
        RECT 659.830 3.670 674.630 4.280 ;
        RECT 675.470 3.670 690.730 4.280 ;
        RECT 691.570 3.670 706.370 4.280 ;
        RECT 707.210 3.670 722.470 4.280 ;
        RECT 723.310 3.670 738.110 4.280 ;
        RECT 738.950 3.670 754.210 4.280 ;
        RECT 755.050 3.670 770.310 4.280 ;
        RECT 771.150 3.670 785.950 4.280 ;
        RECT 786.790 3.670 802.050 4.280 ;
        RECT 802.890 3.670 817.690 4.280 ;
        RECT 818.530 3.670 833.790 4.280 ;
        RECT 834.630 3.670 849.430 4.280 ;
        RECT 850.270 3.670 865.530 4.280 ;
        RECT 866.370 3.670 881.170 4.280 ;
        RECT 882.010 3.670 897.270 4.280 ;
        RECT 898.110 3.670 912.910 4.280 ;
        RECT 913.750 3.670 929.010 4.280 ;
        RECT 929.850 3.670 944.650 4.280 ;
        RECT 945.490 3.670 960.750 4.280 ;
        RECT 961.590 3.670 976.850 4.280 ;
        RECT 977.690 3.670 992.490 4.280 ;
        RECT 993.330 3.670 1008.590 4.280 ;
        RECT 1009.430 3.670 1024.230 4.280 ;
        RECT 1025.070 3.670 1040.330 4.280 ;
        RECT 1041.170 3.670 1055.970 4.280 ;
        RECT 1056.810 3.670 1072.070 4.280 ;
        RECT 1072.910 3.670 1087.710 4.280 ;
        RECT 1088.550 3.670 1103.810 4.280 ;
        RECT 1104.650 3.670 1119.450 4.280 ;
        RECT 1120.290 3.670 1135.550 4.280 ;
        RECT 1136.390 3.670 1151.650 4.280 ;
        RECT 1152.490 3.670 1167.290 4.280 ;
        RECT 1168.130 3.670 1183.390 4.280 ;
        RECT 1184.230 3.670 1199.030 4.280 ;
        RECT 1199.870 3.670 1215.130 4.280 ;
        RECT 1215.970 3.670 1230.770 4.280 ;
        RECT 1231.610 3.670 1246.870 4.280 ;
        RECT 1247.710 3.670 1262.510 4.280 ;
        RECT 1263.350 3.670 1278.610 4.280 ;
        RECT 1279.450 3.670 1294.250 4.280 ;
        RECT 1295.090 3.670 1310.350 4.280 ;
        RECT 1311.190 3.670 1325.990 4.280 ;
        RECT 1326.830 3.670 1342.090 4.280 ;
        RECT 1342.930 3.670 1358.190 4.280 ;
        RECT 1359.030 3.670 1373.830 4.280 ;
        RECT 1374.670 3.670 1389.930 4.280 ;
        RECT 1390.770 3.670 1405.570 4.280 ;
        RECT 1406.410 3.670 1421.670 4.280 ;
        RECT 1422.510 3.670 1437.310 4.280 ;
        RECT 1438.150 3.670 1453.410 4.280 ;
        RECT 1454.250 3.670 1469.050 4.280 ;
        RECT 1469.890 3.670 1485.150 4.280 ;
        RECT 1485.990 3.670 1500.790 4.280 ;
        RECT 1501.630 3.670 1516.890 4.280 ;
        RECT 1517.730 3.670 1532.990 4.280 ;
        RECT 1533.830 3.670 1548.630 4.280 ;
        RECT 1549.470 3.670 1564.730 4.280 ;
        RECT 1565.570 3.670 1580.370 4.280 ;
        RECT 1581.210 3.670 1596.470 4.280 ;
        RECT 1597.310 3.670 1612.110 4.280 ;
        RECT 1612.950 3.670 1628.210 4.280 ;
        RECT 1629.050 3.670 1643.850 4.280 ;
        RECT 1644.690 3.670 1659.950 4.280 ;
        RECT 1660.790 3.670 1675.590 4.280 ;
        RECT 1676.430 3.670 1691.690 4.280 ;
        RECT 1692.530 3.670 1699.140 4.280 ;
      LAYER met3 ;
        RECT 21.040 250.600 1696.000 290.865 ;
        RECT 21.040 249.200 1695.600 250.600 ;
        RECT 21.040 150.640 1696.000 249.200 ;
        RECT 21.040 149.240 1695.600 150.640 ;
        RECT 21.040 50.680 1696.000 149.240 ;
        RECT 21.040 49.280 1695.600 50.680 ;
        RECT 21.040 10.715 1696.000 49.280 ;
      LAYER met4 ;
        RECT 146.575 288.960 1306.105 290.865 ;
        RECT 146.575 74.975 174.240 288.960 ;
        RECT 176.640 74.975 251.040 288.960 ;
        RECT 253.440 74.975 327.840 288.960 ;
        RECT 330.240 74.975 404.640 288.960 ;
        RECT 407.040 74.975 481.440 288.960 ;
        RECT 483.840 74.975 558.240 288.960 ;
        RECT 560.640 74.975 635.040 288.960 ;
        RECT 637.440 74.975 711.840 288.960 ;
        RECT 714.240 74.975 788.640 288.960 ;
        RECT 791.040 74.975 865.440 288.960 ;
        RECT 867.840 74.975 942.240 288.960 ;
        RECT 944.640 74.975 1019.040 288.960 ;
        RECT 1021.440 74.975 1095.840 288.960 ;
        RECT 1098.240 74.975 1172.640 288.960 ;
        RECT 1175.040 74.975 1249.440 288.960 ;
        RECT 1251.840 74.975 1306.105 288.960 ;
  END
END soric_soc
END LIBRARY

