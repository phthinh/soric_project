magic
tech sky130A
magscale 1 2
timestamp 1640357211
<< obsli1 >>
rect 1104 765 239171 237745
<< obsm1 >>
rect 14 756 239186 237924
<< metal2 >>
rect 938 239200 994 240000
rect 2778 239200 2834 240000
rect 4710 239200 4766 240000
rect 6642 239200 6698 240000
rect 8482 239200 8538 240000
rect 10414 239200 10470 240000
rect 12346 239200 12402 240000
rect 14186 239200 14242 240000
rect 16118 239200 16174 240000
rect 18050 239200 18106 240000
rect 19982 239200 20038 240000
rect 21822 239200 21878 240000
rect 23754 239200 23810 240000
rect 25686 239200 25742 240000
rect 27526 239200 27582 240000
rect 29458 239200 29514 240000
rect 31390 239200 31446 240000
rect 33322 239200 33378 240000
rect 35162 239200 35218 240000
rect 37094 239200 37150 240000
rect 39026 239200 39082 240000
rect 40866 239200 40922 240000
rect 42798 239200 42854 240000
rect 44730 239200 44786 240000
rect 46570 239200 46626 240000
rect 48502 239200 48558 240000
rect 50434 239200 50490 240000
rect 52366 239200 52422 240000
rect 54206 239200 54262 240000
rect 56138 239200 56194 240000
rect 58070 239200 58126 240000
rect 59910 239200 59966 240000
rect 61842 239200 61898 240000
rect 63774 239200 63830 240000
rect 65706 239200 65762 240000
rect 67546 239200 67602 240000
rect 69478 239200 69534 240000
rect 71410 239200 71466 240000
rect 73250 239200 73306 240000
rect 75182 239200 75238 240000
rect 77114 239200 77170 240000
rect 78954 239200 79010 240000
rect 80886 239200 80942 240000
rect 82818 239200 82874 240000
rect 84750 239200 84806 240000
rect 86590 239200 86646 240000
rect 88522 239200 88578 240000
rect 90454 239200 90510 240000
rect 92294 239200 92350 240000
rect 94226 239200 94282 240000
rect 96158 239200 96214 240000
rect 98090 239200 98146 240000
rect 99930 239200 99986 240000
rect 101862 239200 101918 240000
rect 103794 239200 103850 240000
rect 105634 239200 105690 240000
rect 107566 239200 107622 240000
rect 109498 239200 109554 240000
rect 111338 239200 111394 240000
rect 113270 239200 113326 240000
rect 115202 239200 115258 240000
rect 117134 239200 117190 240000
rect 118974 239200 119030 240000
rect 120906 239200 120962 240000
rect 122838 239200 122894 240000
rect 124678 239200 124734 240000
rect 126610 239200 126666 240000
rect 128542 239200 128598 240000
rect 130474 239200 130530 240000
rect 132314 239200 132370 240000
rect 134246 239200 134302 240000
rect 136178 239200 136234 240000
rect 138018 239200 138074 240000
rect 139950 239200 140006 240000
rect 141882 239200 141938 240000
rect 143722 239200 143778 240000
rect 145654 239200 145710 240000
rect 147586 239200 147642 240000
rect 149518 239200 149574 240000
rect 151358 239200 151414 240000
rect 153290 239200 153346 240000
rect 155222 239200 155278 240000
rect 157062 239200 157118 240000
rect 158994 239200 159050 240000
rect 160926 239200 160982 240000
rect 162858 239200 162914 240000
rect 164698 239200 164754 240000
rect 166630 239200 166686 240000
rect 168562 239200 168618 240000
rect 170402 239200 170458 240000
rect 172334 239200 172390 240000
rect 174266 239200 174322 240000
rect 176106 239200 176162 240000
rect 178038 239200 178094 240000
rect 179970 239200 180026 240000
rect 181902 239200 181958 240000
rect 183742 239200 183798 240000
rect 185674 239200 185730 240000
rect 187606 239200 187662 240000
rect 189446 239200 189502 240000
rect 191378 239200 191434 240000
rect 193310 239200 193366 240000
rect 195242 239200 195298 240000
rect 197082 239200 197138 240000
rect 199014 239200 199070 240000
rect 200946 239200 201002 240000
rect 202786 239200 202842 240000
rect 204718 239200 204774 240000
rect 206650 239200 206706 240000
rect 208490 239200 208546 240000
rect 210422 239200 210478 240000
rect 212354 239200 212410 240000
rect 214286 239200 214342 240000
rect 216126 239200 216182 240000
rect 218058 239200 218114 240000
rect 219990 239200 220046 240000
rect 221830 239200 221886 240000
rect 223762 239200 223818 240000
rect 225694 239200 225750 240000
rect 227626 239200 227682 240000
rect 229466 239200 229522 240000
rect 231398 239200 231454 240000
rect 233330 239200 233386 240000
rect 235170 239200 235226 240000
rect 237102 239200 237158 240000
rect 239034 239200 239090 240000
rect 846 0 902 800
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5814 0 5870 800
rect 7470 0 7526 800
rect 9126 0 9182 800
rect 10782 0 10838 800
rect 12438 0 12494 800
rect 14094 0 14150 800
rect 15842 0 15898 800
rect 17498 0 17554 800
rect 19154 0 19210 800
rect 20810 0 20866 800
rect 22466 0 22522 800
rect 24122 0 24178 800
rect 25778 0 25834 800
rect 27434 0 27490 800
rect 29182 0 29238 800
rect 30838 0 30894 800
rect 32494 0 32550 800
rect 34150 0 34206 800
rect 35806 0 35862 800
rect 37462 0 37518 800
rect 39118 0 39174 800
rect 40774 0 40830 800
rect 42430 0 42486 800
rect 44178 0 44234 800
rect 45834 0 45890 800
rect 47490 0 47546 800
rect 49146 0 49202 800
rect 50802 0 50858 800
rect 52458 0 52514 800
rect 54114 0 54170 800
rect 55770 0 55826 800
rect 57518 0 57574 800
rect 59174 0 59230 800
rect 60830 0 60886 800
rect 62486 0 62542 800
rect 64142 0 64198 800
rect 65798 0 65854 800
rect 67454 0 67510 800
rect 69110 0 69166 800
rect 70766 0 70822 800
rect 72514 0 72570 800
rect 74170 0 74226 800
rect 75826 0 75882 800
rect 77482 0 77538 800
rect 79138 0 79194 800
rect 80794 0 80850 800
rect 82450 0 82506 800
rect 84106 0 84162 800
rect 85854 0 85910 800
rect 87510 0 87566 800
rect 89166 0 89222 800
rect 90822 0 90878 800
rect 92478 0 92534 800
rect 94134 0 94190 800
rect 95790 0 95846 800
rect 97446 0 97502 800
rect 99102 0 99158 800
rect 100850 0 100906 800
rect 102506 0 102562 800
rect 104162 0 104218 800
rect 105818 0 105874 800
rect 107474 0 107530 800
rect 109130 0 109186 800
rect 110786 0 110842 800
rect 112442 0 112498 800
rect 114190 0 114246 800
rect 115846 0 115902 800
rect 117502 0 117558 800
rect 119158 0 119214 800
rect 120814 0 120870 800
rect 122470 0 122526 800
rect 124126 0 124182 800
rect 125782 0 125838 800
rect 127438 0 127494 800
rect 129186 0 129242 800
rect 130842 0 130898 800
rect 132498 0 132554 800
rect 134154 0 134210 800
rect 135810 0 135866 800
rect 137466 0 137522 800
rect 139122 0 139178 800
rect 140778 0 140834 800
rect 142526 0 142582 800
rect 144182 0 144238 800
rect 145838 0 145894 800
rect 147494 0 147550 800
rect 149150 0 149206 800
rect 150806 0 150862 800
rect 152462 0 152518 800
rect 154118 0 154174 800
rect 155774 0 155830 800
rect 157522 0 157578 800
rect 159178 0 159234 800
rect 160834 0 160890 800
rect 162490 0 162546 800
rect 164146 0 164202 800
rect 165802 0 165858 800
rect 167458 0 167514 800
rect 169114 0 169170 800
rect 170862 0 170918 800
rect 172518 0 172574 800
rect 174174 0 174230 800
rect 175830 0 175886 800
rect 177486 0 177542 800
rect 179142 0 179198 800
rect 180798 0 180854 800
rect 182454 0 182510 800
rect 184110 0 184166 800
rect 185858 0 185914 800
rect 187514 0 187570 800
rect 189170 0 189226 800
rect 190826 0 190882 800
rect 192482 0 192538 800
rect 194138 0 194194 800
rect 195794 0 195850 800
rect 197450 0 197506 800
rect 199198 0 199254 800
rect 200854 0 200910 800
rect 202510 0 202566 800
rect 204166 0 204222 800
rect 205822 0 205878 800
rect 207478 0 207534 800
rect 209134 0 209190 800
rect 210790 0 210846 800
rect 212446 0 212502 800
rect 214194 0 214250 800
rect 215850 0 215906 800
rect 217506 0 217562 800
rect 219162 0 219218 800
rect 220818 0 220874 800
rect 222474 0 222530 800
rect 224130 0 224186 800
rect 225786 0 225842 800
rect 227534 0 227590 800
rect 229190 0 229246 800
rect 230846 0 230902 800
rect 232502 0 232558 800
rect 234158 0 234214 800
rect 235814 0 235870 800
rect 237470 0 237526 800
rect 239126 0 239182 800
<< obsm2 >>
rect 20 239144 882 239329
rect 1050 239144 2722 239329
rect 2890 239144 4654 239329
rect 4822 239144 6586 239329
rect 6754 239144 8426 239329
rect 8594 239144 10358 239329
rect 10526 239144 12290 239329
rect 12458 239144 14130 239329
rect 14298 239144 16062 239329
rect 16230 239144 17994 239329
rect 18162 239144 19926 239329
rect 20094 239144 21766 239329
rect 21934 239144 23698 239329
rect 23866 239144 25630 239329
rect 25798 239144 27470 239329
rect 27638 239144 29402 239329
rect 29570 239144 31334 239329
rect 31502 239144 33266 239329
rect 33434 239144 35106 239329
rect 35274 239144 37038 239329
rect 37206 239144 38970 239329
rect 39138 239144 40810 239329
rect 40978 239144 42742 239329
rect 42910 239144 44674 239329
rect 44842 239144 46514 239329
rect 46682 239144 48446 239329
rect 48614 239144 50378 239329
rect 50546 239144 52310 239329
rect 52478 239144 54150 239329
rect 54318 239144 56082 239329
rect 56250 239144 58014 239329
rect 58182 239144 59854 239329
rect 60022 239144 61786 239329
rect 61954 239144 63718 239329
rect 63886 239144 65650 239329
rect 65818 239144 67490 239329
rect 67658 239144 69422 239329
rect 69590 239144 71354 239329
rect 71522 239144 73194 239329
rect 73362 239144 75126 239329
rect 75294 239144 77058 239329
rect 77226 239144 78898 239329
rect 79066 239144 80830 239329
rect 80998 239144 82762 239329
rect 82930 239144 84694 239329
rect 84862 239144 86534 239329
rect 86702 239144 88466 239329
rect 88634 239144 90398 239329
rect 90566 239144 92238 239329
rect 92406 239144 94170 239329
rect 94338 239144 96102 239329
rect 96270 239144 98034 239329
rect 98202 239144 99874 239329
rect 100042 239144 101806 239329
rect 101974 239144 103738 239329
rect 103906 239144 105578 239329
rect 105746 239144 107510 239329
rect 107678 239144 109442 239329
rect 109610 239144 111282 239329
rect 111450 239144 113214 239329
rect 113382 239144 115146 239329
rect 115314 239144 117078 239329
rect 117246 239144 118918 239329
rect 119086 239144 120850 239329
rect 121018 239144 122782 239329
rect 122950 239144 124622 239329
rect 124790 239144 126554 239329
rect 126722 239144 128486 239329
rect 128654 239144 130418 239329
rect 130586 239144 132258 239329
rect 132426 239144 134190 239329
rect 134358 239144 136122 239329
rect 136290 239144 137962 239329
rect 138130 239144 139894 239329
rect 140062 239144 141826 239329
rect 141994 239144 143666 239329
rect 143834 239144 145598 239329
rect 145766 239144 147530 239329
rect 147698 239144 149462 239329
rect 149630 239144 151302 239329
rect 151470 239144 153234 239329
rect 153402 239144 155166 239329
rect 155334 239144 157006 239329
rect 157174 239144 158938 239329
rect 159106 239144 160870 239329
rect 161038 239144 162802 239329
rect 162970 239144 164642 239329
rect 164810 239144 166574 239329
rect 166742 239144 168506 239329
rect 168674 239144 170346 239329
rect 170514 239144 172278 239329
rect 172446 239144 174210 239329
rect 174378 239144 176050 239329
rect 176218 239144 177982 239329
rect 178150 239144 179914 239329
rect 180082 239144 181846 239329
rect 182014 239144 183686 239329
rect 183854 239144 185618 239329
rect 185786 239144 187550 239329
rect 187718 239144 189390 239329
rect 189558 239144 191322 239329
rect 191490 239144 193254 239329
rect 193422 239144 195186 239329
rect 195354 239144 197026 239329
rect 197194 239144 198958 239329
rect 199126 239144 200890 239329
rect 201058 239144 202730 239329
rect 202898 239144 204662 239329
rect 204830 239144 206594 239329
rect 206762 239144 208434 239329
rect 208602 239144 210366 239329
rect 210534 239144 212298 239329
rect 212466 239144 214230 239329
rect 214398 239144 216070 239329
rect 216238 239144 218002 239329
rect 218170 239144 219934 239329
rect 220102 239144 221774 239329
rect 221942 239144 223706 239329
rect 223874 239144 225638 239329
rect 225806 239144 227570 239329
rect 227738 239144 229410 239329
rect 229578 239144 231342 239329
rect 231510 239144 233274 239329
rect 233442 239144 235114 239329
rect 235282 239144 237046 239329
rect 237214 239144 238978 239329
rect 239146 239144 239180 239329
rect 20 856 239180 239144
rect 20 711 790 856
rect 958 711 2446 856
rect 2614 711 4102 856
rect 4270 711 5758 856
rect 5926 711 7414 856
rect 7582 711 9070 856
rect 9238 711 10726 856
rect 10894 711 12382 856
rect 12550 711 14038 856
rect 14206 711 15786 856
rect 15954 711 17442 856
rect 17610 711 19098 856
rect 19266 711 20754 856
rect 20922 711 22410 856
rect 22578 711 24066 856
rect 24234 711 25722 856
rect 25890 711 27378 856
rect 27546 711 29126 856
rect 29294 711 30782 856
rect 30950 711 32438 856
rect 32606 711 34094 856
rect 34262 711 35750 856
rect 35918 711 37406 856
rect 37574 711 39062 856
rect 39230 711 40718 856
rect 40886 711 42374 856
rect 42542 711 44122 856
rect 44290 711 45778 856
rect 45946 711 47434 856
rect 47602 711 49090 856
rect 49258 711 50746 856
rect 50914 711 52402 856
rect 52570 711 54058 856
rect 54226 711 55714 856
rect 55882 711 57462 856
rect 57630 711 59118 856
rect 59286 711 60774 856
rect 60942 711 62430 856
rect 62598 711 64086 856
rect 64254 711 65742 856
rect 65910 711 67398 856
rect 67566 711 69054 856
rect 69222 711 70710 856
rect 70878 711 72458 856
rect 72626 711 74114 856
rect 74282 711 75770 856
rect 75938 711 77426 856
rect 77594 711 79082 856
rect 79250 711 80738 856
rect 80906 711 82394 856
rect 82562 711 84050 856
rect 84218 711 85798 856
rect 85966 711 87454 856
rect 87622 711 89110 856
rect 89278 711 90766 856
rect 90934 711 92422 856
rect 92590 711 94078 856
rect 94246 711 95734 856
rect 95902 711 97390 856
rect 97558 711 99046 856
rect 99214 711 100794 856
rect 100962 711 102450 856
rect 102618 711 104106 856
rect 104274 711 105762 856
rect 105930 711 107418 856
rect 107586 711 109074 856
rect 109242 711 110730 856
rect 110898 711 112386 856
rect 112554 711 114134 856
rect 114302 711 115790 856
rect 115958 711 117446 856
rect 117614 711 119102 856
rect 119270 711 120758 856
rect 120926 711 122414 856
rect 122582 711 124070 856
rect 124238 711 125726 856
rect 125894 711 127382 856
rect 127550 711 129130 856
rect 129298 711 130786 856
rect 130954 711 132442 856
rect 132610 711 134098 856
rect 134266 711 135754 856
rect 135922 711 137410 856
rect 137578 711 139066 856
rect 139234 711 140722 856
rect 140890 711 142470 856
rect 142638 711 144126 856
rect 144294 711 145782 856
rect 145950 711 147438 856
rect 147606 711 149094 856
rect 149262 711 150750 856
rect 150918 711 152406 856
rect 152574 711 154062 856
rect 154230 711 155718 856
rect 155886 711 157466 856
rect 157634 711 159122 856
rect 159290 711 160778 856
rect 160946 711 162434 856
rect 162602 711 164090 856
rect 164258 711 165746 856
rect 165914 711 167402 856
rect 167570 711 169058 856
rect 169226 711 170806 856
rect 170974 711 172462 856
rect 172630 711 174118 856
rect 174286 711 175774 856
rect 175942 711 177430 856
rect 177598 711 179086 856
rect 179254 711 180742 856
rect 180910 711 182398 856
rect 182566 711 184054 856
rect 184222 711 185802 856
rect 185970 711 187458 856
rect 187626 711 189114 856
rect 189282 711 190770 856
rect 190938 711 192426 856
rect 192594 711 194082 856
rect 194250 711 195738 856
rect 195906 711 197394 856
rect 197562 711 199142 856
rect 199310 711 200798 856
rect 200966 711 202454 856
rect 202622 711 204110 856
rect 204278 711 205766 856
rect 205934 711 207422 856
rect 207590 711 209078 856
rect 209246 711 210734 856
rect 210902 711 212390 856
rect 212558 711 214138 856
rect 214306 711 215794 856
rect 215962 711 217450 856
rect 217618 711 219106 856
rect 219274 711 220762 856
rect 220930 711 222418 856
rect 222586 711 224074 856
rect 224242 711 225730 856
rect 225898 711 227478 856
rect 227646 711 229134 856
rect 229302 711 230790 856
rect 230958 711 232446 856
rect 232614 711 234102 856
rect 234270 711 235758 856
rect 235926 711 237414 856
rect 237582 711 239070 856
<< metal3 >>
rect 0 239096 800 239216
rect 239200 239232 240000 239352
rect 239200 237736 240000 237856
rect 0 237464 800 237584
rect 239200 236240 240000 236360
rect 0 235832 800 235952
rect 239200 234880 240000 235000
rect 0 234200 800 234320
rect 239200 233384 240000 233504
rect 0 232568 800 232688
rect 239200 231888 240000 232008
rect 0 230936 800 231056
rect 239200 230528 240000 230648
rect 0 229440 800 229560
rect 239200 229032 240000 229152
rect 0 227808 800 227928
rect 239200 227536 240000 227656
rect 0 226176 800 226296
rect 239200 226176 240000 226296
rect 0 224544 800 224664
rect 239200 224680 240000 224800
rect 239200 223184 240000 223304
rect 0 222912 800 223032
rect 239200 221688 240000 221808
rect 0 221280 800 221400
rect 239200 220328 240000 220448
rect 0 219784 800 219904
rect 239200 218832 240000 218952
rect 0 218152 800 218272
rect 239200 217336 240000 217456
rect 0 216520 800 216640
rect 239200 215976 240000 216096
rect 0 214888 800 215008
rect 239200 214480 240000 214600
rect 0 213256 800 213376
rect 239200 212984 240000 213104
rect 0 211624 800 211744
rect 239200 211624 240000 211744
rect 0 209992 800 210112
rect 239200 210128 240000 210248
rect 0 208496 800 208616
rect 239200 208632 240000 208752
rect 239200 207136 240000 207256
rect 0 206864 800 206984
rect 239200 205776 240000 205896
rect 0 205232 800 205352
rect 239200 204280 240000 204400
rect 0 203600 800 203720
rect 239200 202784 240000 202904
rect 0 201968 800 202088
rect 239200 201424 240000 201544
rect 0 200336 800 200456
rect 239200 199928 240000 200048
rect 0 198840 800 198960
rect 239200 198432 240000 198552
rect 0 197208 800 197328
rect 239200 197072 240000 197192
rect 0 195576 800 195696
rect 239200 195576 240000 195696
rect 0 193944 800 194064
rect 239200 194080 240000 194200
rect 239200 192720 240000 192840
rect 0 192312 800 192432
rect 239200 191224 240000 191344
rect 0 190680 800 190800
rect 239200 189728 240000 189848
rect 0 189048 800 189168
rect 239200 188232 240000 188352
rect 0 187552 800 187672
rect 239200 186872 240000 186992
rect 0 185920 800 186040
rect 239200 185376 240000 185496
rect 0 184288 800 184408
rect 239200 183880 240000 184000
rect 0 182656 800 182776
rect 239200 182520 240000 182640
rect 0 181024 800 181144
rect 239200 181024 240000 181144
rect 0 179392 800 179512
rect 239200 179528 240000 179648
rect 239200 178168 240000 178288
rect 0 177896 800 178016
rect 239200 176672 240000 176792
rect 0 176264 800 176384
rect 239200 175176 240000 175296
rect 0 174632 800 174752
rect 239200 173680 240000 173800
rect 0 173000 800 173120
rect 239200 172320 240000 172440
rect 0 171368 800 171488
rect 239200 170824 240000 170944
rect 0 169736 800 169856
rect 239200 169328 240000 169448
rect 0 168104 800 168224
rect 239200 167968 240000 168088
rect 0 166608 800 166728
rect 239200 166472 240000 166592
rect 0 164976 800 165096
rect 239200 164976 240000 165096
rect 239200 163616 240000 163736
rect 0 163344 800 163464
rect 239200 162120 240000 162240
rect 0 161712 800 161832
rect 239200 160624 240000 160744
rect 0 160080 800 160200
rect 239200 159128 240000 159248
rect 0 158448 800 158568
rect 239200 157768 240000 157888
rect 0 156952 800 157072
rect 239200 156272 240000 156392
rect 0 155320 800 155440
rect 239200 154776 240000 154896
rect 0 153688 800 153808
rect 239200 153416 240000 153536
rect 0 152056 800 152176
rect 239200 151920 240000 152040
rect 0 150424 800 150544
rect 239200 150424 240000 150544
rect 239200 149064 240000 149184
rect 0 148792 800 148912
rect 239200 147568 240000 147688
rect 0 147160 800 147280
rect 239200 146072 240000 146192
rect 0 145664 800 145784
rect 239200 144712 240000 144832
rect 0 144032 800 144152
rect 239200 143216 240000 143336
rect 0 142400 800 142520
rect 239200 141720 240000 141840
rect 0 140768 800 140888
rect 239200 140224 240000 140344
rect 0 139136 800 139256
rect 239200 138864 240000 138984
rect 0 137504 800 137624
rect 239200 137368 240000 137488
rect 0 136008 800 136128
rect 239200 135872 240000 135992
rect 0 134376 800 134496
rect 239200 134512 240000 134632
rect 239200 133016 240000 133136
rect 0 132744 800 132864
rect 239200 131520 240000 131640
rect 0 131112 800 131232
rect 239200 130160 240000 130280
rect 0 129480 800 129600
rect 239200 128664 240000 128784
rect 0 127848 800 127968
rect 239200 127168 240000 127288
rect 0 126216 800 126336
rect 239200 125672 240000 125792
rect 0 124720 800 124840
rect 239200 124312 240000 124432
rect 0 123088 800 123208
rect 239200 122816 240000 122936
rect 0 121456 800 121576
rect 239200 121320 240000 121440
rect 0 119824 800 119944
rect 239200 119960 240000 120080
rect 239200 118464 240000 118584
rect 0 118192 800 118312
rect 239200 116968 240000 117088
rect 0 116560 800 116680
rect 239200 115608 240000 115728
rect 0 115064 800 115184
rect 239200 114112 240000 114232
rect 0 113432 800 113552
rect 239200 112616 240000 112736
rect 0 111800 800 111920
rect 239200 111120 240000 111240
rect 0 110168 800 110288
rect 239200 109760 240000 109880
rect 0 108536 800 108656
rect 239200 108264 240000 108384
rect 0 106904 800 107024
rect 239200 106768 240000 106888
rect 0 105272 800 105392
rect 239200 105408 240000 105528
rect 0 103776 800 103896
rect 239200 103912 240000 104032
rect 239200 102416 240000 102536
rect 0 102144 800 102264
rect 239200 101056 240000 101176
rect 0 100512 800 100632
rect 239200 99560 240000 99680
rect 0 98880 800 99000
rect 239200 98064 240000 98184
rect 0 97248 800 97368
rect 239200 96704 240000 96824
rect 0 95616 800 95736
rect 239200 95208 240000 95328
rect 0 94120 800 94240
rect 239200 93712 240000 93832
rect 0 92488 800 92608
rect 239200 92216 240000 92336
rect 0 90856 800 90976
rect 239200 90856 240000 90976
rect 0 89224 800 89344
rect 239200 89360 240000 89480
rect 239200 87864 240000 87984
rect 0 87592 800 87712
rect 239200 86504 240000 86624
rect 0 85960 800 86080
rect 239200 85008 240000 85128
rect 0 84328 800 84448
rect 239200 83512 240000 83632
rect 0 82832 800 82952
rect 239200 82152 240000 82272
rect 0 81200 800 81320
rect 239200 80656 240000 80776
rect 0 79568 800 79688
rect 239200 79160 240000 79280
rect 0 77936 800 78056
rect 239200 77664 240000 77784
rect 0 76304 800 76424
rect 239200 76304 240000 76424
rect 0 74672 800 74792
rect 239200 74808 240000 74928
rect 0 73176 800 73296
rect 239200 73312 240000 73432
rect 239200 71952 240000 72072
rect 0 71544 800 71664
rect 239200 70456 240000 70576
rect 0 69912 800 70032
rect 239200 68960 240000 69080
rect 0 68280 800 68400
rect 239200 67600 240000 67720
rect 0 66648 800 66768
rect 239200 66104 240000 66224
rect 0 65016 800 65136
rect 239200 64608 240000 64728
rect 0 63384 800 63504
rect 239200 63112 240000 63232
rect 0 61888 800 62008
rect 239200 61752 240000 61872
rect 0 60256 800 60376
rect 239200 60256 240000 60376
rect 0 58624 800 58744
rect 239200 58760 240000 58880
rect 239200 57400 240000 57520
rect 0 56992 800 57112
rect 239200 55904 240000 56024
rect 0 55360 800 55480
rect 239200 54408 240000 54528
rect 0 53728 800 53848
rect 239200 53048 240000 53168
rect 0 52232 800 52352
rect 239200 51552 240000 51672
rect 0 50600 800 50720
rect 239200 50056 240000 50176
rect 0 48968 800 49088
rect 239200 48696 240000 48816
rect 0 47336 800 47456
rect 239200 47200 240000 47320
rect 0 45704 800 45824
rect 239200 45704 240000 45824
rect 0 44072 800 44192
rect 239200 44208 240000 44328
rect 239200 42848 240000 42968
rect 0 42440 800 42560
rect 239200 41352 240000 41472
rect 0 40944 800 41064
rect 239200 39856 240000 39976
rect 0 39312 800 39432
rect 239200 38496 240000 38616
rect 0 37680 800 37800
rect 239200 37000 240000 37120
rect 0 36048 800 36168
rect 239200 35504 240000 35624
rect 0 34416 800 34536
rect 239200 34144 240000 34264
rect 0 32784 800 32904
rect 239200 32648 240000 32768
rect 0 31288 800 31408
rect 239200 31152 240000 31272
rect 0 29656 800 29776
rect 239200 29656 240000 29776
rect 239200 28296 240000 28416
rect 0 28024 800 28144
rect 239200 26800 240000 26920
rect 0 26392 800 26512
rect 239200 25304 240000 25424
rect 0 24760 800 24880
rect 239200 23944 240000 24064
rect 0 23128 800 23248
rect 239200 22448 240000 22568
rect 0 21496 800 21616
rect 239200 20952 240000 21072
rect 0 20000 800 20120
rect 239200 19592 240000 19712
rect 0 18368 800 18488
rect 239200 18096 240000 18216
rect 0 16736 800 16856
rect 239200 16600 240000 16720
rect 0 15104 800 15224
rect 239200 15104 240000 15224
rect 239200 13744 240000 13864
rect 0 13472 800 13592
rect 239200 12248 240000 12368
rect 0 11840 800 11960
rect 239200 10752 240000 10872
rect 0 10344 800 10464
rect 239200 9392 240000 9512
rect 0 8712 800 8832
rect 239200 7896 240000 8016
rect 0 7080 800 7200
rect 239200 6400 240000 6520
rect 0 5448 800 5568
rect 239200 5040 240000 5160
rect 0 3816 800 3936
rect 239200 3544 240000 3664
rect 0 2184 800 2304
rect 239200 2048 240000 2168
rect 0 688 800 808
rect 239200 688 240000 808
<< obsm3 >>
rect 105 239296 239120 239325
rect 880 239152 239120 239296
rect 880 239016 239322 239152
rect 105 237936 239322 239016
rect 105 237664 239120 237936
rect 880 237656 239120 237664
rect 880 237384 239322 237656
rect 105 236440 239322 237384
rect 105 236160 239120 236440
rect 105 236032 239322 236160
rect 880 235752 239322 236032
rect 105 235080 239322 235752
rect 105 234800 239120 235080
rect 105 234400 239322 234800
rect 880 234120 239322 234400
rect 105 233584 239322 234120
rect 105 233304 239120 233584
rect 105 232768 239322 233304
rect 880 232488 239322 232768
rect 105 232088 239322 232488
rect 105 231808 239120 232088
rect 105 231136 239322 231808
rect 880 230856 239322 231136
rect 105 230728 239322 230856
rect 105 230448 239120 230728
rect 105 229640 239322 230448
rect 880 229360 239322 229640
rect 105 229232 239322 229360
rect 105 228952 239120 229232
rect 105 228008 239322 228952
rect 880 227736 239322 228008
rect 880 227728 239120 227736
rect 105 227456 239120 227728
rect 105 226376 239322 227456
rect 880 226096 239120 226376
rect 105 224880 239322 226096
rect 105 224744 239120 224880
rect 880 224600 239120 224744
rect 880 224464 239322 224600
rect 105 223384 239322 224464
rect 105 223112 239120 223384
rect 880 223104 239120 223112
rect 880 222832 239322 223104
rect 105 221888 239322 222832
rect 105 221608 239120 221888
rect 105 221480 239322 221608
rect 880 221200 239322 221480
rect 105 220528 239322 221200
rect 105 220248 239120 220528
rect 105 219984 239322 220248
rect 880 219704 239322 219984
rect 105 219032 239322 219704
rect 105 218752 239120 219032
rect 105 218352 239322 218752
rect 880 218072 239322 218352
rect 105 217536 239322 218072
rect 105 217256 239120 217536
rect 105 216720 239322 217256
rect 880 216440 239322 216720
rect 105 216176 239322 216440
rect 105 215896 239120 216176
rect 105 215088 239322 215896
rect 880 214808 239322 215088
rect 105 214680 239322 214808
rect 105 214400 239120 214680
rect 105 213456 239322 214400
rect 880 213184 239322 213456
rect 880 213176 239120 213184
rect 105 212904 239120 213176
rect 105 211824 239322 212904
rect 880 211544 239120 211824
rect 105 210328 239322 211544
rect 105 210192 239120 210328
rect 880 210048 239120 210192
rect 880 209912 239322 210048
rect 105 208832 239322 209912
rect 105 208696 239120 208832
rect 880 208552 239120 208696
rect 880 208416 239322 208552
rect 105 207336 239322 208416
rect 105 207064 239120 207336
rect 880 207056 239120 207064
rect 880 206784 239322 207056
rect 105 205976 239322 206784
rect 105 205696 239120 205976
rect 105 205432 239322 205696
rect 880 205152 239322 205432
rect 105 204480 239322 205152
rect 105 204200 239120 204480
rect 105 203800 239322 204200
rect 880 203520 239322 203800
rect 105 202984 239322 203520
rect 105 202704 239120 202984
rect 105 202168 239322 202704
rect 880 201888 239322 202168
rect 105 201624 239322 201888
rect 105 201344 239120 201624
rect 105 200536 239322 201344
rect 880 200256 239322 200536
rect 105 200128 239322 200256
rect 105 199848 239120 200128
rect 105 199040 239322 199848
rect 880 198760 239322 199040
rect 105 198632 239322 198760
rect 105 198352 239120 198632
rect 105 197408 239322 198352
rect 880 197272 239322 197408
rect 880 197128 239120 197272
rect 105 196992 239120 197128
rect 105 195776 239322 196992
rect 880 195496 239120 195776
rect 105 194280 239322 195496
rect 105 194144 239120 194280
rect 880 194000 239120 194144
rect 880 193864 239322 194000
rect 105 192920 239322 193864
rect 105 192640 239120 192920
rect 105 192512 239322 192640
rect 880 192232 239322 192512
rect 105 191424 239322 192232
rect 105 191144 239120 191424
rect 105 190880 239322 191144
rect 880 190600 239322 190880
rect 105 189928 239322 190600
rect 105 189648 239120 189928
rect 105 189248 239322 189648
rect 880 188968 239322 189248
rect 105 188432 239322 188968
rect 105 188152 239120 188432
rect 105 187752 239322 188152
rect 880 187472 239322 187752
rect 105 187072 239322 187472
rect 105 186792 239120 187072
rect 105 186120 239322 186792
rect 880 185840 239322 186120
rect 105 185576 239322 185840
rect 105 185296 239120 185576
rect 105 184488 239322 185296
rect 880 184208 239322 184488
rect 105 184080 239322 184208
rect 105 183800 239120 184080
rect 105 182856 239322 183800
rect 880 182720 239322 182856
rect 880 182576 239120 182720
rect 105 182440 239120 182576
rect 105 181224 239322 182440
rect 880 180944 239120 181224
rect 105 179728 239322 180944
rect 105 179592 239120 179728
rect 880 179448 239120 179592
rect 880 179312 239322 179448
rect 105 178368 239322 179312
rect 105 178096 239120 178368
rect 880 178088 239120 178096
rect 880 177816 239322 178088
rect 105 176872 239322 177816
rect 105 176592 239120 176872
rect 105 176464 239322 176592
rect 880 176184 239322 176464
rect 105 175376 239322 176184
rect 105 175096 239120 175376
rect 105 174832 239322 175096
rect 880 174552 239322 174832
rect 105 173880 239322 174552
rect 105 173600 239120 173880
rect 105 173200 239322 173600
rect 880 172920 239322 173200
rect 105 172520 239322 172920
rect 105 172240 239120 172520
rect 105 171568 239322 172240
rect 880 171288 239322 171568
rect 105 171024 239322 171288
rect 105 170744 239120 171024
rect 105 169936 239322 170744
rect 880 169656 239322 169936
rect 105 169528 239322 169656
rect 105 169248 239120 169528
rect 105 168304 239322 169248
rect 880 168168 239322 168304
rect 880 168024 239120 168168
rect 105 167888 239120 168024
rect 105 166808 239322 167888
rect 880 166672 239322 166808
rect 880 166528 239120 166672
rect 105 166392 239120 166528
rect 105 165176 239322 166392
rect 880 164896 239120 165176
rect 105 163816 239322 164896
rect 105 163544 239120 163816
rect 880 163536 239120 163544
rect 880 163264 239322 163536
rect 105 162320 239322 163264
rect 105 162040 239120 162320
rect 105 161912 239322 162040
rect 880 161632 239322 161912
rect 105 160824 239322 161632
rect 105 160544 239120 160824
rect 105 160280 239322 160544
rect 880 160000 239322 160280
rect 105 159328 239322 160000
rect 105 159048 239120 159328
rect 105 158648 239322 159048
rect 880 158368 239322 158648
rect 105 157968 239322 158368
rect 105 157688 239120 157968
rect 105 157152 239322 157688
rect 880 156872 239322 157152
rect 105 156472 239322 156872
rect 105 156192 239120 156472
rect 105 155520 239322 156192
rect 880 155240 239322 155520
rect 105 154976 239322 155240
rect 105 154696 239120 154976
rect 105 153888 239322 154696
rect 880 153616 239322 153888
rect 880 153608 239120 153616
rect 105 153336 239120 153608
rect 105 152256 239322 153336
rect 880 152120 239322 152256
rect 880 151976 239120 152120
rect 105 151840 239120 151976
rect 105 150624 239322 151840
rect 880 150344 239120 150624
rect 105 149264 239322 150344
rect 105 148992 239120 149264
rect 880 148984 239120 148992
rect 880 148712 239322 148984
rect 105 147768 239322 148712
rect 105 147488 239120 147768
rect 105 147360 239322 147488
rect 880 147080 239322 147360
rect 105 146272 239322 147080
rect 105 145992 239120 146272
rect 105 145864 239322 145992
rect 880 145584 239322 145864
rect 105 144912 239322 145584
rect 105 144632 239120 144912
rect 105 144232 239322 144632
rect 880 143952 239322 144232
rect 105 143416 239322 143952
rect 105 143136 239120 143416
rect 105 142600 239322 143136
rect 880 142320 239322 142600
rect 105 141920 239322 142320
rect 105 141640 239120 141920
rect 105 140968 239322 141640
rect 880 140688 239322 140968
rect 105 140424 239322 140688
rect 105 140144 239120 140424
rect 105 139336 239322 140144
rect 880 139064 239322 139336
rect 880 139056 239120 139064
rect 105 138784 239120 139056
rect 105 137704 239322 138784
rect 880 137568 239322 137704
rect 880 137424 239120 137568
rect 105 137288 239120 137424
rect 105 136208 239322 137288
rect 880 136072 239322 136208
rect 880 135928 239120 136072
rect 105 135792 239120 135928
rect 105 134712 239322 135792
rect 105 134576 239120 134712
rect 880 134432 239120 134576
rect 880 134296 239322 134432
rect 105 133216 239322 134296
rect 105 132944 239120 133216
rect 880 132936 239120 132944
rect 880 132664 239322 132936
rect 105 131720 239322 132664
rect 105 131440 239120 131720
rect 105 131312 239322 131440
rect 880 131032 239322 131312
rect 105 130360 239322 131032
rect 105 130080 239120 130360
rect 105 129680 239322 130080
rect 880 129400 239322 129680
rect 105 128864 239322 129400
rect 105 128584 239120 128864
rect 105 128048 239322 128584
rect 880 127768 239322 128048
rect 105 127368 239322 127768
rect 105 127088 239120 127368
rect 105 126416 239322 127088
rect 880 126136 239322 126416
rect 105 125872 239322 126136
rect 105 125592 239120 125872
rect 105 124920 239322 125592
rect 880 124640 239322 124920
rect 105 124512 239322 124640
rect 105 124232 239120 124512
rect 105 123288 239322 124232
rect 880 123016 239322 123288
rect 880 123008 239120 123016
rect 105 122736 239120 123008
rect 105 121656 239322 122736
rect 880 121520 239322 121656
rect 880 121376 239120 121520
rect 105 121240 239120 121376
rect 105 120160 239322 121240
rect 105 120024 239120 120160
rect 880 119880 239120 120024
rect 880 119744 239322 119880
rect 105 118664 239322 119744
rect 105 118392 239120 118664
rect 880 118384 239120 118392
rect 880 118112 239322 118384
rect 105 117168 239322 118112
rect 105 116888 239120 117168
rect 105 116760 239322 116888
rect 880 116480 239322 116760
rect 105 115808 239322 116480
rect 105 115528 239120 115808
rect 105 115264 239322 115528
rect 880 114984 239322 115264
rect 105 114312 239322 114984
rect 105 114032 239120 114312
rect 105 113632 239322 114032
rect 880 113352 239322 113632
rect 105 112816 239322 113352
rect 105 112536 239120 112816
rect 105 112000 239322 112536
rect 880 111720 239322 112000
rect 105 111320 239322 111720
rect 105 111040 239120 111320
rect 105 110368 239322 111040
rect 880 110088 239322 110368
rect 105 109960 239322 110088
rect 105 109680 239120 109960
rect 105 108736 239322 109680
rect 880 108464 239322 108736
rect 880 108456 239120 108464
rect 105 108184 239120 108456
rect 105 107104 239322 108184
rect 880 106968 239322 107104
rect 880 106824 239120 106968
rect 105 106688 239120 106824
rect 105 105608 239322 106688
rect 105 105472 239120 105608
rect 880 105328 239120 105472
rect 880 105192 239322 105328
rect 105 104112 239322 105192
rect 105 103976 239120 104112
rect 880 103832 239120 103976
rect 880 103696 239322 103832
rect 105 102616 239322 103696
rect 105 102344 239120 102616
rect 880 102336 239120 102344
rect 880 102064 239322 102336
rect 105 101256 239322 102064
rect 105 100976 239120 101256
rect 105 100712 239322 100976
rect 880 100432 239322 100712
rect 105 99760 239322 100432
rect 105 99480 239120 99760
rect 105 99080 239322 99480
rect 880 98800 239322 99080
rect 105 98264 239322 98800
rect 105 97984 239120 98264
rect 105 97448 239322 97984
rect 880 97168 239322 97448
rect 105 96904 239322 97168
rect 105 96624 239120 96904
rect 105 95816 239322 96624
rect 880 95536 239322 95816
rect 105 95408 239322 95536
rect 105 95128 239120 95408
rect 105 94320 239322 95128
rect 880 94040 239322 94320
rect 105 93912 239322 94040
rect 105 93632 239120 93912
rect 105 92688 239322 93632
rect 880 92416 239322 92688
rect 880 92408 239120 92416
rect 105 92136 239120 92408
rect 105 91056 239322 92136
rect 880 90776 239120 91056
rect 105 89560 239322 90776
rect 105 89424 239120 89560
rect 880 89280 239120 89424
rect 880 89144 239322 89280
rect 105 88064 239322 89144
rect 105 87792 239120 88064
rect 880 87784 239120 87792
rect 880 87512 239322 87784
rect 105 86704 239322 87512
rect 105 86424 239120 86704
rect 105 86160 239322 86424
rect 880 85880 239322 86160
rect 105 85208 239322 85880
rect 105 84928 239120 85208
rect 105 84528 239322 84928
rect 880 84248 239322 84528
rect 105 83712 239322 84248
rect 105 83432 239120 83712
rect 105 83032 239322 83432
rect 880 82752 239322 83032
rect 105 82352 239322 82752
rect 105 82072 239120 82352
rect 105 81400 239322 82072
rect 880 81120 239322 81400
rect 105 80856 239322 81120
rect 105 80576 239120 80856
rect 105 79768 239322 80576
rect 880 79488 239322 79768
rect 105 79360 239322 79488
rect 105 79080 239120 79360
rect 105 78136 239322 79080
rect 880 77864 239322 78136
rect 880 77856 239120 77864
rect 105 77584 239120 77856
rect 105 76504 239322 77584
rect 880 76224 239120 76504
rect 105 75008 239322 76224
rect 105 74872 239120 75008
rect 880 74728 239120 74872
rect 880 74592 239322 74728
rect 105 73512 239322 74592
rect 105 73376 239120 73512
rect 880 73232 239120 73376
rect 880 73096 239322 73232
rect 105 72152 239322 73096
rect 105 71872 239120 72152
rect 105 71744 239322 71872
rect 880 71464 239322 71744
rect 105 70656 239322 71464
rect 105 70376 239120 70656
rect 105 70112 239322 70376
rect 880 69832 239322 70112
rect 105 69160 239322 69832
rect 105 68880 239120 69160
rect 105 68480 239322 68880
rect 880 68200 239322 68480
rect 105 67800 239322 68200
rect 105 67520 239120 67800
rect 105 66848 239322 67520
rect 880 66568 239322 66848
rect 105 66304 239322 66568
rect 105 66024 239120 66304
rect 105 65216 239322 66024
rect 880 64936 239322 65216
rect 105 64808 239322 64936
rect 105 64528 239120 64808
rect 105 63584 239322 64528
rect 880 63312 239322 63584
rect 880 63304 239120 63312
rect 105 63032 239120 63304
rect 105 62088 239322 63032
rect 880 61952 239322 62088
rect 880 61808 239120 61952
rect 105 61672 239120 61808
rect 105 60456 239322 61672
rect 880 60176 239120 60456
rect 105 58960 239322 60176
rect 105 58824 239120 58960
rect 880 58680 239120 58824
rect 880 58544 239322 58680
rect 105 57600 239322 58544
rect 105 57320 239120 57600
rect 105 57192 239322 57320
rect 880 56912 239322 57192
rect 105 56104 239322 56912
rect 105 55824 239120 56104
rect 105 55560 239322 55824
rect 880 55280 239322 55560
rect 105 54608 239322 55280
rect 105 54328 239120 54608
rect 105 53928 239322 54328
rect 880 53648 239322 53928
rect 105 53248 239322 53648
rect 105 52968 239120 53248
rect 105 52432 239322 52968
rect 880 52152 239322 52432
rect 105 51752 239322 52152
rect 105 51472 239120 51752
rect 105 50800 239322 51472
rect 880 50520 239322 50800
rect 105 50256 239322 50520
rect 105 49976 239120 50256
rect 105 49168 239322 49976
rect 880 48896 239322 49168
rect 880 48888 239120 48896
rect 105 48616 239120 48888
rect 105 47536 239322 48616
rect 880 47400 239322 47536
rect 880 47256 239120 47400
rect 105 47120 239120 47256
rect 105 45904 239322 47120
rect 880 45624 239120 45904
rect 105 44408 239322 45624
rect 105 44272 239120 44408
rect 880 44128 239120 44272
rect 880 43992 239322 44128
rect 105 43048 239322 43992
rect 105 42768 239120 43048
rect 105 42640 239322 42768
rect 880 42360 239322 42640
rect 105 41552 239322 42360
rect 105 41272 239120 41552
rect 105 41144 239322 41272
rect 880 40864 239322 41144
rect 105 40056 239322 40864
rect 105 39776 239120 40056
rect 105 39512 239322 39776
rect 880 39232 239322 39512
rect 105 38696 239322 39232
rect 105 38416 239120 38696
rect 105 37880 239322 38416
rect 880 37600 239322 37880
rect 105 37200 239322 37600
rect 105 36920 239120 37200
rect 105 36248 239322 36920
rect 880 35968 239322 36248
rect 105 35704 239322 35968
rect 105 35424 239120 35704
rect 105 34616 239322 35424
rect 880 34344 239322 34616
rect 880 34336 239120 34344
rect 105 34064 239120 34336
rect 105 32984 239322 34064
rect 880 32848 239322 32984
rect 880 32704 239120 32848
rect 105 32568 239120 32704
rect 105 31488 239322 32568
rect 880 31352 239322 31488
rect 880 31208 239120 31352
rect 105 31072 239120 31208
rect 105 29856 239322 31072
rect 880 29576 239120 29856
rect 105 28496 239322 29576
rect 105 28224 239120 28496
rect 880 28216 239120 28224
rect 880 27944 239322 28216
rect 105 27000 239322 27944
rect 105 26720 239120 27000
rect 105 26592 239322 26720
rect 880 26312 239322 26592
rect 105 25504 239322 26312
rect 105 25224 239120 25504
rect 105 24960 239322 25224
rect 880 24680 239322 24960
rect 105 24144 239322 24680
rect 105 23864 239120 24144
rect 105 23328 239322 23864
rect 880 23048 239322 23328
rect 105 22648 239322 23048
rect 105 22368 239120 22648
rect 105 21696 239322 22368
rect 880 21416 239322 21696
rect 105 21152 239322 21416
rect 105 20872 239120 21152
rect 105 20200 239322 20872
rect 880 19920 239322 20200
rect 105 19792 239322 19920
rect 105 19512 239120 19792
rect 105 18568 239322 19512
rect 880 18296 239322 18568
rect 880 18288 239120 18296
rect 105 18016 239120 18288
rect 105 16936 239322 18016
rect 880 16800 239322 16936
rect 880 16656 239120 16800
rect 105 16520 239120 16656
rect 105 15304 239322 16520
rect 880 15024 239120 15304
rect 105 13944 239322 15024
rect 105 13672 239120 13944
rect 880 13664 239120 13672
rect 880 13392 239322 13664
rect 105 12448 239322 13392
rect 105 12168 239120 12448
rect 105 12040 239322 12168
rect 880 11760 239322 12040
rect 105 10952 239322 11760
rect 105 10672 239120 10952
rect 105 10544 239322 10672
rect 880 10264 239322 10544
rect 105 9592 239322 10264
rect 105 9312 239120 9592
rect 105 8912 239322 9312
rect 880 8632 239322 8912
rect 105 8096 239322 8632
rect 105 7816 239120 8096
rect 105 7280 239322 7816
rect 880 7000 239322 7280
rect 105 6600 239322 7000
rect 105 6320 239120 6600
rect 105 5648 239322 6320
rect 880 5368 239322 5648
rect 105 5240 239322 5368
rect 105 4960 239120 5240
rect 105 4016 239322 4960
rect 880 3744 239322 4016
rect 880 3736 239120 3744
rect 105 3464 239120 3736
rect 105 2384 239322 3464
rect 880 2248 239322 2384
rect 880 2104 239120 2248
rect 105 1968 239120 2104
rect 105 888 239322 1968
rect 880 715 239120 888
<< metal4 >>
rect 4208 2128 4528 237776
rect 9208 2128 9528 237776
rect 14208 2128 14528 237776
rect 19208 2128 19528 237776
rect 24208 2128 24528 237776
rect 29208 2128 29528 237776
rect 34208 2128 34528 237776
rect 39208 2128 39528 237776
rect 44208 2128 44528 237776
rect 49208 2128 49528 237776
rect 54208 2128 54528 237776
rect 59208 2128 59528 237776
rect 64208 2128 64528 237776
rect 69208 2128 69528 237776
rect 74208 2128 74528 237776
rect 79208 2128 79528 237776
rect 84208 2128 84528 237776
rect 89208 2128 89528 237776
rect 94208 2128 94528 237776
rect 99208 2128 99528 237776
rect 104208 2128 104528 237776
rect 109208 2128 109528 237776
rect 114208 2128 114528 237776
rect 119208 2128 119528 237776
rect 124208 2128 124528 237776
rect 129208 2128 129528 237776
rect 134208 2128 134528 237776
rect 139208 2128 139528 237776
rect 144208 2128 144528 237776
rect 149208 2128 149528 237776
rect 154208 2128 154528 237776
rect 159208 2128 159528 237776
rect 164208 2128 164528 237776
rect 169208 2128 169528 237776
rect 174208 2128 174528 237776
rect 179208 2128 179528 237776
rect 184208 2128 184528 237776
rect 189208 2128 189528 237776
rect 194208 2128 194528 237776
rect 199208 2128 199528 237776
rect 204208 2128 204528 237776
rect 209208 2128 209528 237776
rect 214208 2128 214528 237776
rect 219208 2128 219528 237776
rect 224208 2128 224528 237776
rect 229208 2128 229528 237776
rect 234208 2128 234528 237776
<< obsm4 >>
rect 23059 3299 24128 235381
rect 24608 3299 29128 235381
rect 29608 3299 34128 235381
rect 34608 3299 39128 235381
rect 39608 3299 44128 235381
rect 44608 3299 49128 235381
rect 49608 3299 54128 235381
rect 54608 3299 59128 235381
rect 59608 3299 64128 235381
rect 64608 3299 69128 235381
rect 69608 3299 74128 235381
rect 74608 3299 79128 235381
rect 79608 3299 84128 235381
rect 84608 3299 89128 235381
rect 89608 3299 94128 235381
rect 94608 3299 99128 235381
rect 99608 3299 104128 235381
rect 104608 3299 109128 235381
rect 109608 3299 114128 235381
rect 114608 3299 119128 235381
rect 119608 3299 124128 235381
rect 124608 3299 129128 235381
rect 129608 3299 134128 235381
rect 134608 3299 139128 235381
rect 139608 3299 144128 235381
rect 144608 3299 149128 235381
rect 149608 3299 154128 235381
rect 154608 3299 159128 235381
rect 159608 3299 164128 235381
rect 164608 3299 169128 235381
rect 169608 3299 174128 235381
rect 174608 3299 179128 235381
rect 179608 3299 184128 235381
rect 184608 3299 189128 235381
rect 189608 3299 194128 235381
rect 194608 3299 199128 235381
rect 199608 3299 203813 235381
<< labels >>
rlabel metal3 s 0 688 800 808 6 alert_major_o
port 1 nsew signal output
rlabel metal3 s 239200 688 240000 808 6 alert_minor_o
port 2 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 boot_addr_i[0]
port 3 nsew signal input
rlabel metal3 s 239200 80656 240000 80776 6 boot_addr_i[10]
port 4 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 boot_addr_i[11]
port 5 nsew signal input
rlabel metal3 s 239200 90856 240000 90976 6 boot_addr_i[12]
port 6 nsew signal input
rlabel metal2 s 82818 239200 82874 240000 6 boot_addr_i[13]
port 7 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 boot_addr_i[14]
port 8 nsew signal input
rlabel metal2 s 92294 239200 92350 240000 6 boot_addr_i[15]
port 9 nsew signal input
rlabel metal3 s 0 124720 800 124840 6 boot_addr_i[16]
port 10 nsew signal input
rlabel metal3 s 0 129480 800 129600 6 boot_addr_i[17]
port 11 nsew signal input
rlabel metal3 s 239200 121320 240000 121440 6 boot_addr_i[18]
port 12 nsew signal input
rlabel metal3 s 239200 127168 240000 127288 6 boot_addr_i[19]
port 13 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 boot_addr_i[1]
port 14 nsew signal input
rlabel metal3 s 239200 134512 240000 134632 6 boot_addr_i[20]
port 15 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 boot_addr_i[21]
port 16 nsew signal input
rlabel metal3 s 0 150424 800 150544 6 boot_addr_i[22]
port 17 nsew signal input
rlabel metal3 s 239200 150424 240000 150544 6 boot_addr_i[23]
port 18 nsew signal input
rlabel metal3 s 0 164976 800 165096 6 boot_addr_i[24]
port 19 nsew signal input
rlabel metal3 s 0 174632 800 174752 6 boot_addr_i[25]
port 20 nsew signal input
rlabel metal2 s 155222 239200 155278 240000 6 boot_addr_i[26]
port 21 nsew signal input
rlabel metal3 s 0 182656 800 182776 6 boot_addr_i[27]
port 22 nsew signal input
rlabel metal2 s 168562 239200 168618 240000 6 boot_addr_i[28]
port 23 nsew signal input
rlabel metal2 s 187514 0 187570 800 6 boot_addr_i[29]
port 24 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 boot_addr_i[2]
port 25 nsew signal input
rlabel metal3 s 0 193944 800 194064 6 boot_addr_i[30]
port 26 nsew signal input
rlabel metal3 s 239200 195576 240000 195696 6 boot_addr_i[31]
port 27 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 boot_addr_i[3]
port 28 nsew signal input
rlabel metal2 s 33322 239200 33378 240000 6 boot_addr_i[4]
port 29 nsew signal input
rlabel metal2 s 42798 239200 42854 240000 6 boot_addr_i[5]
port 30 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 boot_addr_i[6]
port 31 nsew signal input
rlabel metal3 s 239200 64608 240000 64728 6 boot_addr_i[7]
port 32 nsew signal input
rlabel metal3 s 239200 73312 240000 73432 6 boot_addr_i[8]
port 33 nsew signal input
rlabel metal2 s 50434 239200 50490 240000 6 boot_addr_i[9]
port 34 nsew signal input
rlabel metal3 s 239200 2048 240000 2168 6 clk_i
port 35 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 core_sleep_o
port 36 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 crash_dump_o[0]
port 37 nsew signal output
rlabel metal3 s 0 229440 800 229560 6 crash_dump_o[100]
port 38 nsew signal output
rlabel metal3 s 239200 226176 240000 226296 6 crash_dump_o[101]
port 39 nsew signal output
rlabel metal3 s 0 230936 800 231056 6 crash_dump_o[102]
port 40 nsew signal output
rlabel metal2 s 230846 0 230902 800 6 crash_dump_o[103]
port 41 nsew signal output
rlabel metal3 s 0 232568 800 232688 6 crash_dump_o[104]
port 42 nsew signal output
rlabel metal2 s 232502 0 232558 800 6 crash_dump_o[105]
port 43 nsew signal output
rlabel metal3 s 0 234200 800 234320 6 crash_dump_o[106]
port 44 nsew signal output
rlabel metal3 s 239200 227536 240000 227656 6 crash_dump_o[107]
port 45 nsew signal output
rlabel metal3 s 0 235832 800 235952 6 crash_dump_o[108]
port 46 nsew signal output
rlabel metal3 s 239200 229032 240000 229152 6 crash_dump_o[109]
port 47 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 crash_dump_o[10]
port 48 nsew signal output
rlabel metal3 s 239200 230528 240000 230648 6 crash_dump_o[110]
port 49 nsew signal output
rlabel metal3 s 239200 231888 240000 232008 6 crash_dump_o[111]
port 50 nsew signal output
rlabel metal3 s 239200 233384 240000 233504 6 crash_dump_o[112]
port 51 nsew signal output
rlabel metal2 s 234158 0 234214 800 6 crash_dump_o[113]
port 52 nsew signal output
rlabel metal2 s 235814 0 235870 800 6 crash_dump_o[114]
port 53 nsew signal output
rlabel metal3 s 239200 234880 240000 235000 6 crash_dump_o[115]
port 54 nsew signal output
rlabel metal3 s 239200 236240 240000 236360 6 crash_dump_o[116]
port 55 nsew signal output
rlabel metal3 s 0 237464 800 237584 6 crash_dump_o[117]
port 56 nsew signal output
rlabel metal2 s 231398 239200 231454 240000 6 crash_dump_o[118]
port 57 nsew signal output
rlabel metal2 s 237470 0 237526 800 6 crash_dump_o[119]
port 58 nsew signal output
rlabel metal3 s 239200 86504 240000 86624 6 crash_dump_o[11]
port 59 nsew signal output
rlabel metal3 s 239200 237736 240000 237856 6 crash_dump_o[120]
port 60 nsew signal output
rlabel metal2 s 233330 239200 233386 240000 6 crash_dump_o[121]
port 61 nsew signal output
rlabel metal2 s 235170 239200 235226 240000 6 crash_dump_o[122]
port 62 nsew signal output
rlabel metal3 s 239200 239232 240000 239352 6 crash_dump_o[123]
port 63 nsew signal output
rlabel metal2 s 237102 239200 237158 240000 6 crash_dump_o[124]
port 64 nsew signal output
rlabel metal2 s 239126 0 239182 800 6 crash_dump_o[125]
port 65 nsew signal output
rlabel metal3 s 0 239096 800 239216 6 crash_dump_o[126]
port 66 nsew signal output
rlabel metal2 s 239034 239200 239090 240000 6 crash_dump_o[127]
port 67 nsew signal output
rlabel metal2 s 75182 239200 75238 240000 6 crash_dump_o[12]
port 68 nsew signal output
rlabel metal2 s 112442 0 112498 800 6 crash_dump_o[13]
port 69 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 crash_dump_o[14]
port 70 nsew signal output
rlabel metal3 s 239200 105408 240000 105528 6 crash_dump_o[15]
port 71 nsew signal output
rlabel metal2 s 96158 239200 96214 240000 6 crash_dump_o[16]
port 72 nsew signal output
rlabel metal3 s 0 131112 800 131232 6 crash_dump_o[17]
port 73 nsew signal output
rlabel metal3 s 0 137504 800 137624 6 crash_dump_o[18]
port 74 nsew signal output
rlabel metal3 s 239200 128664 240000 128784 6 crash_dump_o[19]
port 75 nsew signal output
rlabel metal2 s 14186 239200 14242 240000 6 crash_dump_o[1]
port 76 nsew signal output
rlabel metal3 s 239200 135872 240000 135992 6 crash_dump_o[20]
port 77 nsew signal output
rlabel metal2 s 124678 239200 124734 240000 6 crash_dump_o[21]
port 78 nsew signal output
rlabel metal2 s 130474 239200 130530 240000 6 crash_dump_o[22]
port 79 nsew signal output
rlabel metal2 s 138018 239200 138074 240000 6 crash_dump_o[23]
port 80 nsew signal output
rlabel metal2 s 143722 239200 143778 240000 6 crash_dump_o[24]
port 81 nsew signal output
rlabel metal2 s 149518 239200 149574 240000 6 crash_dump_o[25]
port 82 nsew signal output
rlabel metal2 s 157062 239200 157118 240000 6 crash_dump_o[26]
port 83 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 crash_dump_o[27]
port 84 nsew signal output
rlabel metal2 s 170402 239200 170458 240000 6 crash_dump_o[28]
port 85 nsew signal output
rlabel metal3 s 239200 185376 240000 185496 6 crash_dump_o[29]
port 86 nsew signal output
rlabel metal3 s 239200 22448 240000 22568 6 crash_dump_o[2]
port 87 nsew signal output
rlabel metal3 s 239200 189728 240000 189848 6 crash_dump_o[30]
port 88 nsew signal output
rlabel metal3 s 0 198840 800 198960 6 crash_dump_o[31]
port 89 nsew signal output
rlabel metal3 s 0 205232 800 205352 6 crash_dump_o[32]
port 90 nsew signal output
rlabel metal3 s 239200 201424 240000 201544 6 crash_dump_o[33]
port 91 nsew signal output
rlabel metal2 s 205822 0 205878 800 6 crash_dump_o[34]
port 92 nsew signal output
rlabel metal2 s 191378 239200 191434 240000 6 crash_dump_o[35]
port 93 nsew signal output
rlabel metal3 s 239200 202784 240000 202904 6 crash_dump_o[36]
port 94 nsew signal output
rlabel metal2 s 193310 239200 193366 240000 6 crash_dump_o[37]
port 95 nsew signal output
rlabel metal2 s 195242 239200 195298 240000 6 crash_dump_o[38]
port 96 nsew signal output
rlabel metal3 s 0 206864 800 206984 6 crash_dump_o[39]
port 97 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 crash_dump_o[3]
port 98 nsew signal output
rlabel metal3 s 239200 204280 240000 204400 6 crash_dump_o[40]
port 99 nsew signal output
rlabel metal2 s 207478 0 207534 800 6 crash_dump_o[41]
port 100 nsew signal output
rlabel metal2 s 197082 239200 197138 240000 6 crash_dump_o[42]
port 101 nsew signal output
rlabel metal3 s 239200 205776 240000 205896 6 crash_dump_o[43]
port 102 nsew signal output
rlabel metal3 s 0 208496 800 208616 6 crash_dump_o[44]
port 103 nsew signal output
rlabel metal2 s 199014 239200 199070 240000 6 crash_dump_o[45]
port 104 nsew signal output
rlabel metal2 s 209134 0 209190 800 6 crash_dump_o[46]
port 105 nsew signal output
rlabel metal2 s 210790 0 210846 800 6 crash_dump_o[47]
port 106 nsew signal output
rlabel metal2 s 200946 239200 201002 240000 6 crash_dump_o[48]
port 107 nsew signal output
rlabel metal3 s 0 209992 800 210112 6 crash_dump_o[49]
port 108 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 crash_dump_o[4]
port 109 nsew signal output
rlabel metal2 s 202786 239200 202842 240000 6 crash_dump_o[50]
port 110 nsew signal output
rlabel metal2 s 204718 239200 204774 240000 6 crash_dump_o[51]
port 111 nsew signal output
rlabel metal3 s 0 211624 800 211744 6 crash_dump_o[52]
port 112 nsew signal output
rlabel metal2 s 206650 239200 206706 240000 6 crash_dump_o[53]
port 113 nsew signal output
rlabel metal2 s 212446 0 212502 800 6 crash_dump_o[54]
port 114 nsew signal output
rlabel metal3 s 0 213256 800 213376 6 crash_dump_o[55]
port 115 nsew signal output
rlabel metal3 s 239200 207136 240000 207256 6 crash_dump_o[56]
port 116 nsew signal output
rlabel metal2 s 208490 239200 208546 240000 6 crash_dump_o[57]
port 117 nsew signal output
rlabel metal3 s 0 214888 800 215008 6 crash_dump_o[58]
port 118 nsew signal output
rlabel metal2 s 210422 239200 210478 240000 6 crash_dump_o[59]
port 119 nsew signal output
rlabel metal3 s 239200 44208 240000 44328 6 crash_dump_o[5]
port 120 nsew signal output
rlabel metal3 s 239200 208632 240000 208752 6 crash_dump_o[60]
port 121 nsew signal output
rlabel metal2 s 212354 239200 212410 240000 6 crash_dump_o[61]
port 122 nsew signal output
rlabel metal2 s 214194 0 214250 800 6 crash_dump_o[62]
port 123 nsew signal output
rlabel metal3 s 0 216520 800 216640 6 crash_dump_o[63]
port 124 nsew signal output
rlabel metal3 s 0 218152 800 218272 6 crash_dump_o[64]
port 125 nsew signal output
rlabel metal2 s 215850 0 215906 800 6 crash_dump_o[65]
port 126 nsew signal output
rlabel metal3 s 239200 210128 240000 210248 6 crash_dump_o[66]
port 127 nsew signal output
rlabel metal2 s 214286 239200 214342 240000 6 crash_dump_o[67]
port 128 nsew signal output
rlabel metal2 s 216126 239200 216182 240000 6 crash_dump_o[68]
port 129 nsew signal output
rlabel metal2 s 218058 239200 218114 240000 6 crash_dump_o[69]
port 130 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 crash_dump_o[6]
port 131 nsew signal output
rlabel metal3 s 0 219784 800 219904 6 crash_dump_o[70]
port 132 nsew signal output
rlabel metal3 s 0 221280 800 221400 6 crash_dump_o[71]
port 133 nsew signal output
rlabel metal2 s 217506 0 217562 800 6 crash_dump_o[72]
port 134 nsew signal output
rlabel metal3 s 0 222912 800 223032 6 crash_dump_o[73]
port 135 nsew signal output
rlabel metal2 s 219990 239200 220046 240000 6 crash_dump_o[74]
port 136 nsew signal output
rlabel metal3 s 239200 211624 240000 211744 6 crash_dump_o[75]
port 137 nsew signal output
rlabel metal3 s 239200 212984 240000 213104 6 crash_dump_o[76]
port 138 nsew signal output
rlabel metal3 s 239200 214480 240000 214600 6 crash_dump_o[77]
port 139 nsew signal output
rlabel metal2 s 221830 239200 221886 240000 6 crash_dump_o[78]
port 140 nsew signal output
rlabel metal2 s 219162 0 219218 800 6 crash_dump_o[79]
port 141 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 crash_dump_o[7]
port 142 nsew signal output
rlabel metal3 s 239200 215976 240000 216096 6 crash_dump_o[80]
port 143 nsew signal output
rlabel metal2 s 223762 239200 223818 240000 6 crash_dump_o[81]
port 144 nsew signal output
rlabel metal2 s 220818 0 220874 800 6 crash_dump_o[82]
port 145 nsew signal output
rlabel metal3 s 239200 217336 240000 217456 6 crash_dump_o[83]
port 146 nsew signal output
rlabel metal3 s 239200 218832 240000 218952 6 crash_dump_o[84]
port 147 nsew signal output
rlabel metal2 s 225694 239200 225750 240000 6 crash_dump_o[85]
port 148 nsew signal output
rlabel metal3 s 0 224544 800 224664 6 crash_dump_o[86]
port 149 nsew signal output
rlabel metal2 s 222474 0 222530 800 6 crash_dump_o[87]
port 150 nsew signal output
rlabel metal3 s 0 226176 800 226296 6 crash_dump_o[88]
port 151 nsew signal output
rlabel metal2 s 224130 0 224186 800 6 crash_dump_o[89]
port 152 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 crash_dump_o[8]
port 153 nsew signal output
rlabel metal3 s 239200 220328 240000 220448 6 crash_dump_o[90]
port 154 nsew signal output
rlabel metal3 s 239200 221688 240000 221808 6 crash_dump_o[91]
port 155 nsew signal output
rlabel metal3 s 239200 223184 240000 223304 6 crash_dump_o[92]
port 156 nsew signal output
rlabel metal2 s 227626 239200 227682 240000 6 crash_dump_o[93]
port 157 nsew signal output
rlabel metal2 s 225786 0 225842 800 6 crash_dump_o[94]
port 158 nsew signal output
rlabel metal3 s 239200 224680 240000 224800 6 crash_dump_o[95]
port 159 nsew signal output
rlabel metal2 s 229466 239200 229522 240000 6 crash_dump_o[96]
port 160 nsew signal output
rlabel metal3 s 0 227808 800 227928 6 crash_dump_o[97]
port 161 nsew signal output
rlabel metal2 s 227534 0 227590 800 6 crash_dump_o[98]
port 162 nsew signal output
rlabel metal2 s 229190 0 229246 800 6 crash_dump_o[99]
port 163 nsew signal output
rlabel metal3 s 239200 79160 240000 79280 6 crash_dump_o[9]
port 164 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 data_addr_o[0]
port 165 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 data_addr_o[10]
port 166 nsew signal output
rlabel metal3 s 0 98880 800 99000 6 data_addr_o[11]
port 167 nsew signal output
rlabel metal3 s 239200 92216 240000 92336 6 data_addr_o[12]
port 168 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 data_addr_o[13]
port 169 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 data_addr_o[14]
port 170 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 data_addr_o[15]
port 171 nsew signal output
rlabel metal2 s 98090 239200 98146 240000 6 data_addr_o[16]
port 172 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 data_addr_o[17]
port 173 nsew signal output
rlabel metal2 s 105634 239200 105690 240000 6 data_addr_o[18]
port 174 nsew signal output
rlabel metal2 s 142526 0 142582 800 6 data_addr_o[19]
port 175 nsew signal output
rlabel metal2 s 16118 239200 16174 240000 6 data_addr_o[1]
port 176 nsew signal output
rlabel metal2 s 117134 239200 117190 240000 6 data_addr_o[20]
port 177 nsew signal output
rlabel metal3 s 239200 141720 240000 141840 6 data_addr_o[21]
port 178 nsew signal output
rlabel metal2 s 160834 0 160890 800 6 data_addr_o[22]
port 179 nsew signal output
rlabel metal2 s 139950 239200 140006 240000 6 data_addr_o[23]
port 180 nsew signal output
rlabel metal2 s 145654 239200 145710 240000 6 data_addr_o[24]
port 181 nsew signal output
rlabel metal3 s 239200 162120 240000 162240 6 data_addr_o[25]
port 182 nsew signal output
rlabel metal3 s 239200 167968 240000 168088 6 data_addr_o[26]
port 183 nsew signal output
rlabel metal2 s 162858 239200 162914 240000 6 data_addr_o[27]
port 184 nsew signal output
rlabel metal2 s 182454 0 182510 800 6 data_addr_o[28]
port 185 nsew signal output
rlabel metal3 s 0 190680 800 190800 6 data_addr_o[29]
port 186 nsew signal output
rlabel metal2 s 19982 239200 20038 240000 6 data_addr_o[2]
port 187 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 data_addr_o[30]
port 188 nsew signal output
rlabel metal2 s 183742 239200 183798 240000 6 data_addr_o[31]
port 189 nsew signal output
rlabel metal3 s 239200 35504 240000 35624 6 data_addr_o[3]
port 190 nsew signal output
rlabel metal3 s 239200 39856 240000 39976 6 data_addr_o[4]
port 191 nsew signal output
rlabel metal3 s 239200 45704 240000 45824 6 data_addr_o[5]
port 192 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 data_addr_o[6]
port 193 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 data_addr_o[7]
port 194 nsew signal output
rlabel metal3 s 239200 74808 240000 74928 6 data_addr_o[8]
port 195 nsew signal output
rlabel metal2 s 94134 0 94190 800 6 data_addr_o[9]
port 196 nsew signal output
rlabel metal3 s 239200 9392 240000 9512 6 data_be_o[0]
port 197 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 data_be_o[1]
port 198 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 data_be_o[2]
port 199 nsew signal output
rlabel metal3 s 239200 37000 240000 37120 6 data_be_o[3]
port 200 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 data_err_i
port 201 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 data_gnt_i
port 202 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 data_rdata_i[0]
port 203 nsew signal input
rlabel metal3 s 239200 82152 240000 82272 6 data_rdata_i[10]
port 204 nsew signal input
rlabel metal3 s 239200 87864 240000 87984 6 data_rdata_i[11]
port 205 nsew signal input
rlabel metal3 s 239200 93712 240000 93832 6 data_rdata_i[12]
port 206 nsew signal input
rlabel metal2 s 84750 239200 84806 240000 6 data_rdata_i[13]
port 207 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 data_rdata_i[14]
port 208 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 data_rdata_i[15]
port 209 nsew signal input
rlabel metal2 s 99930 239200 99986 240000 6 data_rdata_i[16]
port 210 nsew signal input
rlabel metal3 s 239200 114112 240000 114232 6 data_rdata_i[17]
port 211 nsew signal input
rlabel metal3 s 0 139136 800 139256 6 data_rdata_i[18]
port 212 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 data_rdata_i[19]
port 213 nsew signal input
rlabel metal2 s 18050 239200 18106 240000 6 data_rdata_i[1]
port 214 nsew signal input
rlabel metal3 s 239200 137368 240000 137488 6 data_rdata_i[20]
port 215 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 data_rdata_i[21]
port 216 nsew signal input
rlabel metal3 s 0 152056 800 152176 6 data_rdata_i[22]
port 217 nsew signal input
rlabel metal3 s 0 156952 800 157072 6 data_rdata_i[23]
port 218 nsew signal input
rlabel metal3 s 239200 157768 240000 157888 6 data_rdata_i[24]
port 219 nsew signal input
rlabel metal2 s 151358 239200 151414 240000 6 data_rdata_i[25]
port 220 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 data_rdata_i[26]
port 221 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 data_rdata_i[27]
port 222 nsew signal input
rlabel metal3 s 239200 181024 240000 181144 6 data_rdata_i[28]
port 223 nsew signal input
rlabel metal3 s 239200 186872 240000 186992 6 data_rdata_i[29]
port 224 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 data_rdata_i[2]
port 225 nsew signal input
rlabel metal3 s 0 195576 800 195696 6 data_rdata_i[30]
port 226 nsew signal input
rlabel metal2 s 204166 0 204222 800 6 data_rdata_i[31]
port 227 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 data_rdata_i[3]
port 228 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 data_rdata_i[4]
port 229 nsew signal input
rlabel metal3 s 0 60256 800 60376 6 data_rdata_i[5]
port 230 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 data_rdata_i[6]
port 231 nsew signal input
rlabel metal3 s 239200 66104 240000 66224 6 data_rdata_i[7]
port 232 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 data_rdata_i[8]
port 233 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 data_rdata_i[9]
port 234 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 data_rdata_intg_i[0]
port 235 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 data_rdata_intg_i[1]
port 236 nsew signal input
rlabel metal2 s 21822 239200 21878 240000 6 data_rdata_intg_i[2]
port 237 nsew signal input
rlabel metal2 s 25686 239200 25742 240000 6 data_rdata_intg_i[3]
port 238 nsew signal input
rlabel metal3 s 239200 41352 240000 41472 6 data_rdata_intg_i[4]
port 239 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 data_rdata_intg_i[5]
port 240 nsew signal input
rlabel metal3 s 239200 53048 240000 53168 6 data_rdata_intg_i[6]
port 241 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 data_req_o
port 242 nsew signal output
rlabel metal2 s 938 239200 994 240000 6 data_rvalid_i
port 243 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 data_wdata_intg_o[0]
port 244 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 data_wdata_intg_o[1]
port 245 nsew signal output
rlabel metal3 s 239200 23944 240000 24064 6 data_wdata_intg_o[2]
port 246 nsew signal output
rlabel metal2 s 27526 239200 27582 240000 6 data_wdata_intg_o[3]
port 247 nsew signal output
rlabel metal2 s 35162 239200 35218 240000 6 data_wdata_intg_o[4]
port 248 nsew signal output
rlabel metal3 s 239200 47200 240000 47320 6 data_wdata_intg_o[5]
port 249 nsew signal output
rlabel metal3 s 239200 54408 240000 54528 6 data_wdata_intg_o[6]
port 250 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 data_wdata_o[0]
port 251 nsew signal output
rlabel metal3 s 0 94120 800 94240 6 data_wdata_o[10]
port 252 nsew signal output
rlabel metal2 s 65706 239200 65762 240000 6 data_wdata_o[11]
port 253 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 data_wdata_o[12]
port 254 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 data_wdata_o[13]
port 255 nsew signal output
rlabel metal2 s 88522 239200 88578 240000 6 data_wdata_o[14]
port 256 nsew signal output
rlabel metal3 s 239200 106768 240000 106888 6 data_wdata_o[15]
port 257 nsew signal output
rlabel metal3 s 0 126216 800 126336 6 data_wdata_o[16]
port 258 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 data_wdata_o[17]
port 259 nsew signal output
rlabel metal3 s 239200 122816 240000 122936 6 data_wdata_o[18]
port 260 nsew signal output
rlabel metal2 s 113270 239200 113326 240000 6 data_wdata_o[19]
port 261 nsew signal output
rlabel metal3 s 239200 13744 240000 13864 6 data_wdata_o[1]
port 262 nsew signal output
rlabel metal2 s 118974 239200 119030 240000 6 data_wdata_o[20]
port 263 nsew signal output
rlabel metal2 s 155774 0 155830 800 6 data_wdata_o[21]
port 264 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 data_wdata_o[22]
port 265 nsew signal output
rlabel metal3 s 239200 151920 240000 152040 6 data_wdata_o[23]
port 266 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 data_wdata_o[24]
port 267 nsew signal output
rlabel metal3 s 239200 163616 240000 163736 6 data_wdata_o[25]
port 268 nsew signal output
rlabel metal3 s 0 179392 800 179512 6 data_wdata_o[26]
port 269 nsew signal output
rlabel metal3 s 0 184288 800 184408 6 data_wdata_o[27]
port 270 nsew signal output
rlabel metal2 s 172334 239200 172390 240000 6 data_wdata_o[28]
port 271 nsew signal output
rlabel metal2 s 176106 239200 176162 240000 6 data_wdata_o[29]
port 272 nsew signal output
rlabel metal3 s 239200 25304 240000 25424 6 data_wdata_o[2]
port 273 nsew signal output
rlabel metal2 s 197450 0 197506 800 6 data_wdata_o[30]
port 274 nsew signal output
rlabel metal3 s 239200 197072 240000 197192 6 data_wdata_o[31]
port 275 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 data_wdata_o[3]
port 276 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 data_wdata_o[4]
port 277 nsew signal output
rlabel metal2 s 44730 239200 44786 240000 6 data_wdata_o[5]
port 278 nsew signal output
rlabel metal3 s 239200 55904 240000 56024 6 data_wdata_o[6]
port 279 nsew signal output
rlabel metal3 s 239200 67600 240000 67720 6 data_wdata_o[7]
port 280 nsew signal output
rlabel metal2 s 87510 0 87566 800 6 data_wdata_o[8]
port 281 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 data_wdata_o[9]
port 282 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 data_we_o
port 283 nsew signal output
rlabel metal2 s 2778 239200 2834 240000 6 debug_req_i
port 284 nsew signal input
rlabel metal2 s 10414 239200 10470 240000 6 eFPGA_delay_o[0]
port 285 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 eFPGA_delay_o[1]
port 286 nsew signal output
rlabel metal3 s 239200 26800 240000 26920 6 eFPGA_delay_o[2]
port 287 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 eFPGA_delay_o[3]
port 288 nsew signal output
rlabel metal3 s 239200 3544 240000 3664 6 eFPGA_en_o
port 289 nsew signal output
rlabel metal2 s 4710 239200 4766 240000 6 eFPGA_fpga_done_i
port 290 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 eFPGA_operand_a_o[0]
port 291 nsew signal output
rlabel metal3 s 239200 83512 240000 83632 6 eFPGA_operand_a_o[10]
port 292 nsew signal output
rlabel metal2 s 67546 239200 67602 240000 6 eFPGA_operand_a_o[11]
port 293 nsew signal output
rlabel metal3 s 239200 95208 240000 95328 6 eFPGA_operand_a_o[12]
port 294 nsew signal output
rlabel metal3 s 0 105272 800 105392 6 eFPGA_operand_a_o[13]
port 295 nsew signal output
rlabel metal3 s 0 113432 800 113552 6 eFPGA_operand_a_o[14]
port 296 nsew signal output
rlabel metal3 s 0 118192 800 118312 6 eFPGA_operand_a_o[15]
port 297 nsew signal output
rlabel metal2 s 101862 239200 101918 240000 6 eFPGA_operand_a_o[16]
port 298 nsew signal output
rlabel metal3 s 239200 115608 240000 115728 6 eFPGA_operand_a_o[17]
port 299 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 eFPGA_operand_a_o[18]
port 300 nsew signal output
rlabel metal3 s 239200 130160 240000 130280 6 eFPGA_operand_a_o[19]
port 301 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 eFPGA_operand_a_o[1]
port 302 nsew signal output
rlabel metal3 s 239200 138864 240000 138984 6 eFPGA_operand_a_o[20]
port 303 nsew signal output
rlabel metal2 s 157522 0 157578 800 6 eFPGA_operand_a_o[21]
port 304 nsew signal output
rlabel metal2 s 132314 239200 132370 240000 6 eFPGA_operand_a_o[22]
port 305 nsew signal output
rlabel metal3 s 239200 153416 240000 153536 6 eFPGA_operand_a_o[23]
port 306 nsew signal output
rlabel metal3 s 0 166608 800 166728 6 eFPGA_operand_a_o[24]
port 307 nsew signal output
rlabel metal3 s 0 176264 800 176384 6 eFPGA_operand_a_o[25]
port 308 nsew signal output
rlabel metal3 s 239200 169328 240000 169448 6 eFPGA_operand_a_o[26]
port 309 nsew signal output
rlabel metal3 s 239200 175176 240000 175296 6 eFPGA_operand_a_o[27]
port 310 nsew signal output
rlabel metal3 s 0 185920 800 186040 6 eFPGA_operand_a_o[28]
port 311 nsew signal output
rlabel metal2 s 178038 239200 178094 240000 6 eFPGA_operand_a_o[29]
port 312 nsew signal output
rlabel metal3 s 239200 28296 240000 28416 6 eFPGA_operand_a_o[2]
port 313 nsew signal output
rlabel metal2 s 181902 239200 181958 240000 6 eFPGA_operand_a_o[30]
port 314 nsew signal output
rlabel metal3 s 239200 198432 240000 198552 6 eFPGA_operand_a_o[31]
port 315 nsew signal output
rlabel metal2 s 29458 239200 29514 240000 6 eFPGA_operand_a_o[3]
port 316 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 eFPGA_operand_a_o[4]
port 317 nsew signal output
rlabel metal3 s 239200 48696 240000 48816 6 eFPGA_operand_a_o[5]
port 318 nsew signal output
rlabel metal3 s 239200 57400 240000 57520 6 eFPGA_operand_a_o[6]
port 319 nsew signal output
rlabel metal3 s 0 73176 800 73296 6 eFPGA_operand_a_o[7]
port 320 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 eFPGA_operand_a_o[8]
port 321 nsew signal output
rlabel metal2 s 52366 239200 52422 240000 6 eFPGA_operand_a_o[9]
port 322 nsew signal output
rlabel metal3 s 239200 10752 240000 10872 6 eFPGA_operand_b_o[0]
port 323 nsew signal output
rlabel metal3 s 0 95616 800 95736 6 eFPGA_operand_b_o[10]
port 324 nsew signal output
rlabel metal3 s 0 100512 800 100632 6 eFPGA_operand_b_o[11]
port 325 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 eFPGA_operand_b_o[12]
port 326 nsew signal output
rlabel metal3 s 239200 96704 240000 96824 6 eFPGA_operand_b_o[13]
port 327 nsew signal output
rlabel metal3 s 239200 101056 240000 101176 6 eFPGA_operand_b_o[14]
port 328 nsew signal output
rlabel metal3 s 0 119824 800 119944 6 eFPGA_operand_b_o[15]
port 329 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 eFPGA_operand_b_o[16]
port 330 nsew signal output
rlabel metal3 s 239200 116968 240000 117088 6 eFPGA_operand_b_o[17]
port 331 nsew signal output
rlabel metal3 s 239200 124312 240000 124432 6 eFPGA_operand_b_o[18]
port 332 nsew signal output
rlabel metal3 s 0 142400 800 142520 6 eFPGA_operand_b_o[19]
port 333 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 eFPGA_operand_b_o[1]
port 334 nsew signal output
rlabel metal3 s 0 145664 800 145784 6 eFPGA_operand_b_o[20]
port 335 nsew signal output
rlabel metal3 s 0 148792 800 148912 6 eFPGA_operand_b_o[21]
port 336 nsew signal output
rlabel metal3 s 0 155320 800 155440 6 eFPGA_operand_b_o[22]
port 337 nsew signal output
rlabel metal3 s 0 158448 800 158568 6 eFPGA_operand_b_o[23]
port 338 nsew signal output
rlabel metal3 s 0 168104 800 168224 6 eFPGA_operand_b_o[24]
port 339 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 eFPGA_operand_b_o[25]
port 340 nsew signal output
rlabel metal3 s 239200 170824 240000 170944 6 eFPGA_operand_b_o[26]
port 341 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 eFPGA_operand_b_o[27]
port 342 nsew signal output
rlabel metal2 s 184110 0 184166 800 6 eFPGA_operand_b_o[28]
port 343 nsew signal output
rlabel metal2 s 189170 0 189226 800 6 eFPGA_operand_b_o[29]
port 344 nsew signal output
rlabel metal3 s 239200 29656 240000 29776 6 eFPGA_operand_b_o[2]
port 345 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 eFPGA_operand_b_o[30]
port 346 nsew signal output
rlabel metal3 s 0 200336 800 200456 6 eFPGA_operand_b_o[31]
port 347 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 eFPGA_operand_b_o[3]
port 348 nsew signal output
rlabel metal2 s 37094 239200 37150 240000 6 eFPGA_operand_b_o[4]
port 349 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 eFPGA_operand_b_o[5]
port 350 nsew signal output
rlabel metal3 s 239200 58760 240000 58880 6 eFPGA_operand_b_o[6]
port 351 nsew signal output
rlabel metal3 s 239200 68960 240000 69080 6 eFPGA_operand_b_o[7]
port 352 nsew signal output
rlabel metal3 s 0 81200 800 81320 6 eFPGA_operand_b_o[8]
port 353 nsew signal output
rlabel metal2 s 54206 239200 54262 240000 6 eFPGA_operand_b_o[9]
port 354 nsew signal output
rlabel metal2 s 12346 239200 12402 240000 6 eFPGA_operator_o[0]
port 355 nsew signal output
rlabel metal3 s 239200 15104 240000 15224 6 eFPGA_operator_o[1]
port 356 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 eFPGA_result_a_i[0]
port 357 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 eFPGA_result_a_i[10]
port 358 nsew signal input
rlabel metal3 s 0 102144 800 102264 6 eFPGA_result_a_i[11]
port 359 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 eFPGA_result_a_i[12]
port 360 nsew signal input
rlabel metal3 s 239200 98064 240000 98184 6 eFPGA_result_a_i[13]
port 361 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 eFPGA_result_a_i[14]
port 362 nsew signal input
rlabel metal3 s 0 121456 800 121576 6 eFPGA_result_a_i[15]
port 363 nsew signal input
rlabel metal3 s 239200 112616 240000 112736 6 eFPGA_result_a_i[16]
port 364 nsew signal input
rlabel metal3 s 0 132744 800 132864 6 eFPGA_result_a_i[17]
port 365 nsew signal input
rlabel metal2 s 107566 239200 107622 240000 6 eFPGA_result_a_i[18]
port 366 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 eFPGA_result_a_i[19]
port 367 nsew signal input
rlabel metal3 s 239200 16600 240000 16720 6 eFPGA_result_a_i[1]
port 368 nsew signal input
rlabel metal3 s 0 147160 800 147280 6 eFPGA_result_a_i[20]
port 369 nsew signal input
rlabel metal3 s 239200 143216 240000 143336 6 eFPGA_result_a_i[21]
port 370 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 eFPGA_result_a_i[22]
port 371 nsew signal input
rlabel metal2 s 141882 239200 141938 240000 6 eFPGA_result_a_i[23]
port 372 nsew signal input
rlabel metal3 s 239200 159128 240000 159248 6 eFPGA_result_a_i[24]
port 373 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 eFPGA_result_a_i[25]
port 374 nsew signal input
rlabel metal2 s 158994 239200 159050 240000 6 eFPGA_result_a_i[26]
port 375 nsew signal input
rlabel metal3 s 239200 176672 240000 176792 6 eFPGA_result_a_i[27]
port 376 nsew signal input
rlabel metal2 s 174266 239200 174322 240000 6 eFPGA_result_a_i[28]
port 377 nsew signal input
rlabel metal3 s 239200 188232 240000 188352 6 eFPGA_result_a_i[29]
port 378 nsew signal input
rlabel metal3 s 239200 31152 240000 31272 6 eFPGA_result_a_i[2]
port 379 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 eFPGA_result_a_i[30]
port 380 nsew signal input
rlabel metal2 s 185674 239200 185730 240000 6 eFPGA_result_a_i[31]
port 381 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 eFPGA_result_a_i[3]
port 382 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 eFPGA_result_a_i[4]
port 383 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 eFPGA_result_a_i[5]
port 384 nsew signal input
rlabel metal2 s 46570 239200 46626 240000 6 eFPGA_result_a_i[6]
port 385 nsew signal input
rlabel metal3 s 0 74672 800 74792 6 eFPGA_result_a_i[7]
port 386 nsew signal input
rlabel metal3 s 239200 76304 240000 76424 6 eFPGA_result_a_i[8]
port 387 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 eFPGA_result_a_i[9]
port 388 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 eFPGA_result_b_i[0]
port 389 nsew signal input
rlabel metal2 s 58070 239200 58126 240000 6 eFPGA_result_b_i[10]
port 390 nsew signal input
rlabel metal2 s 69478 239200 69534 240000 6 eFPGA_result_b_i[11]
port 391 nsew signal input
rlabel metal2 s 77114 239200 77170 240000 6 eFPGA_result_b_i[12]
port 392 nsew signal input
rlabel metal2 s 86590 239200 86646 240000 6 eFPGA_result_b_i[13]
port 393 nsew signal input
rlabel metal2 s 90454 239200 90510 240000 6 eFPGA_result_b_i[14]
port 394 nsew signal input
rlabel metal3 s 239200 108264 240000 108384 6 eFPGA_result_b_i[15]
port 395 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 eFPGA_result_b_i[16]
port 396 nsew signal input
rlabel metal3 s 0 134376 800 134496 6 eFPGA_result_b_i[17]
port 397 nsew signal input
rlabel metal2 s 109498 239200 109554 240000 6 eFPGA_result_b_i[18]
port 398 nsew signal input
rlabel metal2 s 115202 239200 115258 240000 6 eFPGA_result_b_i[19]
port 399 nsew signal input
rlabel metal3 s 239200 18096 240000 18216 6 eFPGA_result_b_i[1]
port 400 nsew signal input
rlabel metal2 s 120906 239200 120962 240000 6 eFPGA_result_b_i[20]
port 401 nsew signal input
rlabel metal2 s 126610 239200 126666 240000 6 eFPGA_result_b_i[21]
port 402 nsew signal input
rlabel metal3 s 239200 147568 240000 147688 6 eFPGA_result_b_i[22]
port 403 nsew signal input
rlabel metal3 s 0 160080 800 160200 6 eFPGA_result_b_i[23]
port 404 nsew signal input
rlabel metal3 s 239200 160624 240000 160744 6 eFPGA_result_b_i[24]
port 405 nsew signal input
rlabel metal3 s 239200 164976 240000 165096 6 eFPGA_result_b_i[25]
port 406 nsew signal input
rlabel metal2 s 160926 239200 160982 240000 6 eFPGA_result_b_i[26]
port 407 nsew signal input
rlabel metal3 s 239200 178168 240000 178288 6 eFPGA_result_b_i[27]
port 408 nsew signal input
rlabel metal3 s 0 187552 800 187672 6 eFPGA_result_b_i[28]
port 409 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 eFPGA_result_b_i[29]
port 410 nsew signal input
rlabel metal3 s 239200 32648 240000 32768 6 eFPGA_result_b_i[2]
port 411 nsew signal input
rlabel metal3 s 0 197208 800 197328 6 eFPGA_result_b_i[30]
port 412 nsew signal input
rlabel metal2 s 187606 239200 187662 240000 6 eFPGA_result_b_i[31]
port 413 nsew signal input
rlabel metal2 s 31390 239200 31446 240000 6 eFPGA_result_b_i[3]
port 414 nsew signal input
rlabel metal2 s 39026 239200 39082 240000 6 eFPGA_result_b_i[4]
port 415 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 eFPGA_result_b_i[5]
port 416 nsew signal input
rlabel metal3 s 239200 60256 240000 60376 6 eFPGA_result_b_i[6]
port 417 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 eFPGA_result_b_i[7]
port 418 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 eFPGA_result_b_i[8]
port 419 nsew signal input
rlabel metal2 s 56138 239200 56194 240000 6 eFPGA_result_b_i[9]
port 420 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 eFPGA_result_c_i[0]
port 421 nsew signal input
rlabel metal3 s 239200 85008 240000 85128 6 eFPGA_result_c_i[10]
port 422 nsew signal input
rlabel metal3 s 0 103776 800 103896 6 eFPGA_result_c_i[11]
port 423 nsew signal input
rlabel metal2 s 78954 239200 79010 240000 6 eFPGA_result_c_i[12]
port 424 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 eFPGA_result_c_i[13]
port 425 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 eFPGA_result_c_i[14]
port 426 nsew signal input
rlabel metal3 s 239200 109760 240000 109880 6 eFPGA_result_c_i[15]
port 427 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 eFPGA_result_c_i[16]
port 428 nsew signal input
rlabel metal3 s 239200 118464 240000 118584 6 eFPGA_result_c_i[17]
port 429 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 eFPGA_result_c_i[18]
port 430 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 eFPGA_result_c_i[19]
port 431 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 eFPGA_result_c_i[1]
port 432 nsew signal input
rlabel metal3 s 239200 140224 240000 140344 6 eFPGA_result_c_i[20]
port 433 nsew signal input
rlabel metal3 s 239200 144712 240000 144832 6 eFPGA_result_c_i[21]
port 434 nsew signal input
rlabel metal2 s 134246 239200 134302 240000 6 eFPGA_result_c_i[22]
port 435 nsew signal input
rlabel metal3 s 239200 154776 240000 154896 6 eFPGA_result_c_i[23]
port 436 nsew signal input
rlabel metal3 s 0 169736 800 169856 6 eFPGA_result_c_i[24]
port 437 nsew signal input
rlabel metal3 s 0 177896 800 178016 6 eFPGA_result_c_i[25]
port 438 nsew signal input
rlabel metal3 s 239200 172320 240000 172440 6 eFPGA_result_c_i[26]
port 439 nsew signal input
rlabel metal2 s 164698 239200 164754 240000 6 eFPGA_result_c_i[27]
port 440 nsew signal input
rlabel metal3 s 239200 182520 240000 182640 6 eFPGA_result_c_i[28]
port 441 nsew signal input
rlabel metal2 s 192482 0 192538 800 6 eFPGA_result_c_i[29]
port 442 nsew signal input
rlabel metal3 s 239200 34144 240000 34264 6 eFPGA_result_c_i[2]
port 443 nsew signal input
rlabel metal3 s 239200 191224 240000 191344 6 eFPGA_result_c_i[30]
port 444 nsew signal input
rlabel metal3 s 0 201968 800 202088 6 eFPGA_result_c_i[31]
port 445 nsew signal input
rlabel metal3 s 239200 38496 240000 38616 6 eFPGA_result_c_i[3]
port 446 nsew signal input
rlabel metal3 s 239200 42848 240000 42968 6 eFPGA_result_c_i[4]
port 447 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 eFPGA_result_c_i[5]
port 448 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 eFPGA_result_c_i[6]
port 449 nsew signal input
rlabel metal3 s 239200 70456 240000 70576 6 eFPGA_result_c_i[7]
port 450 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 eFPGA_result_c_i[8]
port 451 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 eFPGA_result_c_i[9]
port 452 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 eFPGA_write_strobe_o
port 453 nsew signal output
rlabel metal2 s 6642 239200 6698 240000 6 fetch_enable_i
port 454 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 hart_id_i[0]
port 455 nsew signal input
rlabel metal2 s 59910 239200 59966 240000 6 hart_id_i[10]
port 456 nsew signal input
rlabel metal2 s 71410 239200 71466 240000 6 hart_id_i[11]
port 457 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 hart_id_i[12]
port 458 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 hart_id_i[13]
port 459 nsew signal input
rlabel metal3 s 239200 102416 240000 102536 6 hart_id_i[14]
port 460 nsew signal input
rlabel metal3 s 239200 111120 240000 111240 6 hart_id_i[15]
port 461 nsew signal input
rlabel metal2 s 103794 239200 103850 240000 6 hart_id_i[16]
port 462 nsew signal input
rlabel metal3 s 239200 119960 240000 120080 6 hart_id_i[17]
port 463 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 hart_id_i[18]
port 464 nsew signal input
rlabel metal3 s 239200 131520 240000 131640 6 hart_id_i[19]
port 465 nsew signal input
rlabel metal3 s 239200 19592 240000 19712 6 hart_id_i[1]
port 466 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 hart_id_i[20]
port 467 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 hart_id_i[21]
port 468 nsew signal input
rlabel metal3 s 239200 149064 240000 149184 6 hart_id_i[22]
port 469 nsew signal input
rlabel metal3 s 0 161712 800 161832 6 hart_id_i[23]
port 470 nsew signal input
rlabel metal3 s 0 171368 800 171488 6 hart_id_i[24]
port 471 nsew signal input
rlabel metal3 s 239200 166472 240000 166592 6 hart_id_i[25]
port 472 nsew signal input
rlabel metal3 s 239200 173680 240000 173800 6 hart_id_i[26]
port 473 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 hart_id_i[27]
port 474 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 hart_id_i[28]
port 475 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 hart_id_i[29]
port 476 nsew signal input
rlabel metal2 s 23754 239200 23810 240000 6 hart_id_i[2]
port 477 nsew signal input
rlabel metal3 s 239200 192720 240000 192840 6 hart_id_i[30]
port 478 nsew signal input
rlabel metal3 s 239200 199928 240000 200048 6 hart_id_i[31]
port 479 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 hart_id_i[3]
port 480 nsew signal input
rlabel metal2 s 40866 239200 40922 240000 6 hart_id_i[4]
port 481 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 hart_id_i[5]
port 482 nsew signal input
rlabel metal3 s 239200 61752 240000 61872 6 hart_id_i[6]
port 483 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 hart_id_i[7]
port 484 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 hart_id_i[8]
port 485 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 hart_id_i[9]
port 486 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 instr_addr_o[0]
port 487 nsew signal output
rlabel metal2 s 61842 239200 61898 240000 6 instr_addr_o[10]
port 488 nsew signal output
rlabel metal3 s 239200 89360 240000 89480 6 instr_addr_o[11]
port 489 nsew signal output
rlabel metal2 s 80886 239200 80942 240000 6 instr_addr_o[12]
port 490 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 instr_addr_o[13]
port 491 nsew signal output
rlabel metal3 s 0 116560 800 116680 6 instr_addr_o[14]
port 492 nsew signal output
rlabel metal3 s 0 123088 800 123208 6 instr_addr_o[15]
port 493 nsew signal output
rlabel metal2 s 130842 0 130898 800 6 instr_addr_o[16]
port 494 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 instr_addr_o[17]
port 495 nsew signal output
rlabel metal2 s 111338 239200 111394 240000 6 instr_addr_o[18]
port 496 nsew signal output
rlabel metal3 s 239200 133016 240000 133136 6 instr_addr_o[19]
port 497 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 instr_addr_o[1]
port 498 nsew signal output
rlabel metal2 s 150806 0 150862 800 6 instr_addr_o[20]
port 499 nsew signal output
rlabel metal2 s 128542 239200 128598 240000 6 instr_addr_o[21]
port 500 nsew signal output
rlabel metal2 s 164146 0 164202 800 6 instr_addr_o[22]
port 501 nsew signal output
rlabel metal3 s 239200 156272 240000 156392 6 instr_addr_o[23]
port 502 nsew signal output
rlabel metal3 s 0 173000 800 173120 6 instr_addr_o[24]
port 503 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 instr_addr_o[25]
port 504 nsew signal output
rlabel metal3 s 0 181024 800 181144 6 instr_addr_o[26]
port 505 nsew signal output
rlabel metal3 s 239200 179528 240000 179648 6 instr_addr_o[27]
port 506 nsew signal output
rlabel metal3 s 0 189048 800 189168 6 instr_addr_o[28]
port 507 nsew signal output
rlabel metal2 s 179970 239200 180026 240000 6 instr_addr_o[29]
port 508 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 instr_addr_o[2]
port 509 nsew signal output
rlabel metal2 s 202510 0 202566 800 6 instr_addr_o[30]
port 510 nsew signal output
rlabel metal3 s 0 203600 800 203720 6 instr_addr_o[31]
port 511 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 instr_addr_o[3]
port 512 nsew signal output
rlabel metal3 s 0 56992 800 57112 6 instr_addr_o[4]
port 513 nsew signal output
rlabel metal3 s 239200 50056 240000 50176 6 instr_addr_o[5]
port 514 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 instr_addr_o[6]
port 515 nsew signal output
rlabel metal3 s 0 77936 800 78056 6 instr_addr_o[7]
port 516 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 instr_addr_o[8]
port 517 nsew signal output
rlabel metal3 s 0 90856 800 90976 6 instr_addr_o[9]
port 518 nsew signal output
rlabel metal3 s 239200 5040 240000 5160 6 instr_err_i
port 519 nsew signal input
rlabel metal2 s 8482 239200 8538 240000 6 instr_gnt_i
port 520 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 instr_rdata_i[0]
port 521 nsew signal input
rlabel metal2 s 63774 239200 63830 240000 6 instr_rdata_i[10]
port 522 nsew signal input
rlabel metal2 s 73250 239200 73306 240000 6 instr_rdata_i[11]
port 523 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 instr_rdata_i[12]
port 524 nsew signal input
rlabel metal3 s 239200 99560 240000 99680 6 instr_rdata_i[13]
port 525 nsew signal input
rlabel metal3 s 239200 103912 240000 104032 6 instr_rdata_i[14]
port 526 nsew signal input
rlabel metal2 s 94226 239200 94282 240000 6 instr_rdata_i[15]
port 527 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 instr_rdata_i[16]
port 528 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 instr_rdata_i[17]
port 529 nsew signal input
rlabel metal3 s 239200 125672 240000 125792 6 instr_rdata_i[18]
port 530 nsew signal input
rlabel metal3 s 0 144032 800 144152 6 instr_rdata_i[19]
port 531 nsew signal input
rlabel metal3 s 239200 20952 240000 21072 6 instr_rdata_i[1]
port 532 nsew signal input
rlabel metal2 s 122838 239200 122894 240000 6 instr_rdata_i[20]
port 533 nsew signal input
rlabel metal3 s 239200 146072 240000 146192 6 instr_rdata_i[21]
port 534 nsew signal input
rlabel metal2 s 136178 239200 136234 240000 6 instr_rdata_i[22]
port 535 nsew signal input
rlabel metal3 s 0 163344 800 163464 6 instr_rdata_i[23]
port 536 nsew signal input
rlabel metal2 s 147586 239200 147642 240000 6 instr_rdata_i[24]
port 537 nsew signal input
rlabel metal2 s 153290 239200 153346 240000 6 instr_rdata_i[25]
port 538 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 instr_rdata_i[26]
port 539 nsew signal input
rlabel metal2 s 166630 239200 166686 240000 6 instr_rdata_i[27]
port 540 nsew signal input
rlabel metal3 s 239200 183880 240000 184000 6 instr_rdata_i[28]
port 541 nsew signal input
rlabel metal3 s 0 192312 800 192432 6 instr_rdata_i[29]
port 542 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 instr_rdata_i[2]
port 543 nsew signal input
rlabel metal3 s 239200 194080 240000 194200 6 instr_rdata_i[30]
port 544 nsew signal input
rlabel metal2 s 189446 239200 189502 240000 6 instr_rdata_i[31]
port 545 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 instr_rdata_i[3]
port 546 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 instr_rdata_i[4]
port 547 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 instr_rdata_i[5]
port 548 nsew signal input
rlabel metal2 s 48502 239200 48558 240000 6 instr_rdata_i[6]
port 549 nsew signal input
rlabel metal3 s 239200 71952 240000 72072 6 instr_rdata_i[7]
port 550 nsew signal input
rlabel metal3 s 239200 77664 240000 77784 6 instr_rdata_i[8]
port 551 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 instr_rdata_i[9]
port 552 nsew signal input
rlabel metal3 s 239200 12248 240000 12368 6 instr_rdata_intg_i[0]
port 553 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 instr_rdata_intg_i[1]
port 554 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 instr_rdata_intg_i[2]
port 555 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 instr_rdata_intg_i[3]
port 556 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 instr_rdata_intg_i[4]
port 557 nsew signal input
rlabel metal3 s 239200 51552 240000 51672 6 instr_rdata_intg_i[5]
port 558 nsew signal input
rlabel metal3 s 239200 63112 240000 63232 6 instr_rdata_intg_i[6]
port 559 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 instr_req_o
port 560 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 instr_rvalid_i
port 561 nsew signal input
rlabel metal2 s 846 0 902 800 6 irq_external_i
port 562 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 irq_fast_i[0]
port 563 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 irq_fast_i[10]
port 564 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 irq_fast_i[11]
port 565 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 irq_fast_i[12]
port 566 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 irq_fast_i[13]
port 567 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 irq_fast_i[14]
port 568 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 irq_fast_i[1]
port 569 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 irq_fast_i[2]
port 570 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 irq_fast_i[3]
port 571 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 irq_fast_i[4]
port 572 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 irq_fast_i[5]
port 573 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 irq_fast_i[6]
port 574 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 irq_fast_i[7]
port 575 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 irq_fast_i[8]
port 576 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 irq_fast_i[9]
port 577 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 irq_nm_i
port 578 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 irq_software_i
port 579 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 irq_timer_i
port 580 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 ram_cfg_i
port 581 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 rst_ni
port 582 nsew signal input
rlabel metal3 s 239200 6400 240000 6520 6 scan_rst_ni
port 583 nsew signal input
rlabel metal3 s 239200 7896 240000 8016 6 test_en_i
port 584 nsew signal input
rlabel metal4 s 4208 2128 4528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 14208 2128 14528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 24208 2128 24528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 34208 2128 34528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 44208 2128 44528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 54208 2128 54528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 64208 2128 64528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 74208 2128 74528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 84208 2128 84528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 94208 2128 94528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 104208 2128 104528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 114208 2128 114528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 124208 2128 124528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 134208 2128 134528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 144208 2128 144528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 154208 2128 154528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 164208 2128 164528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 174208 2128 174528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 184208 2128 184528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 194208 2128 194528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 204208 2128 204528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 214208 2128 214528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 224208 2128 224528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 234208 2128 234528 237776 6 vccd1
port 585 nsew power input
rlabel metal4 s 9208 2128 9528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 19208 2128 19528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 29208 2128 29528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 39208 2128 39528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 49208 2128 49528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 59208 2128 59528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 69208 2128 69528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 79208 2128 79528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 89208 2128 89528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 99208 2128 99528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 109208 2128 109528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 119208 2128 119528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 129208 2128 129528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 139208 2128 139528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 149208 2128 149528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 159208 2128 159528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 169208 2128 169528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 179208 2128 179528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 189208 2128 189528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 199208 2128 199528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 209208 2128 209528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 219208 2128 219528 237776 6 vssd1
port 586 nsew ground input
rlabel metal4 s 229208 2128 229528 237776 6 vssd1
port 586 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 240000 240000
string LEFview TRUE
string GDS_FILE /project/openlane/ibex_top/runs/ibex_top/results/magic/ibex_top.gds
string GDS_END 112073372
string GDS_START 721754
<< end >>

