magic
tech sky130A
magscale 1 2
timestamp 1640350729
<< locali >>
rect 26249 25823 26283 28441
rect 19073 24055 19107 24361
rect 9873 20791 9907 21097
rect 4353 20247 4387 20417
rect 21833 16031 21867 16133
rect 14749 15351 14783 15657
rect 14105 14263 14139 14501
rect 11805 12767 11839 12937
rect 20085 12291 20119 12393
rect 8493 11135 8527 11305
rect 6193 10455 6227 10557
rect 8769 9911 8803 10217
rect 13737 9027 13771 9129
rect 8769 7871 8803 8041
rect 17877 7259 17911 7429
rect 4629 6103 4663 6409
<< viali >>
rect 26249 28441 26283 28475
rect 12817 26537 12851 26571
rect 15117 26401 15151 26435
rect 11805 26333 11839 26367
rect 11897 26333 11931 26367
rect 12264 26333 12298 26367
rect 12541 26333 12575 26367
rect 14105 26333 14139 26367
rect 14289 26333 14323 26367
rect 14807 26333 14841 26367
rect 15209 26333 15243 26367
rect 15301 26333 15335 26367
rect 12725 26265 12759 26299
rect 14473 26265 14507 26299
rect 14565 26265 14599 26299
rect 15485 26265 15519 26299
rect 15669 26265 15703 26299
rect 16313 26265 16347 26299
rect 16497 26265 16531 26299
rect 16681 26265 16715 26299
rect 12357 26197 12391 26231
rect 12909 25993 12943 26027
rect 16037 25993 16071 26027
rect 7932 25857 7966 25891
rect 11069 25857 11103 25891
rect 11161 25857 11195 25891
rect 11529 25857 11563 25891
rect 11785 25857 11819 25891
rect 13093 25857 13127 25891
rect 13349 25857 13383 25891
rect 14924 25857 14958 25891
rect 16681 25857 16715 25891
rect 21833 25857 21867 25891
rect 23121 25857 23155 25891
rect 25053 25857 25087 25891
rect 7665 25789 7699 25823
rect 14657 25789 14691 25823
rect 16773 25789 16807 25823
rect 25329 25789 25363 25823
rect 26249 25789 26283 25823
rect 11345 25721 11379 25755
rect 7481 25653 7515 25687
rect 9045 25653 9079 25687
rect 10885 25653 10919 25687
rect 14473 25653 14507 25687
rect 16681 25653 16715 25687
rect 17049 25653 17083 25687
rect 13001 25449 13035 25483
rect 14381 25449 14415 25483
rect 16681 25449 16715 25483
rect 11805 25381 11839 25415
rect 8585 25313 8619 25347
rect 10425 25313 10459 25347
rect 12449 25313 12483 25347
rect 12633 25313 12667 25347
rect 13737 25313 13771 25347
rect 15301 25313 15335 25347
rect 25053 25313 25087 25347
rect 6745 25245 6779 25279
rect 7021 25245 7055 25279
rect 7481 25245 7515 25279
rect 7665 25245 7699 25279
rect 8033 25245 8067 25279
rect 8309 25245 8343 25279
rect 8953 25245 8987 25279
rect 10333 25245 10367 25279
rect 10692 25245 10726 25279
rect 12817 25245 12851 25279
rect 13427 25245 13461 25279
rect 13829 25245 13863 25279
rect 14105 25245 14139 25279
rect 15025 25245 15059 25279
rect 18337 25245 18371 25279
rect 7205 25177 7239 25211
rect 7389 25177 7423 25211
rect 7941 25177 7975 25211
rect 8125 25177 8159 25211
rect 8493 25177 8527 25211
rect 13185 25177 13219 25211
rect 14749 25177 14783 25211
rect 15546 25177 15580 25211
rect 18070 25177 18104 25211
rect 6929 25109 6963 25143
rect 10241 25109 10275 25143
rect 11989 25109 12023 25143
rect 12357 25109 12391 25143
rect 14372 25109 14406 25143
rect 14841 25109 14875 25143
rect 15209 25109 15243 25143
rect 16957 25109 16991 25143
rect 7205 24905 7239 24939
rect 8033 24905 8067 24939
rect 8585 24905 8619 24939
rect 10333 24905 10367 24939
rect 13001 24905 13035 24939
rect 13369 24905 13403 24939
rect 14657 24905 14691 24939
rect 15761 24905 15795 24939
rect 10968 24837 11002 24871
rect 11897 24837 11931 24871
rect 14289 24837 14323 24871
rect 15117 24837 15151 24871
rect 6653 24769 6687 24803
rect 6745 24769 6779 24803
rect 7113 24769 7147 24803
rect 7297 24769 7331 24803
rect 7389 24769 7423 24803
rect 7554 24769 7588 24803
rect 7662 24769 7696 24803
rect 7941 24769 7975 24803
rect 9229 24769 9263 24803
rect 10425 24769 10459 24803
rect 10701 24769 10735 24803
rect 11345 24769 11379 24803
rect 11989 24769 12023 24803
rect 12909 24769 12943 24803
rect 13553 24769 13587 24803
rect 13645 24769 13679 24803
rect 14197 24769 14231 24803
rect 15577 24769 15611 24803
rect 16095 24769 16129 24803
rect 16405 24769 16439 24803
rect 17083 24769 17117 24803
rect 7757 24701 7791 24735
rect 8677 24701 8711 24735
rect 8861 24701 8895 24735
rect 12173 24701 12207 24735
rect 12449 24701 12483 24735
rect 13185 24701 13219 24735
rect 14013 24701 14047 24735
rect 15209 24701 15243 24735
rect 15393 24701 15427 24735
rect 16497 24701 16531 24735
rect 16681 24701 16715 24735
rect 16773 24701 16807 24735
rect 8217 24633 8251 24667
rect 9045 24633 9079 24667
rect 10609 24633 10643 24667
rect 13829 24633 13863 24667
rect 17325 24633 17359 24667
rect 6745 24565 6779 24599
rect 9321 24565 9355 24599
rect 9597 24565 9631 24599
rect 10977 24565 11011 24599
rect 11529 24565 11563 24599
rect 12541 24565 12575 24599
rect 14749 24565 14783 24599
rect 15945 24565 15979 24599
rect 2145 24361 2179 24395
rect 6193 24361 6227 24395
rect 11437 24361 11471 24395
rect 11621 24361 11655 24395
rect 12541 24361 12575 24395
rect 12725 24361 12759 24395
rect 13001 24361 13035 24395
rect 13829 24361 13863 24395
rect 14565 24361 14599 24395
rect 14749 24361 14783 24395
rect 15485 24361 15519 24395
rect 15669 24361 15703 24395
rect 19073 24361 19107 24395
rect 19257 24361 19291 24395
rect 15853 24293 15887 24327
rect 8401 24225 8435 24259
rect 8585 24225 8619 24259
rect 10425 24225 10459 24259
rect 10793 24225 10827 24259
rect 11161 24225 11195 24259
rect 16313 24225 16347 24259
rect 16405 24225 16439 24259
rect 4813 24157 4847 24191
rect 6377 24157 6411 24191
rect 8309 24157 8343 24191
rect 10977 24157 11011 24191
rect 11989 24157 12023 24191
rect 12173 24157 12207 24191
rect 15117 24157 15151 24191
rect 17509 24157 17543 24191
rect 5080 24089 5114 24123
rect 6622 24089 6656 24123
rect 10158 24089 10192 24123
rect 12587 24089 12621 24123
rect 14197 24089 14231 24123
rect 14574 24089 14608 24123
rect 17754 24089 17788 24123
rect 19257 24157 19291 24191
rect 19441 24157 19475 24191
rect 7757 24021 7791 24055
rect 7941 24021 7975 24055
rect 9045 24021 9079 24055
rect 10609 24021 10643 24055
rect 11612 24021 11646 24055
rect 15494 24021 15528 24055
rect 16221 24021 16255 24055
rect 18889 24021 18923 24055
rect 19073 24021 19107 24055
rect 19625 24021 19659 24055
rect 5273 23817 5307 23851
rect 5917 23817 5951 23851
rect 8033 23817 8067 23851
rect 10149 23817 10183 23851
rect 11713 23817 11747 23851
rect 11989 23817 12023 23851
rect 12265 23817 12299 23851
rect 13277 23817 13311 23851
rect 17049 23817 17083 23851
rect 4905 23749 4939 23783
rect 5089 23749 5123 23783
rect 9965 23749 9999 23783
rect 12909 23749 12943 23783
rect 15853 23749 15887 23783
rect 16267 23749 16301 23783
rect 20637 23749 20671 23783
rect 20821 23749 20855 23783
rect 5365 23681 5399 23715
rect 5549 23681 5583 23715
rect 5733 23681 5767 23715
rect 5917 23681 5951 23715
rect 6469 23681 6503 23715
rect 6653 23681 6687 23715
rect 7021 23681 7055 23715
rect 7389 23681 7423 23715
rect 7481 23681 7515 23715
rect 7849 23681 7883 23715
rect 8405 23681 8439 23715
rect 8677 23681 8711 23715
rect 8769 23681 8803 23715
rect 8953 23681 8987 23715
rect 9045 23681 9079 23715
rect 9597 23681 9631 23715
rect 10149 23681 10183 23715
rect 10425 23681 10459 23715
rect 10517 23681 10551 23715
rect 11069 23681 11103 23715
rect 11529 23681 11563 23715
rect 12173 23681 12207 23715
rect 12449 23681 12483 23715
rect 16497 23681 16531 23715
rect 16865 23681 16899 23715
rect 17509 23681 17543 23715
rect 17601 23681 17635 23715
rect 18153 23681 18187 23715
rect 18395 23681 18429 23715
rect 18797 23681 18831 23715
rect 19156 23681 19190 23715
rect 20453 23681 20487 23715
rect 7205 23613 7239 23647
rect 7573 23613 7607 23647
rect 7665 23613 7699 23647
rect 8221 23613 8255 23647
rect 8309 23613 8343 23647
rect 8493 23613 8527 23647
rect 9413 23613 9447 23647
rect 9873 23613 9907 23647
rect 12633 23613 12667 23647
rect 12817 23613 12851 23647
rect 16681 23613 16715 23647
rect 17693 23613 17727 23647
rect 18705 23613 18739 23647
rect 18889 23613 18923 23647
rect 6193 23545 6227 23579
rect 17141 23545 17175 23579
rect 6745 23477 6779 23511
rect 8861 23477 8895 23511
rect 9229 23477 9263 23511
rect 10609 23477 10643 23511
rect 10885 23477 10919 23511
rect 11253 23477 11287 23511
rect 15669 23477 15703 23511
rect 16221 23477 16255 23511
rect 20269 23477 20303 23511
rect 7205 23273 7239 23307
rect 8493 23273 8527 23307
rect 14197 23273 14231 23307
rect 16589 23273 16623 23307
rect 18705 23273 18739 23307
rect 19257 23273 19291 23307
rect 6745 23205 6779 23239
rect 8033 23205 8067 23239
rect 10241 23205 10275 23239
rect 13461 23205 13495 23239
rect 7481 23137 7515 23171
rect 7573 23137 7607 23171
rect 15301 23137 15335 23171
rect 15761 23137 15795 23171
rect 15945 23137 15979 23171
rect 17325 23137 17359 23171
rect 19809 23137 19843 23171
rect 2145 23069 2179 23103
rect 6837 23069 6871 23103
rect 7389 23069 7423 23103
rect 7665 23069 7699 23103
rect 7849 23069 7883 23103
rect 7941 23069 7975 23103
rect 8953 23069 8987 23103
rect 9137 23069 9171 23103
rect 9505 23069 9539 23103
rect 9781 23069 9815 23103
rect 9873 23069 9907 23103
rect 13277 23069 13311 23103
rect 14381 23069 14415 23103
rect 18153 23069 18187 23103
rect 18429 23069 18463 23103
rect 20269 23069 20303 23103
rect 20545 23069 20579 23103
rect 22109 23069 22143 23103
rect 8309 23001 8343 23035
rect 8493 23001 8527 23035
rect 9689 23001 9723 23035
rect 10057 23001 10091 23035
rect 14657 23001 14691 23035
rect 14841 23001 14875 23035
rect 18696 23001 18730 23035
rect 19073 23001 19107 23035
rect 19625 23001 19659 23035
rect 20790 23001 20824 23035
rect 22354 23001 22388 23035
rect 6469 22933 6503 22967
rect 7021 22933 7055 22967
rect 8677 22933 8711 22967
rect 9137 22933 9171 22967
rect 12449 22933 12483 22967
rect 14565 22933 14599 22967
rect 16129 22933 16163 22967
rect 16221 22933 16255 22967
rect 18337 22933 18371 22967
rect 19717 22933 19751 22967
rect 20177 22933 20211 22967
rect 20453 22933 20487 22967
rect 21925 22933 21959 22967
rect 23489 22933 23523 22967
rect 7205 22729 7239 22763
rect 7665 22729 7699 22763
rect 8309 22729 8343 22763
rect 9045 22729 9079 22763
rect 14473 22729 14507 22763
rect 15301 22729 15335 22763
rect 15761 22729 15795 22763
rect 17049 22729 17083 22763
rect 17509 22729 17543 22763
rect 17877 22729 17911 22763
rect 19533 22729 19567 22763
rect 20094 22729 20128 22763
rect 22201 22729 22235 22763
rect 22753 22729 22787 22763
rect 7297 22661 7331 22695
rect 8861 22661 8895 22695
rect 10057 22661 10091 22695
rect 10517 22661 10551 22695
rect 18429 22661 18463 22695
rect 20913 22661 20947 22695
rect 23765 22661 23799 22695
rect 4077 22593 4111 22627
rect 7849 22593 7883 22627
rect 8401 22593 8435 22627
rect 8585 22593 8619 22627
rect 8769 22593 8803 22627
rect 9229 22593 9263 22627
rect 9321 22593 9355 22627
rect 10701 22593 10735 22627
rect 11897 22593 11931 22627
rect 14105 22593 14139 22627
rect 14933 22593 14967 22627
rect 18705 22593 18739 22627
rect 18981 22593 19015 22627
rect 19440 22593 19474 22627
rect 19717 22593 19751 22627
rect 20361 22593 20395 22627
rect 20821 22593 20855 22627
rect 22017 22593 22051 22627
rect 22661 22593 22695 22627
rect 23213 22593 23247 22627
rect 23580 22593 23614 22627
rect 23857 22593 23891 22627
rect 24225 22593 24259 22627
rect 4261 22525 4295 22559
rect 7113 22525 7147 22559
rect 9597 22525 9631 22559
rect 10149 22525 10183 22559
rect 10333 22525 10367 22559
rect 11253 22525 11287 22559
rect 13645 22525 13679 22559
rect 13829 22525 13863 22559
rect 14013 22525 14047 22559
rect 14657 22525 14691 22559
rect 14841 22525 14875 22559
rect 15853 22525 15887 22559
rect 16037 22525 16071 22559
rect 16773 22525 16807 22559
rect 16957 22525 16991 22559
rect 17969 22525 18003 22559
rect 18061 22525 18095 22559
rect 19073 22525 19107 22559
rect 21097 22525 21131 22559
rect 21925 22525 21959 22559
rect 22845 22525 22879 22559
rect 23121 22525 23155 22559
rect 24409 22525 24443 22559
rect 11069 22457 11103 22491
rect 15393 22457 15427 22491
rect 17417 22457 17451 22491
rect 18889 22457 18923 22491
rect 3893 22389 3927 22423
rect 7941 22389 7975 22423
rect 9505 22389 9539 22423
rect 9689 22389 9723 22423
rect 10793 22389 10827 22423
rect 12081 22389 12115 22423
rect 16405 22389 16439 22423
rect 18521 22389 18555 22423
rect 20085 22389 20119 22423
rect 20453 22389 20487 22423
rect 22293 22389 22327 22423
rect 23949 22389 23983 22423
rect 8033 22185 8067 22219
rect 9505 22185 9539 22219
rect 10241 22185 10275 22219
rect 13461 22185 13495 22219
rect 14105 22185 14139 22219
rect 16221 22185 16255 22219
rect 17233 22185 17267 22219
rect 20361 22185 20395 22219
rect 22109 22185 22143 22219
rect 22845 22185 22879 22219
rect 23397 22185 23431 22219
rect 24869 22185 24903 22219
rect 5917 22117 5951 22151
rect 22293 22117 22327 22151
rect 23213 22117 23247 22151
rect 6009 22049 6043 22083
rect 8953 22049 8987 22083
rect 13829 22049 13863 22083
rect 14749 22049 14783 22083
rect 15669 22049 15703 22083
rect 16865 22049 16899 22083
rect 23857 22049 23891 22083
rect 23949 22049 23983 22083
rect 1961 21981 1995 22015
rect 3801 21981 3835 22015
rect 5641 21981 5675 22015
rect 5733 21981 5767 22015
rect 8125 21981 8159 22015
rect 8769 21981 8803 22015
rect 9137 21981 9171 22015
rect 9689 21981 9723 22015
rect 9873 21981 9907 22015
rect 9965 21981 9999 22015
rect 10425 21981 10459 22015
rect 11253 21981 11287 22015
rect 13093 21981 13127 22015
rect 13369 21981 13403 22015
rect 15209 21981 15243 22015
rect 15393 21981 15427 22015
rect 16313 21981 16347 22015
rect 16497 21981 16531 22015
rect 16681 21981 16715 22015
rect 17417 21981 17451 22015
rect 21741 21981 21775 22015
rect 22477 21981 22511 22015
rect 23121 21981 23155 22015
rect 24685 21981 24719 22015
rect 25237 21981 25271 22015
rect 2228 21913 2262 21947
rect 4068 21913 4102 21947
rect 11520 21913 11554 21947
rect 12909 21913 12943 21947
rect 13277 21913 13311 21947
rect 15853 21913 15887 21947
rect 17049 21913 17083 21947
rect 17509 21913 17543 21947
rect 22155 21913 22189 21947
rect 22854 21913 22888 21947
rect 24409 21913 24443 21947
rect 3341 21845 3375 21879
rect 5181 21845 5215 21879
rect 5457 21845 5491 21879
rect 7849 21845 7883 21879
rect 8677 21845 8711 21879
rect 9229 21845 9263 21879
rect 10149 21845 10183 21879
rect 12633 21845 12667 21879
rect 14473 21845 14507 21879
rect 14565 21845 14599 21879
rect 15025 21845 15059 21879
rect 15761 21845 15795 21879
rect 23765 21845 23799 21879
rect 24501 21845 24535 21879
rect 25053 21845 25087 21879
rect 3249 21641 3283 21675
rect 4261 21641 4295 21675
rect 5825 21641 5859 21675
rect 7481 21641 7515 21675
rect 8401 21641 8435 21675
rect 10609 21641 10643 21675
rect 11161 21641 11195 21675
rect 11621 21641 11655 21675
rect 12633 21641 12667 21675
rect 13829 21641 13863 21675
rect 14749 21641 14783 21675
rect 15853 21641 15887 21675
rect 23213 21641 23247 21675
rect 21833 21573 21867 21607
rect 22017 21573 22051 21607
rect 23664 21573 23698 21607
rect 3433 21505 3467 21539
rect 3525 21505 3559 21539
rect 5374 21505 5408 21539
rect 6009 21505 6043 21539
rect 6561 21505 6595 21539
rect 7021 21505 7055 21539
rect 7665 21505 7699 21539
rect 8217 21505 8251 21539
rect 9045 21505 9079 21539
rect 9413 21505 9447 21539
rect 9689 21505 9723 21539
rect 10057 21505 10091 21539
rect 10149 21505 10183 21539
rect 10425 21505 10459 21539
rect 11345 21505 11379 21539
rect 11805 21505 11839 21539
rect 11989 21505 12023 21539
rect 12081 21505 12115 21539
rect 12265 21505 12299 21539
rect 12817 21505 12851 21539
rect 13093 21505 13127 21539
rect 13553 21505 13587 21539
rect 13829 21505 13863 21539
rect 14565 21505 14599 21539
rect 15209 21505 15243 21539
rect 15301 21505 15335 21539
rect 15485 21505 15519 21539
rect 15669 21505 15703 21539
rect 18337 21505 18371 21539
rect 18521 21505 18555 21539
rect 23121 21505 23155 21539
rect 23213 21505 23247 21539
rect 23397 21505 23431 21539
rect 3709 21437 3743 21471
rect 3801 21437 3835 21471
rect 5641 21437 5675 21471
rect 6193 21437 6227 21471
rect 6377 21437 6411 21471
rect 9229 21437 9263 21471
rect 9873 21437 9907 21471
rect 11897 21437 11931 21471
rect 13369 21437 13403 21471
rect 22201 21437 22235 21471
rect 7389 21369 7423 21403
rect 9689 21369 9723 21403
rect 16037 21369 16071 21403
rect 6745 21301 6779 21335
rect 7113 21301 7147 21335
rect 9321 21301 9355 21335
rect 10333 21301 10367 21335
rect 13277 21301 13311 21335
rect 14105 21301 14139 21335
rect 18245 21301 18279 21335
rect 24777 21301 24811 21335
rect 3985 21097 4019 21131
rect 4169 21097 4203 21131
rect 4629 21097 4663 21131
rect 8401 21097 8435 21131
rect 9229 21097 9263 21131
rect 9873 21097 9907 21131
rect 10333 21097 10367 21131
rect 17693 21097 17727 21131
rect 22477 21097 22511 21131
rect 22661 21097 22695 21131
rect 23121 21097 23155 21131
rect 23765 21097 23799 21131
rect 23949 21097 23983 21131
rect 24501 21097 24535 21131
rect 7849 21029 7883 21063
rect 4721 20961 4755 20995
rect 7021 20961 7055 20995
rect 7297 20961 7331 20995
rect 8585 20961 8619 20995
rect 9321 20961 9355 20995
rect 3249 20893 3283 20927
rect 3341 20893 3375 20927
rect 3801 20893 3835 20927
rect 4353 20893 4387 20927
rect 4445 20893 4479 20927
rect 6377 20893 6411 20927
rect 6745 20893 6779 20927
rect 6837 20893 6871 20927
rect 7113 20893 7147 20927
rect 7481 20893 7515 20927
rect 7665 20893 7699 20927
rect 8033 20893 8067 20927
rect 8401 20893 8435 20927
rect 9413 20893 9447 20927
rect 9689 20893 9723 20927
rect 6132 20825 6166 20859
rect 6561 20825 6595 20859
rect 8677 20825 8711 20859
rect 15117 20961 15151 20995
rect 17417 20961 17451 20995
rect 19809 20961 19843 20995
rect 23029 20961 23063 20995
rect 9965 20893 9999 20927
rect 10149 20893 10183 20927
rect 11345 20893 11379 20927
rect 14841 20893 14875 20927
rect 15485 20893 15519 20927
rect 17050 20893 17084 20927
rect 17509 20893 17543 20927
rect 19073 20893 19107 20927
rect 19349 20893 19383 20927
rect 22385 20893 22419 20927
rect 22477 20893 22511 20927
rect 22845 20893 22879 20927
rect 23581 20893 23615 20927
rect 23765 20893 23799 20927
rect 24593 20893 24627 20927
rect 10609 20825 10643 20859
rect 11069 20825 11103 20859
rect 15301 20825 15335 20859
rect 18828 20825 18862 20859
rect 20076 20825 20110 20859
rect 23121 20825 23155 20859
rect 3525 20757 3559 20791
rect 4997 20757 5031 20791
rect 8217 20757 8251 20791
rect 9045 20757 9079 20791
rect 9505 20757 9539 20791
rect 9873 20757 9907 20791
rect 10885 20757 10919 20791
rect 10977 20757 11011 20791
rect 14657 20757 14691 20791
rect 16957 20757 16991 20791
rect 19533 20757 19567 20791
rect 19717 20757 19751 20791
rect 21189 20757 21223 20791
rect 22109 20757 22143 20791
rect 4445 20553 4479 20587
rect 5273 20553 5307 20587
rect 7757 20553 7791 20587
rect 8769 20553 8803 20587
rect 9965 20553 9999 20587
rect 11345 20553 11379 20587
rect 15577 20553 15611 20587
rect 16221 20553 16255 20587
rect 18061 20553 18095 20587
rect 22569 20553 22603 20587
rect 3985 20485 4019 20519
rect 5825 20485 5859 20519
rect 16313 20485 16347 20519
rect 23029 20485 23063 20519
rect 1685 20417 1719 20451
rect 1952 20417 1986 20451
rect 3341 20417 3375 20451
rect 3525 20417 3559 20451
rect 3617 20417 3651 20451
rect 3893 20417 3927 20451
rect 4169 20417 4203 20451
rect 4353 20417 4387 20451
rect 4629 20417 4663 20451
rect 4905 20417 4939 20451
rect 5089 20417 5123 20451
rect 5181 20417 5215 20451
rect 5457 20417 5491 20451
rect 5549 20417 5583 20451
rect 5733 20417 5767 20451
rect 5922 20417 5956 20451
rect 6633 20417 6667 20451
rect 9873 20417 9907 20451
rect 10885 20417 10919 20451
rect 11161 20417 11195 20451
rect 11529 20417 11563 20451
rect 11785 20417 11819 20451
rect 14197 20417 14231 20451
rect 14464 20417 14498 20451
rect 16037 20417 16071 20451
rect 16681 20417 16715 20451
rect 16937 20417 16971 20451
rect 18613 20417 18647 20451
rect 19073 20417 19107 20451
rect 19165 20417 19199 20451
rect 20085 20417 20119 20451
rect 20177 20417 20211 20451
rect 20913 20417 20947 20451
rect 21098 20417 21132 20451
rect 21465 20417 21499 20451
rect 22753 20417 22787 20451
rect 24317 20417 24351 20451
rect 24501 20417 24535 20451
rect 24777 20417 24811 20451
rect 3801 20349 3835 20383
rect 6377 20349 6411 20383
rect 18705 20349 18739 20383
rect 18797 20349 18831 20383
rect 20361 20349 20395 20383
rect 21557 20349 21591 20383
rect 22937 20349 22971 20383
rect 4721 20281 4755 20315
rect 6101 20281 6135 20315
rect 11069 20281 11103 20315
rect 19441 20281 19475 20315
rect 3065 20213 3099 20247
rect 4353 20213 4387 20247
rect 8033 20213 8067 20247
rect 12909 20213 12943 20247
rect 15853 20213 15887 20247
rect 18245 20213 18279 20247
rect 19073 20213 19107 20247
rect 19717 20213 19751 20247
rect 23029 20213 23063 20247
rect 24225 20213 24259 20247
rect 24593 20213 24627 20247
rect 6285 20009 6319 20043
rect 11713 20009 11747 20043
rect 14749 20009 14783 20043
rect 14933 20009 14967 20043
rect 16313 20009 16347 20043
rect 18429 20009 18463 20043
rect 18981 20009 19015 20043
rect 19625 20009 19659 20043
rect 20177 20009 20211 20043
rect 11621 19941 11655 19975
rect 12817 19941 12851 19975
rect 15117 19941 15151 19975
rect 22201 19941 22235 19975
rect 1501 19873 1535 19907
rect 3433 19873 3467 19907
rect 4353 19873 4387 19907
rect 4445 19873 4479 19907
rect 12357 19873 12391 19907
rect 15577 19873 15611 19907
rect 15761 19873 15795 19907
rect 17049 19873 17083 19907
rect 17233 19873 17267 19907
rect 17877 19873 17911 19907
rect 22937 19873 22971 19907
rect 24133 19873 24167 19907
rect 25513 19873 25547 19907
rect 3157 19805 3191 19839
rect 3249 19805 3283 19839
rect 4077 19805 4111 19839
rect 4169 19805 4203 19839
rect 4537 19805 4571 19839
rect 4721 19805 4755 19839
rect 7113 19805 7147 19839
rect 11161 19805 11195 19839
rect 11253 19805 11287 19839
rect 11437 19805 11471 19839
rect 11897 19805 11931 19839
rect 11989 19805 12023 19839
rect 12154 19805 12188 19839
rect 12265 19805 12299 19839
rect 12541 19805 12575 19839
rect 13001 19805 13035 19839
rect 14381 19805 14415 19839
rect 16129 19805 16163 19839
rect 16497 19805 16531 19839
rect 18705 19805 18739 19839
rect 18797 19805 18831 19839
rect 19901 19805 19935 19839
rect 19993 19805 20027 19839
rect 20821 19805 20855 19839
rect 22570 19805 22604 19839
rect 23029 19805 23063 19839
rect 23305 19805 23339 19839
rect 23489 19805 23523 19839
rect 23823 19805 23857 19839
rect 24225 19805 24259 19839
rect 24651 19805 24685 19839
rect 24961 19805 24995 19839
rect 25053 19805 25087 19839
rect 25145 19805 25179 19839
rect 1768 19737 1802 19771
rect 3893 19737 3927 19771
rect 14758 19737 14792 19771
rect 15485 19737 15519 19771
rect 18061 19737 18095 19771
rect 19257 19737 19291 19771
rect 21088 19737 21122 19771
rect 22385 19737 22419 19771
rect 23121 19737 23155 19771
rect 24409 19737 24443 19771
rect 25329 19737 25363 19771
rect 2881 19669 2915 19703
rect 4905 19669 4939 19703
rect 6929 19669 6963 19703
rect 7297 19669 7331 19703
rect 11069 19669 11103 19703
rect 12633 19669 12667 19703
rect 16589 19669 16623 19703
rect 16957 19669 16991 19703
rect 18438 19669 18472 19703
rect 19634 19669 19668 19703
rect 20545 19669 20579 19703
rect 23673 19669 23707 19703
rect 3525 19465 3559 19499
rect 4445 19465 4479 19499
rect 8769 19465 8803 19499
rect 10241 19465 10275 19499
rect 10885 19465 10919 19499
rect 14105 19465 14139 19499
rect 15770 19465 15804 19499
rect 18705 19465 18739 19499
rect 19533 19465 19567 19499
rect 20278 19465 20312 19499
rect 21097 19465 21131 19499
rect 21465 19465 21499 19499
rect 22753 19465 22787 19499
rect 25513 19465 25547 19499
rect 9106 19397 9140 19431
rect 12970 19397 13004 19431
rect 15393 19397 15427 19431
rect 19901 19397 19935 19431
rect 23590 19397 23624 19431
rect 2145 19329 2179 19363
rect 2412 19329 2446 19363
rect 3801 19329 3835 19363
rect 3985 19329 4019 19363
rect 4077 19329 4111 19363
rect 4353 19329 4387 19363
rect 4629 19329 4663 19363
rect 6561 19329 6595 19363
rect 6930 19329 6964 19363
rect 7113 19329 7147 19363
rect 7205 19329 7239 19363
rect 7389 19329 7423 19363
rect 7849 19329 7883 19363
rect 8585 19329 8619 19363
rect 8861 19329 8895 19363
rect 11069 19329 11103 19363
rect 11345 19329 11379 19363
rect 11529 19329 11563 19363
rect 11712 19329 11746 19363
rect 11805 19329 11839 19363
rect 11897 19329 11931 19363
rect 12081 19329 12115 19363
rect 16037 19329 16071 19363
rect 18245 19329 18279 19363
rect 18555 19329 18589 19363
rect 19717 19329 19751 19363
rect 20545 19329 20579 19363
rect 21005 19329 21039 19363
rect 21649 19329 21683 19363
rect 22167 19329 22201 19363
rect 23121 19329 23155 19363
rect 23213 19329 23247 19363
rect 23857 19329 23891 19363
rect 24400 19329 24434 19363
rect 4261 19261 4295 19295
rect 6745 19261 6779 19295
rect 6837 19261 6871 19295
rect 12725 19261 12759 19295
rect 15025 19261 15059 19295
rect 18153 19261 18187 19295
rect 21281 19261 21315 19295
rect 22477 19261 22511 19295
rect 22569 19261 22603 19295
rect 23029 19261 23063 19295
rect 24133 19261 24167 19295
rect 7481 19193 7515 19227
rect 11161 19193 11195 19227
rect 12357 19193 12391 19227
rect 20637 19193 20671 19227
rect 6469 19125 6503 19159
rect 7757 19125 7791 19159
rect 10793 19125 10827 19159
rect 12173 19125 12207 19159
rect 15761 19125 15795 19159
rect 20269 19125 20303 19159
rect 22017 19125 22051 19159
rect 23121 19125 23155 19159
rect 23581 19125 23615 19159
rect 5549 18921 5583 18955
rect 9045 18921 9079 18955
rect 15669 18921 15703 18955
rect 20453 18921 20487 18955
rect 22201 18921 22235 18955
rect 23121 18921 23155 18955
rect 23305 18921 23339 18955
rect 25237 18921 25271 18955
rect 11253 18853 11287 18887
rect 17141 18853 17175 18887
rect 20637 18853 20671 18887
rect 24409 18853 24443 18887
rect 17877 18785 17911 18819
rect 23949 18785 23983 18819
rect 24133 18785 24167 18819
rect 24869 18785 24903 18819
rect 25053 18785 25087 18819
rect 25513 18785 25547 18819
rect 5365 18717 5399 18751
rect 5641 18717 5675 18751
rect 5908 18717 5942 18751
rect 7205 18717 7239 18751
rect 10425 18717 10459 18751
rect 11069 18717 11103 18751
rect 11529 18717 11563 18751
rect 11805 18717 11839 18751
rect 14289 18717 14323 18751
rect 20085 18717 20119 18751
rect 20821 18717 20855 18751
rect 22753 18717 22787 18751
rect 25421 18717 25455 18751
rect 7472 18649 7506 18683
rect 10180 18649 10214 18683
rect 12072 18649 12106 18683
rect 14556 18649 14590 18683
rect 16497 18649 16531 18683
rect 20462 18649 20496 18683
rect 21088 18649 21122 18683
rect 23167 18649 23201 18683
rect 24777 18649 24811 18683
rect 4169 18581 4203 18615
rect 7021 18581 7055 18615
rect 8585 18581 8619 18615
rect 11345 18581 11379 18615
rect 13185 18581 13219 18615
rect 16129 18581 16163 18615
rect 16405 18581 16439 18615
rect 17325 18581 17359 18615
rect 17693 18581 17727 18615
rect 17785 18581 17819 18615
rect 23489 18581 23523 18615
rect 23857 18581 23891 18615
rect 4353 18377 4387 18411
rect 8493 18377 8527 18411
rect 14749 18377 14783 18411
rect 15577 18377 15611 18411
rect 18981 18377 19015 18411
rect 21005 18377 21039 18411
rect 21373 18377 21407 18411
rect 21833 18377 21867 18411
rect 22293 18377 22327 18411
rect 23397 18377 23431 18411
rect 25421 18377 25455 18411
rect 8125 18309 8159 18343
rect 8309 18309 8343 18343
rect 9689 18309 9723 18343
rect 11345 18309 11379 18343
rect 15945 18309 15979 18343
rect 18889 18309 18923 18343
rect 21649 18309 21683 18343
rect 24308 18309 24342 18343
rect 3065 18241 3099 18275
rect 3434 18241 3468 18275
rect 3617 18241 3651 18275
rect 3801 18241 3835 18275
rect 4261 18241 4295 18275
rect 4537 18241 4571 18275
rect 4629 18241 4663 18275
rect 4812 18241 4846 18275
rect 4905 18241 4939 18275
rect 5181 18241 5215 18275
rect 5463 18241 5497 18275
rect 5622 18247 5656 18281
rect 5733 18241 5767 18275
rect 6009 18241 6043 18275
rect 6377 18241 6411 18275
rect 6633 18241 6667 18275
rect 11529 18241 11563 18275
rect 11712 18241 11746 18275
rect 11897 18241 11931 18275
rect 12081 18241 12115 18275
rect 13369 18241 13403 18275
rect 13625 18241 13659 18275
rect 14933 18241 14967 18275
rect 15116 18247 15150 18281
rect 15209 18241 15243 18275
rect 15485 18241 15519 18275
rect 16773 18241 16807 18275
rect 16957 18241 16991 18275
rect 17325 18241 17359 18275
rect 17785 18241 17819 18275
rect 18245 18241 18279 18275
rect 18429 18241 18463 18275
rect 20821 18241 20855 18275
rect 21189 18241 21223 18275
rect 22201 18241 22235 18275
rect 3249 18173 3283 18207
rect 3341 18173 3375 18207
rect 4997 18173 5031 18207
rect 5825 18173 5859 18207
rect 6193 18173 6227 18207
rect 11805 18173 11839 18207
rect 15301 18173 15335 18207
rect 17233 18173 17267 18207
rect 17877 18173 17911 18207
rect 17969 18173 18003 18207
rect 22477 18173 22511 18207
rect 24041 18173 24075 18207
rect 2881 18105 2915 18139
rect 3985 18105 4019 18139
rect 15761 18105 15795 18139
rect 17417 18105 17451 18139
rect 19165 18105 19199 18139
rect 4077 18037 4111 18071
rect 5273 18037 5307 18071
rect 7757 18037 7791 18071
rect 8309 18037 8343 18071
rect 12173 18037 12207 18071
rect 18613 18037 18647 18071
rect 5365 17833 5399 17867
rect 12909 17833 12943 17867
rect 13737 17833 13771 17867
rect 16773 17833 16807 17867
rect 18061 17833 18095 17867
rect 19257 17833 19291 17867
rect 10517 17765 10551 17799
rect 4629 17697 4663 17731
rect 4721 17697 4755 17731
rect 10977 17697 11011 17731
rect 13369 17697 13403 17731
rect 13461 17697 13495 17731
rect 14657 17697 14691 17731
rect 15117 17697 15151 17731
rect 17325 17697 17359 17731
rect 18613 17697 18647 17731
rect 19809 17697 19843 17731
rect 2053 17629 2087 17663
rect 4353 17629 4387 17663
rect 4536 17629 4570 17663
rect 4905 17629 4939 17663
rect 5549 17629 5583 17663
rect 5733 17629 5767 17663
rect 5989 17629 6023 17663
rect 8953 17629 8987 17663
rect 10701 17629 10735 17663
rect 10885 17629 10919 17663
rect 11070 17623 11104 17657
rect 11253 17629 11287 17663
rect 11529 17629 11563 17663
rect 11796 17629 11830 17663
rect 13093 17629 13127 17663
rect 13276 17629 13310 17663
rect 13645 17629 13679 17663
rect 14381 17629 14415 17663
rect 14546 17629 14580 17663
rect 14749 17629 14783 17663
rect 14933 17629 14967 17663
rect 15209 17629 15243 17663
rect 15465 17629 15499 17663
rect 17141 17629 17175 17663
rect 17601 17629 17635 17663
rect 17877 17629 17911 17663
rect 19073 17629 19107 17663
rect 2320 17561 2354 17595
rect 3985 17561 4019 17595
rect 4169 17561 4203 17595
rect 9220 17561 9254 17595
rect 19717 17561 19751 17595
rect 3433 17493 3467 17527
rect 4997 17493 5031 17527
rect 7113 17493 7147 17527
rect 10333 17493 10367 17527
rect 16589 17493 16623 17527
rect 17233 17493 17267 17527
rect 17693 17493 17727 17527
rect 18429 17493 18463 17527
rect 18521 17493 18555 17527
rect 18889 17493 18923 17527
rect 19625 17493 19659 17527
rect 3249 17289 3283 17323
rect 6561 17289 6595 17323
rect 9689 17289 9723 17323
rect 9873 17289 9907 17323
rect 12909 17289 12943 17323
rect 15301 17289 15335 17323
rect 18061 17289 18095 17323
rect 19993 17289 20027 17323
rect 20269 17289 20303 17323
rect 8401 17221 8435 17255
rect 11345 17221 11379 17255
rect 11774 17221 11808 17255
rect 18245 17221 18279 17255
rect 21097 17221 21131 17255
rect 23949 17221 23983 17255
rect 1869 17153 1903 17187
rect 2136 17153 2170 17187
rect 3792 17153 3826 17187
rect 5089 17153 5123 17187
rect 5273 17153 5307 17187
rect 5457 17153 5491 17187
rect 5677 17156 5711 17190
rect 5825 17153 5859 17187
rect 6101 17153 6135 17187
rect 6653 17153 6687 17187
rect 8861 17153 8895 17187
rect 9045 17153 9079 17187
rect 9230 17153 9264 17187
rect 9413 17153 9447 17187
rect 9965 17153 9999 17187
rect 10103 17153 10137 17187
rect 10241 17153 10275 17187
rect 10351 17153 10385 17187
rect 10517 17153 10551 17187
rect 10609 17153 10643 17187
rect 10792 17153 10826 17187
rect 10885 17153 10919 17187
rect 11161 17153 11195 17187
rect 16937 17153 16971 17187
rect 18337 17153 18371 17187
rect 18521 17153 18555 17187
rect 18889 17153 18923 17187
rect 19625 17153 19659 17187
rect 20085 17153 20119 17187
rect 20729 17153 20763 17187
rect 24225 17153 24259 17187
rect 3525 17085 3559 17119
rect 5549 17085 5583 17119
rect 6837 17085 6871 17119
rect 8217 17085 8251 17119
rect 9137 17085 9171 17119
rect 10977 17085 11011 17119
rect 11529 17085 11563 17119
rect 16681 17085 16715 17119
rect 18705 17085 18739 17119
rect 19441 17085 19475 17119
rect 19533 17085 19567 17119
rect 20545 17085 20579 17119
rect 5917 17017 5951 17051
rect 8585 17017 8619 17051
rect 24409 17017 24443 17051
rect 4905 16949 4939 16983
rect 7113 16949 7147 16983
rect 8769 16949 8803 16983
rect 19073 16949 19107 16983
rect 20913 16949 20947 16983
rect 21833 16949 21867 16983
rect 22477 16949 22511 16983
rect 23121 16949 23155 16983
rect 23305 16949 23339 16983
rect 24501 16949 24535 16983
rect 3893 16745 3927 16779
rect 8769 16745 8803 16779
rect 10517 16745 10551 16779
rect 16773 16745 16807 16779
rect 17969 16745 18003 16779
rect 18705 16745 18739 16779
rect 19441 16745 19475 16779
rect 19625 16745 19659 16779
rect 25605 16745 25639 16779
rect 20913 16677 20947 16711
rect 2145 16609 2179 16643
rect 4629 16609 4663 16643
rect 8217 16609 8251 16643
rect 8953 16609 8987 16643
rect 12449 16609 12483 16643
rect 14565 16609 14599 16643
rect 16497 16609 16531 16643
rect 17325 16609 17359 16643
rect 17877 16609 17911 16643
rect 20361 16609 20395 16643
rect 20453 16609 20487 16643
rect 21465 16609 21499 16643
rect 21557 16609 21591 16643
rect 21925 16609 21959 16643
rect 23213 16609 23247 16643
rect 24041 16609 24075 16643
rect 24501 16609 24535 16643
rect 24685 16609 24719 16643
rect 2412 16541 2446 16575
rect 3985 16541 4019 16575
rect 4123 16541 4157 16575
rect 4242 16541 4276 16575
rect 4354 16541 4388 16575
rect 4549 16541 4583 16575
rect 4896 16541 4930 16575
rect 9209 16541 9243 16575
rect 10701 16541 10735 16575
rect 16129 16541 16163 16575
rect 16312 16535 16346 16569
rect 16405 16541 16439 16575
rect 16681 16541 16715 16575
rect 17417 16541 17451 16575
rect 17693 16541 17727 16575
rect 19809 16541 19843 16575
rect 20729 16541 20763 16575
rect 22201 16541 22235 16575
rect 25329 16541 25363 16575
rect 25421 16541 25455 16575
rect 8401 16473 8435 16507
rect 12716 16473 12750 16507
rect 14832 16473 14866 16507
rect 21373 16473 21407 16507
rect 22109 16473 22143 16507
rect 23121 16473 23155 16507
rect 23857 16473 23891 16507
rect 3525 16405 3559 16439
rect 6009 16405 6043 16439
rect 8309 16405 8343 16439
rect 10333 16405 10367 16439
rect 13829 16405 13863 16439
rect 15945 16405 15979 16439
rect 19349 16405 19383 16439
rect 19901 16405 19935 16439
rect 20269 16405 20303 16439
rect 21005 16405 21039 16439
rect 22569 16405 22603 16439
rect 22661 16405 22695 16439
rect 23029 16405 23063 16439
rect 23489 16405 23523 16439
rect 23949 16405 23983 16439
rect 24777 16405 24811 16439
rect 25145 16405 25179 16439
rect 9781 16201 9815 16235
rect 9965 16201 9999 16235
rect 10609 16201 10643 16235
rect 13093 16201 13127 16235
rect 14013 16201 14047 16235
rect 14841 16201 14875 16235
rect 20729 16201 20763 16235
rect 21189 16201 21223 16235
rect 21281 16201 21315 16235
rect 23213 16201 23247 16235
rect 24041 16201 24075 16235
rect 24869 16201 24903 16235
rect 24961 16201 24995 16235
rect 25421 16201 25455 16235
rect 2881 16133 2915 16167
rect 16405 16133 16439 16167
rect 16926 16133 16960 16167
rect 21833 16133 21867 16167
rect 23581 16133 23615 16167
rect 24501 16133 24535 16167
rect 3065 16065 3099 16099
rect 3249 16065 3283 16099
rect 3434 16065 3468 16099
rect 3617 16065 3651 16099
rect 8116 16065 8150 16099
rect 9597 16065 9631 16099
rect 9689 16065 9723 16099
rect 10241 16065 10275 16099
rect 10793 16065 10827 16099
rect 12449 16065 12483 16099
rect 12632 16065 12666 16099
rect 13001 16065 13035 16099
rect 14197 16065 14231 16099
rect 14380 16065 14414 16099
rect 14473 16065 14507 16099
rect 14749 16065 14783 16099
rect 15669 16065 15703 16099
rect 15817 16071 15851 16105
rect 15945 16065 15979 16099
rect 16221 16065 16255 16099
rect 20361 16065 20395 16099
rect 22109 16065 22143 16099
rect 22845 16065 22879 16099
rect 23673 16065 23707 16099
rect 25329 16065 25363 16099
rect 3341 15997 3375 16031
rect 7849 15997 7883 16031
rect 12725 15997 12759 16031
rect 12817 15997 12851 16031
rect 14565 15997 14599 16031
rect 16037 15997 16071 16031
rect 16681 15997 16715 16031
rect 19717 15997 19751 16031
rect 19901 15997 19935 16031
rect 20177 15997 20211 16031
rect 20269 15997 20303 16031
rect 21373 15997 21407 16031
rect 21833 15997 21867 16031
rect 21925 15997 21959 16031
rect 22569 15997 22603 16031
rect 22753 15997 22787 16031
rect 23397 15997 23431 16031
rect 24225 15997 24259 16031
rect 24409 15997 24443 16031
rect 25513 15997 25547 16031
rect 9229 15929 9263 15963
rect 10425 15929 10459 15963
rect 20821 15929 20855 15963
rect 9505 15861 9539 15895
rect 13369 15861 13403 15895
rect 18061 15861 18095 15895
rect 22293 15861 22327 15895
rect 3893 15657 3927 15691
rect 7021 15657 7055 15691
rect 9505 15657 9539 15691
rect 12081 15657 12115 15691
rect 12357 15657 12391 15691
rect 13553 15657 13587 15691
rect 14749 15657 14783 15691
rect 19073 15657 19107 15691
rect 19993 15657 20027 15691
rect 20453 15657 20487 15691
rect 21281 15657 21315 15691
rect 22845 15657 22879 15691
rect 22937 15657 22971 15691
rect 24133 15657 24167 15691
rect 24409 15657 24443 15691
rect 25237 15657 25271 15691
rect 11897 15589 11931 15623
rect 14289 15589 14323 15623
rect 3157 15521 3191 15555
rect 5641 15521 5675 15555
rect 8217 15521 8251 15555
rect 9045 15521 9079 15555
rect 10149 15521 10183 15555
rect 2973 15453 3007 15487
rect 3249 15453 3283 15487
rect 3342 15453 3376 15487
rect 3525 15453 3559 15487
rect 7389 15453 7423 15487
rect 8401 15453 8435 15487
rect 8493 15453 8527 15487
rect 9229 15453 9263 15487
rect 9321 15453 9355 15487
rect 9597 15453 9631 15487
rect 11713 15453 11747 15487
rect 12265 15453 12299 15487
rect 12541 15453 12575 15487
rect 13369 15453 13403 15487
rect 13645 15453 13679 15487
rect 14105 15453 14139 15487
rect 2789 15385 2823 15419
rect 5908 15385 5942 15419
rect 10416 15385 10450 15419
rect 25513 15589 25547 15623
rect 19349 15521 19383 15555
rect 19533 15521 19567 15555
rect 20913 15521 20947 15555
rect 21097 15521 21131 15555
rect 21833 15521 21867 15555
rect 22109 15521 22143 15555
rect 22293 15521 22327 15555
rect 22477 15521 22511 15555
rect 23489 15521 23523 15555
rect 23765 15521 23799 15555
rect 24961 15521 24995 15555
rect 18705 15453 18739 15487
rect 20177 15453 20211 15487
rect 20821 15453 20855 15487
rect 22661 15453 22695 15487
rect 23949 15453 23983 15487
rect 24777 15453 24811 15487
rect 25421 15453 25455 15487
rect 18245 15385 18279 15419
rect 18429 15385 18463 15419
rect 18613 15385 18647 15419
rect 21741 15385 21775 15419
rect 23305 15385 23339 15419
rect 24869 15385 24903 15419
rect 8033 15317 8067 15351
rect 11529 15317 11563 15351
rect 13829 15317 13863 15351
rect 14749 15317 14783 15351
rect 14933 15317 14967 15351
rect 18889 15317 18923 15351
rect 19625 15317 19659 15351
rect 20361 15317 20395 15351
rect 21649 15317 21683 15351
rect 23397 15317 23431 15351
rect 1593 15113 1627 15147
rect 4261 15113 4295 15147
rect 4721 15113 4755 15147
rect 8769 15113 8803 15147
rect 10609 15113 10643 15147
rect 18245 15113 18279 15147
rect 18797 15113 18831 15147
rect 19165 15113 19199 15147
rect 20269 15113 20303 15147
rect 20821 15113 20855 15147
rect 21281 15113 21315 15147
rect 23305 15113 23339 15147
rect 24317 15113 24351 15147
rect 24777 15045 24811 15079
rect 2717 14977 2751 15011
rect 2973 14977 3007 15011
rect 3433 14977 3467 15011
rect 3616 14977 3650 15011
rect 3985 14977 4019 15011
rect 4629 14977 4663 15011
rect 5089 14977 5123 15011
rect 6561 14977 6595 15011
rect 6653 14977 6687 15011
rect 6920 14977 6954 15011
rect 8953 14977 8987 15011
rect 9965 14977 9999 15011
rect 10148 14977 10182 15011
rect 10333 14977 10367 15011
rect 10517 14977 10551 15011
rect 12909 14977 12943 15011
rect 14933 14977 14967 15011
rect 15281 14977 15315 15011
rect 16681 14977 16715 15011
rect 16937 14977 16971 15011
rect 19533 14977 19567 15011
rect 20453 14977 20487 15011
rect 20821 14977 20855 15011
rect 21097 14977 21131 15011
rect 21189 14977 21223 15011
rect 23305 14977 23339 15011
rect 23581 14977 23615 15011
rect 23949 14977 23983 15011
rect 24133 14977 24167 15011
rect 3709 14909 3743 14943
rect 3801 14909 3835 14943
rect 4813 14909 4847 14943
rect 10241 14909 10275 14943
rect 15025 14909 15059 14943
rect 18521 14909 18555 14943
rect 18705 14909 18739 14943
rect 19993 14909 20027 14943
rect 20637 14909 20671 14943
rect 14749 14841 14783 14875
rect 4077 14773 4111 14807
rect 8033 14773 8067 14807
rect 9137 14773 9171 14807
rect 10885 14773 10919 14807
rect 12817 14773 12851 14807
rect 14197 14773 14231 14807
rect 16405 14773 16439 14807
rect 18061 14773 18095 14807
rect 19625 14773 19659 14807
rect 21557 14773 21591 14807
rect 23673 14773 23707 14807
rect 24501 14773 24535 14807
rect 5181 14569 5215 14603
rect 6285 14569 6319 14603
rect 7113 14569 7147 14603
rect 7297 14569 7331 14603
rect 8125 14569 8159 14603
rect 8677 14569 8711 14603
rect 11437 14569 11471 14603
rect 14841 14569 14875 14603
rect 16497 14569 16531 14603
rect 14105 14501 14139 14535
rect 18705 14501 18739 14535
rect 20177 14501 20211 14535
rect 3070 14433 3104 14467
rect 3801 14433 3835 14467
rect 5917 14433 5951 14467
rect 6745 14433 6779 14467
rect 6837 14433 6871 14467
rect 7757 14433 7791 14467
rect 7849 14433 7883 14467
rect 11989 14433 12023 14467
rect 2789 14365 2823 14399
rect 2973 14365 3007 14399
rect 3158 14365 3192 14399
rect 3341 14365 3375 14399
rect 4068 14365 4102 14399
rect 5641 14365 5675 14399
rect 5824 14365 5858 14399
rect 6009 14365 6043 14399
rect 6193 14365 6227 14399
rect 6469 14365 6503 14399
rect 6652 14365 6686 14399
rect 7021 14365 7055 14399
rect 8585 14365 8619 14399
rect 8763 14365 8797 14399
rect 8953 14365 8987 14399
rect 9229 14365 9263 14399
rect 9413 14365 9447 14399
rect 11621 14365 11655 14399
rect 11786 14365 11820 14399
rect 11897 14365 11931 14399
rect 12173 14365 12207 14399
rect 12449 14365 12483 14399
rect 7665 14297 7699 14331
rect 12357 14297 12391 14331
rect 12694 14297 12728 14331
rect 14473 14433 14507 14467
rect 14565 14433 14599 14467
rect 15301 14433 15335 14467
rect 15393 14433 15427 14467
rect 15761 14433 15795 14467
rect 16129 14433 16163 14467
rect 16221 14433 16255 14467
rect 18153 14433 18187 14467
rect 19625 14433 19659 14467
rect 20637 14433 20671 14467
rect 24225 14433 24259 14467
rect 14197 14365 14231 14399
rect 14380 14365 14414 14399
rect 14749 14365 14783 14399
rect 15025 14365 15059 14399
rect 15208 14365 15242 14399
rect 15577 14365 15611 14399
rect 15853 14365 15887 14399
rect 16036 14365 16070 14399
rect 16405 14365 16439 14399
rect 18061 14365 18095 14399
rect 18463 14365 18497 14399
rect 19809 14365 19843 14399
rect 20085 14365 20119 14399
rect 20453 14365 20487 14399
rect 23489 14365 23523 14399
rect 23581 14365 23615 14399
rect 23857 14365 23891 14399
rect 24133 14365 24167 14399
rect 24409 14365 24443 14399
rect 19441 14297 19475 14331
rect 19533 14297 19567 14331
rect 2697 14229 2731 14263
rect 8401 14229 8435 14263
rect 9045 14229 9079 14263
rect 9781 14229 9815 14263
rect 13829 14229 13863 14263
rect 14105 14229 14139 14263
rect 16681 14229 16715 14263
rect 23397 14229 23431 14263
rect 24501 14229 24535 14263
rect 3709 14025 3743 14059
rect 4813 14025 4847 14059
rect 5457 14025 5491 14059
rect 5917 14025 5951 14059
rect 6377 14025 6411 14059
rect 6837 14025 6871 14059
rect 7665 14025 7699 14059
rect 8125 14025 8159 14059
rect 11161 14025 11195 14059
rect 12909 14025 12943 14059
rect 14841 14025 14875 14059
rect 16405 14025 16439 14059
rect 17785 14025 17819 14059
rect 18613 14025 18647 14059
rect 19073 14025 19107 14059
rect 19717 14025 19751 14059
rect 20269 14025 20303 14059
rect 23305 14025 23339 14059
rect 24409 14025 24443 14059
rect 4077 13957 4111 13991
rect 8217 13957 8251 13991
rect 9781 13957 9815 13991
rect 15292 13957 15326 13991
rect 2973 13889 3007 13923
rect 3157 13889 3191 13923
rect 3342 13889 3376 13923
rect 3525 13889 3559 13923
rect 4169 13889 4203 13923
rect 4721 13889 4755 13923
rect 4997 13889 5031 13923
rect 5089 13889 5123 13923
rect 5632 13889 5666 13923
rect 5725 13889 5759 13923
rect 6009 13889 6043 13923
rect 6745 13889 6779 13923
rect 7573 13889 7607 13923
rect 8677 13889 8711 13923
rect 9137 13889 9171 13923
rect 9321 13889 9355 13923
rect 9597 13889 9631 13923
rect 11796 13889 11830 13923
rect 13093 13889 13127 13923
rect 13349 13889 13383 13923
rect 14657 13889 14691 13923
rect 15025 13889 15059 13923
rect 17693 13889 17727 13923
rect 18521 13889 18555 13923
rect 19073 13889 19107 13923
rect 19349 13889 19383 13923
rect 19441 13889 19475 13923
rect 19901 13889 19935 13923
rect 20085 13889 20119 13923
rect 20361 13889 20395 13923
rect 20453 13889 20487 13923
rect 20821 13889 20855 13923
rect 21097 13889 21131 13923
rect 21281 13889 21315 13923
rect 21833 13889 21867 13923
rect 22201 13889 22235 13923
rect 23213 13889 23247 13923
rect 23581 13889 23615 13923
rect 23949 13889 23983 13923
rect 24133 13889 24167 13923
rect 24317 13889 24351 13923
rect 3249 13821 3283 13855
rect 4353 13821 4387 13855
rect 4629 13821 4663 13855
rect 6929 13821 6963 13855
rect 7757 13821 7791 13855
rect 8953 13821 8987 13855
rect 11529 13821 11563 13855
rect 17877 13821 17911 13855
rect 18705 13821 18739 13855
rect 20913 13821 20947 13855
rect 22017 13821 22051 13855
rect 23765 13821 23799 13855
rect 2789 13753 2823 13787
rect 5273 13753 5307 13787
rect 8769 13753 8803 13787
rect 9413 13753 9447 13787
rect 17049 13753 17083 13787
rect 17233 13753 17267 13787
rect 21465 13753 21499 13787
rect 22201 13753 22235 13787
rect 23949 13753 23983 13787
rect 6193 13685 6227 13719
rect 7205 13685 7239 13719
rect 9965 13685 9999 13719
rect 10057 13685 10091 13719
rect 10241 13685 10275 13719
rect 14473 13685 14507 13719
rect 17325 13685 17359 13719
rect 18153 13685 18187 13719
rect 19901 13685 19935 13719
rect 3801 13481 3835 13515
rect 4629 13481 4663 13515
rect 9781 13481 9815 13515
rect 11989 13481 12023 13515
rect 14657 13481 14691 13515
rect 17049 13481 17083 13515
rect 21465 13481 21499 13515
rect 21649 13481 21683 13515
rect 23121 13481 23155 13515
rect 24501 13481 24535 13515
rect 8953 13413 8987 13447
rect 12909 13413 12943 13447
rect 14105 13413 14139 13447
rect 4261 13345 4295 13379
rect 4353 13345 4387 13379
rect 5917 13345 5951 13379
rect 7665 13345 7699 13379
rect 10885 13345 10919 13379
rect 11713 13345 11747 13379
rect 12449 13345 12483 13379
rect 13369 13345 13403 13379
rect 13921 13345 13955 13379
rect 17601 13345 17635 13379
rect 17693 13345 17727 13379
rect 18429 13345 18463 13379
rect 18613 13345 18647 13379
rect 20545 13345 20579 13379
rect 21741 13345 21775 13379
rect 23489 13345 23523 13379
rect 24041 13345 24075 13379
rect 24961 13345 24995 13379
rect 25145 13345 25179 13379
rect 2973 13277 3007 13311
rect 4813 13277 4847 13311
rect 5641 13277 5675 13311
rect 5825 13277 5859 13311
rect 6027 13277 6061 13311
rect 6193 13277 6227 13311
rect 6469 13277 6503 13311
rect 6653 13277 6687 13311
rect 6745 13277 6779 13311
rect 6873 13277 6907 13311
rect 7021 13277 7055 13311
rect 7573 13277 7607 13311
rect 9195 13277 9229 13311
rect 9321 13277 9355 13311
rect 9450 13277 9484 13311
rect 9597 13277 9631 13311
rect 9689 13277 9723 13311
rect 9873 13277 9907 13311
rect 10241 13277 10275 13311
rect 10701 13277 10735 13311
rect 10977 13277 11011 13311
rect 11105 13274 11139 13308
rect 11253 13251 11287 13285
rect 11351 13277 11385 13311
rect 11528 13277 11562 13311
rect 11621 13277 11655 13311
rect 11897 13277 11931 13311
rect 12173 13277 12207 13311
rect 12338 13274 12372 13308
rect 12541 13277 12575 13311
rect 12725 13277 12759 13311
rect 13001 13277 13035 13311
rect 13184 13277 13218 13311
rect 13277 13277 13311 13311
rect 13553 13277 13587 13311
rect 14473 13277 14507 13311
rect 14749 13277 14783 13311
rect 17509 13277 17543 13311
rect 18337 13277 18371 13311
rect 20729 13277 20763 13311
rect 20821 13277 20855 13311
rect 21649 13277 21683 13311
rect 21925 13277 21959 13311
rect 22385 13277 22419 13311
rect 22937 13277 22971 13311
rect 23029 13277 23063 13311
rect 23673 13277 23707 13311
rect 24777 13277 24811 13311
rect 25053 13277 25087 13311
rect 2706 13209 2740 13243
rect 4169 13209 4203 13243
rect 7481 13209 7515 13243
rect 14289 13209 14323 13243
rect 22017 13209 22051 13243
rect 22201 13209 22235 13243
rect 23949 13209 23983 13243
rect 24409 13209 24443 13243
rect 1593 13141 1627 13175
rect 5549 13141 5583 13175
rect 6377 13141 6411 13175
rect 7113 13141 7147 13175
rect 10057 13141 10091 13175
rect 10609 13141 10643 13175
rect 13645 13141 13679 13175
rect 14933 13141 14967 13175
rect 17141 13141 17175 13175
rect 17969 13141 18003 13175
rect 20361 13141 20395 13175
rect 21189 13141 21223 13175
rect 23305 13141 23339 13175
rect 3249 12937 3283 12971
rect 3433 12937 3467 12971
rect 3801 12937 3835 12971
rect 6101 12937 6135 12971
rect 7757 12937 7791 12971
rect 9689 12937 9723 12971
rect 9965 12937 9999 12971
rect 11529 12937 11563 12971
rect 11805 12937 11839 12971
rect 16405 12937 16439 12971
rect 18337 12937 18371 12971
rect 20913 12937 20947 12971
rect 21005 12937 21039 12971
rect 21557 12937 21591 12971
rect 22017 12937 22051 12971
rect 23397 12937 23431 12971
rect 23857 12937 23891 12971
rect 24225 12937 24259 12971
rect 2136 12869 2170 12903
rect 3893 12869 3927 12903
rect 8953 12869 8987 12903
rect 11078 12869 11112 12903
rect 4721 12801 4755 12835
rect 4988 12801 5022 12835
rect 6377 12801 6411 12835
rect 6633 12801 6667 12835
rect 9045 12801 9079 12835
rect 9321 12801 9355 12835
rect 9505 12801 9539 12835
rect 11345 12801 11379 12835
rect 11713 12801 11747 12835
rect 24317 12869 24351 12903
rect 11897 12801 11931 12835
rect 12173 12801 12207 12835
rect 12633 12801 12667 12835
rect 14114 12801 14148 12835
rect 14381 12801 14415 12835
rect 15025 12801 15059 12835
rect 15292 12801 15326 12835
rect 18429 12801 18463 12835
rect 21373 12801 21407 12835
rect 21833 12801 21867 12835
rect 22568 12801 22602 12835
rect 1869 12733 1903 12767
rect 4077 12733 4111 12767
rect 11805 12733 11839 12767
rect 17877 12733 17911 12767
rect 19165 12733 19199 12767
rect 20361 12733 20395 12767
rect 21097 12733 21131 12767
rect 22109 12733 22143 12767
rect 22201 12733 22235 12767
rect 23121 12733 23155 12767
rect 23305 12733 23339 12767
rect 24409 12733 24443 12767
rect 9137 12665 9171 12699
rect 12357 12665 12391 12699
rect 13001 12665 13035 12699
rect 12081 12597 12115 12631
rect 12541 12597 12575 12631
rect 20545 12597 20579 12631
rect 22661 12597 22695 12631
rect 22845 12597 22879 12631
rect 23765 12597 23799 12631
rect 10425 12393 10459 12427
rect 12357 12393 12391 12427
rect 20085 12393 20119 12427
rect 22753 12393 22787 12427
rect 9781 12325 9815 12359
rect 10057 12325 10091 12359
rect 12909 12325 12943 12359
rect 17325 12325 17359 12359
rect 18429 12325 18463 12359
rect 20821 12325 20855 12359
rect 9413 12257 9447 12291
rect 11345 12257 11379 12291
rect 15301 12257 15335 12291
rect 15669 12257 15703 12291
rect 16129 12257 16163 12291
rect 17601 12257 17635 12291
rect 18889 12257 18923 12291
rect 19717 12257 19751 12291
rect 19809 12257 19843 12291
rect 20085 12257 20119 12291
rect 20269 12257 20303 12291
rect 21465 12257 21499 12291
rect 24869 12257 24903 12291
rect 24961 12257 24995 12291
rect 6929 12189 6963 12223
rect 8769 12189 8803 12223
rect 9137 12189 9171 12223
rect 9321 12189 9355 12223
rect 9506 12189 9540 12223
rect 9689 12189 9723 12223
rect 9965 12189 9999 12223
rect 10241 12189 10275 12223
rect 11069 12189 11103 12223
rect 11234 12189 11268 12223
rect 11437 12189 11471 12223
rect 11621 12189 11655 12223
rect 12541 12189 12575 12223
rect 12725 12189 12759 12223
rect 13001 12189 13035 12223
rect 14933 12189 14967 12223
rect 15116 12189 15150 12223
rect 15209 12189 15243 12223
rect 15485 12189 15519 12223
rect 16037 12189 16071 12223
rect 16496 12189 16530 12223
rect 16957 12189 16991 12223
rect 17969 12189 18003 12223
rect 18153 12189 18187 12223
rect 18521 12189 18555 12223
rect 18613 12189 18647 12223
rect 20177 12189 20211 12223
rect 20636 12189 20670 12223
rect 22109 12189 22143 12223
rect 22569 12189 22603 12223
rect 24777 12189 24811 12223
rect 16773 12121 16807 12155
rect 17141 12121 17175 12155
rect 21741 12121 21775 12155
rect 21925 12121 21959 12155
rect 7021 12053 7055 12087
rect 8585 12053 8619 12087
rect 9045 12053 9079 12087
rect 10885 12053 10919 12087
rect 11713 12053 11747 12087
rect 13185 12053 13219 12087
rect 16589 12053 16623 12087
rect 18705 12053 18739 12087
rect 19257 12053 19291 12087
rect 19625 12053 19659 12087
rect 20913 12053 20947 12087
rect 21281 12053 21315 12087
rect 21373 12053 21407 12087
rect 22201 12053 22235 12087
rect 23673 12053 23707 12087
rect 24133 12053 24167 12087
rect 24409 12053 24443 12087
rect 3249 11849 3283 11883
rect 10701 11849 10735 11883
rect 16865 11849 16899 11883
rect 17325 11849 17359 11883
rect 17785 11849 17819 11883
rect 18153 11849 18187 11883
rect 18889 11849 18923 11883
rect 19349 11849 19383 11883
rect 19809 11849 19843 11883
rect 20637 11849 20671 11883
rect 21189 11849 21223 11883
rect 21833 11849 21867 11883
rect 22293 11849 22327 11883
rect 23305 11849 23339 11883
rect 24133 11849 24167 11883
rect 5181 11781 5215 11815
rect 5365 11781 5399 11815
rect 9045 11781 9079 11815
rect 17417 11781 17451 11815
rect 18245 11781 18279 11815
rect 19441 11781 19475 11815
rect 20361 11781 20395 11815
rect 21281 11781 21315 11815
rect 22201 11781 22235 11815
rect 24225 11781 24259 11815
rect 2697 11713 2731 11747
rect 2973 11713 3007 11747
rect 3157 11713 3191 11747
rect 6561 11713 6595 11747
rect 7941 11713 7975 11747
rect 8106 11713 8140 11747
rect 8217 11713 8251 11747
rect 8493 11713 8527 11747
rect 9229 11713 9263 11747
rect 9321 11713 9355 11747
rect 9577 11713 9611 11747
rect 11796 11713 11830 11747
rect 15292 11713 15326 11747
rect 16681 11713 16715 11747
rect 18613 11713 18647 11747
rect 18797 11713 18831 11747
rect 19901 11713 19935 11747
rect 20085 11713 20119 11747
rect 20453 11713 20487 11747
rect 2789 11645 2823 11679
rect 8309 11645 8343 11679
rect 11529 11645 11563 11679
rect 15025 11645 15059 11679
rect 17509 11645 17543 11679
rect 18337 11645 18371 11679
rect 19165 11645 19199 11679
rect 21465 11645 21499 11679
rect 22385 11645 22419 11679
rect 22753 11645 22787 11679
rect 23397 11645 23431 11679
rect 23489 11645 23523 11679
rect 24317 11645 24351 11679
rect 2881 11577 2915 11611
rect 2513 11509 2547 11543
rect 6377 11509 6411 11543
rect 7757 11509 7791 11543
rect 8585 11509 8619 11543
rect 12909 11509 12943 11543
rect 14473 11509 14507 11543
rect 16405 11509 16439 11543
rect 16957 11509 16991 11543
rect 20821 11509 20855 11543
rect 22937 11509 22971 11543
rect 23765 11509 23799 11543
rect 1777 11305 1811 11339
rect 8493 11305 8527 11339
rect 8769 11305 8803 11339
rect 10333 11305 10367 11339
rect 15669 11305 15703 11339
rect 18337 11305 18371 11339
rect 18705 11305 18739 11339
rect 21005 11305 21039 11339
rect 22661 11305 22695 11339
rect 6745 11237 6779 11271
rect 8309 11237 8343 11271
rect 5365 11169 5399 11203
rect 13829 11237 13863 11271
rect 14473 11237 14507 11271
rect 17049 11237 17083 11271
rect 18981 11237 19015 11271
rect 19257 11237 19291 11271
rect 24409 11237 24443 11271
rect 8953 11169 8987 11203
rect 12541 11169 12575 11203
rect 12633 11169 12667 11203
rect 13369 11169 13403 11203
rect 15393 11169 15427 11203
rect 16405 11169 16439 11203
rect 17693 11169 17727 11203
rect 19809 11169 19843 11203
rect 20821 11169 20855 11203
rect 21465 11169 21499 11203
rect 21557 11169 21591 11203
rect 21833 11169 21867 11203
rect 23397 11169 23431 11203
rect 23673 11169 23707 11203
rect 24133 11169 24167 11203
rect 24869 11169 24903 11203
rect 24961 11169 24995 11203
rect 3157 11101 3191 11135
rect 3341 11101 3375 11135
rect 3525 11101 3559 11135
rect 3801 11101 3835 11135
rect 6929 11101 6963 11135
rect 8493 11101 8527 11135
rect 8585 11101 8619 11135
rect 9209 11101 9243 11135
rect 12357 11101 12391 11135
rect 12726 11101 12760 11135
rect 12909 11101 12943 11135
rect 13001 11101 13035 11135
rect 13184 11101 13218 11135
rect 13277 11101 13311 11135
rect 13507 11101 13541 11135
rect 15025 11101 15059 11135
rect 15208 11101 15242 11135
rect 15301 11101 15335 11135
rect 15577 11101 15611 11135
rect 16221 11101 16255 11135
rect 16589 11101 16623 11135
rect 16681 11101 16715 11135
rect 17509 11101 17543 11135
rect 18337 11101 18371 11135
rect 18429 11101 18463 11135
rect 19625 11101 19659 11135
rect 21373 11101 21407 11135
rect 23213 11101 23247 11135
rect 23305 11101 23339 11135
rect 2912 11033 2946 11067
rect 3249 11033 3283 11067
rect 5089 11033 5123 11067
rect 5632 11033 5666 11067
rect 7174 11033 7208 11067
rect 12173 11033 12207 11067
rect 13737 11033 13771 11067
rect 14105 11033 14139 11067
rect 14289 11033 14323 11067
rect 14657 11033 14691 11067
rect 14841 11033 14875 11067
rect 17601 11033 17635 11067
rect 19717 11033 19751 11067
rect 17141 10965 17175 10999
rect 22845 10965 22879 10999
rect 24777 10965 24811 10999
rect 5273 10761 5307 10795
rect 7205 10761 7239 10795
rect 10793 10761 10827 10795
rect 15853 10761 15887 10795
rect 17049 10761 17083 10795
rect 18797 10761 18831 10795
rect 19349 10761 19383 10795
rect 23765 10761 23799 10795
rect 24225 10761 24259 10795
rect 2136 10693 2170 10727
rect 3525 10693 3559 10727
rect 5089 10693 5123 10727
rect 13194 10693 13228 10727
rect 14758 10693 14792 10727
rect 19257 10693 19291 10727
rect 23397 10693 23431 10727
rect 23857 10693 23891 10727
rect 3433 10625 3467 10659
rect 3801 10625 3835 10659
rect 4077 10625 4111 10659
rect 4353 10625 4387 10659
rect 4536 10625 4570 10659
rect 4629 10625 4663 10659
rect 4905 10625 4939 10659
rect 5365 10625 5399 10659
rect 5734 10625 5768 10659
rect 5917 10625 5951 10659
rect 6561 10625 6595 10659
rect 7297 10625 7331 10659
rect 7573 10625 7607 10659
rect 7849 10625 7883 10659
rect 8116 10625 8150 10659
rect 9413 10625 9447 10659
rect 9680 10625 9714 10659
rect 13461 10625 13495 10659
rect 15117 10625 15151 10659
rect 15519 10625 15553 10659
rect 15761 10625 15795 10659
rect 16037 10625 16071 10659
rect 1869 10557 1903 10591
rect 3617 10557 3651 10591
rect 4721 10557 4755 10591
rect 5549 10557 5583 10591
rect 5641 10557 5675 10591
rect 6101 10557 6135 10591
rect 6193 10557 6227 10591
rect 15025 10557 15059 10591
rect 15209 10557 15243 10591
rect 19073 10557 19107 10591
rect 23581 10557 23615 10591
rect 4169 10489 4203 10523
rect 6377 10489 6411 10523
rect 3249 10421 3283 10455
rect 6193 10421 6227 10455
rect 9229 10421 9263 10455
rect 12081 10421 12115 10455
rect 13645 10421 13679 10455
rect 19717 10421 19751 10455
rect 2421 10217 2455 10251
rect 8033 10217 8067 10251
rect 8769 10217 8803 10251
rect 9597 10217 9631 10251
rect 13553 10217 13587 10251
rect 13921 10217 13955 10251
rect 15209 10217 15243 10251
rect 3249 10149 3283 10183
rect 2697 10081 2731 10115
rect 2789 10081 2823 10115
rect 2881 10081 2915 10115
rect 3525 10081 3559 10115
rect 4353 10081 4387 10115
rect 4813 10081 4847 10115
rect 8309 10081 8343 10115
rect 2605 10013 2639 10047
rect 3065 10013 3099 10047
rect 3341 10013 3375 10047
rect 3617 10013 3651 10047
rect 3985 10013 4019 10047
rect 4150 10013 4184 10047
rect 4261 10013 4295 10047
rect 4537 10013 4571 10047
rect 6377 10013 6411 10047
rect 8125 10013 8159 10047
rect 8401 10013 8435 10047
rect 8494 10013 8528 10047
rect 8677 10013 8711 10047
rect 4721 9945 4755 9979
rect 5058 9945 5092 9979
rect 6622 9945 6656 9979
rect 23121 10149 23155 10183
rect 9321 10081 9355 10115
rect 9873 10081 9907 10115
rect 14197 10081 14231 10115
rect 21465 10081 21499 10115
rect 8953 10013 8987 10047
rect 9136 10013 9170 10047
rect 9229 10013 9263 10047
rect 9505 10013 9539 10047
rect 13737 10013 13771 10047
rect 14105 10013 14139 10047
rect 14564 10013 14598 10047
rect 14933 10013 14967 10047
rect 20729 10013 20763 10047
rect 21189 10013 21223 10047
rect 24594 10013 24628 10047
rect 24961 10013 24995 10047
rect 25053 10013 25087 10047
rect 14749 9945 14783 9979
rect 15117 9945 15151 9979
rect 22845 9945 22879 9979
rect 24409 9945 24443 9979
rect 3801 9877 3835 9911
rect 6193 9877 6227 9911
rect 7757 9877 7791 9911
rect 8769 9877 8803 9911
rect 20545 9877 20579 9911
rect 20821 9877 20855 9911
rect 21281 9877 21315 9911
rect 23305 9877 23339 9911
rect 3341 9673 3375 9707
rect 5641 9673 5675 9707
rect 13185 9673 13219 9707
rect 14565 9673 14599 9707
rect 15393 9673 15427 9707
rect 22845 9673 22879 9707
rect 25053 9673 25087 9707
rect 5457 9605 5491 9639
rect 17969 9605 18003 9639
rect 20821 9605 20855 9639
rect 21649 9605 21683 9639
rect 23305 9605 23339 9639
rect 25421 9605 25455 9639
rect 2513 9537 2547 9571
rect 2697 9537 2731 9571
rect 2881 9537 2915 9571
rect 3157 9537 3191 9571
rect 3709 9537 3743 9571
rect 4721 9537 4755 9571
rect 4904 9537 4938 9571
rect 5089 9537 5123 9571
rect 5273 9537 5307 9571
rect 8033 9537 8067 9571
rect 8309 9537 8343 9571
rect 9689 9537 9723 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 13277 9537 13311 9571
rect 14657 9537 14691 9571
rect 15485 9537 15519 9571
rect 17325 9537 17359 9571
rect 21465 9537 21499 9571
rect 23213 9537 23247 9571
rect 23929 9537 23963 9571
rect 25605 9537 25639 9571
rect 2237 9469 2271 9503
rect 3617 9469 3651 9503
rect 4997 9469 5031 9503
rect 8401 9469 8435 9503
rect 13829 9469 13863 9503
rect 14105 9469 14139 9503
rect 14841 9469 14875 9503
rect 15669 9469 15703 9503
rect 18061 9469 18095 9503
rect 18153 9469 18187 9503
rect 19809 9469 19843 9503
rect 20913 9469 20947 9503
rect 21097 9469 21131 9503
rect 23397 9469 23431 9503
rect 23673 9469 23707 9503
rect 2421 9401 2455 9435
rect 3065 9401 3099 9435
rect 7849 9401 7883 9435
rect 9873 9401 9907 9435
rect 10241 9401 10275 9435
rect 13369 9401 13403 9435
rect 17601 9401 17635 9435
rect 20177 9401 20211 9435
rect 20453 9401 20487 9435
rect 25237 9401 25271 9435
rect 2053 9333 2087 9367
rect 3709 9333 3743 9367
rect 4537 9333 4571 9367
rect 8125 9333 8159 9367
rect 9965 9333 9999 9367
rect 11621 9333 11655 9367
rect 14197 9333 14231 9367
rect 15025 9333 15059 9367
rect 17509 9333 17543 9367
rect 20269 9333 20303 9367
rect 21373 9333 21407 9367
rect 3801 9129 3835 9163
rect 4261 9129 4295 9163
rect 12725 9129 12759 9163
rect 13645 9129 13679 9163
rect 13737 9129 13771 9163
rect 20085 9129 20119 9163
rect 23397 9129 23431 9163
rect 3065 9061 3099 9095
rect 10609 9061 10643 9095
rect 14841 9061 14875 9095
rect 22109 9061 22143 9095
rect 22293 9061 22327 9095
rect 1685 8993 1719 9027
rect 3893 8993 3927 9027
rect 12817 8993 12851 9027
rect 12909 8993 12943 9027
rect 13737 8993 13771 9027
rect 13829 8993 13863 9027
rect 14197 8993 14231 9027
rect 14381 8993 14415 9027
rect 15117 8993 15151 9027
rect 18705 8993 18739 9027
rect 19809 8993 19843 9027
rect 20545 8993 20579 9027
rect 22845 8993 22879 9027
rect 24041 8993 24075 9027
rect 24961 8993 24995 9027
rect 1952 8925 1986 8959
rect 3801 8925 3835 8959
rect 4077 8925 4111 8959
rect 7297 8925 7331 8959
rect 9137 8925 9171 8959
rect 9321 8925 9355 8959
rect 10241 8925 10275 8959
rect 11989 8925 12023 8959
rect 12265 8925 12299 8959
rect 13093 8925 13127 8959
rect 13185 8925 13219 8959
rect 14473 8925 14507 8959
rect 16405 8925 16439 8959
rect 18521 8925 18555 8959
rect 19499 8925 19533 8959
rect 19901 8925 19935 8959
rect 20235 8925 20269 8959
rect 20637 8925 20671 8959
rect 20729 8925 20763 8959
rect 22478 8925 22512 8959
rect 22937 8925 22971 8959
rect 23213 8925 23247 8959
rect 23857 8925 23891 8959
rect 24651 8925 24685 8959
rect 25053 8925 25087 8959
rect 25145 8925 25179 8959
rect 25329 8925 25363 8959
rect 7564 8857 7598 8891
rect 8953 8857 8987 8891
rect 9873 8857 9907 8891
rect 10057 8857 10091 8891
rect 11722 8857 11756 8891
rect 15301 8857 15335 8891
rect 16650 8857 16684 8891
rect 18613 8857 18647 8891
rect 19257 8857 19291 8891
rect 20996 8857 21030 8891
rect 23949 8857 23983 8891
rect 24409 8857 24443 8891
rect 25513 8857 25547 8891
rect 8677 8789 8711 8823
rect 12081 8789 12115 8823
rect 12541 8789 12575 8823
rect 13369 8789 13403 8823
rect 15209 8789 15243 8823
rect 15669 8789 15703 8823
rect 17785 8789 17819 8823
rect 18153 8789 18187 8823
rect 23489 8789 23523 8823
rect 2605 8585 2639 8619
rect 6101 8585 6135 8619
rect 7113 8585 7147 8619
rect 8033 8585 8067 8619
rect 9045 8585 9079 8619
rect 11161 8585 11195 8619
rect 11621 8585 11655 8619
rect 12817 8585 12851 8619
rect 13369 8585 13403 8619
rect 14013 8585 14047 8619
rect 14105 8585 14139 8619
rect 15025 8585 15059 8619
rect 15853 8585 15887 8619
rect 16037 8585 16071 8619
rect 17049 8585 17083 8619
rect 17877 8585 17911 8619
rect 19441 8585 19475 8619
rect 21557 8585 21591 8619
rect 25237 8585 25271 8619
rect 7665 8517 7699 8551
rect 11897 8517 11931 8551
rect 13277 8517 13311 8551
rect 14933 8517 14967 8551
rect 20444 8517 20478 8551
rect 21833 8517 21867 8551
rect 22017 8517 22051 8551
rect 22201 8517 22235 8551
rect 2789 8449 2823 8483
rect 3065 8449 3099 8483
rect 3157 8449 3191 8483
rect 3249 8449 3283 8483
rect 3893 8449 3927 8483
rect 5273 8449 5307 8483
rect 5456 8452 5490 8486
rect 5825 8449 5859 8483
rect 6837 8449 6871 8483
rect 7297 8449 7331 8483
rect 8125 8449 8159 8483
rect 8494 8449 8528 8483
rect 8677 8449 8711 8483
rect 8953 8449 8987 8483
rect 10793 8449 10827 8483
rect 11069 8449 11103 8483
rect 12311 8449 12345 8483
rect 12437 8449 12471 8483
rect 12633 8449 12667 8483
rect 15669 8449 15703 8483
rect 17693 8449 17727 8483
rect 18990 8449 19024 8483
rect 19534 8449 19568 8483
rect 20177 8449 20211 8483
rect 23857 8449 23891 8483
rect 24113 8449 24147 8483
rect 5549 8381 5583 8415
rect 5641 8381 5675 8415
rect 8309 8381 8343 8415
rect 8401 8381 8435 8415
rect 10241 8381 10275 8415
rect 10885 8381 10919 8415
rect 11805 8381 11839 8415
rect 12081 8381 12115 8415
rect 13185 8381 13219 8415
rect 16497 8381 16531 8415
rect 17141 8381 17175 8415
rect 17233 8381 17267 8415
rect 19257 8381 19291 8415
rect 19901 8381 19935 8415
rect 19993 8381 20027 8415
rect 23029 8381 23063 8415
rect 2973 8313 3007 8347
rect 3709 8313 3743 8347
rect 6009 8313 6043 8347
rect 6929 8313 6963 8347
rect 7481 8313 7515 8347
rect 8769 8313 8803 8347
rect 10517 8313 10551 8347
rect 12173 8313 12207 8347
rect 13737 8313 13771 8347
rect 16221 8313 16255 8347
rect 16681 8313 16715 8347
rect 17509 8313 17543 8347
rect 23397 8313 23431 8347
rect 3157 8245 3191 8279
rect 3525 8245 3559 8279
rect 12541 8245 12575 8279
rect 23489 8245 23523 8279
rect 2973 8041 3007 8075
rect 6469 8041 6503 8075
rect 6745 8041 6779 8075
rect 8769 8041 8803 8075
rect 9873 8041 9907 8075
rect 16313 8041 16347 8075
rect 17325 8041 17359 8075
rect 19533 8041 19567 8075
rect 19901 8041 19935 8075
rect 21097 8041 21131 8075
rect 23857 8041 23891 8075
rect 4353 7905 4387 7939
rect 4445 7905 4479 7939
rect 7297 7905 7331 7939
rect 7389 7905 7423 7939
rect 8217 7905 8251 7939
rect 11713 7973 11747 8007
rect 14197 7973 14231 8007
rect 17233 7973 17267 8007
rect 18889 7973 18923 8007
rect 20821 7973 20855 8007
rect 9321 7905 9355 7939
rect 11897 7905 11931 7939
rect 12357 7905 12391 7939
rect 13369 7905 13403 7939
rect 13921 7905 13955 7939
rect 17509 7905 17543 7939
rect 19625 7905 19659 7939
rect 1593 7837 1627 7871
rect 3341 7837 3375 7871
rect 4077 7837 4111 7871
rect 4242 7837 4276 7871
rect 4629 7837 4663 7871
rect 6377 7837 6411 7871
rect 6653 7837 6687 7871
rect 6929 7837 6963 7871
rect 7021 7837 7055 7871
rect 7204 7837 7238 7871
rect 7573 7837 7607 7871
rect 7849 7837 7883 7871
rect 8032 7837 8066 7871
rect 8125 7837 8159 7871
rect 8401 7837 8435 7871
rect 8769 7837 8803 7871
rect 8953 7837 8987 7871
rect 9136 7837 9170 7871
rect 9229 7837 9263 7871
rect 9505 7837 9539 7871
rect 10333 7837 10367 7871
rect 10600 7837 10634 7871
rect 12081 7837 12115 7871
rect 12449 7837 12483 7871
rect 12909 7837 12943 7871
rect 13553 7837 13587 7871
rect 15577 7837 15611 7871
rect 16497 7837 16531 7871
rect 16681 7837 16715 7871
rect 19717 7837 19751 7871
rect 19993 7837 20027 7871
rect 20177 7837 20211 7871
rect 21281 7837 21315 7871
rect 23305 7837 23339 7871
rect 23673 7837 23707 7871
rect 1860 7769 1894 7803
rect 6110 7769 6144 7803
rect 7757 7769 7791 7803
rect 12541 7769 12575 7803
rect 13093 7769 13127 7803
rect 15310 7769 15344 7803
rect 16773 7769 16807 7803
rect 16865 7769 16899 7803
rect 17754 7769 17788 7803
rect 20453 7769 20487 7803
rect 3249 7701 3283 7735
rect 3893 7701 3927 7735
rect 4721 7701 4755 7735
rect 4997 7701 5031 7735
rect 8493 7701 8527 7735
rect 9597 7701 9631 7735
rect 12725 7701 12759 7735
rect 12817 7701 12851 7735
rect 13185 7701 13219 7735
rect 13829 7701 13863 7735
rect 19349 7701 19383 7735
rect 20913 7701 20947 7735
rect 23121 7701 23155 7735
rect 2145 7497 2179 7531
rect 5733 7497 5767 7531
rect 11621 7497 11655 7531
rect 12541 7497 12575 7531
rect 13461 7497 13495 7531
rect 13553 7497 13587 7531
rect 14013 7497 14047 7531
rect 18613 7497 18647 7531
rect 19901 7497 19935 7531
rect 22845 7497 22879 7531
rect 23673 7497 23707 7531
rect 3433 7429 3467 7463
rect 4620 7429 4654 7463
rect 11253 7429 11287 7463
rect 14197 7429 14231 7463
rect 17141 7429 17175 7463
rect 17877 7429 17911 7463
rect 2237 7361 2271 7395
rect 2329 7361 2363 7395
rect 2789 7361 2823 7395
rect 2881 7361 2915 7395
rect 3157 7361 3191 7395
rect 3249 7361 3283 7395
rect 4353 7361 4387 7395
rect 7582 7361 7616 7395
rect 9514 7361 9548 7395
rect 11161 7361 11195 7395
rect 11713 7361 11747 7395
rect 12449 7361 12483 7395
rect 12909 7361 12943 7395
rect 13277 7361 13311 7395
rect 13737 7361 13771 7395
rect 13921 7361 13955 7395
rect 16681 7361 16715 7395
rect 16957 7361 16991 7395
rect 2605 7293 2639 7327
rect 7849 7293 7883 7327
rect 9781 7293 9815 7327
rect 12679 7293 12713 7327
rect 17233 7293 17267 7327
rect 17969 7361 18003 7395
rect 18153 7361 18187 7395
rect 18337 7361 18371 7395
rect 18429 7361 18463 7395
rect 19349 7361 19383 7395
rect 19717 7361 19751 7395
rect 20545 7361 20579 7395
rect 22937 7361 22971 7395
rect 24225 7361 24259 7395
rect 24409 7361 24443 7395
rect 23121 7293 23155 7327
rect 23765 7293 23799 7327
rect 23857 7293 23891 7327
rect 3065 7225 3099 7259
rect 3617 7225 3651 7259
rect 13093 7225 13127 7259
rect 17601 7225 17635 7259
rect 17693 7225 17727 7259
rect 17877 7225 17911 7259
rect 19533 7225 19567 7259
rect 1869 7157 1903 7191
rect 5917 7157 5951 7191
rect 6469 7157 6503 7191
rect 8401 7157 8435 7191
rect 12081 7157 12115 7191
rect 20361 7157 20395 7191
rect 22477 7157 22511 7191
rect 23305 7157 23339 7191
rect 24501 7157 24535 7191
rect 12173 6953 12207 6987
rect 20361 6953 20395 6987
rect 24961 6953 24995 6987
rect 13369 6885 13403 6919
rect 13553 6885 13587 6919
rect 20177 6885 20211 6919
rect 22477 6885 22511 6919
rect 24133 6885 24167 6919
rect 4537 6817 4571 6851
rect 6469 6817 6503 6851
rect 6837 6817 6871 6851
rect 8033 6817 8067 6851
rect 15485 6817 15519 6851
rect 16313 6817 16347 6851
rect 22753 6817 22787 6851
rect 24501 6817 24535 6851
rect 6101 6749 6135 6783
rect 6266 6749 6300 6783
rect 6377 6749 6411 6783
rect 6653 6749 6687 6783
rect 7849 6749 7883 6783
rect 10158 6749 10192 6783
rect 10425 6749 10459 6783
rect 12081 6749 12115 6783
rect 13185 6749 13219 6783
rect 13277 6749 13311 6783
rect 14657 6749 14691 6783
rect 15301 6749 15335 6783
rect 16129 6749 16163 6783
rect 16773 6749 16807 6783
rect 20971 6749 21005 6783
rect 21281 6749 21315 6783
rect 21373 6749 21407 6783
rect 23020 6749 23054 6783
rect 24409 6749 24443 6783
rect 24868 6749 24902 6783
rect 4804 6681 4838 6715
rect 16589 6681 16623 6715
rect 19901 6681 19935 6715
rect 22109 6681 22143 6715
rect 5917 6613 5951 6647
rect 7757 6613 7791 6647
rect 9045 6613 9079 6647
rect 13001 6613 13035 6647
rect 14841 6613 14875 6647
rect 14933 6613 14967 6647
rect 15393 6613 15427 6647
rect 15761 6613 15795 6647
rect 16221 6613 16255 6647
rect 20821 6613 20855 6647
rect 22569 6613 22603 6647
rect 3341 6409 3375 6443
rect 4169 6409 4203 6443
rect 4629 6409 4663 6443
rect 5549 6409 5583 6443
rect 9413 6409 9447 6443
rect 14197 6409 14231 6443
rect 16773 6409 16807 6443
rect 18981 6409 19015 6443
rect 19441 6409 19475 6443
rect 20361 6409 20395 6443
rect 20821 6409 20855 6443
rect 22109 6409 22143 6443
rect 24317 6409 24351 6443
rect 1869 6341 1903 6375
rect 3893 6341 3927 6375
rect 1961 6273 1995 6307
rect 2145 6273 2179 6307
rect 2697 6273 2731 6307
rect 2881 6273 2915 6307
rect 3065 6273 3099 6307
rect 3341 6273 3375 6307
rect 3985 6273 4019 6307
rect 3249 6205 3283 6239
rect 2697 6137 2731 6171
rect 4721 6341 4755 6375
rect 8300 6341 8334 6375
rect 20085 6341 20119 6375
rect 20729 6341 20763 6375
rect 21373 6341 21407 6375
rect 21557 6341 21591 6375
rect 22446 6341 22480 6375
rect 4905 6273 4939 6307
rect 5070 6273 5104 6307
rect 5181 6273 5215 6307
rect 5457 6273 5491 6307
rect 5917 6273 5951 6307
rect 11621 6273 11655 6307
rect 11989 6273 12023 6307
rect 12173 6273 12207 6307
rect 14749 6273 14783 6307
rect 15005 6273 15039 6307
rect 16497 6273 16531 6307
rect 16866 6273 16900 6307
rect 18797 6273 18831 6307
rect 19901 6273 19935 6307
rect 21189 6273 21223 6307
rect 21925 6273 21959 6307
rect 22201 6273 22235 6307
rect 24167 6273 24201 6307
rect 5273 6205 5307 6239
rect 8033 6205 8067 6239
rect 14657 6205 14691 6239
rect 17233 6205 17267 6239
rect 17325 6205 17359 6239
rect 19533 6205 19567 6239
rect 19625 6205 19659 6239
rect 20913 6205 20947 6239
rect 23765 6205 23799 6239
rect 23857 6205 23891 6239
rect 5733 6137 5767 6171
rect 14381 6137 14415 6171
rect 16129 6137 16163 6171
rect 2329 6069 2363 6103
rect 4629 6069 4663 6103
rect 11805 6069 11839 6103
rect 12173 6069 12207 6103
rect 16313 6069 16347 6103
rect 19073 6069 19107 6103
rect 20177 6069 20211 6103
rect 23581 6069 23615 6103
rect 3157 5865 3191 5899
rect 8677 5865 8711 5899
rect 12725 5865 12759 5899
rect 15209 5865 15243 5899
rect 19349 5865 19383 5899
rect 21373 5865 21407 5899
rect 22385 5865 22419 5899
rect 11713 5797 11747 5831
rect 18613 5797 18647 5831
rect 18797 5797 18831 5831
rect 22293 5797 22327 5831
rect 23673 5797 23707 5831
rect 2973 5729 3007 5763
rect 12265 5729 12299 5763
rect 15669 5729 15703 5763
rect 15761 5729 15795 5763
rect 19993 5729 20027 5763
rect 21925 5729 21959 5763
rect 2706 5661 2740 5695
rect 5457 5661 5491 5695
rect 8217 5661 8251 5695
rect 8401 5661 8435 5695
rect 8493 5661 8527 5695
rect 8769 5661 8803 5695
rect 11437 5661 11471 5695
rect 12081 5661 12115 5695
rect 12909 5661 12943 5695
rect 13001 5661 13035 5695
rect 14841 5661 14875 5695
rect 15359 5661 15393 5695
rect 15853 5661 15887 5695
rect 17785 5661 17819 5695
rect 18245 5661 18279 5695
rect 19073 5661 19107 5695
rect 19499 5661 19533 5695
rect 19809 5661 19843 5695
rect 19901 5661 19935 5695
rect 20260 5661 20294 5695
rect 23305 5661 23339 5695
rect 23489 5661 23523 5695
rect 9229 5593 9263 5627
rect 9413 5593 9447 5627
rect 12173 5593 12207 5627
rect 13093 5593 13127 5627
rect 16120 5593 16154 5627
rect 17417 5593 17451 5627
rect 17601 5593 17635 5627
rect 1593 5525 1627 5559
rect 5273 5525 5307 5559
rect 5917 5525 5951 5559
rect 11621 5525 11655 5559
rect 14657 5525 14691 5559
rect 17233 5525 17267 5559
rect 18429 5525 18463 5559
rect 2789 5321 2823 5355
rect 4997 5321 5031 5355
rect 9321 5321 9355 5355
rect 9873 5321 9907 5355
rect 11253 5321 11287 5355
rect 15669 5321 15703 5355
rect 16405 5321 16439 5355
rect 17141 5321 17175 5355
rect 17233 5321 17267 5355
rect 20269 5321 20303 5355
rect 4629 5253 4663 5287
rect 4721 5253 4755 5287
rect 5365 5253 5399 5287
rect 8208 5253 8242 5287
rect 9965 5253 9999 5287
rect 10793 5253 10827 5287
rect 11774 5253 11808 5287
rect 13277 5253 13311 5287
rect 19134 5253 19168 5287
rect 3902 5185 3936 5219
rect 4169 5185 4203 5219
rect 4532 5185 4566 5219
rect 4905 5185 4939 5219
rect 6009 5185 6043 5219
rect 6377 5185 6411 5219
rect 6644 5185 6678 5219
rect 7941 5185 7975 5219
rect 11529 5185 11563 5219
rect 13093 5185 13127 5219
rect 16037 5185 16071 5219
rect 16221 5185 16255 5219
rect 17601 5185 17635 5219
rect 17877 5185 17911 5219
rect 5457 5117 5491 5151
rect 5641 5117 5675 5151
rect 10149 5117 10183 5151
rect 15209 5117 15243 5151
rect 17325 5117 17359 5151
rect 17693 5117 17727 5151
rect 18889 5117 18923 5151
rect 11161 5049 11195 5083
rect 13461 5049 13495 5083
rect 15577 5049 15611 5083
rect 4353 4981 4387 5015
rect 5825 4981 5859 5015
rect 6193 4981 6227 5015
rect 7757 4981 7791 5015
rect 9505 4981 9539 5015
rect 10425 4981 10459 5015
rect 12909 4981 12943 5015
rect 16221 4981 16255 5015
rect 16773 4981 16807 5015
rect 17601 4981 17635 5015
rect 18061 4981 18095 5015
rect 5273 4777 5307 4811
rect 6377 4777 6411 4811
rect 6837 4777 6871 4811
rect 7849 4777 7883 4811
rect 8769 4777 8803 4811
rect 10609 4777 10643 4811
rect 14105 4777 14139 4811
rect 17601 4777 17635 4811
rect 9045 4709 9079 4743
rect 11069 4709 11103 4743
rect 11345 4709 11379 4743
rect 16129 4709 16163 4743
rect 16957 4709 16991 4743
rect 3893 4641 3927 4675
rect 5917 4641 5951 4675
rect 6101 4641 6135 4675
rect 7941 4641 7975 4675
rect 8217 4641 8251 4675
rect 8309 4641 8343 4675
rect 10701 4641 10735 4675
rect 11989 4641 12023 4675
rect 12725 4641 12759 4675
rect 13553 4641 13587 4675
rect 15393 4641 15427 4675
rect 17049 4641 17083 4675
rect 2053 4573 2087 4607
rect 6285 4573 6319 4607
rect 6561 4573 6595 4607
rect 6653 4573 6687 4607
rect 7021 4573 7055 4607
rect 7573 4573 7607 4607
rect 7665 4573 7699 4607
rect 8401 4573 8435 4607
rect 10425 4573 10459 4607
rect 11713 4573 11747 4607
rect 12541 4573 12575 4607
rect 13369 4573 13403 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 15209 4573 15243 4607
rect 17141 4573 17175 4607
rect 17508 4573 17542 4607
rect 4160 4505 4194 4539
rect 7389 4505 7423 4539
rect 10158 4505 10192 4539
rect 12633 4505 12667 4539
rect 15761 4505 15795 4539
rect 16589 4505 16623 4539
rect 16773 4505 16807 4539
rect 5457 4437 5491 4471
rect 5825 4437 5859 4471
rect 7113 4437 7147 4471
rect 11161 4437 11195 4471
rect 11805 4437 11839 4471
rect 12173 4437 12207 4471
rect 13001 4437 13035 4471
rect 13461 4437 13495 4471
rect 14473 4437 14507 4471
rect 14841 4437 14875 4471
rect 15301 4437 15335 4471
rect 16221 4437 16255 4471
rect 4813 4233 4847 4267
rect 5917 4233 5951 4267
rect 7757 4233 7791 4267
rect 9229 4233 9263 4267
rect 9781 4233 9815 4267
rect 9965 4233 9999 4267
rect 14289 4233 14323 4267
rect 6745 4165 6779 4199
rect 10701 4165 10735 4199
rect 10793 4165 10827 4199
rect 12081 4165 12115 4199
rect 15209 4165 15243 4199
rect 15761 4165 15795 4199
rect 16865 4165 16899 4199
rect 4997 4097 5031 4131
rect 5089 4097 5123 4131
rect 5365 4097 5399 4131
rect 5825 4097 5859 4131
rect 7205 4097 7239 4131
rect 7941 4097 7975 4131
rect 8401 4097 8435 4131
rect 9321 4097 9355 4131
rect 11529 4097 11563 4131
rect 12323 4097 12357 4131
rect 12633 4097 12667 4131
rect 12725 4097 12759 4131
rect 13176 4097 13210 4131
rect 14473 4097 14507 4131
rect 14715 4097 14749 4131
rect 15025 4097 15059 4131
rect 15393 4097 15427 4131
rect 16003 4097 16037 4131
rect 16313 4097 16347 4131
rect 16681 4097 16715 4131
rect 17141 4097 17175 4131
rect 22017 4097 22051 4131
rect 22284 4097 22318 4131
rect 5273 4029 5307 4063
rect 6009 4029 6043 4063
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 7573 4029 7607 4063
rect 8493 4029 8527 4063
rect 8677 4029 8711 4063
rect 9505 4029 9539 4063
rect 12909 4029 12943 4063
rect 15117 4029 15151 4063
rect 16405 4029 16439 4063
rect 7389 3961 7423 3995
rect 10425 3961 10459 3995
rect 11161 3961 11195 3995
rect 15577 3961 15611 3995
rect 23397 3961 23431 3995
rect 5457 3893 5491 3927
rect 6377 3893 6411 3927
rect 8033 3893 8067 3927
rect 8861 3893 8895 3927
rect 10241 3893 10275 3927
rect 11253 3893 11287 3927
rect 11713 3893 11747 3927
rect 16957 3893 16991 3927
rect 17325 3893 17359 3927
rect 5825 3689 5859 3723
rect 7665 3689 7699 3723
rect 11897 3689 11931 3723
rect 13737 3689 13771 3723
rect 22293 3689 22327 3723
rect 2145 3621 2179 3655
rect 9045 3621 9079 3655
rect 14105 3621 14139 3655
rect 16497 3621 16531 3655
rect 16773 3621 16807 3655
rect 4445 3553 4479 3587
rect 7481 3553 7515 3587
rect 8125 3553 8159 3587
rect 8217 3553 8251 3587
rect 15117 3553 15151 3587
rect 18153 3553 18187 3587
rect 2329 3485 2363 3519
rect 2513 3485 2547 3519
rect 8401 3485 8435 3519
rect 8493 3485 8527 3519
rect 10425 3485 10459 3519
rect 10517 3485 10551 3519
rect 10784 3485 10818 3519
rect 12081 3485 12115 3519
rect 12357 3485 12391 3519
rect 14347 3485 14381 3519
rect 14637 3485 14671 3519
rect 14742 3485 14776 3519
rect 14841 3485 14875 3519
rect 17886 3485 17920 3519
rect 21833 3485 21867 3519
rect 22477 3485 22511 3519
rect 23121 3485 23155 3519
rect 24409 3485 24443 3519
rect 25053 3485 25087 3519
rect 4712 3417 4746 3451
rect 7214 3417 7248 3451
rect 8677 3417 8711 3451
rect 10158 3417 10192 3451
rect 12602 3417 12636 3451
rect 15362 3417 15396 3451
rect 22017 3417 22051 3451
rect 22201 3417 22235 3451
rect 6101 3349 6135 3383
rect 12265 3349 12299 3383
rect 15025 3349 15059 3383
rect 21649 3349 21683 3383
rect 22661 3349 22695 3383
rect 4813 3145 4847 3179
rect 6009 3145 6043 3179
rect 6377 3145 6411 3179
rect 7481 3145 7515 3179
rect 12909 3145 12943 3179
rect 13277 3145 13311 3179
rect 14841 3145 14875 3179
rect 15301 3077 15335 3111
rect 4997 3009 5031 3043
rect 5089 3009 5123 3043
rect 5365 3009 5399 3043
rect 5733 3009 5767 3043
rect 5825 3009 5859 3043
rect 8594 3009 8628 3043
rect 8861 3009 8895 3043
rect 11529 3009 11563 3043
rect 11796 3009 11830 3043
rect 13093 3009 13127 3043
rect 5457 2941 5491 2975
rect 14933 2873 14967 2907
rect 5273 2805 5307 2839
rect 5549 2805 5583 2839
rect 8033 2601 8067 2635
rect 8493 2601 8527 2635
rect 7941 2465 7975 2499
rect 8217 2397 8251 2431
rect 8309 2397 8343 2431
<< metal1 >>
rect 26234 28472 26240 28484
rect 26195 28444 26240 28472
rect 26234 28432 26240 28444
rect 26292 28432 26298 28484
rect 1104 27226 26128 27248
rect 1104 27174 9291 27226
rect 9343 27174 9355 27226
rect 9407 27174 9419 27226
rect 9471 27174 9483 27226
rect 9535 27174 9547 27226
rect 9599 27174 17632 27226
rect 17684 27174 17696 27226
rect 17748 27174 17760 27226
rect 17812 27174 17824 27226
rect 17876 27174 17888 27226
rect 17940 27174 26128 27226
rect 1104 27152 26128 27174
rect 1104 26682 26128 26704
rect 1104 26630 5120 26682
rect 5172 26630 5184 26682
rect 5236 26630 5248 26682
rect 5300 26630 5312 26682
rect 5364 26630 5376 26682
rect 5428 26630 13462 26682
rect 13514 26630 13526 26682
rect 13578 26630 13590 26682
rect 13642 26630 13654 26682
rect 13706 26630 13718 26682
rect 13770 26630 21803 26682
rect 21855 26630 21867 26682
rect 21919 26630 21931 26682
rect 21983 26630 21995 26682
rect 22047 26630 22059 26682
rect 22111 26630 26128 26682
rect 1104 26608 26128 26630
rect 12342 26528 12348 26580
rect 12400 26568 12406 26580
rect 12805 26571 12863 26577
rect 12805 26568 12817 26571
rect 12400 26540 12817 26568
rect 12400 26528 12406 26540
rect 12805 26537 12817 26540
rect 12851 26537 12863 26571
rect 12805 26531 12863 26537
rect 11808 26472 12572 26500
rect 11808 26376 11836 26472
rect 11790 26364 11796 26376
rect 11751 26336 11796 26364
rect 11790 26324 11796 26336
rect 11848 26324 11854 26376
rect 11885 26367 11943 26373
rect 11885 26333 11897 26367
rect 11931 26333 11943 26367
rect 11885 26327 11943 26333
rect 12252 26367 12310 26373
rect 12252 26333 12264 26367
rect 12298 26364 12310 26367
rect 12342 26364 12348 26376
rect 12298 26336 12348 26364
rect 12298 26333 12310 26336
rect 12252 26327 12310 26333
rect 11900 26296 11928 26327
rect 12342 26324 12348 26336
rect 12400 26324 12406 26376
rect 12544 26373 12572 26472
rect 12529 26367 12587 26373
rect 12529 26333 12541 26367
rect 12575 26333 12587 26367
rect 12820 26364 12848 26531
rect 15105 26435 15163 26441
rect 14476 26404 14964 26432
rect 13814 26364 13820 26376
rect 12820 26336 13820 26364
rect 12529 26327 12587 26333
rect 13814 26324 13820 26336
rect 13872 26364 13878 26376
rect 14093 26367 14151 26373
rect 14093 26364 14105 26367
rect 13872 26336 14105 26364
rect 13872 26324 13878 26336
rect 14093 26333 14105 26336
rect 14139 26333 14151 26367
rect 14093 26327 14151 26333
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26364 14335 26367
rect 14366 26364 14372 26376
rect 14323 26336 14372 26364
rect 14323 26333 14335 26336
rect 14277 26327 14335 26333
rect 14366 26324 14372 26336
rect 14424 26324 14430 26376
rect 12710 26296 12716 26308
rect 11900 26268 12716 26296
rect 12710 26256 12716 26268
rect 12768 26256 12774 26308
rect 14182 26256 14188 26308
rect 14240 26296 14246 26308
rect 14476 26305 14504 26404
rect 14795 26367 14853 26373
rect 14795 26333 14807 26367
rect 14841 26364 14853 26367
rect 14936 26364 14964 26404
rect 15105 26401 15117 26435
rect 15151 26432 15163 26435
rect 15151 26404 15516 26432
rect 15151 26401 15163 26404
rect 15105 26395 15163 26401
rect 15197 26367 15255 26373
rect 15197 26364 15209 26367
rect 14841 26333 14872 26364
rect 14936 26336 15209 26364
rect 14795 26327 14872 26333
rect 15197 26333 15209 26336
rect 15243 26364 15255 26367
rect 15289 26367 15347 26373
rect 15289 26364 15301 26367
rect 15243 26336 15301 26364
rect 15243 26333 15255 26336
rect 15197 26327 15255 26333
rect 15289 26333 15301 26336
rect 15335 26333 15347 26367
rect 15289 26327 15347 26333
rect 14461 26299 14519 26305
rect 14461 26296 14473 26299
rect 14240 26268 14473 26296
rect 14240 26256 14246 26268
rect 14461 26265 14473 26268
rect 14507 26265 14519 26299
rect 14461 26259 14519 26265
rect 14550 26256 14556 26308
rect 14608 26296 14614 26308
rect 14608 26268 14653 26296
rect 14608 26256 14614 26268
rect 12342 26228 12348 26240
rect 12303 26200 12348 26228
rect 12342 26188 12348 26200
rect 12400 26188 12406 26240
rect 14844 26228 14872 26327
rect 15488 26308 15516 26404
rect 15470 26296 15476 26308
rect 15431 26268 15476 26296
rect 15470 26256 15476 26268
rect 15528 26256 15534 26308
rect 15657 26299 15715 26305
rect 15657 26265 15669 26299
rect 15703 26296 15715 26299
rect 16301 26299 16359 26305
rect 16301 26296 16313 26299
rect 15703 26268 16313 26296
rect 15703 26265 15715 26268
rect 15657 26259 15715 26265
rect 16301 26265 16313 26268
rect 16347 26296 16359 26299
rect 16390 26296 16396 26308
rect 16347 26268 16396 26296
rect 16347 26265 16359 26268
rect 16301 26259 16359 26265
rect 15672 26228 15700 26259
rect 16390 26256 16396 26268
rect 16448 26256 16454 26308
rect 16485 26299 16543 26305
rect 16485 26265 16497 26299
rect 16531 26296 16543 26299
rect 16574 26296 16580 26308
rect 16531 26268 16580 26296
rect 16531 26265 16543 26268
rect 16485 26259 16543 26265
rect 16574 26256 16580 26268
rect 16632 26256 16638 26308
rect 16666 26256 16672 26308
rect 16724 26296 16730 26308
rect 16724 26268 16769 26296
rect 16724 26256 16730 26268
rect 14844 26200 15700 26228
rect 1104 26138 26128 26160
rect 1104 26086 9291 26138
rect 9343 26086 9355 26138
rect 9407 26086 9419 26138
rect 9471 26086 9483 26138
rect 9535 26086 9547 26138
rect 9599 26086 17632 26138
rect 17684 26086 17696 26138
rect 17748 26086 17760 26138
rect 17812 26086 17824 26138
rect 17876 26086 17888 26138
rect 17940 26086 26128 26138
rect 1104 26064 26128 26086
rect 566 25984 572 26036
rect 624 26024 630 26036
rect 11606 26024 11612 26036
rect 624 25996 11612 26024
rect 624 25984 630 25996
rect 11606 25984 11612 25996
rect 11664 25984 11670 26036
rect 12710 25984 12716 26036
rect 12768 26024 12774 26036
rect 12897 26027 12955 26033
rect 12897 26024 12909 26027
rect 12768 25996 12909 26024
rect 12768 25984 12774 25996
rect 12897 25993 12909 25996
rect 12943 25993 12955 26027
rect 12897 25987 12955 25993
rect 15470 25984 15476 26036
rect 15528 26024 15534 26036
rect 16025 26027 16083 26033
rect 16025 26024 16037 26027
rect 15528 25996 16037 26024
rect 15528 25984 15534 25996
rect 16025 25993 16037 25996
rect 16071 25993 16083 26027
rect 16025 25987 16083 25993
rect 11532 25928 14688 25956
rect 7926 25897 7932 25900
rect 7920 25851 7932 25897
rect 7984 25888 7990 25900
rect 11054 25888 11060 25900
rect 7984 25860 8020 25888
rect 11015 25860 11060 25888
rect 7926 25848 7932 25851
rect 7984 25848 7990 25860
rect 11054 25848 11060 25860
rect 11112 25848 11118 25900
rect 11146 25848 11152 25900
rect 11204 25888 11210 25900
rect 11532 25897 11560 25928
rect 13096 25897 13124 25928
rect 11517 25891 11575 25897
rect 11204 25860 11249 25888
rect 11204 25848 11210 25860
rect 11517 25857 11529 25891
rect 11563 25857 11575 25891
rect 11773 25891 11831 25897
rect 11773 25888 11785 25891
rect 11517 25851 11575 25857
rect 11624 25860 11785 25888
rect 6914 25780 6920 25832
rect 6972 25820 6978 25832
rect 7653 25823 7711 25829
rect 7653 25820 7665 25823
rect 6972 25792 7665 25820
rect 6972 25780 6978 25792
rect 7653 25789 7665 25792
rect 7699 25789 7711 25823
rect 11624 25820 11652 25860
rect 11773 25857 11785 25860
rect 11819 25857 11831 25891
rect 11773 25851 11831 25857
rect 13081 25891 13139 25897
rect 13081 25857 13093 25891
rect 13127 25857 13139 25891
rect 13081 25851 13139 25857
rect 13170 25848 13176 25900
rect 13228 25888 13234 25900
rect 13337 25891 13395 25897
rect 13337 25888 13349 25891
rect 13228 25860 13349 25888
rect 13228 25848 13234 25860
rect 13337 25857 13349 25860
rect 13383 25857 13395 25891
rect 13337 25851 13395 25857
rect 14660 25832 14688 25928
rect 14918 25897 14924 25900
rect 14912 25851 14924 25897
rect 14976 25888 14982 25900
rect 14976 25860 15012 25888
rect 14918 25848 14924 25851
rect 14976 25848 14982 25860
rect 16482 25848 16488 25900
rect 16540 25888 16546 25900
rect 16669 25891 16727 25897
rect 16669 25888 16681 25891
rect 16540 25860 16681 25888
rect 16540 25848 16546 25860
rect 16669 25857 16681 25860
rect 16715 25857 16727 25891
rect 16669 25851 16727 25857
rect 21726 25848 21732 25900
rect 21784 25888 21790 25900
rect 21821 25891 21879 25897
rect 21821 25888 21833 25891
rect 21784 25860 21833 25888
rect 21784 25848 21790 25860
rect 21821 25857 21833 25860
rect 21867 25857 21879 25891
rect 23106 25888 23112 25900
rect 23067 25860 23112 25888
rect 21821 25851 21879 25857
rect 23106 25848 23112 25860
rect 23164 25848 23170 25900
rect 25041 25891 25099 25897
rect 25041 25857 25053 25891
rect 25087 25888 25099 25891
rect 25498 25888 25504 25900
rect 25087 25860 25504 25888
rect 25087 25857 25099 25860
rect 25041 25851 25099 25857
rect 25498 25848 25504 25860
rect 25556 25848 25562 25900
rect 14642 25820 14648 25832
rect 7653 25783 7711 25789
rect 11348 25792 11652 25820
rect 14603 25792 14648 25820
rect 11348 25761 11376 25792
rect 14642 25780 14648 25792
rect 14700 25780 14706 25832
rect 16390 25780 16396 25832
rect 16448 25820 16454 25832
rect 16761 25823 16819 25829
rect 16761 25820 16773 25823
rect 16448 25792 16773 25820
rect 16448 25780 16454 25792
rect 16761 25789 16773 25792
rect 16807 25789 16819 25823
rect 16761 25783 16819 25789
rect 25317 25823 25375 25829
rect 25317 25789 25329 25823
rect 25363 25820 25375 25823
rect 26237 25823 26295 25829
rect 26237 25820 26249 25823
rect 25363 25792 26249 25820
rect 25363 25789 25375 25792
rect 25317 25783 25375 25789
rect 26237 25789 26249 25792
rect 26283 25789 26295 25823
rect 26237 25783 26295 25789
rect 11333 25755 11391 25761
rect 11333 25721 11345 25755
rect 11379 25721 11391 25755
rect 11333 25715 11391 25721
rect 16114 25712 16120 25764
rect 16172 25752 16178 25764
rect 16172 25724 17080 25752
rect 16172 25712 16178 25724
rect 7190 25644 7196 25696
rect 7248 25684 7254 25696
rect 7469 25687 7527 25693
rect 7469 25684 7481 25687
rect 7248 25656 7481 25684
rect 7248 25644 7254 25656
rect 7469 25653 7481 25656
rect 7515 25653 7527 25687
rect 7469 25647 7527 25653
rect 7558 25644 7564 25696
rect 7616 25684 7622 25696
rect 8846 25684 8852 25696
rect 7616 25656 8852 25684
rect 7616 25644 7622 25656
rect 8846 25644 8852 25656
rect 8904 25684 8910 25696
rect 9033 25687 9091 25693
rect 9033 25684 9045 25687
rect 8904 25656 9045 25684
rect 8904 25644 8910 25656
rect 9033 25653 9045 25656
rect 9079 25653 9091 25687
rect 9033 25647 9091 25653
rect 10686 25644 10692 25696
rect 10744 25684 10750 25696
rect 10873 25687 10931 25693
rect 10873 25684 10885 25687
rect 10744 25656 10885 25684
rect 10744 25644 10750 25656
rect 10873 25653 10885 25656
rect 10919 25653 10931 25687
rect 14458 25684 14464 25696
rect 14419 25656 14464 25684
rect 10873 25647 10931 25653
rect 14458 25644 14464 25656
rect 14516 25644 14522 25696
rect 16574 25644 16580 25696
rect 16632 25684 16638 25696
rect 17052 25693 17080 25724
rect 16669 25687 16727 25693
rect 16669 25684 16681 25687
rect 16632 25656 16681 25684
rect 16632 25644 16638 25656
rect 16669 25653 16681 25656
rect 16715 25653 16727 25687
rect 16669 25647 16727 25653
rect 17037 25687 17095 25693
rect 17037 25653 17049 25687
rect 17083 25684 17095 25687
rect 19242 25684 19248 25696
rect 17083 25656 19248 25684
rect 17083 25653 17095 25656
rect 17037 25647 17095 25653
rect 19242 25644 19248 25656
rect 19300 25644 19306 25696
rect 1104 25594 26128 25616
rect 1104 25542 5120 25594
rect 5172 25542 5184 25594
rect 5236 25542 5248 25594
rect 5300 25542 5312 25594
rect 5364 25542 5376 25594
rect 5428 25542 13462 25594
rect 13514 25542 13526 25594
rect 13578 25542 13590 25594
rect 13642 25542 13654 25594
rect 13706 25542 13718 25594
rect 13770 25542 21803 25594
rect 21855 25542 21867 25594
rect 21919 25542 21931 25594
rect 21983 25542 21995 25594
rect 22047 25542 22059 25594
rect 22111 25542 26128 25594
rect 1104 25520 26128 25542
rect 6914 25440 6920 25492
rect 6972 25480 6978 25492
rect 12989 25483 13047 25489
rect 6972 25452 10364 25480
rect 6972 25440 6978 25452
rect 7190 25372 7196 25424
rect 7248 25412 7254 25424
rect 7248 25384 8156 25412
rect 7248 25372 7254 25384
rect 7282 25304 7288 25356
rect 7340 25344 7346 25356
rect 7340 25316 7604 25344
rect 7340 25304 7346 25316
rect 7576 25288 7604 25316
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25276 6791 25279
rect 7009 25279 7067 25285
rect 7009 25276 7021 25279
rect 6779 25248 7021 25276
rect 6779 25245 6791 25248
rect 6733 25239 6791 25245
rect 7009 25245 7021 25248
rect 7055 25245 7067 25279
rect 7009 25239 7067 25245
rect 7098 25236 7104 25288
rect 7156 25276 7162 25288
rect 7469 25279 7527 25285
rect 7469 25276 7481 25279
rect 7156 25248 7481 25276
rect 7156 25236 7162 25248
rect 7469 25245 7481 25248
rect 7515 25245 7527 25279
rect 7469 25239 7527 25245
rect 7558 25236 7564 25288
rect 7616 25276 7622 25288
rect 7653 25279 7711 25285
rect 7653 25276 7665 25279
rect 7616 25248 7665 25276
rect 7616 25236 7622 25248
rect 7653 25245 7665 25248
rect 7699 25245 7711 25279
rect 7653 25239 7711 25245
rect 7834 25236 7840 25288
rect 7892 25276 7898 25288
rect 8021 25279 8079 25285
rect 8021 25276 8033 25279
rect 7892 25248 8033 25276
rect 7892 25236 7898 25248
rect 8021 25245 8033 25248
rect 8067 25245 8079 25279
rect 8128 25276 8156 25384
rect 8202 25304 8208 25356
rect 8260 25344 8266 25356
rect 8573 25347 8631 25353
rect 8573 25344 8585 25347
rect 8260 25316 8585 25344
rect 8260 25304 8266 25316
rect 8573 25313 8585 25316
rect 8619 25313 8631 25347
rect 10336 25344 10364 25452
rect 12989 25449 13001 25483
rect 13035 25480 13047 25483
rect 13170 25480 13176 25492
rect 13035 25452 13176 25480
rect 13035 25449 13047 25452
rect 12989 25443 13047 25449
rect 13170 25440 13176 25452
rect 13228 25440 13234 25492
rect 14366 25480 14372 25492
rect 14327 25452 14372 25480
rect 14366 25440 14372 25452
rect 14424 25440 14430 25492
rect 16574 25440 16580 25492
rect 16632 25480 16638 25492
rect 16669 25483 16727 25489
rect 16669 25480 16681 25483
rect 16632 25452 16681 25480
rect 16632 25440 16638 25452
rect 16669 25449 16681 25452
rect 16715 25480 16727 25483
rect 16758 25480 16764 25492
rect 16715 25452 16764 25480
rect 16715 25449 16727 25452
rect 16669 25443 16727 25449
rect 16758 25440 16764 25452
rect 16816 25440 16822 25492
rect 11790 25412 11796 25424
rect 11624 25384 11796 25412
rect 10410 25344 10416 25356
rect 10323 25316 10416 25344
rect 8573 25307 8631 25313
rect 10410 25304 10416 25316
rect 10468 25304 10474 25356
rect 10686 25285 10692 25288
rect 8297 25279 8355 25285
rect 8297 25276 8309 25279
rect 8128 25248 8309 25276
rect 8021 25239 8079 25245
rect 8297 25245 8309 25248
rect 8343 25276 8355 25279
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8343 25248 8953 25276
rect 8343 25245 8355 25248
rect 8297 25239 8355 25245
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 10321 25279 10379 25285
rect 10321 25245 10333 25279
rect 10367 25245 10379 25279
rect 10680 25276 10692 25285
rect 10647 25248 10692 25276
rect 10321 25239 10379 25245
rect 10680 25239 10692 25248
rect 6638 25168 6644 25220
rect 6696 25208 6702 25220
rect 7190 25208 7196 25220
rect 6696 25180 7196 25208
rect 6696 25168 6702 25180
rect 7190 25168 7196 25180
rect 7248 25168 7254 25220
rect 7374 25208 7380 25220
rect 7335 25180 7380 25208
rect 7374 25168 7380 25180
rect 7432 25168 7438 25220
rect 7929 25211 7987 25217
rect 7929 25177 7941 25211
rect 7975 25208 7987 25211
rect 8110 25208 8116 25220
rect 7975 25180 8116 25208
rect 7975 25177 7987 25180
rect 7929 25171 7987 25177
rect 8110 25168 8116 25180
rect 8168 25168 8174 25220
rect 8481 25211 8539 25217
rect 8481 25177 8493 25211
rect 8527 25208 8539 25211
rect 9214 25208 9220 25220
rect 8527 25180 9220 25208
rect 8527 25177 8539 25180
rect 8481 25171 8539 25177
rect 9214 25168 9220 25180
rect 9272 25168 9278 25220
rect 10336 25208 10364 25239
rect 10686 25236 10692 25239
rect 10744 25236 10750 25288
rect 11624 25208 11652 25384
rect 11790 25372 11796 25384
rect 11848 25372 11854 25424
rect 14182 25412 14188 25424
rect 13648 25384 14188 25412
rect 12342 25304 12348 25356
rect 12400 25344 12406 25356
rect 12437 25347 12495 25353
rect 12437 25344 12449 25347
rect 12400 25316 12449 25344
rect 12400 25304 12406 25316
rect 12437 25313 12449 25316
rect 12483 25313 12495 25347
rect 12618 25344 12624 25356
rect 12579 25316 12624 25344
rect 12437 25307 12495 25313
rect 12618 25304 12624 25316
rect 12676 25304 12682 25356
rect 12802 25276 12808 25288
rect 12763 25248 12808 25276
rect 12802 25236 12808 25248
rect 12860 25236 12866 25288
rect 13415 25279 13473 25285
rect 13415 25245 13427 25279
rect 13461 25276 13473 25279
rect 13648 25276 13676 25384
rect 14182 25372 14188 25384
rect 14240 25372 14246 25424
rect 13725 25347 13783 25353
rect 13725 25313 13737 25347
rect 13771 25344 13783 25347
rect 14458 25344 14464 25356
rect 13771 25316 14464 25344
rect 13771 25313 13783 25316
rect 13725 25307 13783 25313
rect 14458 25304 14464 25316
rect 14516 25304 14522 25356
rect 14642 25304 14648 25356
rect 14700 25344 14706 25356
rect 15289 25347 15347 25353
rect 15289 25344 15301 25347
rect 14700 25316 15301 25344
rect 14700 25304 14706 25316
rect 15289 25313 15301 25316
rect 15335 25313 15347 25347
rect 25038 25344 25044 25356
rect 24999 25316 25044 25344
rect 15289 25307 15347 25313
rect 25038 25304 25044 25316
rect 25096 25304 25102 25356
rect 13814 25276 13820 25288
rect 13461 25248 13676 25276
rect 13775 25248 13820 25276
rect 13461 25245 13473 25248
rect 13415 25239 13473 25245
rect 13814 25236 13820 25248
rect 13872 25236 13878 25288
rect 14090 25276 14096 25288
rect 14051 25248 14096 25276
rect 14090 25236 14096 25248
rect 14148 25236 14154 25288
rect 15010 25276 15016 25288
rect 14971 25248 15016 25276
rect 15010 25236 15016 25248
rect 15068 25236 15074 25288
rect 18322 25276 18328 25288
rect 18283 25248 18328 25276
rect 18322 25236 18328 25248
rect 18380 25236 18386 25288
rect 13170 25208 13176 25220
rect 10336 25180 11652 25208
rect 13131 25180 13176 25208
rect 13170 25168 13176 25180
rect 13228 25168 13234 25220
rect 14737 25211 14795 25217
rect 14737 25177 14749 25211
rect 14783 25208 14795 25211
rect 15102 25208 15108 25220
rect 14783 25180 15108 25208
rect 14783 25177 14795 25180
rect 14737 25171 14795 25177
rect 15102 25168 15108 25180
rect 15160 25168 15166 25220
rect 15534 25211 15592 25217
rect 15534 25208 15546 25211
rect 15212 25180 15546 25208
rect 6917 25143 6975 25149
rect 6917 25109 6929 25143
rect 6963 25140 6975 25143
rect 8386 25140 8392 25152
rect 6963 25112 8392 25140
rect 6963 25109 6975 25112
rect 6917 25103 6975 25109
rect 8386 25100 8392 25112
rect 8444 25100 8450 25152
rect 10229 25143 10287 25149
rect 10229 25109 10241 25143
rect 10275 25140 10287 25143
rect 11698 25140 11704 25152
rect 10275 25112 11704 25140
rect 10275 25109 10287 25112
rect 10229 25103 10287 25109
rect 11698 25100 11704 25112
rect 11756 25100 11762 25152
rect 11974 25140 11980 25152
rect 11935 25112 11980 25140
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 12342 25140 12348 25152
rect 12303 25112 12348 25140
rect 12342 25100 12348 25112
rect 12400 25100 12406 25152
rect 14360 25143 14418 25149
rect 14360 25109 14372 25143
rect 14406 25140 14418 25143
rect 14458 25140 14464 25152
rect 14406 25112 14464 25140
rect 14406 25109 14418 25112
rect 14360 25103 14418 25109
rect 14458 25100 14464 25112
rect 14516 25100 14522 25152
rect 14826 25140 14832 25152
rect 14787 25112 14832 25140
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 15212 25149 15240 25180
rect 15534 25177 15546 25180
rect 15580 25177 15592 25211
rect 15534 25171 15592 25177
rect 16850 25168 16856 25220
rect 16908 25208 16914 25220
rect 18058 25211 18116 25217
rect 18058 25208 18070 25211
rect 16908 25180 18070 25208
rect 16908 25168 16914 25180
rect 18058 25177 18070 25180
rect 18104 25177 18116 25211
rect 18058 25171 18116 25177
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25109 15255 25143
rect 15197 25103 15255 25109
rect 16390 25100 16396 25152
rect 16448 25140 16454 25152
rect 16945 25143 17003 25149
rect 16945 25140 16957 25143
rect 16448 25112 16957 25140
rect 16448 25100 16454 25112
rect 16945 25109 16957 25112
rect 16991 25109 17003 25143
rect 16945 25103 17003 25109
rect 1104 25050 26128 25072
rect 1104 24998 9291 25050
rect 9343 24998 9355 25050
rect 9407 24998 9419 25050
rect 9471 24998 9483 25050
rect 9535 24998 9547 25050
rect 9599 24998 17632 25050
rect 17684 24998 17696 25050
rect 17748 24998 17760 25050
rect 17812 24998 17824 25050
rect 17876 24998 17888 25050
rect 17940 24998 26128 25050
rect 1104 24976 26128 24998
rect 7193 24939 7251 24945
rect 7193 24905 7205 24939
rect 7239 24936 7251 24939
rect 7834 24936 7840 24948
rect 7239 24908 7840 24936
rect 7239 24905 7251 24908
rect 7193 24899 7251 24905
rect 7834 24896 7840 24908
rect 7892 24896 7898 24948
rect 7926 24896 7932 24948
rect 7984 24936 7990 24948
rect 8021 24939 8079 24945
rect 8021 24936 8033 24939
rect 7984 24908 8033 24936
rect 7984 24896 7990 24908
rect 8021 24905 8033 24908
rect 8067 24905 8079 24939
rect 8021 24899 8079 24905
rect 8110 24896 8116 24948
rect 8168 24936 8174 24948
rect 8573 24939 8631 24945
rect 8573 24936 8585 24939
rect 8168 24908 8585 24936
rect 8168 24896 8174 24908
rect 8573 24905 8585 24908
rect 8619 24905 8631 24939
rect 10321 24939 10379 24945
rect 10321 24936 10333 24939
rect 8573 24899 8631 24905
rect 8680 24908 10333 24936
rect 1670 24828 1676 24880
rect 1728 24868 1734 24880
rect 2682 24868 2688 24880
rect 1728 24840 2688 24868
rect 1728 24828 1734 24840
rect 2682 24828 2688 24840
rect 2740 24828 2746 24880
rect 7742 24868 7748 24880
rect 7300 24840 7512 24868
rect 7300 24812 7328 24840
rect 6641 24803 6699 24809
rect 6641 24769 6653 24803
rect 6687 24769 6699 24803
rect 6641 24763 6699 24769
rect 6656 24732 6684 24763
rect 6730 24760 6736 24812
rect 6788 24800 6794 24812
rect 7098 24800 7104 24812
rect 6788 24772 6833 24800
rect 7059 24772 7104 24800
rect 6788 24760 6794 24772
rect 7098 24760 7104 24772
rect 7156 24760 7162 24812
rect 7282 24800 7288 24812
rect 7243 24772 7288 24800
rect 7282 24760 7288 24772
rect 7340 24760 7346 24812
rect 7377 24803 7435 24809
rect 7377 24769 7389 24803
rect 7423 24769 7435 24803
rect 7484 24800 7512 24840
rect 7668 24840 7748 24868
rect 7668 24809 7696 24840
rect 7742 24828 7748 24840
rect 7800 24828 7806 24880
rect 7852 24868 7880 24896
rect 8478 24868 8484 24880
rect 7852 24840 8484 24868
rect 8478 24828 8484 24840
rect 8536 24828 8542 24880
rect 7542 24803 7600 24809
rect 7542 24800 7554 24803
rect 7484 24772 7554 24800
rect 7377 24763 7435 24769
rect 7542 24769 7554 24772
rect 7588 24769 7600 24803
rect 7542 24763 7600 24769
rect 7650 24803 7708 24809
rect 7650 24769 7662 24803
rect 7696 24769 7708 24803
rect 7650 24763 7708 24769
rect 7929 24803 7987 24809
rect 7929 24769 7941 24803
rect 7975 24800 7987 24803
rect 8202 24800 8208 24812
rect 7975 24772 8208 24800
rect 7975 24769 7987 24772
rect 7929 24763 7987 24769
rect 6656 24704 6776 24732
rect 6748 24664 6776 24704
rect 7190 24692 7196 24744
rect 7248 24732 7254 24744
rect 7392 24732 7420 24763
rect 8202 24760 8208 24772
rect 8260 24800 8266 24812
rect 8680 24800 8708 24908
rect 10321 24905 10333 24908
rect 10367 24936 10379 24939
rect 12158 24936 12164 24948
rect 10367 24908 12164 24936
rect 10367 24905 10379 24908
rect 10321 24899 10379 24905
rect 12158 24896 12164 24908
rect 12216 24896 12222 24948
rect 12989 24939 13047 24945
rect 12989 24905 13001 24939
rect 13035 24936 13047 24939
rect 13170 24936 13176 24948
rect 13035 24908 13176 24936
rect 13035 24905 13047 24908
rect 12989 24899 13047 24905
rect 13170 24896 13176 24908
rect 13228 24896 13234 24948
rect 13357 24939 13415 24945
rect 13357 24905 13369 24939
rect 13403 24905 13415 24939
rect 13357 24899 13415 24905
rect 10962 24877 10968 24880
rect 10956 24868 10968 24877
rect 10923 24840 10968 24868
rect 10956 24831 10968 24840
rect 10962 24828 10968 24831
rect 11020 24828 11026 24880
rect 11885 24871 11943 24877
rect 11885 24837 11897 24871
rect 11931 24868 11943 24871
rect 13372 24868 13400 24899
rect 14366 24896 14372 24948
rect 14424 24936 14430 24948
rect 14645 24939 14703 24945
rect 14645 24936 14657 24939
rect 14424 24908 14657 24936
rect 14424 24896 14430 24908
rect 14645 24905 14657 24908
rect 14691 24905 14703 24939
rect 14645 24899 14703 24905
rect 15749 24939 15807 24945
rect 15749 24905 15761 24939
rect 15795 24936 15807 24939
rect 16850 24936 16856 24948
rect 15795 24908 16856 24936
rect 15795 24905 15807 24908
rect 15749 24899 15807 24905
rect 16850 24896 16856 24908
rect 16908 24896 16914 24948
rect 14274 24868 14280 24880
rect 11931 24840 13400 24868
rect 14235 24840 14280 24868
rect 11931 24837 11943 24840
rect 11885 24831 11943 24837
rect 14274 24828 14280 24840
rect 14332 24828 14338 24880
rect 15105 24871 15163 24877
rect 15105 24837 15117 24871
rect 15151 24868 15163 24871
rect 15378 24868 15384 24880
rect 15151 24840 15384 24868
rect 15151 24837 15163 24840
rect 15105 24831 15163 24837
rect 15378 24828 15384 24840
rect 15436 24828 15442 24880
rect 16482 24828 16488 24880
rect 16540 24868 16546 24880
rect 16540 24840 16712 24868
rect 16540 24828 16546 24840
rect 9214 24800 9220 24812
rect 8260 24772 8708 24800
rect 9175 24772 9220 24800
rect 8260 24760 8266 24772
rect 9214 24760 9220 24772
rect 9272 24760 9278 24812
rect 10413 24803 10471 24809
rect 10413 24769 10425 24803
rect 10459 24769 10471 24803
rect 10413 24763 10471 24769
rect 10689 24803 10747 24809
rect 10689 24769 10701 24803
rect 10735 24800 10747 24803
rect 11054 24800 11060 24812
rect 10735 24772 11060 24800
rect 10735 24769 10747 24772
rect 10689 24763 10747 24769
rect 7248 24704 7420 24732
rect 7745 24735 7803 24741
rect 7248 24692 7254 24704
rect 7745 24701 7757 24735
rect 7791 24732 7803 24735
rect 7834 24732 7840 24744
rect 7791 24704 7840 24732
rect 7791 24701 7803 24704
rect 7745 24695 7803 24701
rect 7834 24692 7840 24704
rect 7892 24692 7898 24744
rect 8665 24735 8723 24741
rect 8665 24701 8677 24735
rect 8711 24701 8723 24735
rect 8665 24695 8723 24701
rect 8205 24667 8263 24673
rect 8205 24664 8217 24667
rect 6748 24636 8217 24664
rect 8205 24633 8217 24636
rect 8251 24633 8263 24667
rect 8680 24664 8708 24695
rect 8754 24692 8760 24744
rect 8812 24732 8818 24744
rect 8849 24735 8907 24741
rect 8849 24732 8861 24735
rect 8812 24704 8861 24732
rect 8812 24692 8818 24704
rect 8849 24701 8861 24704
rect 8895 24732 8907 24735
rect 10428 24732 10456 24763
rect 11054 24760 11060 24772
rect 11112 24760 11118 24812
rect 11330 24800 11336 24812
rect 11291 24772 11336 24800
rect 11330 24760 11336 24772
rect 11388 24760 11394 24812
rect 11698 24760 11704 24812
rect 11756 24800 11762 24812
rect 11977 24803 12035 24809
rect 11977 24800 11989 24803
rect 11756 24772 11989 24800
rect 11756 24760 11762 24772
rect 11977 24769 11989 24772
rect 12023 24769 12035 24803
rect 11977 24763 12035 24769
rect 12897 24803 12955 24809
rect 12897 24769 12909 24803
rect 12943 24800 12955 24803
rect 13262 24800 13268 24812
rect 12943 24772 13268 24800
rect 12943 24769 12955 24772
rect 12897 24763 12955 24769
rect 13262 24760 13268 24772
rect 13320 24760 13326 24812
rect 13354 24760 13360 24812
rect 13412 24800 13418 24812
rect 13541 24803 13599 24809
rect 13541 24800 13553 24803
rect 13412 24772 13553 24800
rect 13412 24760 13418 24772
rect 13541 24769 13553 24772
rect 13587 24769 13599 24803
rect 13541 24763 13599 24769
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24800 13691 24803
rect 14090 24800 14096 24812
rect 13679 24772 14096 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 14090 24760 14096 24772
rect 14148 24760 14154 24812
rect 14185 24803 14243 24809
rect 14185 24769 14197 24803
rect 14231 24800 14243 24803
rect 14550 24800 14556 24812
rect 14231 24772 14556 24800
rect 14231 24769 14243 24772
rect 14185 24763 14243 24769
rect 14550 24760 14556 24772
rect 14608 24760 14614 24812
rect 14826 24760 14832 24812
rect 14884 24800 14890 24812
rect 15562 24800 15568 24812
rect 14884 24772 15424 24800
rect 15523 24772 15568 24800
rect 14884 24760 14890 24772
rect 11882 24732 11888 24744
rect 8895 24704 9628 24732
rect 10428 24704 11888 24732
rect 8895 24701 8907 24704
rect 8849 24695 8907 24701
rect 9033 24667 9091 24673
rect 9033 24664 9045 24667
rect 8680 24636 9045 24664
rect 8205 24627 8263 24633
rect 9033 24633 9045 24636
rect 9079 24633 9091 24667
rect 9033 24627 9091 24633
rect 6733 24599 6791 24605
rect 6733 24565 6745 24599
rect 6779 24596 6791 24599
rect 7834 24596 7840 24608
rect 6779 24568 7840 24596
rect 6779 24565 6791 24568
rect 6733 24559 6791 24565
rect 7834 24556 7840 24568
rect 7892 24556 7898 24608
rect 8110 24556 8116 24608
rect 8168 24596 8174 24608
rect 9600 24605 9628 24704
rect 11882 24692 11888 24704
rect 11940 24692 11946 24744
rect 12158 24732 12164 24744
rect 12071 24704 12164 24732
rect 12158 24692 12164 24704
rect 12216 24732 12222 24744
rect 12437 24735 12495 24741
rect 12437 24732 12449 24735
rect 12216 24704 12449 24732
rect 12216 24692 12222 24704
rect 12437 24701 12449 24704
rect 12483 24732 12495 24735
rect 12618 24732 12624 24744
rect 12483 24704 12624 24732
rect 12483 24701 12495 24704
rect 12437 24695 12495 24701
rect 12618 24692 12624 24704
rect 12676 24732 12682 24744
rect 13173 24735 13231 24741
rect 13173 24732 13185 24735
rect 12676 24704 13185 24732
rect 12676 24692 12682 24704
rect 13173 24701 13185 24704
rect 13219 24732 13231 24735
rect 13998 24732 14004 24744
rect 13219 24704 14004 24732
rect 13219 24701 13231 24704
rect 13173 24695 13231 24701
rect 13998 24692 14004 24704
rect 14056 24732 14062 24744
rect 14844 24732 14872 24760
rect 15396 24741 15424 24772
rect 15562 24760 15568 24772
rect 15620 24760 15626 24812
rect 16114 24809 16120 24812
rect 16083 24803 16120 24809
rect 16083 24769 16095 24803
rect 16083 24763 16120 24769
rect 16114 24760 16120 24763
rect 16172 24760 16178 24812
rect 16390 24800 16396 24812
rect 16351 24772 16396 24800
rect 16390 24760 16396 24772
rect 16448 24760 16454 24812
rect 14056 24704 14872 24732
rect 15197 24735 15255 24741
rect 14056 24692 14062 24704
rect 15197 24701 15209 24735
rect 15243 24701 15255 24735
rect 15197 24695 15255 24701
rect 15381 24735 15439 24741
rect 15381 24701 15393 24735
rect 15427 24732 15439 24735
rect 15654 24732 15660 24744
rect 15427 24704 15660 24732
rect 15427 24701 15439 24704
rect 15381 24695 15439 24701
rect 10597 24667 10655 24673
rect 10597 24633 10609 24667
rect 10643 24664 10655 24667
rect 12342 24664 12348 24676
rect 10643 24636 12348 24664
rect 10643 24633 10655 24636
rect 10597 24627 10655 24633
rect 12342 24624 12348 24636
rect 12400 24624 12406 24676
rect 13817 24667 13875 24673
rect 13817 24633 13829 24667
rect 13863 24664 13875 24667
rect 14918 24664 14924 24676
rect 13863 24636 14924 24664
rect 13863 24633 13875 24636
rect 13817 24627 13875 24633
rect 14918 24624 14924 24636
rect 14976 24624 14982 24676
rect 15212 24664 15240 24695
rect 15654 24692 15660 24704
rect 15712 24692 15718 24744
rect 16485 24735 16543 24741
rect 16485 24701 16497 24735
rect 16531 24732 16543 24735
rect 16574 24732 16580 24744
rect 16531 24704 16580 24732
rect 16531 24701 16543 24704
rect 16485 24695 16543 24701
rect 16574 24692 16580 24704
rect 16632 24692 16638 24744
rect 16684 24741 16712 24840
rect 17034 24760 17040 24812
rect 17092 24809 17098 24812
rect 17092 24803 17129 24809
rect 17117 24769 17129 24803
rect 17092 24763 17129 24769
rect 17092 24760 17098 24763
rect 16669 24735 16727 24741
rect 16669 24701 16681 24735
rect 16715 24701 16727 24735
rect 16669 24695 16727 24701
rect 16758 24692 16764 24744
rect 16816 24732 16822 24744
rect 16816 24704 16861 24732
rect 16816 24692 16822 24704
rect 17313 24667 17371 24673
rect 17313 24664 17325 24667
rect 15212 24636 17325 24664
rect 17313 24633 17325 24636
rect 17359 24633 17371 24667
rect 17313 24627 17371 24633
rect 9309 24599 9367 24605
rect 9309 24596 9321 24599
rect 8168 24568 9321 24596
rect 8168 24556 8174 24568
rect 9309 24565 9321 24568
rect 9355 24565 9367 24599
rect 9309 24559 9367 24565
rect 9585 24599 9643 24605
rect 9585 24565 9597 24599
rect 9631 24596 9643 24599
rect 10502 24596 10508 24608
rect 9631 24568 10508 24596
rect 9631 24565 9643 24568
rect 9585 24559 9643 24565
rect 10502 24556 10508 24568
rect 10560 24556 10566 24608
rect 10965 24599 11023 24605
rect 10965 24565 10977 24599
rect 11011 24596 11023 24599
rect 11517 24599 11575 24605
rect 11517 24596 11529 24599
rect 11011 24568 11529 24596
rect 11011 24565 11023 24568
rect 10965 24559 11023 24565
rect 11517 24565 11529 24568
rect 11563 24565 11575 24599
rect 11517 24559 11575 24565
rect 12526 24556 12532 24608
rect 12584 24596 12590 24608
rect 12584 24568 12629 24596
rect 12584 24556 12590 24568
rect 14550 24556 14556 24608
rect 14608 24596 14614 24608
rect 14737 24599 14795 24605
rect 14737 24596 14749 24599
rect 14608 24568 14749 24596
rect 14608 24556 14614 24568
rect 14737 24565 14749 24568
rect 14783 24565 14795 24599
rect 14737 24559 14795 24565
rect 15933 24599 15991 24605
rect 15933 24565 15945 24599
rect 15979 24596 15991 24599
rect 16298 24596 16304 24608
rect 15979 24568 16304 24596
rect 15979 24565 15991 24568
rect 15933 24559 15991 24565
rect 16298 24556 16304 24568
rect 16356 24556 16362 24608
rect 1104 24506 26128 24528
rect 1104 24454 5120 24506
rect 5172 24454 5184 24506
rect 5236 24454 5248 24506
rect 5300 24454 5312 24506
rect 5364 24454 5376 24506
rect 5428 24454 13462 24506
rect 13514 24454 13526 24506
rect 13578 24454 13590 24506
rect 13642 24454 13654 24506
rect 13706 24454 13718 24506
rect 13770 24454 21803 24506
rect 21855 24454 21867 24506
rect 21919 24454 21931 24506
rect 21983 24454 21995 24506
rect 22047 24454 22059 24506
rect 22111 24454 26128 24506
rect 1104 24432 26128 24454
rect 2130 24392 2136 24404
rect 2091 24364 2136 24392
rect 2130 24352 2136 24364
rect 2188 24352 2194 24404
rect 6181 24395 6239 24401
rect 6181 24361 6193 24395
rect 6227 24392 6239 24395
rect 6362 24392 6368 24404
rect 6227 24364 6368 24392
rect 6227 24361 6239 24364
rect 6181 24355 6239 24361
rect 6362 24352 6368 24364
rect 6420 24392 6426 24404
rect 7098 24392 7104 24404
rect 6420 24364 7104 24392
rect 6420 24352 6426 24364
rect 7098 24352 7104 24364
rect 7156 24352 7162 24404
rect 7282 24352 7288 24404
rect 7340 24352 7346 24404
rect 7558 24352 7564 24404
rect 7616 24392 7622 24404
rect 7616 24364 10824 24392
rect 7616 24352 7622 24364
rect 7300 24324 7328 24352
rect 7834 24324 7840 24336
rect 7300 24296 7840 24324
rect 7834 24284 7840 24296
rect 7892 24324 7898 24336
rect 8110 24324 8116 24336
rect 7892 24296 8116 24324
rect 7892 24284 7898 24296
rect 8110 24284 8116 24296
rect 8168 24324 8174 24336
rect 8168 24296 9444 24324
rect 8168 24284 8174 24296
rect 8386 24256 8392 24268
rect 8347 24228 8392 24256
rect 8386 24216 8392 24228
rect 8444 24216 8450 24268
rect 8573 24259 8631 24265
rect 8573 24225 8585 24259
rect 8619 24256 8631 24259
rect 8754 24256 8760 24268
rect 8619 24228 8760 24256
rect 8619 24225 8631 24228
rect 8573 24219 8631 24225
rect 8754 24216 8760 24228
rect 8812 24216 8818 24268
rect 3786 24148 3792 24200
rect 3844 24188 3850 24200
rect 4801 24191 4859 24197
rect 4801 24188 4813 24191
rect 3844 24160 4813 24188
rect 3844 24148 3850 24160
rect 4801 24157 4813 24160
rect 4847 24157 4859 24191
rect 4801 24151 4859 24157
rect 6365 24191 6423 24197
rect 6365 24157 6377 24191
rect 6411 24188 6423 24191
rect 6411 24160 6868 24188
rect 6411 24157 6423 24160
rect 6365 24151 6423 24157
rect 6840 24132 6868 24160
rect 7374 24148 7380 24200
rect 7432 24188 7438 24200
rect 8018 24188 8024 24200
rect 7432 24160 8024 24188
rect 7432 24148 7438 24160
rect 8018 24148 8024 24160
rect 8076 24188 8082 24200
rect 8297 24191 8355 24197
rect 8297 24188 8309 24191
rect 8076 24160 8309 24188
rect 8076 24148 8082 24160
rect 8297 24157 8309 24160
rect 8343 24157 8355 24191
rect 9416 24188 9444 24296
rect 10410 24256 10416 24268
rect 10371 24228 10416 24256
rect 10410 24216 10416 24228
rect 10468 24216 10474 24268
rect 10796 24265 10824 24364
rect 11146 24352 11152 24404
rect 11204 24392 11210 24404
rect 11425 24395 11483 24401
rect 11425 24392 11437 24395
rect 11204 24364 11437 24392
rect 11204 24352 11210 24364
rect 11425 24361 11437 24364
rect 11471 24361 11483 24395
rect 11425 24355 11483 24361
rect 11609 24395 11667 24401
rect 11609 24361 11621 24395
rect 11655 24392 11667 24395
rect 11974 24392 11980 24404
rect 11655 24364 11980 24392
rect 11655 24361 11667 24364
rect 11609 24355 11667 24361
rect 11974 24352 11980 24364
rect 12032 24352 12038 24404
rect 12526 24392 12532 24404
rect 12487 24364 12532 24392
rect 12526 24352 12532 24364
rect 12584 24352 12590 24404
rect 12713 24395 12771 24401
rect 12713 24361 12725 24395
rect 12759 24392 12771 24395
rect 12802 24392 12808 24404
rect 12759 24364 12808 24392
rect 12759 24361 12771 24364
rect 12713 24355 12771 24361
rect 12802 24352 12808 24364
rect 12860 24352 12866 24404
rect 12989 24395 13047 24401
rect 12989 24361 13001 24395
rect 13035 24392 13047 24395
rect 13817 24395 13875 24401
rect 13817 24392 13829 24395
rect 13035 24364 13829 24392
rect 13035 24361 13047 24364
rect 12989 24355 13047 24361
rect 13817 24361 13829 24364
rect 13863 24392 13875 24395
rect 13998 24392 14004 24404
rect 13863 24364 14004 24392
rect 13863 24361 13875 24364
rect 13817 24355 13875 24361
rect 13998 24352 14004 24364
rect 14056 24352 14062 24404
rect 14550 24392 14556 24404
rect 14511 24364 14556 24392
rect 14550 24352 14556 24364
rect 14608 24352 14614 24404
rect 14737 24395 14795 24401
rect 14737 24361 14749 24395
rect 14783 24392 14795 24395
rect 15010 24392 15016 24404
rect 14783 24364 15016 24392
rect 14783 24361 14795 24364
rect 14737 24355 14795 24361
rect 15010 24352 15016 24364
rect 15068 24352 15074 24404
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24361 15531 24395
rect 15473 24355 15531 24361
rect 15488 24324 15516 24355
rect 15562 24352 15568 24404
rect 15620 24392 15626 24404
rect 15657 24395 15715 24401
rect 15657 24392 15669 24395
rect 15620 24364 15669 24392
rect 15620 24352 15626 24364
rect 15657 24361 15669 24364
rect 15703 24361 15715 24395
rect 15657 24355 15715 24361
rect 19061 24395 19119 24401
rect 19061 24361 19073 24395
rect 19107 24392 19119 24395
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 19107 24364 19257 24392
rect 19107 24361 19119 24364
rect 19061 24355 19119 24361
rect 19245 24361 19257 24364
rect 19291 24361 19303 24395
rect 19245 24355 19303 24361
rect 15841 24327 15899 24333
rect 15841 24324 15853 24327
rect 15488 24296 15853 24324
rect 15841 24293 15853 24296
rect 15887 24293 15899 24327
rect 15841 24287 15899 24293
rect 10781 24259 10839 24265
rect 10781 24225 10793 24259
rect 10827 24256 10839 24259
rect 10870 24256 10876 24268
rect 10827 24228 10876 24256
rect 10827 24225 10839 24228
rect 10781 24219 10839 24225
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 11149 24259 11207 24265
rect 11149 24225 11161 24259
rect 11195 24256 11207 24259
rect 13354 24256 13360 24268
rect 11195 24228 13360 24256
rect 11195 24225 11207 24228
rect 11149 24219 11207 24225
rect 13354 24216 13360 24228
rect 13412 24216 13418 24268
rect 16298 24256 16304 24268
rect 16259 24228 16304 24256
rect 16298 24216 16304 24228
rect 16356 24216 16362 24268
rect 16390 24216 16396 24268
rect 16448 24256 16454 24268
rect 16448 24228 16493 24256
rect 16448 24216 16454 24228
rect 10965 24191 11023 24197
rect 9416 24160 10916 24188
rect 8297 24151 8355 24157
rect 5068 24123 5126 24129
rect 5068 24089 5080 24123
rect 5114 24120 5126 24123
rect 5258 24120 5264 24132
rect 5114 24092 5264 24120
rect 5114 24089 5126 24092
rect 5068 24083 5126 24089
rect 5258 24080 5264 24092
rect 5316 24080 5322 24132
rect 5902 24080 5908 24132
rect 5960 24120 5966 24132
rect 6610 24123 6668 24129
rect 6610 24120 6622 24123
rect 5960 24092 6622 24120
rect 5960 24080 5966 24092
rect 6610 24089 6622 24092
rect 6656 24089 6668 24123
rect 6610 24083 6668 24089
rect 6822 24080 6828 24132
rect 6880 24080 6886 24132
rect 8386 24120 8392 24132
rect 7760 24092 8392 24120
rect 6730 24012 6736 24064
rect 6788 24052 6794 24064
rect 7558 24052 7564 24064
rect 6788 24024 7564 24052
rect 6788 24012 6794 24024
rect 7558 24012 7564 24024
rect 7616 24012 7622 24064
rect 7760 24061 7788 24092
rect 8386 24080 8392 24092
rect 8444 24080 8450 24132
rect 10134 24120 10140 24132
rect 10192 24129 10198 24132
rect 10104 24092 10140 24120
rect 10134 24080 10140 24092
rect 10192 24083 10204 24129
rect 10888 24120 10916 24160
rect 10965 24157 10977 24191
rect 11011 24188 11023 24191
rect 11238 24188 11244 24200
rect 11011 24160 11244 24188
rect 11011 24157 11023 24160
rect 10965 24151 11023 24157
rect 11238 24148 11244 24160
rect 11296 24148 11302 24200
rect 11330 24148 11336 24200
rect 11388 24188 11394 24200
rect 11977 24191 12035 24197
rect 11977 24188 11989 24191
rect 11388 24160 11989 24188
rect 11388 24148 11394 24160
rect 11977 24157 11989 24160
rect 12023 24188 12035 24191
rect 12161 24191 12219 24197
rect 12161 24188 12173 24191
rect 12023 24160 12173 24188
rect 12023 24157 12035 24160
rect 11977 24151 12035 24157
rect 12161 24157 12173 24160
rect 12207 24188 12219 24191
rect 12342 24188 12348 24200
rect 12207 24160 12348 24188
rect 12207 24157 12219 24160
rect 12161 24151 12219 24157
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 15102 24188 15108 24200
rect 13464 24160 14504 24188
rect 11146 24120 11152 24132
rect 10888 24092 11152 24120
rect 10192 24080 10198 24083
rect 11146 24080 11152 24092
rect 11204 24080 11210 24132
rect 12575 24123 12633 24129
rect 12575 24120 12587 24123
rect 12406 24092 12587 24120
rect 7745 24055 7803 24061
rect 7745 24021 7757 24055
rect 7791 24021 7803 24055
rect 7926 24052 7932 24064
rect 7887 24024 7932 24052
rect 7745 24015 7803 24021
rect 7926 24012 7932 24024
rect 7984 24012 7990 24064
rect 8938 24012 8944 24064
rect 8996 24052 9002 24064
rect 9033 24055 9091 24061
rect 9033 24052 9045 24055
rect 8996 24024 9045 24052
rect 8996 24012 9002 24024
rect 9033 24021 9045 24024
rect 9079 24021 9091 24055
rect 10594 24052 10600 24064
rect 10555 24024 10600 24052
rect 9033 24015 9091 24021
rect 10594 24012 10600 24024
rect 10652 24012 10658 24064
rect 11600 24055 11658 24061
rect 11600 24021 11612 24055
rect 11646 24052 11658 24055
rect 12250 24052 12256 24064
rect 11646 24024 12256 24052
rect 11646 24021 11658 24024
rect 11600 24015 11658 24021
rect 12250 24012 12256 24024
rect 12308 24052 12314 24064
rect 12406 24052 12434 24092
rect 12575 24089 12587 24092
rect 12621 24120 12633 24123
rect 13464 24120 13492 24160
rect 14476 24132 14504 24160
rect 14844 24160 15108 24188
rect 14182 24120 14188 24132
rect 12621 24092 13492 24120
rect 14143 24092 14188 24120
rect 12621 24089 12633 24092
rect 12575 24083 12633 24089
rect 14182 24080 14188 24092
rect 14240 24080 14246 24132
rect 14458 24080 14464 24132
rect 14516 24120 14522 24132
rect 14562 24123 14620 24129
rect 14562 24120 14574 24123
rect 14516 24092 14574 24120
rect 14516 24080 14522 24092
rect 14562 24089 14574 24092
rect 14608 24089 14620 24123
rect 14562 24083 14620 24089
rect 12308 24024 12434 24052
rect 14200 24052 14228 24080
rect 14844 24052 14872 24160
rect 15102 24148 15108 24160
rect 15160 24148 15166 24200
rect 17497 24191 17555 24197
rect 17497 24157 17509 24191
rect 17543 24188 17555 24191
rect 18322 24188 18328 24200
rect 17543 24160 18328 24188
rect 17543 24157 17555 24160
rect 17497 24151 17555 24157
rect 18322 24148 18328 24160
rect 18380 24188 18386 24200
rect 18874 24188 18880 24200
rect 18380 24160 18880 24188
rect 18380 24148 18386 24160
rect 18874 24148 18880 24160
rect 18932 24148 18938 24200
rect 19242 24188 19248 24200
rect 19203 24160 19248 24188
rect 19242 24148 19248 24160
rect 19300 24188 19306 24200
rect 19429 24191 19487 24197
rect 19300 24148 19334 24188
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 19518 24188 19524 24200
rect 19475 24160 19524 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 17034 24080 17040 24132
rect 17092 24120 17098 24132
rect 17742 24123 17800 24129
rect 17742 24120 17754 24123
rect 17092 24092 17754 24120
rect 17092 24080 17098 24092
rect 17742 24089 17754 24092
rect 17788 24089 17800 24123
rect 17742 24083 17800 24089
rect 18598 24080 18604 24132
rect 18656 24120 18662 24132
rect 19306 24120 19334 24148
rect 20438 24120 20444 24132
rect 18656 24092 20444 24120
rect 18656 24080 18662 24092
rect 20438 24080 20444 24092
rect 20496 24080 20502 24132
rect 14200 24024 14872 24052
rect 15482 24055 15540 24061
rect 12308 24012 12314 24024
rect 15482 24021 15494 24055
rect 15528 24052 15540 24055
rect 16022 24052 16028 24064
rect 15528 24024 16028 24052
rect 15528 24021 15540 24024
rect 15482 24015 15540 24021
rect 16022 24012 16028 24024
rect 16080 24012 16086 24064
rect 16209 24055 16267 24061
rect 16209 24021 16221 24055
rect 16255 24052 16267 24055
rect 16574 24052 16580 24064
rect 16255 24024 16580 24052
rect 16255 24021 16267 24024
rect 16209 24015 16267 24021
rect 16574 24012 16580 24024
rect 16632 24012 16638 24064
rect 18506 24012 18512 24064
rect 18564 24052 18570 24064
rect 18877 24055 18935 24061
rect 18877 24052 18889 24055
rect 18564 24024 18889 24052
rect 18564 24012 18570 24024
rect 18877 24021 18889 24024
rect 18923 24052 18935 24055
rect 19061 24055 19119 24061
rect 19061 24052 19073 24055
rect 18923 24024 19073 24052
rect 18923 24021 18935 24024
rect 18877 24015 18935 24021
rect 19061 24021 19073 24024
rect 19107 24021 19119 24055
rect 19610 24052 19616 24064
rect 19571 24024 19616 24052
rect 19061 24015 19119 24021
rect 19610 24012 19616 24024
rect 19668 24012 19674 24064
rect 1104 23962 26128 23984
rect 1104 23910 9291 23962
rect 9343 23910 9355 23962
rect 9407 23910 9419 23962
rect 9471 23910 9483 23962
rect 9535 23910 9547 23962
rect 9599 23910 17632 23962
rect 17684 23910 17696 23962
rect 17748 23910 17760 23962
rect 17812 23910 17824 23962
rect 17876 23910 17888 23962
rect 17940 23910 26128 23962
rect 1104 23888 26128 23910
rect 5258 23848 5264 23860
rect 5219 23820 5264 23848
rect 5258 23808 5264 23820
rect 5316 23808 5322 23860
rect 5902 23848 5908 23860
rect 5863 23820 5908 23848
rect 5902 23808 5908 23820
rect 5960 23808 5966 23860
rect 8018 23848 8024 23860
rect 7979 23820 8024 23848
rect 8018 23808 8024 23820
rect 8076 23808 8082 23860
rect 8202 23808 8208 23860
rect 8260 23848 8266 23860
rect 8260 23820 8340 23848
rect 8260 23808 8266 23820
rect 4893 23783 4951 23789
rect 4893 23749 4905 23783
rect 4939 23780 4951 23783
rect 5077 23783 5135 23789
rect 5077 23780 5089 23783
rect 4939 23752 5089 23780
rect 4939 23749 4951 23752
rect 4893 23743 4951 23749
rect 5077 23749 5089 23752
rect 5123 23780 5135 23783
rect 7282 23780 7288 23792
rect 5123 23752 7288 23780
rect 5123 23749 5135 23752
rect 5077 23743 5135 23749
rect 5736 23721 5764 23752
rect 7282 23740 7288 23752
rect 7340 23740 7346 23792
rect 7926 23780 7932 23792
rect 7392 23752 7932 23780
rect 5353 23715 5411 23721
rect 5353 23681 5365 23715
rect 5399 23681 5411 23715
rect 5353 23675 5411 23681
rect 5537 23715 5595 23721
rect 5537 23681 5549 23715
rect 5583 23712 5595 23715
rect 5721 23715 5779 23721
rect 5721 23712 5733 23715
rect 5583 23684 5733 23712
rect 5583 23681 5595 23684
rect 5537 23675 5595 23681
rect 5721 23681 5733 23684
rect 5767 23681 5779 23715
rect 5721 23675 5779 23681
rect 5905 23715 5963 23721
rect 5905 23681 5917 23715
rect 5951 23681 5963 23715
rect 5905 23675 5963 23681
rect 5368 23644 5396 23675
rect 5810 23644 5816 23656
rect 5368 23616 5816 23644
rect 5810 23604 5816 23616
rect 5868 23604 5874 23656
rect 5920 23644 5948 23675
rect 6362 23672 6368 23724
rect 6420 23712 6426 23724
rect 6457 23715 6515 23721
rect 6457 23712 6469 23715
rect 6420 23684 6469 23712
rect 6420 23672 6426 23684
rect 6457 23681 6469 23684
rect 6503 23681 6515 23715
rect 6638 23712 6644 23724
rect 6599 23684 6644 23712
rect 6457 23675 6515 23681
rect 6638 23672 6644 23684
rect 6696 23672 6702 23724
rect 7392 23721 7420 23752
rect 7926 23740 7932 23752
rect 7984 23740 7990 23792
rect 7009 23715 7067 23721
rect 7009 23681 7021 23715
rect 7055 23712 7067 23715
rect 7377 23715 7435 23721
rect 7055 23684 7328 23712
rect 7055 23681 7067 23684
rect 7009 23675 7067 23681
rect 7193 23647 7251 23653
rect 7193 23644 7205 23647
rect 5920 23616 7205 23644
rect 7193 23613 7205 23616
rect 7239 23613 7251 23647
rect 7300 23644 7328 23684
rect 7377 23681 7389 23715
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 7469 23715 7527 23721
rect 7469 23681 7481 23715
rect 7515 23712 7527 23715
rect 7742 23712 7748 23724
rect 7515 23684 7748 23712
rect 7515 23681 7527 23684
rect 7469 23675 7527 23681
rect 7484 23644 7512 23675
rect 7742 23672 7748 23684
rect 7800 23672 7806 23724
rect 7837 23715 7895 23721
rect 7837 23681 7849 23715
rect 7883 23712 7895 23715
rect 8018 23712 8024 23724
rect 7883 23684 8024 23712
rect 7883 23681 7895 23684
rect 7837 23675 7895 23681
rect 8018 23672 8024 23684
rect 8076 23672 8082 23724
rect 7300 23616 7512 23644
rect 7561 23647 7619 23653
rect 7193 23607 7251 23613
rect 7561 23613 7573 23647
rect 7607 23613 7619 23647
rect 7561 23607 7619 23613
rect 6181 23579 6239 23585
rect 6181 23545 6193 23579
rect 6227 23576 6239 23579
rect 7576 23576 7604 23607
rect 7650 23604 7656 23656
rect 7708 23644 7714 23656
rect 8312 23653 8340 23820
rect 8386 23808 8392 23860
rect 8444 23808 8450 23860
rect 10134 23848 10140 23860
rect 10095 23820 10140 23848
rect 10134 23808 10140 23820
rect 10192 23808 10198 23860
rect 11238 23808 11244 23860
rect 11296 23848 11302 23860
rect 11701 23851 11759 23857
rect 11701 23848 11713 23851
rect 11296 23820 11713 23848
rect 11296 23808 11302 23820
rect 11701 23817 11713 23820
rect 11747 23817 11759 23851
rect 11701 23811 11759 23817
rect 8404 23721 8432 23808
rect 9766 23780 9772 23792
rect 8956 23752 9772 23780
rect 8956 23724 8984 23752
rect 9766 23740 9772 23752
rect 9824 23780 9830 23792
rect 9953 23783 10011 23789
rect 9953 23780 9965 23783
rect 9824 23752 9965 23780
rect 9824 23740 9830 23752
rect 9953 23749 9965 23752
rect 9999 23749 10011 23783
rect 10962 23780 10968 23792
rect 9953 23743 10011 23749
rect 10428 23752 10968 23780
rect 8393 23715 8451 23721
rect 8393 23681 8405 23715
rect 8439 23681 8451 23715
rect 8662 23712 8668 23724
rect 8623 23684 8668 23712
rect 8393 23675 8451 23681
rect 8209 23647 8267 23653
rect 8209 23644 8221 23647
rect 7708 23616 7753 23644
rect 8128 23616 8221 23644
rect 7708 23604 7714 23616
rect 8018 23576 8024 23588
rect 6227 23548 8024 23576
rect 6227 23545 6239 23548
rect 6181 23539 6239 23545
rect 8018 23536 8024 23548
rect 8076 23536 8082 23588
rect 6730 23508 6736 23520
rect 6691 23480 6736 23508
rect 6730 23468 6736 23480
rect 6788 23468 6794 23520
rect 8128 23508 8156 23616
rect 8209 23613 8221 23616
rect 8255 23613 8267 23647
rect 8209 23607 8267 23613
rect 8297 23647 8355 23653
rect 8297 23613 8309 23647
rect 8343 23613 8355 23647
rect 8297 23607 8355 23613
rect 8404 23576 8432 23675
rect 8662 23672 8668 23684
rect 8720 23672 8726 23724
rect 8754 23672 8760 23724
rect 8812 23712 8818 23724
rect 8938 23712 8944 23724
rect 8812 23684 8857 23712
rect 8899 23684 8944 23712
rect 8812 23672 8818 23684
rect 8938 23672 8944 23684
rect 8996 23672 9002 23724
rect 9033 23715 9091 23721
rect 9033 23681 9045 23715
rect 9079 23681 9091 23715
rect 9033 23675 9091 23681
rect 8478 23604 8484 23656
rect 8536 23644 8542 23656
rect 9048 23644 9076 23675
rect 9122 23672 9128 23724
rect 9180 23712 9186 23724
rect 9585 23715 9643 23721
rect 9585 23712 9597 23715
rect 9180 23684 9597 23712
rect 9180 23672 9186 23684
rect 9585 23681 9597 23684
rect 9631 23681 9643 23715
rect 10134 23712 10140 23724
rect 10095 23684 10140 23712
rect 9585 23675 9643 23681
rect 10134 23672 10140 23684
rect 10192 23672 10198 23724
rect 10428 23721 10456 23752
rect 10962 23740 10968 23752
rect 11020 23740 11026 23792
rect 10413 23715 10471 23721
rect 10413 23681 10425 23715
rect 10459 23681 10471 23715
rect 10413 23675 10471 23681
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23681 10563 23715
rect 11054 23712 11060 23724
rect 11015 23684 11060 23712
rect 10505 23675 10563 23681
rect 9401 23647 9459 23653
rect 9401 23644 9413 23647
rect 8536 23616 8581 23644
rect 8956 23616 9413 23644
rect 8536 23604 8542 23616
rect 8956 23576 8984 23616
rect 9401 23613 9413 23616
rect 9447 23613 9459 23647
rect 9858 23644 9864 23656
rect 9771 23616 9864 23644
rect 9401 23607 9459 23613
rect 9858 23604 9864 23616
rect 9916 23644 9922 23656
rect 10520 23644 10548 23675
rect 11054 23672 11060 23684
rect 11112 23672 11118 23724
rect 11514 23712 11520 23724
rect 11475 23684 11520 23712
rect 11514 23672 11520 23684
rect 11572 23672 11578 23724
rect 11716 23712 11744 23811
rect 11882 23808 11888 23860
rect 11940 23848 11946 23860
rect 11977 23851 12035 23857
rect 11977 23848 11989 23851
rect 11940 23820 11989 23848
rect 11940 23808 11946 23820
rect 11977 23817 11989 23820
rect 12023 23817 12035 23851
rect 12250 23848 12256 23860
rect 12211 23820 12256 23848
rect 11977 23811 12035 23817
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 13262 23848 13268 23860
rect 13223 23820 13268 23848
rect 13262 23808 13268 23820
rect 13320 23808 13326 23860
rect 17034 23848 17040 23860
rect 16995 23820 17040 23848
rect 17034 23808 17040 23820
rect 17092 23808 17098 23860
rect 18966 23848 18972 23860
rect 18432 23820 18972 23848
rect 12897 23783 12955 23789
rect 12897 23780 12909 23783
rect 12176 23752 12909 23780
rect 12176 23721 12204 23752
rect 12897 23749 12909 23752
rect 12943 23749 12955 23783
rect 12897 23743 12955 23749
rect 15102 23740 15108 23792
rect 15160 23780 15166 23792
rect 15841 23783 15899 23789
rect 15841 23780 15853 23783
rect 15160 23752 15853 23780
rect 15160 23740 15166 23752
rect 15841 23749 15853 23752
rect 15887 23749 15899 23783
rect 15841 23743 15899 23749
rect 16022 23740 16028 23792
rect 16080 23780 16086 23792
rect 16255 23783 16313 23789
rect 16255 23780 16267 23783
rect 16080 23752 16267 23780
rect 16080 23740 16086 23752
rect 16255 23749 16267 23752
rect 16301 23780 16313 23783
rect 18046 23780 18052 23792
rect 16301 23752 18052 23780
rect 16301 23749 16313 23752
rect 16255 23743 16313 23749
rect 18046 23740 18052 23752
rect 18104 23740 18110 23792
rect 12161 23715 12219 23721
rect 12161 23712 12173 23715
rect 11716 23684 12173 23712
rect 12161 23681 12173 23684
rect 12207 23681 12219 23715
rect 12161 23675 12219 23681
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23712 12495 23715
rect 13262 23712 13268 23724
rect 12483 23684 13268 23712
rect 12483 23681 12495 23684
rect 12437 23675 12495 23681
rect 13262 23672 13268 23684
rect 13320 23672 13326 23724
rect 16485 23715 16543 23721
rect 16485 23681 16497 23715
rect 16531 23712 16543 23715
rect 16853 23715 16911 23721
rect 16853 23712 16865 23715
rect 16531 23684 16865 23712
rect 16531 23681 16543 23684
rect 16485 23675 16543 23681
rect 16853 23681 16865 23684
rect 16899 23681 16911 23715
rect 17494 23712 17500 23724
rect 17455 23684 17500 23712
rect 16853 23675 16911 23681
rect 17494 23672 17500 23684
rect 17552 23672 17558 23724
rect 18432 23721 18460 23820
rect 18966 23808 18972 23820
rect 19024 23848 19030 23860
rect 19024 23820 20852 23848
rect 19024 23808 19030 23820
rect 18506 23740 18512 23792
rect 18564 23780 18570 23792
rect 20824 23789 20852 23820
rect 20625 23783 20683 23789
rect 20625 23780 20637 23783
rect 18564 23752 20637 23780
rect 18564 23740 18570 23752
rect 20625 23749 20637 23752
rect 20671 23749 20683 23783
rect 20625 23743 20683 23749
rect 20809 23783 20867 23789
rect 20809 23749 20821 23783
rect 20855 23749 20867 23783
rect 20809 23743 20867 23749
rect 17589 23715 17647 23721
rect 17589 23681 17601 23715
rect 17635 23712 17647 23715
rect 18141 23715 18199 23721
rect 18141 23712 18153 23715
rect 17635 23684 18153 23712
rect 17635 23681 17647 23684
rect 17589 23675 17647 23681
rect 18141 23681 18153 23684
rect 18187 23681 18199 23715
rect 18141 23675 18199 23681
rect 18383 23715 18460 23721
rect 18383 23681 18395 23715
rect 18429 23684 18460 23715
rect 18429 23681 18441 23684
rect 18383 23675 18441 23681
rect 18598 23672 18604 23724
rect 18656 23712 18662 23724
rect 19150 23721 19156 23724
rect 18785 23715 18843 23721
rect 18785 23712 18797 23715
rect 18656 23684 18797 23712
rect 18656 23672 18662 23684
rect 18699 23682 18736 23684
rect 18785 23681 18797 23684
rect 18831 23681 18843 23715
rect 18785 23675 18843 23681
rect 19144 23675 19156 23721
rect 19208 23712 19214 23724
rect 20438 23712 20444 23724
rect 19208 23684 19244 23712
rect 20399 23684 20444 23712
rect 19150 23672 19156 23675
rect 19208 23672 19214 23684
rect 20438 23672 20444 23684
rect 20496 23672 20502 23724
rect 12618 23644 12624 23656
rect 9916 23616 10548 23644
rect 12579 23616 12624 23644
rect 9916 23604 9922 23616
rect 12618 23604 12624 23616
rect 12676 23604 12682 23656
rect 12805 23647 12863 23653
rect 12805 23613 12817 23647
rect 12851 23644 12863 23647
rect 14458 23644 14464 23656
rect 12851 23616 14464 23644
rect 12851 23613 12863 23616
rect 12805 23607 12863 23613
rect 14458 23604 14464 23616
rect 14516 23604 14522 23656
rect 16390 23644 16396 23656
rect 15672 23616 16396 23644
rect 8404 23548 8984 23576
rect 15672 23520 15700 23616
rect 16390 23604 16396 23616
rect 16448 23644 16454 23656
rect 16669 23647 16727 23653
rect 16669 23644 16681 23647
rect 16448 23616 16681 23644
rect 16448 23604 16454 23616
rect 16669 23613 16681 23616
rect 16715 23644 16727 23647
rect 17681 23647 17739 23653
rect 17681 23644 17693 23647
rect 16715 23616 17693 23644
rect 16715 23613 16727 23616
rect 16669 23607 16727 23613
rect 17681 23613 17693 23616
rect 17727 23613 17739 23647
rect 17681 23607 17739 23613
rect 17129 23579 17187 23585
rect 17129 23576 17141 23579
rect 16224 23548 17141 23576
rect 8846 23508 8852 23520
rect 8128 23480 8852 23508
rect 8846 23468 8852 23480
rect 8904 23468 8910 23520
rect 8938 23468 8944 23520
rect 8996 23508 9002 23520
rect 9217 23511 9275 23517
rect 9217 23508 9229 23511
rect 8996 23480 9229 23508
rect 8996 23468 9002 23480
rect 9217 23477 9229 23480
rect 9263 23477 9275 23511
rect 10594 23508 10600 23520
rect 10555 23480 10600 23508
rect 9217 23471 9275 23477
rect 10594 23468 10600 23480
rect 10652 23468 10658 23520
rect 10873 23511 10931 23517
rect 10873 23477 10885 23511
rect 10919 23508 10931 23511
rect 10962 23508 10968 23520
rect 10919 23480 10968 23508
rect 10919 23477 10931 23480
rect 10873 23471 10931 23477
rect 10962 23468 10968 23480
rect 11020 23468 11026 23520
rect 11146 23468 11152 23520
rect 11204 23508 11210 23520
rect 11241 23511 11299 23517
rect 11241 23508 11253 23511
rect 11204 23480 11253 23508
rect 11204 23468 11210 23480
rect 11241 23477 11253 23480
rect 11287 23477 11299 23511
rect 15654 23508 15660 23520
rect 15615 23480 15660 23508
rect 11241 23471 11299 23477
rect 15654 23468 15660 23480
rect 15712 23468 15718 23520
rect 16224 23517 16252 23548
rect 17129 23545 17141 23548
rect 17175 23545 17187 23579
rect 17129 23539 17187 23545
rect 16209 23511 16267 23517
rect 16209 23477 16221 23511
rect 16255 23477 16267 23511
rect 17696 23508 17724 23607
rect 18506 23604 18512 23656
rect 18564 23644 18570 23656
rect 18693 23647 18751 23653
rect 18693 23644 18705 23647
rect 18564 23616 18705 23644
rect 18564 23604 18570 23616
rect 18693 23613 18705 23616
rect 18739 23613 18751 23647
rect 18874 23644 18880 23656
rect 18835 23616 18880 23644
rect 18693 23607 18751 23613
rect 18874 23604 18880 23616
rect 18932 23604 18938 23656
rect 19242 23508 19248 23520
rect 17696 23480 19248 23508
rect 16209 23471 16267 23477
rect 19242 23468 19248 23480
rect 19300 23468 19306 23520
rect 19518 23468 19524 23520
rect 19576 23508 19582 23520
rect 20257 23511 20315 23517
rect 20257 23508 20269 23511
rect 19576 23480 20269 23508
rect 19576 23468 19582 23480
rect 20257 23477 20269 23480
rect 20303 23477 20315 23511
rect 20257 23471 20315 23477
rect 1104 23418 26128 23440
rect 1104 23366 5120 23418
rect 5172 23366 5184 23418
rect 5236 23366 5248 23418
rect 5300 23366 5312 23418
rect 5364 23366 5376 23418
rect 5428 23366 13462 23418
rect 13514 23366 13526 23418
rect 13578 23366 13590 23418
rect 13642 23366 13654 23418
rect 13706 23366 13718 23418
rect 13770 23366 21803 23418
rect 21855 23366 21867 23418
rect 21919 23366 21931 23418
rect 21983 23366 21995 23418
rect 22047 23366 22059 23418
rect 22111 23366 26128 23418
rect 1104 23344 26128 23366
rect 5810 23264 5816 23316
rect 5868 23304 5874 23316
rect 7193 23307 7251 23313
rect 7193 23304 7205 23307
rect 5868 23276 7205 23304
rect 5868 23264 5874 23276
rect 7193 23273 7205 23276
rect 7239 23273 7251 23307
rect 7742 23304 7748 23316
rect 7193 23267 7251 23273
rect 7484 23276 7748 23304
rect 6733 23239 6791 23245
rect 6733 23205 6745 23239
rect 6779 23236 6791 23239
rect 7484 23236 7512 23276
rect 7742 23264 7748 23276
rect 7800 23304 7806 23316
rect 8110 23304 8116 23316
rect 7800 23276 8116 23304
rect 7800 23264 7806 23276
rect 8110 23264 8116 23276
rect 8168 23264 8174 23316
rect 8478 23304 8484 23316
rect 8439 23276 8484 23304
rect 8478 23264 8484 23276
rect 8536 23264 8542 23316
rect 14182 23304 14188 23316
rect 14143 23276 14188 23304
rect 14182 23264 14188 23276
rect 14240 23264 14246 23316
rect 16574 23304 16580 23316
rect 16535 23276 16580 23304
rect 16574 23264 16580 23276
rect 16632 23264 16638 23316
rect 18693 23307 18751 23313
rect 18693 23273 18705 23307
rect 18739 23304 18751 23307
rect 19245 23307 19303 23313
rect 19245 23304 19257 23307
rect 18739 23276 19257 23304
rect 18739 23273 18751 23276
rect 18693 23267 18751 23273
rect 19245 23273 19257 23276
rect 19291 23273 19303 23307
rect 19245 23267 19303 23273
rect 6779 23208 7512 23236
rect 6779 23205 6791 23208
rect 6733 23199 6791 23205
rect 7484 23177 7512 23208
rect 8021 23239 8079 23245
rect 8021 23205 8033 23239
rect 8067 23236 8079 23239
rect 8754 23236 8760 23248
rect 8067 23208 8760 23236
rect 8067 23205 8079 23208
rect 8021 23199 8079 23205
rect 7469 23171 7527 23177
rect 7469 23137 7481 23171
rect 7515 23137 7527 23171
rect 7469 23131 7527 23137
rect 7561 23171 7619 23177
rect 7561 23137 7573 23171
rect 7607 23168 7619 23171
rect 7742 23168 7748 23180
rect 7607 23140 7748 23168
rect 7607 23137 7619 23140
rect 7561 23131 7619 23137
rect 7742 23128 7748 23140
rect 7800 23128 7806 23180
rect 8036 23168 8064 23199
rect 8754 23196 8760 23208
rect 8812 23196 8818 23248
rect 10229 23239 10287 23245
rect 10229 23205 10241 23239
rect 10275 23236 10287 23239
rect 11514 23236 11520 23248
rect 10275 23208 11520 23236
rect 10275 23205 10287 23208
rect 10229 23199 10287 23205
rect 11514 23196 11520 23208
rect 11572 23196 11578 23248
rect 13449 23239 13507 23245
rect 13449 23205 13461 23239
rect 13495 23236 13507 23239
rect 16022 23236 16028 23248
rect 13495 23208 16028 23236
rect 13495 23205 13507 23208
rect 13449 23199 13507 23205
rect 16022 23196 16028 23208
rect 16080 23196 16086 23248
rect 18506 23196 18512 23248
rect 18564 23236 18570 23248
rect 18874 23236 18880 23248
rect 18564 23208 18880 23236
rect 18564 23196 18570 23208
rect 18874 23196 18880 23208
rect 18932 23236 18938 23248
rect 18932 23208 20576 23236
rect 18932 23196 18938 23208
rect 7852 23140 8064 23168
rect 2130 23100 2136 23112
rect 2091 23072 2136 23100
rect 2130 23060 2136 23072
rect 2188 23060 2194 23112
rect 6730 23060 6736 23112
rect 6788 23100 6794 23112
rect 6825 23103 6883 23109
rect 6825 23100 6837 23103
rect 6788 23072 6837 23100
rect 6788 23060 6794 23072
rect 6825 23069 6837 23072
rect 6871 23069 6883 23103
rect 7374 23100 7380 23112
rect 7335 23072 7380 23100
rect 6825 23063 6883 23069
rect 7374 23060 7380 23072
rect 7432 23060 7438 23112
rect 7650 23100 7656 23112
rect 7611 23072 7656 23100
rect 7650 23060 7656 23072
rect 7708 23060 7714 23112
rect 7852 23109 7880 23140
rect 8294 23128 8300 23180
rect 8352 23168 8358 23180
rect 15289 23171 15347 23177
rect 8352 23140 9168 23168
rect 8352 23128 8358 23140
rect 7837 23103 7895 23109
rect 7837 23069 7849 23103
rect 7883 23069 7895 23103
rect 7837 23063 7895 23069
rect 7929 23103 7987 23109
rect 7929 23069 7941 23103
rect 7975 23100 7987 23103
rect 8202 23100 8208 23112
rect 7975 23072 8208 23100
rect 7975 23069 7987 23072
rect 7929 23063 7987 23069
rect 7098 22992 7104 23044
rect 7156 23032 7162 23044
rect 7944 23032 7972 23063
rect 8202 23060 8208 23072
rect 8260 23060 8266 23112
rect 8570 23060 8576 23112
rect 8628 23100 8634 23112
rect 9140 23109 9168 23140
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 15749 23171 15807 23177
rect 15749 23168 15761 23171
rect 15335 23140 15761 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 15749 23137 15761 23140
rect 15795 23168 15807 23171
rect 15933 23171 15991 23177
rect 15933 23168 15945 23171
rect 15795 23140 15945 23168
rect 15795 23137 15807 23140
rect 15749 23131 15807 23137
rect 15933 23137 15945 23140
rect 15979 23168 15991 23171
rect 16666 23168 16672 23180
rect 15979 23140 16672 23168
rect 15979 23137 15991 23140
rect 15933 23131 15991 23137
rect 16666 23128 16672 23140
rect 16724 23168 16730 23180
rect 17313 23171 17371 23177
rect 17313 23168 17325 23171
rect 16724 23140 17325 23168
rect 16724 23128 16730 23140
rect 17313 23137 17325 23140
rect 17359 23137 17371 23171
rect 18690 23168 18696 23180
rect 17313 23131 17371 23137
rect 18064 23140 18696 23168
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8628 23072 8953 23100
rect 8628 23060 8634 23072
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 8941 23063 8999 23069
rect 9125 23103 9183 23109
rect 9125 23069 9137 23103
rect 9171 23069 9183 23103
rect 9125 23063 9183 23069
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23069 9551 23103
rect 9766 23100 9772 23112
rect 9727 23072 9772 23100
rect 9493 23063 9551 23069
rect 8294 23032 8300 23044
rect 7156 23004 7972 23032
rect 8255 23004 8300 23032
rect 7156 22992 7162 23004
rect 8294 22992 8300 23004
rect 8352 22992 8358 23044
rect 8481 23035 8539 23041
rect 8481 23001 8493 23035
rect 8527 23032 8539 23035
rect 9214 23032 9220 23044
rect 8527 23004 9220 23032
rect 8527 23001 8539 23004
rect 8481 22995 8539 23001
rect 9214 22992 9220 23004
rect 9272 23032 9278 23044
rect 9508 23032 9536 23063
rect 9766 23060 9772 23072
rect 9824 23060 9830 23112
rect 9858 23060 9864 23112
rect 9916 23100 9922 23112
rect 13262 23100 13268 23112
rect 9916 23072 9961 23100
rect 13223 23072 13268 23100
rect 9916 23060 9922 23072
rect 13262 23060 13268 23072
rect 13320 23060 13326 23112
rect 14369 23103 14427 23109
rect 14369 23069 14381 23103
rect 14415 23100 14427 23103
rect 18064 23100 18092 23140
rect 18690 23128 18696 23140
rect 18748 23128 18754 23180
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 19797 23171 19855 23177
rect 19797 23168 19809 23171
rect 19392 23140 19809 23168
rect 19392 23128 19398 23140
rect 19797 23137 19809 23140
rect 19843 23168 19855 23171
rect 19843 23140 20208 23168
rect 19843 23137 19855 23140
rect 19797 23131 19855 23137
rect 14415 23072 18092 23100
rect 18141 23103 18199 23109
rect 14415 23069 14427 23072
rect 14369 23063 14427 23069
rect 18141 23069 18153 23103
rect 18187 23100 18199 23103
rect 18417 23103 18475 23109
rect 18417 23100 18429 23103
rect 18187 23072 18429 23100
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 18417 23069 18429 23072
rect 18463 23069 18475 23103
rect 19886 23100 19892 23112
rect 18417 23063 18475 23069
rect 18708 23072 19892 23100
rect 9677 23035 9735 23041
rect 9677 23032 9689 23035
rect 9272 23004 9689 23032
rect 9272 22992 9278 23004
rect 9677 23001 9689 23004
rect 9723 23001 9735 23035
rect 10042 23032 10048 23044
rect 10003 23004 10048 23032
rect 9677 22995 9735 23001
rect 10042 22992 10048 23004
rect 10100 22992 10106 23044
rect 11882 22992 11888 23044
rect 11940 23032 11946 23044
rect 14384 23032 14412 23063
rect 14642 23032 14648 23044
rect 11940 23004 14412 23032
rect 14603 23004 14648 23032
rect 11940 22992 11946 23004
rect 14642 22992 14648 23004
rect 14700 22992 14706 23044
rect 14829 23035 14887 23041
rect 14829 23001 14841 23035
rect 14875 23032 14887 23035
rect 16850 23032 16856 23044
rect 14875 23004 16856 23032
rect 14875 23001 14887 23004
rect 14829 22995 14887 23001
rect 16850 22992 16856 23004
rect 16908 22992 16914 23044
rect 18046 22992 18052 23044
rect 18104 23032 18110 23044
rect 18708 23041 18736 23072
rect 19886 23060 19892 23072
rect 19944 23060 19950 23112
rect 18684 23035 18742 23041
rect 18684 23032 18696 23035
rect 18104 23004 18696 23032
rect 18104 22992 18110 23004
rect 18684 23001 18696 23004
rect 18730 23001 18742 23035
rect 18684 22995 18742 23001
rect 19061 23035 19119 23041
rect 19061 23001 19073 23035
rect 19107 23032 19119 23035
rect 19334 23032 19340 23044
rect 19107 23004 19340 23032
rect 19107 23001 19119 23004
rect 19061 22995 19119 23001
rect 19334 22992 19340 23004
rect 19392 22992 19398 23044
rect 19613 23035 19671 23041
rect 19613 23001 19625 23035
rect 19659 23032 19671 23035
rect 19978 23032 19984 23044
rect 19659 23004 19984 23032
rect 19659 23001 19671 23004
rect 19613 22995 19671 23001
rect 19978 22992 19984 23004
rect 20036 22992 20042 23044
rect 6270 22924 6276 22976
rect 6328 22964 6334 22976
rect 6457 22967 6515 22973
rect 6457 22964 6469 22967
rect 6328 22936 6469 22964
rect 6328 22924 6334 22936
rect 6457 22933 6469 22936
rect 6503 22964 6515 22967
rect 6638 22964 6644 22976
rect 6503 22936 6644 22964
rect 6503 22933 6515 22936
rect 6457 22927 6515 22933
rect 6638 22924 6644 22936
rect 6696 22924 6702 22976
rect 7006 22964 7012 22976
rect 6967 22936 7012 22964
rect 7006 22924 7012 22936
rect 7064 22924 7070 22976
rect 8570 22924 8576 22976
rect 8628 22964 8634 22976
rect 8665 22967 8723 22973
rect 8665 22964 8677 22967
rect 8628 22936 8677 22964
rect 8628 22924 8634 22936
rect 8665 22933 8677 22936
rect 8711 22933 8723 22967
rect 8665 22927 8723 22933
rect 8754 22924 8760 22976
rect 8812 22964 8818 22976
rect 9125 22967 9183 22973
rect 9125 22964 9137 22967
rect 8812 22936 9137 22964
rect 8812 22924 8818 22936
rect 9125 22933 9137 22936
rect 9171 22933 9183 22967
rect 9125 22927 9183 22933
rect 9766 22924 9772 22976
rect 9824 22964 9830 22976
rect 10778 22964 10784 22976
rect 9824 22936 10784 22964
rect 9824 22924 9830 22936
rect 10778 22924 10784 22936
rect 10836 22924 10842 22976
rect 11330 22924 11336 22976
rect 11388 22964 11394 22976
rect 12437 22967 12495 22973
rect 12437 22964 12449 22967
rect 11388 22936 12449 22964
rect 11388 22924 11394 22936
rect 12437 22933 12449 22936
rect 12483 22964 12495 22967
rect 12618 22964 12624 22976
rect 12483 22936 12624 22964
rect 12483 22933 12495 22936
rect 12437 22927 12495 22933
rect 12618 22924 12624 22936
rect 12676 22964 12682 22976
rect 13354 22964 13360 22976
rect 12676 22936 13360 22964
rect 12676 22924 12682 22936
rect 13354 22924 13360 22936
rect 13412 22924 13418 22976
rect 14550 22964 14556 22976
rect 14511 22936 14556 22964
rect 14550 22924 14556 22936
rect 14608 22924 14614 22976
rect 16114 22964 16120 22976
rect 16075 22936 16120 22964
rect 16114 22924 16120 22936
rect 16172 22924 16178 22976
rect 16206 22924 16212 22976
rect 16264 22964 16270 22976
rect 18325 22967 18383 22973
rect 16264 22936 16309 22964
rect 16264 22924 16270 22936
rect 18325 22933 18337 22967
rect 18371 22964 18383 22967
rect 19150 22964 19156 22976
rect 18371 22936 19156 22964
rect 18371 22933 18383 22936
rect 18325 22927 18383 22933
rect 19150 22924 19156 22936
rect 19208 22924 19214 22976
rect 19702 22924 19708 22976
rect 19760 22964 19766 22976
rect 20180 22973 20208 23140
rect 20257 23103 20315 23109
rect 20257 23069 20269 23103
rect 20303 23100 20315 23103
rect 20346 23100 20352 23112
rect 20303 23072 20352 23100
rect 20303 23069 20315 23072
rect 20257 23063 20315 23069
rect 20346 23060 20352 23072
rect 20404 23060 20410 23112
rect 20548 23109 20576 23208
rect 20533 23103 20591 23109
rect 20533 23069 20545 23103
rect 20579 23100 20591 23103
rect 22097 23103 22155 23109
rect 22097 23100 22109 23103
rect 20579 23072 22109 23100
rect 20579 23069 20591 23072
rect 20533 23063 20591 23069
rect 22097 23069 22109 23072
rect 22143 23100 22155 23103
rect 23382 23100 23388 23112
rect 22143 23072 23388 23100
rect 22143 23069 22155 23072
rect 22097 23063 22155 23069
rect 23382 23060 23388 23072
rect 23440 23060 23446 23112
rect 20778 23035 20836 23041
rect 20778 23032 20790 23035
rect 20456 23004 20790 23032
rect 20165 22967 20223 22973
rect 19760 22936 19805 22964
rect 19760 22924 19766 22936
rect 20165 22933 20177 22967
rect 20211 22964 20223 22967
rect 20254 22964 20260 22976
rect 20211 22936 20260 22964
rect 20211 22933 20223 22936
rect 20165 22927 20223 22933
rect 20254 22924 20260 22936
rect 20312 22924 20318 22976
rect 20456 22973 20484 23004
rect 20778 23001 20790 23004
rect 20824 23001 20836 23035
rect 20778 22995 20836 23001
rect 22186 22992 22192 23044
rect 22244 23032 22250 23044
rect 22342 23035 22400 23041
rect 22342 23032 22354 23035
rect 22244 23004 22354 23032
rect 22244 22992 22250 23004
rect 22342 23001 22354 23004
rect 22388 23001 22400 23035
rect 22342 22995 22400 23001
rect 20441 22967 20499 22973
rect 20441 22933 20453 22967
rect 20487 22933 20499 22967
rect 20441 22927 20499 22933
rect 21913 22967 21971 22973
rect 21913 22933 21925 22967
rect 21959 22964 21971 22967
rect 22094 22964 22100 22976
rect 21959 22936 22100 22964
rect 21959 22933 21971 22936
rect 21913 22927 21971 22933
rect 22094 22924 22100 22936
rect 22152 22964 22158 22976
rect 23198 22964 23204 22976
rect 22152 22936 23204 22964
rect 22152 22924 22158 22936
rect 23198 22924 23204 22936
rect 23256 22924 23262 22976
rect 23474 22964 23480 22976
rect 23435 22936 23480 22964
rect 23474 22924 23480 22936
rect 23532 22924 23538 22976
rect 1104 22874 26128 22896
rect 1104 22822 9291 22874
rect 9343 22822 9355 22874
rect 9407 22822 9419 22874
rect 9471 22822 9483 22874
rect 9535 22822 9547 22874
rect 9599 22822 17632 22874
rect 17684 22822 17696 22874
rect 17748 22822 17760 22874
rect 17812 22822 17824 22874
rect 17876 22822 17888 22874
rect 17940 22822 26128 22874
rect 1104 22800 26128 22822
rect 7006 22720 7012 22772
rect 7064 22760 7070 22772
rect 7193 22763 7251 22769
rect 7193 22760 7205 22763
rect 7064 22732 7205 22760
rect 7064 22720 7070 22732
rect 7193 22729 7205 22732
rect 7239 22729 7251 22763
rect 7193 22723 7251 22729
rect 7374 22720 7380 22772
rect 7432 22760 7438 22772
rect 7653 22763 7711 22769
rect 7653 22760 7665 22763
rect 7432 22732 7665 22760
rect 7432 22720 7438 22732
rect 7653 22729 7665 22732
rect 7699 22729 7711 22763
rect 8294 22760 8300 22772
rect 8255 22732 8300 22760
rect 7653 22723 7711 22729
rect 8294 22720 8300 22732
rect 8352 22720 8358 22772
rect 9033 22763 9091 22769
rect 9033 22729 9045 22763
rect 9079 22760 9091 22763
rect 10134 22760 10140 22772
rect 9079 22732 10140 22760
rect 9079 22729 9091 22732
rect 9033 22723 9091 22729
rect 10134 22720 10140 22732
rect 10192 22720 10198 22772
rect 14274 22720 14280 22772
rect 14332 22760 14338 22772
rect 14461 22763 14519 22769
rect 14461 22760 14473 22763
rect 14332 22732 14473 22760
rect 14332 22720 14338 22732
rect 14461 22729 14473 22732
rect 14507 22729 14519 22763
rect 14461 22723 14519 22729
rect 15289 22763 15347 22769
rect 15289 22729 15301 22763
rect 15335 22760 15347 22763
rect 15749 22763 15807 22769
rect 15749 22760 15761 22763
rect 15335 22732 15761 22760
rect 15335 22729 15347 22732
rect 15289 22723 15347 22729
rect 15749 22729 15761 22732
rect 15795 22729 15807 22763
rect 15749 22723 15807 22729
rect 16114 22720 16120 22772
rect 16172 22760 16178 22772
rect 17037 22763 17095 22769
rect 17037 22760 17049 22763
rect 16172 22732 17049 22760
rect 16172 22720 16178 22732
rect 17037 22729 17049 22732
rect 17083 22729 17095 22763
rect 17494 22760 17500 22772
rect 17455 22732 17500 22760
rect 17037 22723 17095 22729
rect 17494 22720 17500 22732
rect 17552 22720 17558 22772
rect 17865 22763 17923 22769
rect 17865 22760 17877 22763
rect 17604 22732 17877 22760
rect 7098 22652 7104 22704
rect 7156 22692 7162 22704
rect 7285 22695 7343 22701
rect 7285 22692 7297 22695
rect 7156 22664 7297 22692
rect 7156 22652 7162 22664
rect 7285 22661 7297 22664
rect 7331 22661 7343 22695
rect 7285 22655 7343 22661
rect 8849 22695 8907 22701
rect 8849 22661 8861 22695
rect 8895 22692 8907 22695
rect 10045 22695 10103 22701
rect 10045 22692 10057 22695
rect 8895 22664 10057 22692
rect 8895 22661 8907 22664
rect 8849 22655 8907 22661
rect 10045 22661 10057 22664
rect 10091 22692 10103 22695
rect 10505 22695 10563 22701
rect 10505 22692 10517 22695
rect 10091 22664 10517 22692
rect 10091 22661 10103 22664
rect 10045 22655 10103 22661
rect 10505 22661 10517 22664
rect 10551 22661 10563 22695
rect 10505 22655 10563 22661
rect 13832 22664 16068 22692
rect 3970 22584 3976 22636
rect 4028 22624 4034 22636
rect 4065 22627 4123 22633
rect 4065 22624 4077 22627
rect 4028 22596 4077 22624
rect 4028 22584 4034 22596
rect 4065 22593 4077 22596
rect 4111 22593 4123 22627
rect 7834 22624 7840 22636
rect 7795 22596 7840 22624
rect 4065 22587 4123 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 8386 22624 8392 22636
rect 8347 22596 8392 22624
rect 8386 22584 8392 22596
rect 8444 22584 8450 22636
rect 8570 22624 8576 22636
rect 8531 22596 8576 22624
rect 8570 22584 8576 22596
rect 8628 22584 8634 22636
rect 8754 22624 8760 22636
rect 8715 22596 8760 22624
rect 8754 22584 8760 22596
rect 8812 22584 8818 22636
rect 9214 22624 9220 22636
rect 9175 22596 9220 22624
rect 9214 22584 9220 22596
rect 9272 22584 9278 22636
rect 9309 22627 9367 22633
rect 9309 22593 9321 22627
rect 9355 22624 9367 22627
rect 9766 22624 9772 22636
rect 9355 22596 9772 22624
rect 9355 22593 9367 22596
rect 9309 22587 9367 22593
rect 9766 22584 9772 22596
rect 9824 22584 9830 22636
rect 10686 22624 10692 22636
rect 10647 22596 10692 22624
rect 10686 22584 10692 22596
rect 10744 22584 10750 22636
rect 11882 22624 11888 22636
rect 11843 22596 11888 22624
rect 11882 22584 11888 22596
rect 11940 22584 11946 22636
rect 13354 22584 13360 22636
rect 13412 22624 13418 22636
rect 13832 22624 13860 22664
rect 14090 22624 14096 22636
rect 13412 22596 13860 22624
rect 14051 22596 14096 22624
rect 13412 22584 13418 22596
rect 4249 22559 4307 22565
rect 4249 22525 4261 22559
rect 4295 22556 4307 22559
rect 4338 22556 4344 22568
rect 4295 22528 4344 22556
rect 4295 22525 4307 22528
rect 4249 22519 4307 22525
rect 4338 22516 4344 22528
rect 4396 22516 4402 22568
rect 7101 22559 7159 22565
rect 7101 22525 7113 22559
rect 7147 22556 7159 22559
rect 7147 22528 8248 22556
rect 7147 22525 7159 22528
rect 7101 22519 7159 22525
rect 8220 22500 8248 22528
rect 9122 22516 9128 22568
rect 9180 22556 9186 22568
rect 9585 22559 9643 22565
rect 9585 22556 9597 22559
rect 9180 22528 9597 22556
rect 9180 22516 9186 22528
rect 9585 22525 9597 22528
rect 9631 22525 9643 22559
rect 10134 22556 10140 22568
rect 10095 22528 10140 22556
rect 9585 22519 9643 22525
rect 10134 22516 10140 22528
rect 10192 22516 10198 22568
rect 10318 22516 10324 22568
rect 10376 22556 10382 22568
rect 10594 22556 10600 22568
rect 10376 22528 10600 22556
rect 10376 22516 10382 22528
rect 10594 22516 10600 22528
rect 10652 22556 10658 22568
rect 13832 22565 13860 22596
rect 14090 22584 14096 22596
rect 14148 22584 14154 22636
rect 14921 22627 14979 22633
rect 14921 22593 14933 22627
rect 14967 22624 14979 22627
rect 15194 22624 15200 22636
rect 14967 22596 15200 22624
rect 14967 22593 14979 22596
rect 14921 22587 14979 22593
rect 15194 22584 15200 22596
rect 15252 22584 15258 22636
rect 16040 22624 16068 22664
rect 17402 22652 17408 22704
rect 17460 22692 17466 22704
rect 17604 22692 17632 22732
rect 17865 22729 17877 22732
rect 17911 22729 17923 22763
rect 17865 22723 17923 22729
rect 19521 22763 19579 22769
rect 19521 22729 19533 22763
rect 19567 22760 19579 22763
rect 19702 22760 19708 22772
rect 19567 22732 19708 22760
rect 19567 22729 19579 22732
rect 19521 22723 19579 22729
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 19886 22720 19892 22772
rect 19944 22760 19950 22772
rect 20082 22763 20140 22769
rect 20082 22760 20094 22763
rect 19944 22732 20094 22760
rect 19944 22720 19950 22732
rect 20082 22729 20094 22732
rect 20128 22729 20140 22763
rect 22186 22760 22192 22772
rect 22147 22732 22192 22760
rect 20082 22723 20140 22729
rect 22186 22720 22192 22732
rect 22244 22720 22250 22772
rect 22741 22763 22799 22769
rect 22741 22729 22753 22763
rect 22787 22760 22799 22763
rect 24854 22760 24860 22772
rect 22787 22732 24860 22760
rect 22787 22729 22799 22732
rect 22741 22723 22799 22729
rect 24854 22720 24860 22732
rect 24912 22720 24918 22772
rect 17460 22664 17632 22692
rect 17460 22652 17466 22664
rect 17770 22652 17776 22704
rect 17828 22692 17834 22704
rect 18417 22695 18475 22701
rect 18417 22692 18429 22695
rect 17828 22664 18429 22692
rect 17828 22652 17834 22664
rect 18417 22661 18429 22664
rect 18463 22661 18475 22695
rect 19610 22692 19616 22704
rect 18417 22655 18475 22661
rect 19536 22664 19616 22692
rect 16666 22624 16672 22636
rect 16040 22596 16672 22624
rect 11241 22559 11299 22565
rect 11241 22556 11253 22559
rect 10652 22528 11253 22556
rect 10652 22516 10658 22528
rect 11241 22525 11253 22528
rect 11287 22556 11299 22559
rect 13633 22559 13691 22565
rect 11287 22528 13492 22556
rect 11287 22525 11299 22528
rect 11241 22519 11299 22525
rect 8202 22448 8208 22500
rect 8260 22488 8266 22500
rect 8260 22460 9904 22488
rect 8260 22448 8266 22460
rect 3694 22380 3700 22432
rect 3752 22420 3758 22432
rect 3881 22423 3939 22429
rect 3881 22420 3893 22423
rect 3752 22392 3893 22420
rect 3752 22380 3758 22392
rect 3881 22389 3893 22392
rect 3927 22389 3939 22423
rect 3881 22383 3939 22389
rect 6822 22380 6828 22432
rect 6880 22420 6886 22432
rect 7929 22423 7987 22429
rect 7929 22420 7941 22423
rect 6880 22392 7941 22420
rect 6880 22380 6886 22392
rect 7929 22389 7941 22392
rect 7975 22389 7987 22423
rect 9490 22420 9496 22432
rect 9451 22392 9496 22420
rect 7929 22383 7987 22389
rect 9490 22380 9496 22392
rect 9548 22380 9554 22432
rect 9677 22423 9735 22429
rect 9677 22389 9689 22423
rect 9723 22420 9735 22423
rect 9766 22420 9772 22432
rect 9723 22392 9772 22420
rect 9723 22389 9735 22392
rect 9677 22383 9735 22389
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 9876 22420 9904 22460
rect 10686 22448 10692 22500
rect 10744 22488 10750 22500
rect 11057 22491 11115 22497
rect 11057 22488 11069 22491
rect 10744 22460 11069 22488
rect 10744 22448 10750 22460
rect 11057 22457 11069 22460
rect 11103 22488 11115 22491
rect 13464 22488 13492 22528
rect 13633 22525 13645 22559
rect 13679 22556 13691 22559
rect 13817 22559 13875 22565
rect 13817 22556 13829 22559
rect 13679 22528 13829 22556
rect 13679 22525 13691 22528
rect 13633 22519 13691 22525
rect 13817 22525 13829 22528
rect 13863 22525 13875 22559
rect 13817 22519 13875 22525
rect 13906 22516 13912 22568
rect 13964 22556 13970 22568
rect 14001 22559 14059 22565
rect 14001 22556 14013 22559
rect 13964 22528 14013 22556
rect 13964 22516 13970 22528
rect 14001 22525 14013 22528
rect 14047 22525 14059 22559
rect 14001 22519 14059 22525
rect 14550 22516 14556 22568
rect 14608 22556 14614 22568
rect 14645 22559 14703 22565
rect 14645 22556 14657 22559
rect 14608 22528 14657 22556
rect 14608 22516 14614 22528
rect 14645 22525 14657 22528
rect 14691 22525 14703 22559
rect 14826 22556 14832 22568
rect 14787 22528 14832 22556
rect 14645 22519 14703 22525
rect 14826 22516 14832 22528
rect 14884 22516 14890 22568
rect 15838 22556 15844 22568
rect 15799 22528 15844 22556
rect 15838 22516 15844 22528
rect 15896 22516 15902 22568
rect 16040 22565 16068 22596
rect 16666 22584 16672 22596
rect 16724 22624 16730 22636
rect 18690 22624 18696 22636
rect 16724 22596 18092 22624
rect 18651 22596 18696 22624
rect 16724 22584 16730 22596
rect 16025 22559 16083 22565
rect 16025 22525 16037 22559
rect 16071 22525 16083 22559
rect 16761 22559 16819 22565
rect 16761 22556 16773 22559
rect 16025 22519 16083 22525
rect 16408 22528 16773 22556
rect 14568 22488 14596 22516
rect 15378 22488 15384 22500
rect 11103 22460 13216 22488
rect 13464 22460 14596 22488
rect 15339 22460 15384 22488
rect 11103 22457 11115 22460
rect 11057 22451 11115 22457
rect 10318 22420 10324 22432
rect 9876 22392 10324 22420
rect 10318 22380 10324 22392
rect 10376 22380 10382 22432
rect 10410 22380 10416 22432
rect 10468 22420 10474 22432
rect 10781 22423 10839 22429
rect 10781 22420 10793 22423
rect 10468 22392 10793 22420
rect 10468 22380 10474 22392
rect 10781 22389 10793 22392
rect 10827 22389 10839 22423
rect 10781 22383 10839 22389
rect 12069 22423 12127 22429
rect 12069 22389 12081 22423
rect 12115 22420 12127 22423
rect 12342 22420 12348 22432
rect 12115 22392 12348 22420
rect 12115 22389 12127 22392
rect 12069 22383 12127 22389
rect 12342 22380 12348 22392
rect 12400 22420 12406 22432
rect 13078 22420 13084 22432
rect 12400 22392 13084 22420
rect 12400 22380 12406 22392
rect 13078 22380 13084 22392
rect 13136 22380 13142 22432
rect 13188 22420 13216 22460
rect 15378 22448 15384 22460
rect 15436 22448 15442 22500
rect 16408 22432 16436 22528
rect 16761 22525 16773 22528
rect 16807 22525 16819 22559
rect 16942 22556 16948 22568
rect 16903 22528 16948 22556
rect 16761 22519 16819 22525
rect 16942 22516 16948 22528
rect 17000 22516 17006 22568
rect 18064 22565 18092 22596
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 18966 22624 18972 22636
rect 18927 22596 18972 22624
rect 18966 22584 18972 22596
rect 19024 22584 19030 22636
rect 19428 22627 19486 22633
rect 19428 22593 19440 22627
rect 19474 22624 19486 22627
rect 19536 22624 19564 22664
rect 19610 22652 19616 22664
rect 19668 22692 19674 22704
rect 20901 22695 20959 22701
rect 19668 22664 20024 22692
rect 19668 22652 19674 22664
rect 19702 22624 19708 22636
rect 19474 22596 19564 22624
rect 19663 22596 19708 22624
rect 19474 22593 19486 22596
rect 19428 22587 19486 22593
rect 19702 22584 19708 22596
rect 19760 22584 19766 22636
rect 17957 22559 18015 22565
rect 17957 22525 17969 22559
rect 18003 22525 18015 22559
rect 17957 22519 18015 22525
rect 18049 22559 18107 22565
rect 18049 22525 18061 22559
rect 18095 22525 18107 22559
rect 18049 22519 18107 22525
rect 19061 22559 19119 22565
rect 19061 22525 19073 22559
rect 19107 22556 19119 22559
rect 19518 22556 19524 22568
rect 19107 22528 19524 22556
rect 19107 22525 19119 22528
rect 19061 22519 19119 22525
rect 17402 22488 17408 22500
rect 17363 22460 17408 22488
rect 17402 22448 17408 22460
rect 17460 22448 17466 22500
rect 17972 22488 18000 22519
rect 19518 22516 19524 22528
rect 19576 22516 19582 22568
rect 19996 22556 20024 22664
rect 20901 22661 20913 22695
rect 20947 22692 20959 22695
rect 23753 22695 23811 22701
rect 23753 22692 23765 22695
rect 20947 22664 23765 22692
rect 20947 22661 20959 22664
rect 20901 22655 20959 22661
rect 23753 22661 23765 22664
rect 23799 22661 23811 22695
rect 23753 22655 23811 22661
rect 20346 22624 20352 22636
rect 20307 22596 20352 22624
rect 20346 22584 20352 22596
rect 20404 22584 20410 22636
rect 20714 22584 20720 22636
rect 20772 22624 20778 22636
rect 20809 22627 20867 22633
rect 20809 22624 20821 22627
rect 20772 22596 20821 22624
rect 20772 22584 20778 22596
rect 20809 22593 20821 22596
rect 20855 22593 20867 22627
rect 20809 22587 20867 22593
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22624 22063 22627
rect 22278 22624 22284 22636
rect 22051 22596 22284 22624
rect 22051 22593 22063 22596
rect 22005 22587 22063 22593
rect 22278 22584 22284 22596
rect 22336 22584 22342 22636
rect 22646 22624 22652 22636
rect 22607 22596 22652 22624
rect 22646 22584 22652 22596
rect 22704 22584 22710 22636
rect 23198 22624 23204 22636
rect 23159 22596 23204 22624
rect 23198 22584 23204 22596
rect 23256 22584 23262 22636
rect 23568 22627 23626 22633
rect 23568 22593 23580 22627
rect 23614 22624 23626 22627
rect 23658 22624 23664 22636
rect 23614 22596 23664 22624
rect 23614 22593 23626 22596
rect 23568 22587 23626 22593
rect 23658 22584 23664 22596
rect 23716 22584 23722 22636
rect 23845 22627 23903 22633
rect 23845 22593 23857 22627
rect 23891 22624 23903 22627
rect 23934 22624 23940 22636
rect 23891 22596 23940 22624
rect 23891 22593 23903 22596
rect 23845 22587 23903 22593
rect 23934 22584 23940 22596
rect 23992 22584 23998 22636
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22624 24271 22627
rect 24670 22624 24676 22636
rect 24259 22596 24676 22624
rect 24259 22593 24271 22596
rect 24213 22587 24271 22593
rect 24670 22584 24676 22596
rect 24728 22584 24734 22636
rect 20898 22556 20904 22568
rect 19996 22528 20904 22556
rect 20898 22516 20904 22528
rect 20956 22516 20962 22568
rect 21082 22516 21088 22568
rect 21140 22556 21146 22568
rect 21913 22559 21971 22565
rect 21913 22556 21925 22559
rect 21140 22528 21925 22556
rect 21140 22516 21146 22528
rect 21913 22525 21925 22528
rect 21959 22556 21971 22559
rect 22833 22559 22891 22565
rect 22833 22556 22845 22559
rect 21959 22528 22845 22556
rect 21959 22525 21971 22528
rect 21913 22519 21971 22525
rect 22833 22525 22845 22528
rect 22879 22556 22891 22559
rect 23014 22556 23020 22568
rect 22879 22528 23020 22556
rect 22879 22525 22891 22528
rect 22833 22519 22891 22525
rect 23014 22516 23020 22528
rect 23072 22516 23078 22568
rect 23109 22559 23167 22565
rect 23109 22525 23121 22559
rect 23155 22525 23167 22559
rect 24394 22556 24400 22568
rect 24355 22528 24400 22556
rect 23109 22519 23167 22525
rect 18782 22488 18788 22500
rect 17972 22460 18788 22488
rect 18782 22448 18788 22460
rect 18840 22448 18846 22500
rect 18877 22491 18935 22497
rect 18877 22457 18889 22491
rect 18923 22488 18935 22491
rect 19334 22488 19340 22500
rect 18923 22460 19340 22488
rect 18923 22457 18935 22460
rect 18877 22451 18935 22457
rect 19334 22448 19340 22460
rect 19392 22488 19398 22500
rect 19702 22488 19708 22500
rect 19392 22460 19708 22488
rect 19392 22448 19398 22460
rect 19702 22448 19708 22460
rect 19760 22448 19766 22500
rect 20916 22488 20944 22516
rect 20916 22460 22692 22488
rect 13814 22420 13820 22432
rect 13188 22392 13820 22420
rect 13814 22380 13820 22392
rect 13872 22380 13878 22432
rect 16390 22420 16396 22432
rect 16351 22392 16396 22420
rect 16390 22380 16396 22392
rect 16448 22380 16454 22432
rect 16850 22380 16856 22432
rect 16908 22420 16914 22432
rect 17770 22420 17776 22432
rect 16908 22392 17776 22420
rect 16908 22380 16914 22392
rect 17770 22380 17776 22392
rect 17828 22380 17834 22432
rect 18506 22420 18512 22432
rect 18467 22392 18512 22420
rect 18506 22380 18512 22392
rect 18564 22380 18570 22432
rect 20073 22423 20131 22429
rect 20073 22389 20085 22423
rect 20119 22420 20131 22423
rect 20441 22423 20499 22429
rect 20441 22420 20453 22423
rect 20119 22392 20453 22420
rect 20119 22389 20131 22392
rect 20073 22383 20131 22389
rect 20441 22389 20453 22392
rect 20487 22389 20499 22423
rect 20441 22383 20499 22389
rect 22281 22423 22339 22429
rect 22281 22389 22293 22423
rect 22327 22420 22339 22423
rect 22370 22420 22376 22432
rect 22327 22392 22376 22420
rect 22327 22389 22339 22392
rect 22281 22383 22339 22389
rect 22370 22380 22376 22392
rect 22428 22380 22434 22432
rect 22664 22420 22692 22460
rect 23124 22420 23152 22519
rect 24394 22516 24400 22528
rect 24452 22516 24458 22568
rect 22664 22392 23152 22420
rect 23842 22380 23848 22432
rect 23900 22420 23906 22432
rect 23937 22423 23995 22429
rect 23937 22420 23949 22423
rect 23900 22392 23949 22420
rect 23900 22380 23906 22392
rect 23937 22389 23949 22392
rect 23983 22389 23995 22423
rect 23937 22383 23995 22389
rect 1104 22330 26128 22352
rect 1104 22278 5120 22330
rect 5172 22278 5184 22330
rect 5236 22278 5248 22330
rect 5300 22278 5312 22330
rect 5364 22278 5376 22330
rect 5428 22278 13462 22330
rect 13514 22278 13526 22330
rect 13578 22278 13590 22330
rect 13642 22278 13654 22330
rect 13706 22278 13718 22330
rect 13770 22278 21803 22330
rect 21855 22278 21867 22330
rect 21919 22278 21931 22330
rect 21983 22278 21995 22330
rect 22047 22278 22059 22330
rect 22111 22278 26128 22330
rect 1104 22256 26128 22278
rect 7650 22176 7656 22228
rect 7708 22216 7714 22228
rect 8021 22219 8079 22225
rect 8021 22216 8033 22219
rect 7708 22188 8033 22216
rect 7708 22176 7714 22188
rect 8021 22185 8033 22188
rect 8067 22185 8079 22219
rect 8021 22179 8079 22185
rect 8110 22176 8116 22228
rect 8168 22216 8174 22228
rect 9490 22216 9496 22228
rect 8168 22188 8984 22216
rect 9451 22188 9496 22216
rect 8168 22176 8174 22188
rect 5810 22108 5816 22160
rect 5868 22148 5874 22160
rect 5905 22151 5963 22157
rect 5905 22148 5917 22151
rect 5868 22120 5917 22148
rect 5868 22108 5874 22120
rect 5905 22117 5917 22120
rect 5951 22117 5963 22151
rect 5905 22111 5963 22117
rect 6270 22108 6276 22160
rect 6328 22148 6334 22160
rect 8956 22148 8984 22188
rect 9490 22176 9496 22188
rect 9548 22176 9554 22228
rect 10134 22176 10140 22228
rect 10192 22216 10198 22228
rect 10229 22219 10287 22225
rect 10229 22216 10241 22219
rect 10192 22188 10241 22216
rect 10192 22176 10198 22188
rect 10229 22185 10241 22188
rect 10275 22185 10287 22219
rect 10229 22179 10287 22185
rect 13354 22176 13360 22228
rect 13412 22216 13418 22228
rect 13449 22219 13507 22225
rect 13449 22216 13461 22219
rect 13412 22188 13461 22216
rect 13412 22176 13418 22188
rect 13449 22185 13461 22188
rect 13495 22185 13507 22219
rect 14090 22216 14096 22228
rect 14051 22188 14096 22216
rect 13449 22179 13507 22185
rect 14090 22176 14096 22188
rect 14148 22176 14154 22228
rect 15194 22216 15200 22228
rect 14200 22188 15200 22216
rect 9950 22148 9956 22160
rect 6328 22120 8892 22148
rect 8956 22120 9956 22148
rect 6328 22108 6334 22120
rect 5997 22083 6055 22089
rect 5997 22049 6009 22083
rect 6043 22080 6055 22083
rect 6914 22080 6920 22092
rect 6043 22052 6920 22080
rect 6043 22049 6055 22052
rect 5997 22043 6055 22049
rect 6914 22040 6920 22052
rect 6972 22040 6978 22092
rect 8864 22080 8892 22120
rect 9950 22108 9956 22120
rect 10008 22108 10014 22160
rect 13906 22108 13912 22160
rect 13964 22148 13970 22160
rect 14200 22148 14228 22188
rect 15194 22176 15200 22188
rect 15252 22176 15258 22228
rect 16206 22216 16212 22228
rect 16167 22188 16212 22216
rect 16206 22176 16212 22188
rect 16264 22176 16270 22228
rect 16942 22176 16948 22228
rect 17000 22216 17006 22228
rect 17221 22219 17279 22225
rect 17221 22216 17233 22219
rect 17000 22188 17233 22216
rect 17000 22176 17006 22188
rect 17221 22185 17233 22188
rect 17267 22185 17279 22219
rect 17221 22179 17279 22185
rect 20254 22176 20260 22228
rect 20312 22216 20318 22228
rect 20349 22219 20407 22225
rect 20349 22216 20361 22219
rect 20312 22188 20361 22216
rect 20312 22176 20318 22188
rect 20349 22185 20361 22188
rect 20395 22216 20407 22219
rect 21082 22216 21088 22228
rect 20395 22188 21088 22216
rect 20395 22185 20407 22188
rect 20349 22179 20407 22185
rect 21082 22176 21088 22188
rect 21140 22176 21146 22228
rect 22097 22219 22155 22225
rect 22097 22185 22109 22219
rect 22143 22216 22155 22219
rect 22370 22216 22376 22228
rect 22143 22188 22376 22216
rect 22143 22185 22155 22188
rect 22097 22179 22155 22185
rect 22370 22176 22376 22188
rect 22428 22176 22434 22228
rect 22833 22219 22891 22225
rect 22833 22185 22845 22219
rect 22879 22216 22891 22219
rect 23385 22219 23443 22225
rect 23385 22216 23397 22219
rect 22879 22188 23397 22216
rect 22879 22185 22891 22188
rect 22833 22179 22891 22185
rect 23385 22185 23397 22188
rect 23431 22185 23443 22219
rect 24854 22216 24860 22228
rect 24815 22188 24860 22216
rect 23385 22179 23443 22185
rect 24854 22176 24860 22188
rect 24912 22176 24918 22228
rect 13964 22120 14228 22148
rect 13964 22108 13970 22120
rect 16114 22108 16120 22160
rect 16172 22148 16178 22160
rect 16758 22148 16764 22160
rect 16172 22120 16764 22148
rect 16172 22108 16178 22120
rect 8941 22083 8999 22089
rect 8941 22080 8953 22083
rect 8864 22052 8953 22080
rect 8941 22049 8953 22052
rect 8987 22080 8999 22083
rect 10686 22080 10692 22092
rect 8987 22052 10692 22080
rect 8987 22049 8999 22052
rect 8941 22043 8999 22049
rect 1949 22015 2007 22021
rect 1949 21981 1961 22015
rect 1995 22012 2007 22015
rect 2774 22012 2780 22024
rect 1995 21984 2780 22012
rect 1995 21981 2007 21984
rect 1949 21975 2007 21981
rect 2774 21972 2780 21984
rect 2832 22012 2838 22024
rect 3786 22012 3792 22024
rect 2832 21984 3792 22012
rect 2832 21972 2838 21984
rect 3786 21972 3792 21984
rect 3844 21972 3850 22024
rect 4798 21972 4804 22024
rect 4856 22012 4862 22024
rect 5629 22015 5687 22021
rect 5629 22012 5641 22015
rect 4856 21984 5641 22012
rect 4856 21972 4862 21984
rect 5629 21981 5641 21984
rect 5675 21981 5687 22015
rect 5629 21975 5687 21981
rect 5721 22015 5779 22021
rect 5721 21981 5733 22015
rect 5767 22012 5779 22015
rect 6638 22012 6644 22024
rect 5767 21984 6644 22012
rect 5767 21981 5779 21984
rect 5721 21975 5779 21981
rect 2216 21947 2274 21953
rect 2216 21913 2228 21947
rect 2262 21944 2274 21947
rect 3234 21944 3240 21956
rect 2262 21916 3240 21944
rect 2262 21913 2274 21916
rect 2216 21907 2274 21913
rect 3234 21904 3240 21916
rect 3292 21904 3298 21956
rect 4056 21947 4114 21953
rect 4056 21913 4068 21947
rect 4102 21944 4114 21947
rect 4154 21944 4160 21956
rect 4102 21916 4160 21944
rect 4102 21913 4114 21916
rect 4056 21907 4114 21913
rect 4154 21904 4160 21916
rect 4212 21904 4218 21956
rect 3326 21876 3332 21888
rect 3287 21848 3332 21876
rect 3326 21836 3332 21848
rect 3384 21836 3390 21888
rect 4338 21836 4344 21888
rect 4396 21876 4402 21888
rect 5169 21879 5227 21885
rect 5169 21876 5181 21879
rect 4396 21848 5181 21876
rect 4396 21836 4402 21848
rect 5169 21845 5181 21848
rect 5215 21845 5227 21879
rect 5169 21839 5227 21845
rect 5350 21836 5356 21888
rect 5408 21876 5414 21888
rect 5445 21879 5503 21885
rect 5445 21876 5457 21879
rect 5408 21848 5457 21876
rect 5408 21836 5414 21848
rect 5445 21845 5457 21848
rect 5491 21845 5503 21879
rect 5644 21876 5672 21975
rect 6638 21972 6644 21984
rect 6696 21972 6702 22024
rect 8113 22015 8171 22021
rect 8113 21981 8125 22015
rect 8159 22012 8171 22015
rect 8294 22012 8300 22024
rect 8159 21984 8300 22012
rect 8159 21981 8171 21984
rect 8113 21975 8171 21981
rect 8294 21972 8300 21984
rect 8352 21972 8358 22024
rect 8570 21972 8576 22024
rect 8628 22012 8634 22024
rect 8757 22015 8815 22021
rect 8757 22012 8769 22015
rect 8628 21984 8769 22012
rect 8628 21972 8634 21984
rect 8757 21981 8769 21984
rect 8803 21981 8815 22015
rect 8956 22012 8984 22043
rect 10686 22040 10692 22052
rect 10744 22040 10750 22092
rect 10778 22040 10784 22092
rect 10836 22080 10842 22092
rect 13817 22083 13875 22089
rect 10836 22052 11376 22080
rect 10836 22040 10842 22052
rect 9125 22015 9183 22021
rect 9125 22012 9137 22015
rect 8956 21984 9137 22012
rect 8757 21975 8815 21981
rect 9125 21981 9137 21984
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 5994 21904 6000 21956
rect 6052 21944 6058 21956
rect 8478 21944 8484 21956
rect 6052 21916 8484 21944
rect 6052 21904 6058 21916
rect 8478 21904 8484 21916
rect 8536 21904 8542 21956
rect 8772 21944 8800 21975
rect 9674 21972 9680 22024
rect 9732 22012 9738 22024
rect 9858 22012 9864 22024
rect 9732 21984 9777 22012
rect 9819 21984 9864 22012
rect 9732 21972 9738 21984
rect 9858 21972 9864 21984
rect 9916 21972 9922 22024
rect 9953 22015 10011 22021
rect 9953 21981 9965 22015
rect 9999 21981 10011 22015
rect 10410 22012 10416 22024
rect 10371 21984 10416 22012
rect 9953 21975 10011 21981
rect 9968 21944 9996 21975
rect 10410 21972 10416 21984
rect 10468 21972 10474 22024
rect 11238 22012 11244 22024
rect 11199 21984 11244 22012
rect 11238 21972 11244 21984
rect 11296 21972 11302 22024
rect 11348 22012 11376 22052
rect 12406 22052 13492 22080
rect 12406 22012 12434 22052
rect 11348 21984 12434 22012
rect 13081 22015 13139 22021
rect 13081 21981 13093 22015
rect 13127 21981 13139 22015
rect 13354 22012 13360 22024
rect 13315 21984 13360 22012
rect 13081 21975 13139 21981
rect 8772 21916 9996 21944
rect 11508 21947 11566 21953
rect 11508 21913 11520 21947
rect 11554 21944 11566 21947
rect 11606 21944 11612 21956
rect 11554 21916 11612 21944
rect 11554 21913 11566 21916
rect 11508 21907 11566 21913
rect 11606 21904 11612 21916
rect 11664 21904 11670 21956
rect 12250 21904 12256 21956
rect 12308 21944 12314 21956
rect 12897 21947 12955 21953
rect 12897 21944 12909 21947
rect 12308 21916 12909 21944
rect 12308 21904 12314 21916
rect 12897 21913 12909 21916
rect 12943 21913 12955 21947
rect 12897 21907 12955 21913
rect 6362 21876 6368 21888
rect 5644 21848 6368 21876
rect 5445 21839 5503 21845
rect 6362 21836 6368 21848
rect 6420 21836 6426 21888
rect 7837 21879 7895 21885
rect 7837 21845 7849 21879
rect 7883 21876 7895 21879
rect 8202 21876 8208 21888
rect 7883 21848 8208 21876
rect 7883 21845 7895 21848
rect 7837 21839 7895 21845
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 8662 21876 8668 21888
rect 8623 21848 8668 21876
rect 8662 21836 8668 21848
rect 8720 21836 8726 21888
rect 9217 21879 9275 21885
rect 9217 21845 9229 21879
rect 9263 21876 9275 21879
rect 9858 21876 9864 21888
rect 9263 21848 9864 21876
rect 9263 21845 9275 21848
rect 9217 21839 9275 21845
rect 9858 21836 9864 21848
rect 9916 21836 9922 21888
rect 9950 21836 9956 21888
rect 10008 21876 10014 21888
rect 10137 21879 10195 21885
rect 10137 21876 10149 21879
rect 10008 21848 10149 21876
rect 10008 21836 10014 21848
rect 10137 21845 10149 21848
rect 10183 21876 10195 21879
rect 11330 21876 11336 21888
rect 10183 21848 11336 21876
rect 10183 21845 10195 21848
rect 10137 21839 10195 21845
rect 11330 21836 11336 21848
rect 11388 21836 11394 21888
rect 12066 21836 12072 21888
rect 12124 21876 12130 21888
rect 12621 21879 12679 21885
rect 12621 21876 12633 21879
rect 12124 21848 12633 21876
rect 12124 21836 12130 21848
rect 12621 21845 12633 21848
rect 12667 21876 12679 21879
rect 13096 21876 13124 21975
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 13265 21947 13323 21953
rect 13265 21913 13277 21947
rect 13311 21944 13323 21947
rect 13464 21944 13492 22052
rect 13817 22049 13829 22083
rect 13863 22080 13875 22083
rect 14550 22080 14556 22092
rect 13863 22052 14556 22080
rect 13863 22049 13875 22052
rect 13817 22043 13875 22049
rect 14550 22040 14556 22052
rect 14608 22080 14614 22092
rect 14737 22083 14795 22089
rect 14737 22080 14749 22083
rect 14608 22052 14749 22080
rect 14608 22040 14614 22052
rect 14737 22049 14749 22052
rect 14783 22080 14795 22083
rect 15657 22083 15715 22089
rect 15657 22080 15669 22083
rect 14783 22052 15669 22080
rect 14783 22049 14795 22052
rect 14737 22043 14795 22049
rect 15657 22049 15669 22052
rect 15703 22080 15715 22083
rect 16390 22080 16396 22092
rect 15703 22052 16396 22080
rect 15703 22049 15715 22052
rect 15657 22043 15715 22049
rect 16390 22040 16396 22052
rect 16448 22040 16454 22092
rect 15194 22012 15200 22024
rect 15155 21984 15200 22012
rect 15194 21972 15200 21984
rect 15252 21972 15258 22024
rect 15378 21972 15384 22024
rect 15436 22012 15442 22024
rect 16500 22021 16528 22120
rect 16758 22108 16764 22120
rect 16816 22108 16822 22160
rect 22278 22148 22284 22160
rect 22239 22120 22284 22148
rect 22278 22108 22284 22120
rect 22336 22108 22342 22160
rect 23014 22108 23020 22160
rect 23072 22148 23078 22160
rect 23201 22151 23259 22157
rect 23201 22148 23213 22151
rect 23072 22120 23213 22148
rect 23072 22108 23078 22120
rect 23201 22117 23213 22120
rect 23247 22148 23259 22151
rect 23247 22120 23980 22148
rect 23247 22117 23259 22120
rect 23201 22111 23259 22117
rect 23952 22094 23980 22120
rect 16850 22080 16856 22092
rect 16811 22052 16856 22080
rect 16850 22040 16856 22052
rect 16908 22040 16914 22092
rect 23842 22080 23848 22092
rect 23803 22052 23848 22080
rect 23842 22040 23848 22052
rect 23900 22040 23906 22092
rect 23952 22089 24017 22094
rect 23937 22083 24017 22089
rect 23937 22049 23949 22083
rect 23983 22066 24017 22083
rect 23983 22049 23995 22066
rect 23937 22043 23995 22049
rect 24136 22052 25268 22080
rect 16301 22015 16359 22021
rect 16301 22012 16313 22015
rect 15436 21984 16313 22012
rect 15436 21972 15442 21984
rect 16301 21981 16313 21984
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 16485 22015 16543 22021
rect 16485 21981 16497 22015
rect 16531 21981 16543 22015
rect 16485 21975 16543 21981
rect 16669 22015 16727 22021
rect 16669 21981 16681 22015
rect 16715 22012 16727 22015
rect 17405 22015 17463 22021
rect 17405 22012 17417 22015
rect 16715 21984 17417 22012
rect 16715 21981 16727 21984
rect 16669 21975 16727 21981
rect 17405 21981 17417 21984
rect 17451 21981 17463 22015
rect 17405 21975 17463 21981
rect 19702 21972 19708 22024
rect 19760 22012 19766 22024
rect 21729 22015 21787 22021
rect 21729 22012 21741 22015
rect 19760 21984 21741 22012
rect 19760 21972 19766 21984
rect 21729 21981 21741 21984
rect 21775 22012 21787 22015
rect 22465 22015 22523 22021
rect 22465 22012 22477 22015
rect 21775 21984 22477 22012
rect 21775 21981 21787 21984
rect 21729 21975 21787 21981
rect 22465 21981 22477 21984
rect 22511 21981 22523 22015
rect 22465 21975 22523 21981
rect 23109 22015 23167 22021
rect 23109 21981 23121 22015
rect 23155 22012 23167 22015
rect 24136 22012 24164 22052
rect 24670 22012 24676 22024
rect 23155 21984 24164 22012
rect 24631 21984 24676 22012
rect 23155 21981 23167 21984
rect 23109 21975 23167 21981
rect 24670 21972 24676 21984
rect 24728 21972 24734 22024
rect 25240 22021 25268 22052
rect 25225 22015 25283 22021
rect 25225 21981 25237 22015
rect 25271 21981 25283 22015
rect 25225 21975 25283 21981
rect 13311 21916 15240 21944
rect 13311 21913 13323 21916
rect 13265 21907 13323 21913
rect 15212 21888 15240 21916
rect 15470 21904 15476 21956
rect 15528 21944 15534 21956
rect 15838 21944 15844 21956
rect 15528 21916 15844 21944
rect 15528 21904 15534 21916
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 17034 21944 17040 21956
rect 16995 21916 17040 21944
rect 17034 21904 17040 21916
rect 17092 21944 17098 21956
rect 17497 21947 17555 21953
rect 17497 21944 17509 21947
rect 17092 21916 17509 21944
rect 17092 21904 17098 21916
rect 17497 21913 17509 21916
rect 17543 21913 17555 21947
rect 17497 21907 17555 21913
rect 22143 21947 22201 21953
rect 22143 21913 22155 21947
rect 22189 21944 22201 21947
rect 22842 21947 22900 21953
rect 22842 21944 22854 21947
rect 22189 21916 22854 21944
rect 22189 21913 22201 21916
rect 22143 21907 22201 21913
rect 22842 21913 22854 21916
rect 22888 21944 22900 21947
rect 22888 21916 23428 21944
rect 22888 21913 22900 21916
rect 22842 21907 22900 21913
rect 14458 21876 14464 21888
rect 12667 21848 13124 21876
rect 14419 21848 14464 21876
rect 12667 21845 12679 21848
rect 12621 21839 12679 21845
rect 14458 21836 14464 21848
rect 14516 21836 14522 21888
rect 14550 21836 14556 21888
rect 14608 21876 14614 21888
rect 15010 21876 15016 21888
rect 14608 21848 14653 21876
rect 14971 21848 15016 21876
rect 14608 21836 14614 21848
rect 15010 21836 15016 21848
rect 15068 21836 15074 21888
rect 15194 21836 15200 21888
rect 15252 21836 15258 21888
rect 15746 21876 15752 21888
rect 15707 21848 15752 21876
rect 15746 21836 15752 21848
rect 15804 21836 15810 21888
rect 23400 21876 23428 21916
rect 23474 21904 23480 21956
rect 23532 21944 23538 21956
rect 23532 21916 23888 21944
rect 23532 21904 23538 21916
rect 23860 21888 23888 21916
rect 24026 21904 24032 21956
rect 24084 21944 24090 21956
rect 24397 21947 24455 21953
rect 24397 21944 24409 21947
rect 24084 21916 24409 21944
rect 24084 21904 24090 21916
rect 24397 21913 24409 21916
rect 24443 21913 24455 21947
rect 24397 21907 24455 21913
rect 23566 21876 23572 21888
rect 23400 21848 23572 21876
rect 23566 21836 23572 21848
rect 23624 21836 23630 21888
rect 23750 21876 23756 21888
rect 23711 21848 23756 21876
rect 23750 21836 23756 21848
rect 23808 21836 23814 21888
rect 23842 21836 23848 21888
rect 23900 21876 23906 21888
rect 24489 21879 24547 21885
rect 24489 21876 24501 21879
rect 23900 21848 24501 21876
rect 23900 21836 23906 21848
rect 24489 21845 24501 21848
rect 24535 21845 24547 21879
rect 25038 21876 25044 21888
rect 24999 21848 25044 21876
rect 24489 21839 24547 21845
rect 25038 21836 25044 21848
rect 25096 21836 25102 21888
rect 1104 21786 26128 21808
rect 1104 21734 9291 21786
rect 9343 21734 9355 21786
rect 9407 21734 9419 21786
rect 9471 21734 9483 21786
rect 9535 21734 9547 21786
rect 9599 21734 17632 21786
rect 17684 21734 17696 21786
rect 17748 21734 17760 21786
rect 17812 21734 17824 21786
rect 17876 21734 17888 21786
rect 17940 21734 26128 21786
rect 1104 21712 26128 21734
rect 3234 21672 3240 21684
rect 3195 21644 3240 21672
rect 3234 21632 3240 21644
rect 3292 21632 3298 21684
rect 4249 21675 4307 21681
rect 4249 21641 4261 21675
rect 4295 21672 4307 21675
rect 4798 21672 4804 21684
rect 4295 21644 4804 21672
rect 4295 21641 4307 21644
rect 4249 21635 4307 21641
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 5810 21672 5816 21684
rect 5771 21644 5816 21672
rect 5810 21632 5816 21644
rect 5868 21632 5874 21684
rect 5902 21632 5908 21684
rect 5960 21672 5966 21684
rect 7469 21675 7527 21681
rect 5960 21644 6684 21672
rect 5960 21632 5966 21644
rect 3970 21564 3976 21616
rect 4028 21604 4034 21616
rect 4028 21576 6592 21604
rect 4028 21564 4034 21576
rect 3234 21496 3240 21548
rect 3292 21536 3298 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 3292 21508 3433 21536
rect 3292 21496 3298 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 3513 21539 3571 21545
rect 3513 21505 3525 21539
rect 3559 21536 3571 21539
rect 4430 21536 4436 21548
rect 3559 21508 4436 21536
rect 3559 21505 3571 21508
rect 3513 21499 3571 21505
rect 4430 21496 4436 21508
rect 4488 21496 4494 21548
rect 5350 21496 5356 21548
rect 5408 21545 5414 21548
rect 6012 21545 6040 21576
rect 5408 21536 5420 21545
rect 5997 21539 6055 21545
rect 5408 21508 5453 21536
rect 5408 21499 5420 21508
rect 5997 21505 6009 21539
rect 6043 21505 6055 21539
rect 6454 21536 6460 21548
rect 5997 21499 6055 21505
rect 6196 21508 6460 21536
rect 5408 21496 5414 21499
rect 3694 21468 3700 21480
rect 3655 21440 3700 21468
rect 3694 21428 3700 21440
rect 3752 21428 3758 21480
rect 3789 21471 3847 21477
rect 3789 21437 3801 21471
rect 3835 21468 3847 21471
rect 3878 21468 3884 21480
rect 3835 21440 3884 21468
rect 3835 21437 3847 21440
rect 3789 21431 3847 21437
rect 3878 21428 3884 21440
rect 3936 21428 3942 21480
rect 5629 21471 5687 21477
rect 5629 21437 5641 21471
rect 5675 21437 5687 21471
rect 5629 21431 5687 21437
rect 5644 21400 5672 21431
rect 5718 21428 5724 21480
rect 5776 21468 5782 21480
rect 6196 21477 6224 21508
rect 6454 21496 6460 21508
rect 6512 21496 6518 21548
rect 6564 21545 6592 21576
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 6181 21471 6239 21477
rect 6181 21468 6193 21471
rect 5776 21440 6193 21468
rect 5776 21428 5782 21440
rect 6181 21437 6193 21440
rect 6227 21437 6239 21471
rect 6362 21468 6368 21480
rect 6323 21440 6368 21468
rect 6181 21431 6239 21437
rect 6362 21428 6368 21440
rect 6420 21428 6426 21480
rect 6656 21468 6684 21644
rect 7469 21641 7481 21675
rect 7515 21672 7527 21675
rect 7558 21672 7564 21684
rect 7515 21644 7564 21672
rect 7515 21641 7527 21644
rect 7469 21635 7527 21641
rect 7558 21632 7564 21644
rect 7616 21632 7622 21684
rect 8389 21675 8447 21681
rect 8389 21641 8401 21675
rect 8435 21672 8447 21675
rect 10597 21675 10655 21681
rect 8435 21644 10548 21672
rect 8435 21641 8447 21644
rect 8389 21635 8447 21641
rect 10520 21604 10548 21644
rect 10597 21641 10609 21675
rect 10643 21672 10655 21675
rect 10778 21672 10784 21684
rect 10643 21644 10784 21672
rect 10643 21641 10655 21644
rect 10597 21635 10655 21641
rect 10778 21632 10784 21644
rect 10836 21632 10842 21684
rect 11146 21672 11152 21684
rect 11107 21644 11152 21672
rect 11146 21632 11152 21644
rect 11204 21632 11210 21684
rect 11606 21672 11612 21684
rect 11567 21644 11612 21672
rect 11606 21632 11612 21644
rect 11664 21632 11670 21684
rect 12158 21672 12164 21684
rect 11900 21644 12164 21672
rect 9048 21576 9674 21604
rect 10520 21576 11376 21604
rect 7006 21536 7012 21548
rect 6967 21508 7012 21536
rect 7006 21496 7012 21508
rect 7064 21496 7070 21548
rect 7650 21536 7656 21548
rect 7611 21508 7656 21536
rect 7650 21496 7656 21508
rect 7708 21496 7714 21548
rect 7742 21496 7748 21548
rect 7800 21536 7806 21548
rect 9048 21545 9076 21576
rect 9646 21548 9674 21576
rect 8205 21539 8263 21545
rect 8205 21536 8217 21539
rect 7800 21508 8217 21536
rect 7800 21496 7806 21508
rect 8205 21505 8217 21508
rect 8251 21505 8263 21539
rect 9033 21539 9091 21545
rect 9033 21536 9045 21539
rect 8205 21499 8263 21505
rect 8864 21508 9045 21536
rect 7668 21468 7696 21496
rect 6656 21440 7696 21468
rect 8018 21428 8024 21480
rect 8076 21468 8082 21480
rect 8662 21468 8668 21480
rect 8076 21440 8668 21468
rect 8076 21428 8082 21440
rect 8662 21428 8668 21440
rect 8720 21468 8726 21480
rect 8864 21468 8892 21508
rect 9033 21505 9045 21508
rect 9079 21505 9091 21539
rect 9401 21539 9459 21545
rect 9401 21536 9413 21539
rect 9033 21499 9091 21505
rect 9140 21508 9413 21536
rect 8720 21440 8892 21468
rect 8720 21428 8726 21440
rect 8938 21428 8944 21480
rect 8996 21468 9002 21480
rect 9140 21468 9168 21508
rect 9401 21505 9413 21508
rect 9447 21505 9459 21539
rect 9646 21508 9680 21548
rect 9401 21499 9459 21505
rect 9674 21496 9680 21508
rect 9732 21536 9738 21548
rect 9732 21508 9777 21536
rect 9732 21496 9738 21508
rect 9950 21496 9956 21548
rect 10008 21536 10014 21548
rect 10045 21539 10103 21545
rect 10045 21536 10057 21539
rect 10008 21508 10057 21536
rect 10008 21496 10014 21508
rect 10045 21505 10057 21508
rect 10091 21505 10103 21539
rect 10045 21499 10103 21505
rect 8996 21440 9168 21468
rect 9217 21471 9275 21477
rect 8996 21428 9002 21440
rect 9217 21437 9229 21471
rect 9263 21468 9275 21471
rect 9766 21468 9772 21480
rect 9263 21440 9772 21468
rect 9263 21437 9275 21440
rect 9217 21431 9275 21437
rect 9766 21428 9772 21440
rect 9824 21428 9830 21480
rect 9861 21471 9919 21477
rect 9861 21437 9873 21471
rect 9907 21437 9919 21471
rect 10060 21468 10088 21499
rect 10134 21496 10140 21548
rect 10192 21536 10198 21548
rect 11348 21545 11376 21576
rect 10413 21539 10471 21545
rect 10192 21508 10237 21536
rect 10192 21496 10198 21508
rect 10413 21505 10425 21539
rect 10459 21505 10471 21539
rect 10413 21499 10471 21505
rect 11333 21539 11391 21545
rect 11333 21505 11345 21539
rect 11379 21536 11391 21539
rect 11793 21539 11851 21545
rect 11793 21536 11805 21539
rect 11379 21508 11805 21536
rect 11379 21505 11391 21508
rect 11333 21499 11391 21505
rect 11793 21505 11805 21508
rect 11839 21536 11851 21539
rect 11900 21536 11928 21644
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 12621 21675 12679 21681
rect 12621 21641 12633 21675
rect 12667 21641 12679 21675
rect 12621 21635 12679 21641
rect 13817 21675 13875 21681
rect 13817 21641 13829 21675
rect 13863 21672 13875 21675
rect 14550 21672 14556 21684
rect 13863 21644 14556 21672
rect 13863 21641 13875 21644
rect 13817 21635 13875 21641
rect 12636 21604 12664 21635
rect 14550 21632 14556 21644
rect 14608 21632 14614 21684
rect 14737 21675 14795 21681
rect 14737 21641 14749 21675
rect 14783 21672 14795 21675
rect 14826 21672 14832 21684
rect 14783 21644 14832 21672
rect 14783 21641 14795 21644
rect 14737 21635 14795 21641
rect 14826 21632 14832 21644
rect 14884 21632 14890 21684
rect 15746 21632 15752 21684
rect 15804 21672 15810 21684
rect 15841 21675 15899 21681
rect 15841 21672 15853 21675
rect 15804 21644 15853 21672
rect 15804 21632 15810 21644
rect 15841 21641 15853 21644
rect 15887 21641 15899 21675
rect 15841 21635 15899 21641
rect 23201 21675 23259 21681
rect 23201 21641 23213 21675
rect 23247 21672 23259 21675
rect 24670 21672 24676 21684
rect 23247 21644 24676 21672
rect 23247 21641 23259 21644
rect 23201 21635 23259 21641
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 15378 21604 15384 21616
rect 11992 21576 15384 21604
rect 11992 21545 12020 21576
rect 11839 21508 11928 21536
rect 11977 21539 12035 21545
rect 11839 21505 11851 21508
rect 11793 21499 11851 21505
rect 11977 21505 11989 21539
rect 12023 21505 12035 21539
rect 11977 21499 12035 21505
rect 12069 21539 12127 21545
rect 12069 21505 12081 21539
rect 12115 21505 12127 21539
rect 12250 21536 12256 21548
rect 12211 21508 12256 21536
rect 12069 21499 12127 21505
rect 10428 21468 10456 21499
rect 10060 21440 10456 21468
rect 9861 21431 9919 21437
rect 6822 21400 6828 21412
rect 5644 21372 6828 21400
rect 6822 21360 6828 21372
rect 6880 21360 6886 21412
rect 7006 21360 7012 21412
rect 7064 21400 7070 21412
rect 7377 21403 7435 21409
rect 7377 21400 7389 21403
rect 7064 21372 7389 21400
rect 7064 21360 7070 21372
rect 7377 21369 7389 21372
rect 7423 21400 7435 21403
rect 7558 21400 7564 21412
rect 7423 21372 7564 21400
rect 7423 21369 7435 21372
rect 7377 21363 7435 21369
rect 7558 21360 7564 21372
rect 7616 21360 7622 21412
rect 8294 21360 8300 21412
rect 8352 21400 8358 21412
rect 9122 21400 9128 21412
rect 8352 21372 9128 21400
rect 8352 21360 8358 21372
rect 9122 21360 9128 21372
rect 9180 21400 9186 21412
rect 9677 21403 9735 21409
rect 9677 21400 9689 21403
rect 9180 21372 9689 21400
rect 9180 21360 9186 21372
rect 9677 21369 9689 21372
rect 9723 21369 9735 21403
rect 9876 21400 9904 21431
rect 10870 21428 10876 21480
rect 10928 21468 10934 21480
rect 11885 21471 11943 21477
rect 11885 21468 11897 21471
rect 10928 21440 11897 21468
rect 10928 21428 10934 21440
rect 11885 21437 11897 21440
rect 11931 21437 11943 21471
rect 11885 21431 11943 21437
rect 9876 21372 10364 21400
rect 9677 21363 9735 21369
rect 4614 21292 4620 21344
rect 4672 21332 4678 21344
rect 6733 21335 6791 21341
rect 6733 21332 6745 21335
rect 4672 21304 6745 21332
rect 4672 21292 4678 21304
rect 6733 21301 6745 21304
rect 6779 21301 6791 21335
rect 7098 21332 7104 21344
rect 7059 21304 7104 21332
rect 6733 21295 6791 21301
rect 7098 21292 7104 21304
rect 7156 21332 7162 21344
rect 7834 21332 7840 21344
rect 7156 21304 7840 21332
rect 7156 21292 7162 21304
rect 7834 21292 7840 21304
rect 7892 21292 7898 21344
rect 8662 21292 8668 21344
rect 8720 21332 8726 21344
rect 9309 21335 9367 21341
rect 9309 21332 9321 21335
rect 8720 21304 9321 21332
rect 8720 21292 8726 21304
rect 9309 21301 9321 21304
rect 9355 21332 9367 21335
rect 10134 21332 10140 21344
rect 9355 21304 10140 21332
rect 9355 21301 9367 21304
rect 9309 21295 9367 21301
rect 10134 21292 10140 21304
rect 10192 21292 10198 21344
rect 10336 21341 10364 21372
rect 11146 21360 11152 21412
rect 11204 21400 11210 21412
rect 12084 21400 12112 21499
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 12805 21539 12863 21545
rect 12805 21505 12817 21539
rect 12851 21536 12863 21539
rect 12894 21536 12900 21548
rect 12851 21508 12900 21536
rect 12851 21505 12863 21508
rect 12805 21499 12863 21505
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 13078 21536 13084 21548
rect 13039 21508 13084 21536
rect 13078 21496 13084 21508
rect 13136 21496 13142 21548
rect 13541 21539 13599 21545
rect 13541 21505 13553 21539
rect 13587 21505 13599 21539
rect 13814 21536 13820 21548
rect 13727 21508 13820 21536
rect 13541 21499 13599 21505
rect 13262 21428 13268 21480
rect 13320 21468 13326 21480
rect 13357 21471 13415 21477
rect 13357 21468 13369 21471
rect 13320 21440 13369 21468
rect 13320 21428 13326 21440
rect 13357 21437 13369 21440
rect 13403 21468 13415 21471
rect 13556 21468 13584 21499
rect 13814 21496 13820 21508
rect 13872 21536 13878 21548
rect 14553 21539 14611 21545
rect 13872 21508 14136 21536
rect 13872 21496 13878 21508
rect 13403 21440 13584 21468
rect 13403 21437 13415 21440
rect 13357 21431 13415 21437
rect 11204 21372 12112 21400
rect 11204 21360 11210 21372
rect 10321 21335 10379 21341
rect 10321 21301 10333 21335
rect 10367 21332 10379 21335
rect 10410 21332 10416 21344
rect 10367 21304 10416 21332
rect 10367 21301 10379 21304
rect 10321 21295 10379 21301
rect 10410 21292 10416 21304
rect 10468 21292 10474 21344
rect 13265 21335 13323 21341
rect 13265 21301 13277 21335
rect 13311 21332 13323 21335
rect 13814 21332 13820 21344
rect 13311 21304 13820 21332
rect 13311 21301 13323 21304
rect 13265 21295 13323 21301
rect 13814 21292 13820 21304
rect 13872 21292 13878 21344
rect 14108 21341 14136 21508
rect 14553 21505 14565 21539
rect 14599 21536 14611 21539
rect 15010 21536 15016 21548
rect 14599 21508 15016 21536
rect 14599 21505 14611 21508
rect 14553 21499 14611 21505
rect 15010 21496 15016 21508
rect 15068 21496 15074 21548
rect 15212 21545 15240 21576
rect 15378 21564 15384 21576
rect 15436 21564 15442 21616
rect 20898 21564 20904 21616
rect 20956 21604 20962 21616
rect 21726 21604 21732 21616
rect 20956 21576 21732 21604
rect 20956 21564 20962 21576
rect 21726 21564 21732 21576
rect 21784 21604 21790 21616
rect 21821 21607 21879 21613
rect 21821 21604 21833 21607
rect 21784 21576 21833 21604
rect 21784 21564 21790 21576
rect 21821 21573 21833 21576
rect 21867 21573 21879 21607
rect 21821 21567 21879 21573
rect 22005 21607 22063 21613
rect 22005 21573 22017 21607
rect 22051 21604 22063 21607
rect 22186 21604 22192 21616
rect 22051 21576 22192 21604
rect 22051 21573 22063 21576
rect 22005 21567 22063 21573
rect 22186 21564 22192 21576
rect 22244 21604 22250 21616
rect 22462 21604 22468 21616
rect 22244 21576 22468 21604
rect 22244 21564 22250 21576
rect 22462 21564 22468 21576
rect 22520 21564 22526 21616
rect 23474 21604 23480 21616
rect 23216 21576 23480 21604
rect 15197 21539 15255 21545
rect 15197 21505 15209 21539
rect 15243 21505 15255 21539
rect 15197 21499 15255 21505
rect 15289 21539 15347 21545
rect 15289 21505 15301 21539
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21536 15531 21539
rect 15657 21539 15715 21545
rect 15657 21536 15669 21539
rect 15519 21508 15669 21536
rect 15519 21505 15531 21508
rect 15473 21499 15531 21505
rect 15657 21505 15669 21508
rect 15703 21505 15715 21539
rect 15657 21499 15715 21505
rect 15304 21468 15332 21499
rect 17678 21496 17684 21548
rect 17736 21536 17742 21548
rect 18325 21539 18383 21545
rect 18325 21536 18337 21539
rect 17736 21508 18337 21536
rect 17736 21496 17742 21508
rect 18325 21505 18337 21508
rect 18371 21505 18383 21539
rect 18325 21499 18383 21505
rect 18509 21539 18567 21545
rect 18509 21505 18521 21539
rect 18555 21536 18567 21539
rect 19150 21536 19156 21548
rect 18555 21508 19156 21536
rect 18555 21505 18567 21508
rect 18509 21499 18567 21505
rect 18340 21468 18368 21499
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 23216 21545 23244 21576
rect 23474 21564 23480 21576
rect 23532 21564 23538 21616
rect 23652 21607 23710 21613
rect 23652 21573 23664 21607
rect 23698 21604 23710 21607
rect 25038 21604 25044 21616
rect 23698 21576 25044 21604
rect 23698 21573 23710 21576
rect 23652 21567 23710 21573
rect 25038 21564 25044 21576
rect 25096 21564 25102 21616
rect 23109 21539 23167 21545
rect 23109 21505 23121 21539
rect 23155 21505 23167 21539
rect 23109 21499 23167 21505
rect 23201 21539 23259 21545
rect 23201 21505 23213 21539
rect 23247 21505 23259 21539
rect 23382 21536 23388 21548
rect 23343 21508 23388 21536
rect 23201 21499 23259 21505
rect 18874 21468 18880 21480
rect 15304 21440 15516 21468
rect 18340 21440 18880 21468
rect 15488 21412 15516 21440
rect 18874 21428 18880 21440
rect 18932 21428 18938 21480
rect 22189 21471 22247 21477
rect 22189 21437 22201 21471
rect 22235 21468 22247 21471
rect 23124 21468 23152 21499
rect 23382 21496 23388 21508
rect 23440 21496 23446 21548
rect 22235 21440 23244 21468
rect 22235 21437 22247 21440
rect 22189 21431 22247 21437
rect 15470 21360 15476 21412
rect 15528 21360 15534 21412
rect 16025 21403 16083 21409
rect 16025 21369 16037 21403
rect 16071 21400 16083 21403
rect 16390 21400 16396 21412
rect 16071 21372 16396 21400
rect 16071 21369 16083 21372
rect 16025 21363 16083 21369
rect 16390 21360 16396 21372
rect 16448 21400 16454 21412
rect 17126 21400 17132 21412
rect 16448 21372 17132 21400
rect 16448 21360 16454 21372
rect 17126 21360 17132 21372
rect 17184 21360 17190 21412
rect 18414 21400 18420 21412
rect 17236 21372 18420 21400
rect 14093 21335 14151 21341
rect 14093 21301 14105 21335
rect 14139 21332 14151 21335
rect 17236 21332 17264 21372
rect 18414 21360 18420 21372
rect 18472 21360 18478 21412
rect 14139 21304 17264 21332
rect 18233 21335 18291 21341
rect 14139 21301 14151 21304
rect 14093 21295 14151 21301
rect 18233 21301 18245 21335
rect 18279 21332 18291 21335
rect 18322 21332 18328 21344
rect 18279 21304 18328 21332
rect 18279 21301 18291 21304
rect 18233 21295 18291 21301
rect 18322 21292 18328 21304
rect 18380 21292 18386 21344
rect 23216 21332 23244 21440
rect 23658 21332 23664 21344
rect 23216 21304 23664 21332
rect 23658 21292 23664 21304
rect 23716 21332 23722 21344
rect 24026 21332 24032 21344
rect 23716 21304 24032 21332
rect 23716 21292 23722 21304
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 24578 21292 24584 21344
rect 24636 21332 24642 21344
rect 24765 21335 24823 21341
rect 24765 21332 24777 21335
rect 24636 21304 24777 21332
rect 24636 21292 24642 21304
rect 24765 21301 24777 21304
rect 24811 21301 24823 21335
rect 24765 21295 24823 21301
rect 1104 21242 26128 21264
rect 1104 21190 5120 21242
rect 5172 21190 5184 21242
rect 5236 21190 5248 21242
rect 5300 21190 5312 21242
rect 5364 21190 5376 21242
rect 5428 21190 13462 21242
rect 13514 21190 13526 21242
rect 13578 21190 13590 21242
rect 13642 21190 13654 21242
rect 13706 21190 13718 21242
rect 13770 21190 21803 21242
rect 21855 21190 21867 21242
rect 21919 21190 21931 21242
rect 21983 21190 21995 21242
rect 22047 21190 22059 21242
rect 22111 21190 26128 21242
rect 1104 21168 26128 21190
rect 3970 21128 3976 21140
rect 3931 21100 3976 21128
rect 3970 21088 3976 21100
rect 4028 21088 4034 21140
rect 4154 21128 4160 21140
rect 4115 21100 4160 21128
rect 4154 21088 4160 21100
rect 4212 21088 4218 21140
rect 4614 21128 4620 21140
rect 4575 21100 4620 21128
rect 4614 21088 4620 21100
rect 4672 21088 4678 21140
rect 6638 21128 6644 21140
rect 4724 21100 6644 21128
rect 3988 20992 4016 21088
rect 4430 21020 4436 21072
rect 4488 21060 4494 21072
rect 4724 21060 4752 21100
rect 6638 21088 6644 21100
rect 6696 21088 6702 21140
rect 7742 21088 7748 21140
rect 7800 21128 7806 21140
rect 8389 21131 8447 21137
rect 8389 21128 8401 21131
rect 7800 21100 8401 21128
rect 7800 21088 7806 21100
rect 8389 21097 8401 21100
rect 8435 21097 8447 21131
rect 8389 21091 8447 21097
rect 6822 21060 6828 21072
rect 4488 21032 4752 21060
rect 6380 21032 6828 21060
rect 4488 21020 4494 21032
rect 3344 20964 4016 20992
rect 4080 20964 4660 20992
rect 3234 20924 3240 20936
rect 3195 20896 3240 20924
rect 3234 20884 3240 20896
rect 3292 20884 3298 20936
rect 3344 20933 3372 20964
rect 4080 20936 4108 20964
rect 3329 20927 3387 20933
rect 3329 20893 3341 20927
rect 3375 20893 3387 20927
rect 3329 20887 3387 20893
rect 3789 20927 3847 20933
rect 3789 20893 3801 20927
rect 3835 20924 3847 20927
rect 4062 20924 4068 20936
rect 3835 20896 4068 20924
rect 3835 20893 3847 20896
rect 3789 20887 3847 20893
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 4338 20924 4344 20936
rect 4251 20896 4344 20924
rect 4338 20884 4344 20896
rect 4396 20884 4402 20936
rect 4430 20884 4436 20936
rect 4488 20924 4494 20936
rect 4632 20924 4660 20964
rect 4706 20952 4712 21004
rect 4764 20992 4770 21004
rect 4764 20964 4809 20992
rect 4764 20952 4770 20964
rect 6380 20936 6408 21032
rect 6822 21020 6828 21032
rect 6880 21020 6886 21072
rect 7650 21020 7656 21072
rect 7708 21060 7714 21072
rect 7837 21063 7895 21069
rect 7837 21060 7849 21063
rect 7708 21032 7849 21060
rect 7708 21020 7714 21032
rect 7837 21029 7849 21032
rect 7883 21029 7895 21063
rect 8404 21060 8432 21091
rect 8938 21088 8944 21140
rect 8996 21128 9002 21140
rect 9217 21131 9275 21137
rect 9217 21128 9229 21131
rect 8996 21100 9229 21128
rect 8996 21088 9002 21100
rect 9217 21097 9229 21100
rect 9263 21128 9275 21131
rect 9861 21131 9919 21137
rect 9861 21128 9873 21131
rect 9263 21100 9873 21128
rect 9263 21097 9275 21100
rect 9217 21091 9275 21097
rect 9861 21097 9873 21100
rect 9907 21097 9919 21131
rect 9861 21091 9919 21097
rect 10321 21131 10379 21137
rect 10321 21097 10333 21131
rect 10367 21128 10379 21131
rect 11882 21128 11888 21140
rect 10367 21100 11888 21128
rect 10367 21097 10379 21100
rect 10321 21091 10379 21097
rect 11882 21088 11888 21100
rect 11940 21088 11946 21140
rect 17678 21128 17684 21140
rect 17639 21100 17684 21128
rect 17678 21088 17684 21100
rect 17736 21088 17742 21140
rect 22465 21131 22523 21137
rect 22465 21097 22477 21131
rect 22511 21128 22523 21131
rect 22649 21131 22707 21137
rect 22649 21128 22661 21131
rect 22511 21100 22661 21128
rect 22511 21097 22523 21100
rect 22465 21091 22523 21097
rect 22649 21097 22661 21100
rect 22695 21097 22707 21131
rect 22649 21091 22707 21097
rect 23109 21131 23167 21137
rect 23109 21097 23121 21131
rect 23155 21128 23167 21131
rect 23290 21128 23296 21140
rect 23155 21100 23296 21128
rect 23155 21097 23167 21100
rect 23109 21091 23167 21097
rect 23290 21088 23296 21100
rect 23348 21088 23354 21140
rect 23753 21131 23811 21137
rect 23753 21097 23765 21131
rect 23799 21128 23811 21131
rect 23842 21128 23848 21140
rect 23799 21100 23848 21128
rect 23799 21097 23811 21100
rect 23753 21091 23811 21097
rect 23842 21088 23848 21100
rect 23900 21088 23906 21140
rect 23934 21088 23940 21140
rect 23992 21128 23998 21140
rect 23992 21100 24037 21128
rect 23992 21088 23998 21100
rect 24394 21088 24400 21140
rect 24452 21128 24458 21140
rect 24489 21131 24547 21137
rect 24489 21128 24501 21131
rect 24452 21100 24501 21128
rect 24452 21088 24458 21100
rect 24489 21097 24501 21100
rect 24535 21097 24547 21131
rect 24489 21091 24547 21097
rect 9766 21060 9772 21072
rect 8404 21032 8708 21060
rect 7837 21023 7895 21029
rect 6638 20952 6644 21004
rect 6696 20992 6702 21004
rect 7009 20995 7067 21001
rect 6696 20964 6868 20992
rect 6696 20952 6702 20964
rect 5810 20924 5816 20936
rect 4488 20896 4533 20924
rect 4632 20896 5816 20924
rect 4488 20884 4494 20896
rect 5810 20884 5816 20896
rect 5868 20884 5874 20936
rect 6362 20924 6368 20936
rect 6323 20896 6368 20924
rect 6362 20884 6368 20896
rect 6420 20884 6426 20936
rect 6454 20884 6460 20936
rect 6512 20924 6518 20936
rect 6840 20933 6868 20964
rect 7009 20961 7021 20995
rect 7055 20992 7067 20995
rect 7285 20995 7343 21001
rect 7285 20992 7297 20995
rect 7055 20964 7297 20992
rect 7055 20961 7067 20964
rect 7009 20955 7067 20961
rect 7285 20961 7297 20964
rect 7331 20961 7343 20995
rect 7285 20955 7343 20961
rect 8202 20952 8208 21004
rect 8260 20992 8266 21004
rect 8570 20992 8576 21004
rect 8260 20964 8576 20992
rect 8260 20952 8266 20964
rect 8570 20952 8576 20964
rect 8628 20952 8634 21004
rect 6733 20927 6791 20933
rect 6733 20924 6745 20927
rect 6512 20896 6745 20924
rect 6512 20884 6518 20896
rect 6733 20893 6745 20896
rect 6779 20893 6791 20927
rect 6733 20887 6791 20893
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20893 6883 20927
rect 6825 20887 6883 20893
rect 6914 20884 6920 20936
rect 6972 20924 6978 20936
rect 7101 20927 7159 20933
rect 7101 20924 7113 20927
rect 6972 20896 7113 20924
rect 6972 20884 6978 20896
rect 7101 20893 7113 20896
rect 7147 20893 7159 20927
rect 7466 20924 7472 20936
rect 7427 20896 7472 20924
rect 7101 20887 7159 20893
rect 7466 20884 7472 20896
rect 7524 20884 7530 20936
rect 7650 20924 7656 20936
rect 7611 20896 7656 20924
rect 7650 20884 7656 20896
rect 7708 20884 7714 20936
rect 8018 20924 8024 20936
rect 7979 20896 8024 20924
rect 8018 20884 8024 20896
rect 8076 20884 8082 20936
rect 8386 20924 8392 20936
rect 8347 20896 8392 20924
rect 8386 20884 8392 20896
rect 8444 20884 8450 20936
rect 8680 20924 8708 21032
rect 9324 21032 9772 21060
rect 9324 21001 9352 21032
rect 9766 21020 9772 21032
rect 9824 21020 9830 21072
rect 10410 21020 10416 21072
rect 10468 21060 10474 21072
rect 11146 21060 11152 21072
rect 10468 21032 11152 21060
rect 10468 21020 10474 21032
rect 11146 21020 11152 21032
rect 11204 21020 11210 21072
rect 14458 21020 14464 21072
rect 14516 21060 14522 21072
rect 14918 21060 14924 21072
rect 14516 21032 14924 21060
rect 14516 21020 14522 21032
rect 14918 21020 14924 21032
rect 14976 21020 14982 21072
rect 23952 21060 23980 21088
rect 25038 21060 25044 21072
rect 23952 21032 25044 21060
rect 25038 21020 25044 21032
rect 25096 21020 25102 21072
rect 9309 20995 9367 21001
rect 9309 20961 9321 20995
rect 9355 20961 9367 20995
rect 9858 20992 9864 21004
rect 9309 20955 9367 20961
rect 9692 20964 9864 20992
rect 9692 20933 9720 20964
rect 9858 20952 9864 20964
rect 9916 20992 9922 21004
rect 15105 20995 15163 21001
rect 15105 20992 15117 20995
rect 9916 20964 15117 20992
rect 9916 20952 9922 20964
rect 15105 20961 15117 20964
rect 15151 20961 15163 20995
rect 15105 20955 15163 20961
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 18046 20992 18052 21004
rect 17451 20964 18052 20992
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 18046 20952 18052 20964
rect 18104 20952 18110 21004
rect 19797 20995 19855 21001
rect 19797 20992 19809 20995
rect 19076 20964 19809 20992
rect 9401 20927 9459 20933
rect 9401 20924 9413 20927
rect 8680 20896 9413 20924
rect 9401 20893 9413 20896
rect 9447 20893 9459 20927
rect 9401 20887 9459 20893
rect 9677 20927 9735 20933
rect 9677 20893 9689 20927
rect 9723 20893 9735 20927
rect 9950 20924 9956 20936
rect 9911 20896 9956 20924
rect 9677 20887 9735 20893
rect 4356 20856 4384 20884
rect 4614 20856 4620 20868
rect 4356 20828 4620 20856
rect 4614 20816 4620 20828
rect 4672 20816 4678 20868
rect 5626 20856 5632 20868
rect 5000 20828 5632 20856
rect 3513 20791 3571 20797
rect 3513 20757 3525 20791
rect 3559 20788 3571 20791
rect 3786 20788 3792 20800
rect 3559 20760 3792 20788
rect 3559 20757 3571 20760
rect 3513 20751 3571 20757
rect 3786 20748 3792 20760
rect 3844 20748 3850 20800
rect 5000 20797 5028 20828
rect 5626 20816 5632 20828
rect 5684 20816 5690 20868
rect 6120 20859 6178 20865
rect 6120 20825 6132 20859
rect 6166 20856 6178 20859
rect 6549 20859 6607 20865
rect 6549 20856 6561 20859
rect 6166 20828 6561 20856
rect 6166 20825 6178 20828
rect 6120 20819 6178 20825
rect 6549 20825 6561 20828
rect 6595 20825 6607 20859
rect 8662 20856 8668 20868
rect 6549 20819 6607 20825
rect 6656 20828 8248 20856
rect 8623 20828 8668 20856
rect 4985 20791 5043 20797
rect 4985 20757 4997 20791
rect 5031 20757 5043 20791
rect 4985 20751 5043 20757
rect 5534 20748 5540 20800
rect 5592 20788 5598 20800
rect 6656 20788 6684 20828
rect 8220 20797 8248 20828
rect 8662 20816 8668 20828
rect 8720 20816 8726 20868
rect 5592 20760 6684 20788
rect 8205 20791 8263 20797
rect 5592 20748 5598 20760
rect 8205 20757 8217 20791
rect 8251 20757 8263 20791
rect 8205 20751 8263 20757
rect 8294 20748 8300 20800
rect 8352 20788 8358 20800
rect 9033 20791 9091 20797
rect 9033 20788 9045 20791
rect 8352 20760 9045 20788
rect 8352 20748 8358 20760
rect 9033 20757 9045 20760
rect 9079 20757 9091 20791
rect 9416 20788 9444 20887
rect 9950 20884 9956 20896
rect 10008 20884 10014 20936
rect 10134 20924 10140 20936
rect 10095 20896 10140 20924
rect 10134 20884 10140 20896
rect 10192 20884 10198 20936
rect 10870 20884 10876 20936
rect 10928 20924 10934 20936
rect 11333 20927 11391 20933
rect 11333 20924 11345 20927
rect 10928 20896 11345 20924
rect 10928 20884 10934 20896
rect 11333 20893 11345 20896
rect 11379 20893 11391 20927
rect 14826 20924 14832 20936
rect 14787 20896 14832 20924
rect 11333 20887 11391 20893
rect 14826 20884 14832 20896
rect 14884 20884 14890 20936
rect 15473 20927 15531 20933
rect 15473 20893 15485 20927
rect 15519 20924 15531 20927
rect 16482 20924 16488 20936
rect 15519 20896 16488 20924
rect 15519 20893 15531 20896
rect 15473 20887 15531 20893
rect 16482 20884 16488 20896
rect 16540 20924 16546 20936
rect 17038 20927 17096 20933
rect 17038 20924 17050 20927
rect 16540 20896 17050 20924
rect 16540 20884 16546 20896
rect 17038 20893 17050 20896
rect 17084 20893 17096 20927
rect 17038 20887 17096 20893
rect 17497 20927 17555 20933
rect 17497 20893 17509 20927
rect 17543 20924 17555 20927
rect 18322 20924 18328 20936
rect 17543 20896 18328 20924
rect 17543 20893 17555 20896
rect 17497 20887 17555 20893
rect 18322 20884 18328 20896
rect 18380 20884 18386 20936
rect 18506 20884 18512 20936
rect 18564 20924 18570 20936
rect 19076 20933 19104 20964
rect 19797 20961 19809 20964
rect 19843 20961 19855 20995
rect 19797 20955 19855 20961
rect 21726 20952 21732 21004
rect 21784 20992 21790 21004
rect 23017 20995 23075 21001
rect 21784 20964 22508 20992
rect 21784 20952 21790 20964
rect 19061 20927 19119 20933
rect 19061 20924 19073 20927
rect 18564 20896 19073 20924
rect 18564 20884 18570 20896
rect 19061 20893 19073 20896
rect 19107 20893 19119 20927
rect 19061 20887 19119 20893
rect 19337 20927 19395 20933
rect 19337 20893 19349 20927
rect 19383 20893 19395 20927
rect 22370 20924 22376 20936
rect 22331 20896 22376 20924
rect 19337 20887 19395 20893
rect 10597 20859 10655 20865
rect 10597 20825 10609 20859
rect 10643 20825 10655 20859
rect 11054 20856 11060 20868
rect 11015 20828 11060 20856
rect 10597 20819 10655 20825
rect 9493 20791 9551 20797
rect 9493 20788 9505 20791
rect 9416 20760 9505 20788
rect 9033 20751 9091 20757
rect 9493 20757 9505 20760
rect 9539 20757 9551 20791
rect 9493 20751 9551 20757
rect 9861 20791 9919 20797
rect 9861 20757 9873 20791
rect 9907 20788 9919 20791
rect 10612 20788 10640 20819
rect 11054 20816 11060 20828
rect 11112 20816 11118 20868
rect 15286 20856 15292 20868
rect 15247 20828 15292 20856
rect 15286 20816 15292 20828
rect 15344 20816 15350 20868
rect 18816 20859 18874 20865
rect 18816 20825 18828 20859
rect 18862 20856 18874 20859
rect 18966 20856 18972 20868
rect 18862 20828 18972 20856
rect 18862 20825 18874 20828
rect 18816 20819 18874 20825
rect 18966 20816 18972 20828
rect 19024 20816 19030 20868
rect 9907 20760 10640 20788
rect 9907 20757 9919 20760
rect 9861 20751 9919 20757
rect 10778 20748 10784 20800
rect 10836 20788 10842 20800
rect 10873 20791 10931 20797
rect 10873 20788 10885 20791
rect 10836 20760 10885 20788
rect 10836 20748 10842 20760
rect 10873 20757 10885 20760
rect 10919 20757 10931 20791
rect 10873 20751 10931 20757
rect 10965 20791 11023 20797
rect 10965 20757 10977 20791
rect 11011 20788 11023 20791
rect 11330 20788 11336 20800
rect 11011 20760 11336 20788
rect 11011 20757 11023 20760
rect 10965 20751 11023 20757
rect 11330 20748 11336 20760
rect 11388 20748 11394 20800
rect 14458 20748 14464 20800
rect 14516 20788 14522 20800
rect 14645 20791 14703 20797
rect 14645 20788 14657 20791
rect 14516 20760 14657 20788
rect 14516 20748 14522 20760
rect 14645 20757 14657 20760
rect 14691 20757 14703 20791
rect 16942 20788 16948 20800
rect 16903 20760 16948 20788
rect 14645 20751 14703 20757
rect 16942 20748 16948 20760
rect 17000 20748 17006 20800
rect 18690 20748 18696 20800
rect 18748 20788 18754 20800
rect 19352 20788 19380 20887
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 22480 20933 22508 20964
rect 23017 20961 23029 20995
rect 23063 20992 23075 20995
rect 23063 20964 23796 20992
rect 23063 20961 23075 20964
rect 23017 20955 23075 20961
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20893 22523 20927
rect 22830 20924 22836 20936
rect 22791 20896 22836 20924
rect 22465 20887 22523 20893
rect 22830 20884 22836 20896
rect 22888 20884 22894 20936
rect 23569 20927 23627 20933
rect 23569 20893 23581 20927
rect 23615 20924 23627 20927
rect 23658 20924 23664 20936
rect 23615 20896 23664 20924
rect 23615 20893 23627 20896
rect 23569 20887 23627 20893
rect 23658 20884 23664 20896
rect 23716 20884 23722 20936
rect 23768 20933 23796 20964
rect 23753 20927 23811 20933
rect 23753 20893 23765 20927
rect 23799 20924 23811 20927
rect 24578 20924 24584 20936
rect 23799 20896 24584 20924
rect 23799 20893 23811 20896
rect 23753 20887 23811 20893
rect 24578 20884 24584 20896
rect 24636 20884 24642 20936
rect 20064 20859 20122 20865
rect 20064 20825 20076 20859
rect 20110 20856 20122 20859
rect 20162 20856 20168 20868
rect 20110 20828 20168 20856
rect 20110 20825 20122 20828
rect 20064 20819 20122 20825
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 23109 20859 23167 20865
rect 23109 20825 23121 20859
rect 23155 20856 23167 20859
rect 23842 20856 23848 20868
rect 23155 20828 23848 20856
rect 23155 20825 23167 20828
rect 23109 20819 23167 20825
rect 23842 20816 23848 20828
rect 23900 20816 23906 20868
rect 19518 20788 19524 20800
rect 18748 20760 19380 20788
rect 19479 20760 19524 20788
rect 18748 20748 18754 20760
rect 19518 20748 19524 20760
rect 19576 20748 19582 20800
rect 19705 20791 19763 20797
rect 19705 20757 19717 20791
rect 19751 20788 19763 20791
rect 20254 20788 20260 20800
rect 19751 20760 20260 20788
rect 19751 20757 19763 20760
rect 19705 20751 19763 20757
rect 20254 20748 20260 20760
rect 20312 20788 20318 20800
rect 20530 20788 20536 20800
rect 20312 20760 20536 20788
rect 20312 20748 20318 20760
rect 20530 20748 20536 20760
rect 20588 20748 20594 20800
rect 21177 20791 21235 20797
rect 21177 20757 21189 20791
rect 21223 20788 21235 20791
rect 21450 20788 21456 20800
rect 21223 20760 21456 20788
rect 21223 20757 21235 20760
rect 21177 20751 21235 20757
rect 21450 20748 21456 20760
rect 21508 20748 21514 20800
rect 21542 20748 21548 20800
rect 21600 20788 21606 20800
rect 22097 20791 22155 20797
rect 22097 20788 22109 20791
rect 21600 20760 22109 20788
rect 21600 20748 21606 20760
rect 22097 20757 22109 20760
rect 22143 20757 22155 20791
rect 22097 20751 22155 20757
rect 1104 20698 26128 20720
rect 1104 20646 9291 20698
rect 9343 20646 9355 20698
rect 9407 20646 9419 20698
rect 9471 20646 9483 20698
rect 9535 20646 9547 20698
rect 9599 20646 17632 20698
rect 17684 20646 17696 20698
rect 17748 20646 17760 20698
rect 17812 20646 17824 20698
rect 17876 20646 17888 20698
rect 17940 20646 26128 20698
rect 1104 20624 26128 20646
rect 4430 20584 4436 20596
rect 4391 20556 4436 20584
rect 4430 20544 4436 20556
rect 4488 20544 4494 20596
rect 4706 20544 4712 20596
rect 4764 20584 4770 20596
rect 5261 20587 5319 20593
rect 5261 20584 5273 20587
rect 4764 20556 5273 20584
rect 4764 20544 4770 20556
rect 5261 20553 5273 20556
rect 5307 20584 5319 20587
rect 7006 20584 7012 20596
rect 5307 20556 5672 20584
rect 5307 20553 5319 20556
rect 5261 20547 5319 20553
rect 2774 20516 2780 20528
rect 1688 20488 2780 20516
rect 1486 20408 1492 20460
rect 1544 20448 1550 20460
rect 1688 20457 1716 20488
rect 2774 20476 2780 20488
rect 2832 20516 2838 20528
rect 3973 20519 4031 20525
rect 3973 20516 3985 20519
rect 2832 20488 3985 20516
rect 2832 20476 2838 20488
rect 3973 20485 3985 20488
rect 4019 20485 4031 20519
rect 3973 20479 4031 20485
rect 1673 20451 1731 20457
rect 1673 20448 1685 20451
rect 1544 20420 1685 20448
rect 1544 20408 1550 20420
rect 1673 20417 1685 20420
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 1940 20451 1998 20457
rect 1940 20417 1952 20451
rect 1986 20448 1998 20451
rect 3329 20451 3387 20457
rect 3329 20448 3341 20451
rect 1986 20420 3341 20448
rect 1986 20417 1998 20420
rect 1940 20411 1998 20417
rect 3329 20417 3341 20420
rect 3375 20417 3387 20451
rect 3329 20411 3387 20417
rect 3513 20451 3571 20457
rect 3513 20417 3525 20451
rect 3559 20417 3571 20451
rect 3513 20411 3571 20417
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20417 3663 20451
rect 3878 20448 3884 20460
rect 3839 20420 3884 20448
rect 3605 20411 3663 20417
rect 3528 20380 3556 20411
rect 3160 20352 3556 20380
rect 3160 20256 3188 20352
rect 3620 20312 3648 20411
rect 3878 20408 3884 20420
rect 3936 20408 3942 20460
rect 4157 20451 4215 20457
rect 4157 20417 4169 20451
rect 4203 20448 4215 20451
rect 4341 20451 4399 20457
rect 4341 20448 4353 20451
rect 4203 20420 4353 20448
rect 4203 20417 4215 20420
rect 4157 20411 4215 20417
rect 4341 20417 4353 20420
rect 4387 20417 4399 20451
rect 4341 20411 4399 20417
rect 4617 20451 4675 20457
rect 4617 20417 4629 20451
rect 4663 20448 4675 20451
rect 4893 20451 4951 20457
rect 4893 20448 4905 20451
rect 4663 20420 4905 20448
rect 4663 20417 4675 20420
rect 4617 20411 4675 20417
rect 4893 20417 4905 20420
rect 4939 20448 4951 20451
rect 5077 20451 5135 20457
rect 5077 20448 5089 20451
rect 4939 20420 5089 20448
rect 4939 20417 4951 20420
rect 4893 20411 4951 20417
rect 5077 20417 5089 20420
rect 5123 20417 5135 20451
rect 5077 20411 5135 20417
rect 5169 20451 5227 20457
rect 5169 20417 5181 20451
rect 5215 20448 5227 20451
rect 5442 20448 5448 20460
rect 5215 20420 5448 20448
rect 5215 20417 5227 20420
rect 5169 20411 5227 20417
rect 5442 20408 5448 20420
rect 5500 20408 5506 20460
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 3786 20380 3792 20392
rect 3747 20352 3792 20380
rect 3786 20340 3792 20352
rect 3844 20340 3850 20392
rect 4154 20312 4160 20324
rect 3620 20284 4160 20312
rect 4154 20272 4160 20284
rect 4212 20312 4218 20324
rect 4709 20315 4767 20321
rect 4709 20312 4721 20315
rect 4212 20284 4721 20312
rect 4212 20272 4218 20284
rect 4709 20281 4721 20284
rect 4755 20312 4767 20315
rect 5552 20312 5580 20411
rect 5644 20380 5672 20556
rect 5925 20556 7012 20584
rect 5813 20519 5871 20525
rect 5813 20485 5825 20519
rect 5859 20516 5871 20519
rect 5925 20516 5953 20556
rect 7006 20544 7012 20556
rect 7064 20584 7070 20596
rect 7650 20584 7656 20596
rect 7064 20556 7656 20584
rect 7064 20544 7070 20556
rect 7650 20544 7656 20556
rect 7708 20584 7714 20596
rect 7745 20587 7803 20593
rect 7745 20584 7757 20587
rect 7708 20556 7757 20584
rect 7708 20544 7714 20556
rect 7745 20553 7757 20556
rect 7791 20553 7803 20587
rect 7745 20547 7803 20553
rect 8570 20544 8576 20596
rect 8628 20584 8634 20596
rect 8757 20587 8815 20593
rect 8757 20584 8769 20587
rect 8628 20556 8769 20584
rect 8628 20544 8634 20556
rect 8757 20553 8769 20556
rect 8803 20553 8815 20587
rect 9950 20584 9956 20596
rect 9911 20556 9956 20584
rect 8757 20547 8815 20553
rect 9950 20544 9956 20556
rect 10008 20544 10014 20596
rect 11330 20584 11336 20596
rect 11291 20556 11336 20584
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 11974 20544 11980 20596
rect 12032 20584 12038 20596
rect 12342 20584 12348 20596
rect 12032 20556 12348 20584
rect 12032 20544 12038 20556
rect 12342 20544 12348 20556
rect 12400 20544 12406 20596
rect 15286 20544 15292 20596
rect 15344 20584 15350 20596
rect 15565 20587 15623 20593
rect 15565 20584 15577 20587
rect 15344 20556 15577 20584
rect 15344 20544 15350 20556
rect 15565 20553 15577 20556
rect 15611 20584 15623 20587
rect 16209 20587 16267 20593
rect 16209 20584 16221 20587
rect 15611 20556 16221 20584
rect 15611 20553 15623 20556
rect 15565 20547 15623 20553
rect 16209 20553 16221 20556
rect 16255 20553 16267 20587
rect 18046 20584 18052 20596
rect 18007 20556 18052 20584
rect 16209 20547 16267 20553
rect 18046 20544 18052 20556
rect 18104 20584 18110 20596
rect 18104 20556 19196 20584
rect 18104 20544 18110 20556
rect 6914 20516 6920 20528
rect 5859 20488 5953 20516
rect 6012 20488 6920 20516
rect 5859 20485 5871 20488
rect 5813 20479 5871 20485
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 5910 20451 5968 20457
rect 5776 20420 5821 20448
rect 5776 20408 5782 20420
rect 5910 20417 5922 20451
rect 5956 20446 5968 20451
rect 6012 20446 6040 20488
rect 6914 20476 6920 20488
rect 6972 20476 6978 20528
rect 14642 20516 14648 20528
rect 11532 20488 14648 20516
rect 6621 20451 6679 20457
rect 6621 20448 6633 20451
rect 5956 20418 6040 20446
rect 6104 20420 6633 20448
rect 5956 20417 5968 20418
rect 5910 20411 5968 20417
rect 5925 20380 5953 20411
rect 5644 20352 5953 20380
rect 6104 20321 6132 20420
rect 6621 20417 6633 20420
rect 6667 20417 6679 20451
rect 9858 20448 9864 20460
rect 9819 20420 9864 20448
rect 6621 20411 6679 20417
rect 9858 20408 9864 20420
rect 9916 20408 9922 20460
rect 10870 20448 10876 20460
rect 10831 20420 10876 20448
rect 10870 20408 10876 20420
rect 10928 20408 10934 20460
rect 11146 20448 11152 20460
rect 11107 20420 11152 20448
rect 11146 20408 11152 20420
rect 11204 20408 11210 20460
rect 11238 20408 11244 20460
rect 11296 20448 11302 20460
rect 11532 20457 11560 20488
rect 14200 20457 14228 20488
rect 14642 20476 14648 20488
rect 14700 20476 14706 20528
rect 16301 20519 16359 20525
rect 16301 20485 16313 20519
rect 16347 20516 16359 20519
rect 16482 20516 16488 20528
rect 16347 20488 16488 20516
rect 16347 20485 16359 20488
rect 16301 20479 16359 20485
rect 16482 20476 16488 20488
rect 16540 20476 16546 20528
rect 18506 20516 18512 20528
rect 16684 20488 18512 20516
rect 14458 20457 14464 20460
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 11296 20420 11529 20448
rect 11296 20408 11302 20420
rect 11517 20417 11529 20420
rect 11563 20417 11575 20451
rect 11773 20451 11831 20457
rect 11773 20448 11785 20451
rect 11517 20411 11575 20417
rect 11624 20420 11785 20448
rect 6362 20380 6368 20392
rect 6323 20352 6368 20380
rect 6362 20340 6368 20352
rect 6420 20340 6426 20392
rect 11624 20380 11652 20420
rect 11773 20417 11785 20420
rect 11819 20417 11831 20451
rect 11773 20411 11831 20417
rect 14185 20451 14243 20457
rect 14185 20417 14197 20451
rect 14231 20417 14243 20451
rect 14452 20448 14464 20457
rect 14419 20420 14464 20448
rect 14185 20411 14243 20417
rect 14452 20411 14464 20420
rect 14458 20408 14464 20411
rect 14516 20408 14522 20460
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 16684 20457 16712 20488
rect 18506 20476 18512 20488
rect 18564 20476 18570 20528
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15252 20420 16037 20448
rect 15252 20408 15258 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20417 16727 20451
rect 16925 20451 16983 20457
rect 16925 20448 16937 20451
rect 16669 20411 16727 20417
rect 16776 20420 16937 20448
rect 11072 20352 11652 20380
rect 11072 20321 11100 20352
rect 16390 20340 16396 20392
rect 16448 20380 16454 20392
rect 16776 20380 16804 20420
rect 16925 20417 16937 20420
rect 16971 20417 16983 20451
rect 18598 20448 18604 20460
rect 18559 20420 18604 20448
rect 16925 20411 16983 20417
rect 18598 20408 18604 20420
rect 18656 20408 18662 20460
rect 19058 20448 19064 20460
rect 19019 20420 19064 20448
rect 19058 20408 19064 20420
rect 19116 20408 19122 20460
rect 19168 20457 19196 20556
rect 22370 20544 22376 20596
rect 22428 20584 22434 20596
rect 22557 20587 22615 20593
rect 22557 20584 22569 20587
rect 22428 20556 22569 20584
rect 22428 20544 22434 20556
rect 22557 20553 22569 20556
rect 22603 20553 22615 20587
rect 22557 20547 22615 20553
rect 19242 20476 19248 20528
rect 19300 20516 19306 20528
rect 21542 20516 21548 20528
rect 19300 20488 21548 20516
rect 19300 20476 19306 20488
rect 19153 20451 19211 20457
rect 19153 20417 19165 20451
rect 19199 20417 19211 20451
rect 19153 20411 19211 20417
rect 19886 20408 19892 20460
rect 19944 20448 19950 20460
rect 20073 20451 20131 20457
rect 20073 20448 20085 20451
rect 19944 20420 20085 20448
rect 19944 20408 19950 20420
rect 20073 20417 20085 20420
rect 20119 20417 20131 20451
rect 20073 20411 20131 20417
rect 20165 20451 20223 20457
rect 20165 20417 20177 20451
rect 20211 20448 20223 20451
rect 20901 20451 20959 20457
rect 20901 20448 20913 20451
rect 20211 20420 20913 20448
rect 20211 20417 20223 20420
rect 20165 20411 20223 20417
rect 20901 20417 20913 20420
rect 20947 20417 20959 20451
rect 21008 20448 21036 20488
rect 21542 20476 21548 20488
rect 21600 20476 21606 20528
rect 22462 20476 22468 20528
rect 22520 20516 22526 20528
rect 23017 20519 23075 20525
rect 23017 20516 23029 20519
rect 22520 20488 23029 20516
rect 22520 20476 22526 20488
rect 23017 20485 23029 20488
rect 23063 20485 23075 20519
rect 23017 20479 23075 20485
rect 23658 20476 23664 20528
rect 23716 20516 23722 20528
rect 23716 20488 24808 20516
rect 23716 20476 23722 20488
rect 21086 20451 21144 20457
rect 21086 20448 21098 20451
rect 21008 20420 21098 20448
rect 20901 20411 20959 20417
rect 21086 20417 21098 20420
rect 21132 20417 21144 20451
rect 21450 20448 21456 20460
rect 21411 20420 21456 20448
rect 21086 20411 21144 20417
rect 21450 20408 21456 20420
rect 21508 20448 21514 20460
rect 22741 20451 22799 20457
rect 22741 20448 22753 20451
rect 21508 20420 22753 20448
rect 21508 20408 21514 20420
rect 22741 20417 22753 20420
rect 22787 20417 22799 20451
rect 24302 20448 24308 20460
rect 24263 20420 24308 20448
rect 22741 20411 22799 20417
rect 24302 20408 24308 20420
rect 24360 20408 24366 20460
rect 24486 20448 24492 20460
rect 24447 20420 24492 20448
rect 24486 20408 24492 20420
rect 24544 20408 24550 20460
rect 24780 20457 24808 20488
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20417 24823 20451
rect 24765 20411 24823 20417
rect 18230 20380 18236 20392
rect 16448 20352 16804 20380
rect 18064 20352 18236 20380
rect 16448 20340 16454 20352
rect 4755 20284 5580 20312
rect 6089 20315 6147 20321
rect 4755 20281 4767 20284
rect 4709 20275 4767 20281
rect 6089 20281 6101 20315
rect 6135 20281 6147 20315
rect 6089 20275 6147 20281
rect 11057 20315 11115 20321
rect 11057 20281 11069 20315
rect 11103 20281 11115 20315
rect 11057 20275 11115 20281
rect 12728 20284 14228 20312
rect 3053 20247 3111 20253
rect 3053 20213 3065 20247
rect 3099 20244 3111 20247
rect 3142 20244 3148 20256
rect 3099 20216 3148 20244
rect 3099 20213 3111 20216
rect 3053 20207 3111 20213
rect 3142 20204 3148 20216
rect 3200 20204 3206 20256
rect 4341 20247 4399 20253
rect 4341 20213 4353 20247
rect 4387 20244 4399 20247
rect 7098 20244 7104 20256
rect 4387 20216 7104 20244
rect 4387 20213 4399 20216
rect 4341 20207 4399 20213
rect 7098 20204 7104 20216
rect 7156 20204 7162 20256
rect 8021 20247 8079 20253
rect 8021 20213 8033 20247
rect 8067 20244 8079 20247
rect 8294 20244 8300 20256
rect 8067 20216 8300 20244
rect 8067 20213 8079 20216
rect 8021 20207 8079 20213
rect 8294 20204 8300 20216
rect 8352 20204 8358 20256
rect 11330 20204 11336 20256
rect 11388 20244 11394 20256
rect 12728 20244 12756 20284
rect 12894 20244 12900 20256
rect 11388 20216 12756 20244
rect 12855 20216 12900 20244
rect 11388 20204 11394 20216
rect 12894 20204 12900 20216
rect 12952 20204 12958 20256
rect 14200 20244 14228 20284
rect 15672 20284 16712 20312
rect 15672 20244 15700 20284
rect 15838 20244 15844 20256
rect 14200 20216 15700 20244
rect 15799 20216 15844 20244
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 16684 20244 16712 20284
rect 18064 20244 18092 20352
rect 18230 20340 18236 20352
rect 18288 20340 18294 20392
rect 18690 20380 18696 20392
rect 18651 20352 18696 20380
rect 18690 20340 18696 20352
rect 18748 20340 18754 20392
rect 18785 20383 18843 20389
rect 18785 20349 18797 20383
rect 18831 20380 18843 20383
rect 20349 20383 20407 20389
rect 18831 20352 19334 20380
rect 18831 20349 18843 20352
rect 18785 20343 18843 20349
rect 16684 20216 18092 20244
rect 18233 20247 18291 20253
rect 18233 20213 18245 20247
rect 18279 20244 18291 20247
rect 18414 20244 18420 20256
rect 18279 20216 18420 20244
rect 18279 20213 18291 20216
rect 18233 20207 18291 20213
rect 18414 20204 18420 20216
rect 18472 20204 18478 20256
rect 18874 20204 18880 20256
rect 18932 20244 18938 20256
rect 19061 20247 19119 20253
rect 19061 20244 19073 20247
rect 18932 20216 19073 20244
rect 18932 20204 18938 20216
rect 19061 20213 19073 20216
rect 19107 20213 19119 20247
rect 19306 20244 19334 20352
rect 20349 20349 20361 20383
rect 20395 20380 20407 20383
rect 20530 20380 20536 20392
rect 20395 20352 20536 20380
rect 20395 20349 20407 20352
rect 20349 20343 20407 20349
rect 19426 20312 19432 20324
rect 19387 20284 19432 20312
rect 19426 20272 19432 20284
rect 19484 20272 19490 20324
rect 20364 20312 20392 20343
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 21542 20340 21548 20392
rect 21600 20380 21606 20392
rect 22925 20383 22983 20389
rect 21600 20352 21645 20380
rect 21600 20340 21606 20352
rect 22925 20349 22937 20383
rect 22971 20380 22983 20383
rect 24946 20380 24952 20392
rect 22971 20352 24952 20380
rect 22971 20349 22983 20352
rect 22925 20343 22983 20349
rect 24946 20340 24952 20352
rect 25004 20340 25010 20392
rect 24302 20312 24308 20324
rect 19536 20284 20392 20312
rect 23032 20284 24308 20312
rect 19536 20244 19564 20284
rect 19306 20216 19564 20244
rect 19061 20207 19119 20213
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 23032 20253 23060 20284
rect 24302 20272 24308 20284
rect 24360 20272 24366 20324
rect 19705 20247 19763 20253
rect 19705 20244 19717 20247
rect 19668 20216 19717 20244
rect 19668 20204 19674 20216
rect 19705 20213 19717 20216
rect 19751 20213 19763 20247
rect 19705 20207 19763 20213
rect 23017 20247 23075 20253
rect 23017 20213 23029 20247
rect 23063 20213 23075 20247
rect 23017 20207 23075 20213
rect 23842 20204 23848 20256
rect 23900 20244 23906 20256
rect 24213 20247 24271 20253
rect 24213 20244 24225 20247
rect 23900 20216 24225 20244
rect 23900 20204 23906 20216
rect 24213 20213 24225 20216
rect 24259 20213 24271 20247
rect 24578 20244 24584 20256
rect 24539 20216 24584 20244
rect 24213 20207 24271 20213
rect 24578 20204 24584 20216
rect 24636 20204 24642 20256
rect 1104 20154 26128 20176
rect 1104 20102 5120 20154
rect 5172 20102 5184 20154
rect 5236 20102 5248 20154
rect 5300 20102 5312 20154
rect 5364 20102 5376 20154
rect 5428 20102 13462 20154
rect 13514 20102 13526 20154
rect 13578 20102 13590 20154
rect 13642 20102 13654 20154
rect 13706 20102 13718 20154
rect 13770 20102 21803 20154
rect 21855 20102 21867 20154
rect 21919 20102 21931 20154
rect 21983 20102 21995 20154
rect 22047 20102 22059 20154
rect 22111 20102 26128 20154
rect 1104 20080 26128 20102
rect 4062 20040 4068 20052
rect 3344 20012 4068 20040
rect 1486 19904 1492 19916
rect 1447 19876 1492 19904
rect 1486 19864 1492 19876
rect 1544 19864 1550 19916
rect 3142 19836 3148 19848
rect 3103 19808 3148 19836
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19836 3295 19839
rect 3344 19836 3372 20012
rect 4062 20000 4068 20012
rect 4120 20040 4126 20052
rect 4120 20012 4660 20040
rect 4120 20000 4126 20012
rect 3878 19932 3884 19984
rect 3936 19972 3942 19984
rect 3936 19944 4476 19972
rect 3936 19932 3942 19944
rect 4448 19913 4476 19944
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19904 3479 19907
rect 4341 19907 4399 19913
rect 4341 19904 4353 19907
rect 3467 19876 4353 19904
rect 3467 19873 3479 19876
rect 3421 19867 3479 19873
rect 4341 19873 4353 19876
rect 4387 19873 4399 19907
rect 4341 19867 4399 19873
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 3283 19808 3372 19836
rect 4065 19839 4123 19845
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 4065 19805 4077 19839
rect 4111 19805 4123 19839
rect 4065 19799 4123 19805
rect 1756 19771 1814 19777
rect 1756 19737 1768 19771
rect 1802 19768 1814 19771
rect 3881 19771 3939 19777
rect 3881 19768 3893 19771
rect 1802 19740 3893 19768
rect 1802 19737 1814 19740
rect 1756 19731 1814 19737
rect 3881 19737 3893 19740
rect 3927 19737 3939 19771
rect 3881 19731 3939 19737
rect 4080 19768 4108 19799
rect 4154 19796 4160 19848
rect 4212 19836 4218 19848
rect 4525 19839 4583 19845
rect 4212 19808 4257 19836
rect 4212 19796 4218 19808
rect 4525 19805 4537 19839
rect 4571 19805 4583 19839
rect 4632 19836 4660 20012
rect 5718 20000 5724 20052
rect 5776 20040 5782 20052
rect 6270 20040 6276 20052
rect 5776 20012 6276 20040
rect 5776 20000 5782 20012
rect 6270 20000 6276 20012
rect 6328 20000 6334 20052
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 11701 20043 11759 20049
rect 11701 20040 11713 20043
rect 11112 20012 11713 20040
rect 11112 20000 11118 20012
rect 11701 20009 11713 20012
rect 11747 20009 11759 20043
rect 11701 20003 11759 20009
rect 14737 20043 14795 20049
rect 14737 20009 14749 20043
rect 14783 20009 14795 20043
rect 14737 20003 14795 20009
rect 11514 19932 11520 19984
rect 11572 19972 11578 19984
rect 11609 19975 11667 19981
rect 11609 19972 11621 19975
rect 11572 19944 11621 19972
rect 11572 19932 11578 19944
rect 11609 19941 11621 19944
rect 11655 19941 11667 19975
rect 12805 19975 12863 19981
rect 12805 19972 12817 19975
rect 11609 19935 11667 19941
rect 12268 19944 12817 19972
rect 8110 19904 8116 19916
rect 7116 19876 8116 19904
rect 7116 19845 7144 19876
rect 8110 19864 8116 19876
rect 8168 19904 8174 19916
rect 12268 19904 12296 19944
rect 12805 19941 12817 19944
rect 12851 19972 12863 19975
rect 14752 19972 14780 20003
rect 14826 20000 14832 20052
rect 14884 20040 14890 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 14884 20012 14933 20040
rect 14884 20000 14890 20012
rect 14921 20009 14933 20012
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 16301 20043 16359 20049
rect 16301 20009 16313 20043
rect 16347 20040 16359 20043
rect 16390 20040 16396 20052
rect 16347 20012 16396 20040
rect 16347 20009 16359 20012
rect 16301 20003 16359 20009
rect 16390 20000 16396 20012
rect 16448 20000 16454 20052
rect 16482 20000 16488 20052
rect 16540 20040 16546 20052
rect 18414 20040 18420 20052
rect 16540 20012 18000 20040
rect 18375 20012 18420 20040
rect 16540 20000 16546 20012
rect 15105 19975 15163 19981
rect 15105 19972 15117 19975
rect 12851 19944 13308 19972
rect 14752 19944 15117 19972
rect 12851 19941 12863 19944
rect 12805 19935 12863 19941
rect 8168 19876 12296 19904
rect 12345 19907 12403 19913
rect 8168 19864 8174 19876
rect 12345 19873 12357 19907
rect 12391 19904 12403 19907
rect 12894 19904 12900 19916
rect 12391 19876 12900 19904
rect 12391 19873 12403 19876
rect 12345 19867 12403 19873
rect 12894 19864 12900 19876
rect 12952 19864 12958 19916
rect 4709 19839 4767 19845
rect 4709 19836 4721 19839
rect 4632 19808 4721 19836
rect 4525 19799 4583 19805
rect 4709 19805 4721 19808
rect 4755 19805 4767 19839
rect 4709 19799 4767 19805
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19805 7159 19839
rect 7101 19799 7159 19805
rect 4430 19768 4436 19780
rect 4080 19740 4436 19768
rect 2869 19703 2927 19709
rect 2869 19669 2881 19703
rect 2915 19700 2927 19703
rect 4080 19700 4108 19740
rect 4430 19728 4436 19740
rect 4488 19768 4494 19780
rect 4540 19768 4568 19799
rect 10962 19796 10968 19848
rect 11020 19836 11026 19848
rect 11149 19839 11207 19845
rect 11149 19836 11161 19839
rect 11020 19808 11161 19836
rect 11020 19796 11026 19808
rect 4488 19740 4568 19768
rect 4488 19728 4494 19740
rect 2915 19672 4108 19700
rect 2915 19669 2927 19672
rect 2869 19663 2927 19669
rect 4246 19660 4252 19712
rect 4304 19700 4310 19712
rect 4893 19703 4951 19709
rect 4893 19700 4905 19703
rect 4304 19672 4905 19700
rect 4304 19660 4310 19672
rect 4893 19669 4905 19672
rect 4939 19669 4951 19703
rect 4893 19663 4951 19669
rect 6917 19703 6975 19709
rect 6917 19669 6929 19703
rect 6963 19700 6975 19703
rect 7098 19700 7104 19712
rect 6963 19672 7104 19700
rect 6963 19669 6975 19672
rect 6917 19663 6975 19669
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 7282 19660 7288 19712
rect 7340 19700 7346 19712
rect 8294 19700 8300 19712
rect 7340 19672 8300 19700
rect 7340 19660 7346 19672
rect 8294 19660 8300 19672
rect 8352 19700 8358 19712
rect 11072 19709 11100 19808
rect 11149 19805 11161 19808
rect 11195 19805 11207 19839
rect 11149 19799 11207 19805
rect 11241 19839 11299 19845
rect 11241 19805 11253 19839
rect 11287 19836 11299 19839
rect 11330 19836 11336 19848
rect 11287 19808 11336 19836
rect 11287 19805 11299 19808
rect 11241 19799 11299 19805
rect 11330 19796 11336 19808
rect 11388 19836 11394 19848
rect 11425 19839 11483 19845
rect 11425 19836 11437 19839
rect 11388 19808 11437 19836
rect 11388 19796 11394 19808
rect 11425 19805 11437 19808
rect 11471 19836 11483 19839
rect 11885 19839 11943 19845
rect 11885 19836 11897 19839
rect 11471 19808 11897 19836
rect 11471 19805 11483 19808
rect 11425 19799 11483 19805
rect 11885 19805 11897 19808
rect 11931 19805 11943 19839
rect 11885 19799 11943 19805
rect 11977 19839 12035 19845
rect 11977 19805 11989 19839
rect 12023 19805 12035 19839
rect 12142 19839 12200 19845
rect 12142 19836 12154 19839
rect 11977 19799 12035 19805
rect 12084 19808 12154 19836
rect 11606 19728 11612 19780
rect 11664 19768 11670 19780
rect 11992 19768 12020 19799
rect 11664 19740 12020 19768
rect 11664 19728 11670 19740
rect 11057 19703 11115 19709
rect 11057 19700 11069 19703
rect 8352 19672 11069 19700
rect 8352 19660 8358 19672
rect 11057 19669 11069 19672
rect 11103 19669 11115 19703
rect 11057 19663 11115 19669
rect 11698 19660 11704 19712
rect 11756 19700 11762 19712
rect 12084 19700 12112 19808
rect 12142 19805 12154 19808
rect 12188 19805 12200 19839
rect 12142 19799 12200 19805
rect 12250 19796 12256 19848
rect 12308 19836 12314 19848
rect 12529 19839 12587 19845
rect 12529 19836 12541 19839
rect 12308 19808 12353 19836
rect 12406 19808 12541 19836
rect 12308 19796 12314 19808
rect 12406 19780 12434 19808
rect 12529 19805 12541 19808
rect 12575 19805 12587 19839
rect 12986 19836 12992 19848
rect 12947 19808 12992 19836
rect 12529 19799 12587 19805
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 12342 19728 12348 19780
rect 12400 19740 12434 19780
rect 13280 19768 13308 19944
rect 15105 19941 15117 19944
rect 15151 19941 15163 19975
rect 15838 19972 15844 19984
rect 15105 19935 15163 19941
rect 15580 19944 15844 19972
rect 15580 19913 15608 19944
rect 15838 19932 15844 19944
rect 15896 19932 15902 19984
rect 17972 19972 18000 20012
rect 18414 20000 18420 20012
rect 18472 20000 18478 20052
rect 18966 20040 18972 20052
rect 18927 20012 18972 20040
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 19610 20040 19616 20052
rect 19571 20012 19616 20040
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 20162 20040 20168 20052
rect 20123 20012 20168 20040
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 19426 19972 19432 19984
rect 17972 19944 19432 19972
rect 19426 19932 19432 19944
rect 19484 19932 19490 19984
rect 22189 19975 22247 19981
rect 22189 19941 22201 19975
rect 22235 19941 22247 19975
rect 24302 19972 24308 19984
rect 22189 19935 22247 19941
rect 24136 19944 24308 19972
rect 15565 19907 15623 19913
rect 15565 19873 15577 19907
rect 15611 19873 15623 19907
rect 15565 19867 15623 19873
rect 15654 19864 15660 19916
rect 15712 19904 15718 19916
rect 15749 19907 15807 19913
rect 15749 19904 15761 19907
rect 15712 19876 15761 19904
rect 15712 19864 15718 19876
rect 15749 19873 15761 19876
rect 15795 19904 15807 19907
rect 15795 19876 16528 19904
rect 15795 19873 15807 19876
rect 15749 19867 15807 19873
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 14366 19836 14372 19848
rect 13872 19808 14372 19836
rect 13872 19796 13878 19808
rect 14366 19796 14372 19808
rect 14424 19796 14430 19848
rect 16022 19796 16028 19848
rect 16080 19836 16086 19848
rect 16500 19845 16528 19876
rect 16942 19864 16948 19916
rect 17000 19904 17006 19916
rect 17037 19907 17095 19913
rect 17037 19904 17049 19907
rect 17000 19876 17049 19904
rect 17000 19864 17006 19876
rect 17037 19873 17049 19876
rect 17083 19873 17095 19907
rect 17037 19867 17095 19873
rect 17221 19907 17279 19913
rect 17221 19873 17233 19907
rect 17267 19904 17279 19907
rect 17865 19907 17923 19913
rect 17865 19904 17877 19907
rect 17267 19876 17877 19904
rect 17267 19873 17279 19876
rect 17221 19867 17279 19873
rect 17865 19873 17877 19876
rect 17911 19873 17923 19907
rect 22204 19904 22232 19935
rect 22830 19904 22836 19916
rect 22204 19876 22836 19904
rect 17865 19867 17923 19873
rect 16117 19839 16175 19845
rect 16117 19836 16129 19839
rect 16080 19808 16129 19836
rect 16080 19796 16086 19808
rect 16117 19805 16129 19808
rect 16163 19805 16175 19839
rect 16117 19799 16175 19805
rect 16485 19839 16543 19845
rect 16485 19805 16497 19839
rect 16531 19836 16543 19839
rect 17236 19836 17264 19867
rect 22830 19864 22836 19876
rect 22888 19904 22894 19916
rect 24136 19913 24164 19944
rect 24302 19932 24308 19944
rect 24360 19972 24366 19984
rect 25314 19972 25320 19984
rect 24360 19944 25320 19972
rect 24360 19932 24366 19944
rect 25314 19932 25320 19944
rect 25372 19932 25378 19984
rect 22925 19907 22983 19913
rect 22925 19904 22937 19907
rect 22888 19876 22937 19904
rect 22888 19864 22894 19876
rect 22925 19873 22937 19876
rect 22971 19873 22983 19907
rect 22925 19867 22983 19873
rect 24121 19907 24179 19913
rect 24121 19873 24133 19907
rect 24167 19873 24179 19907
rect 25501 19907 25559 19913
rect 25501 19904 25513 19907
rect 24121 19867 24179 19873
rect 24688 19876 25513 19904
rect 16531 19808 17264 19836
rect 18693 19839 18751 19845
rect 16531 19805 16543 19808
rect 16485 19799 16543 19805
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 18785 19839 18843 19845
rect 18785 19836 18797 19839
rect 18739 19808 18797 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 18785 19805 18797 19808
rect 18831 19805 18843 19839
rect 18785 19799 18843 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 19981 19839 20039 19845
rect 19981 19836 19993 19839
rect 19935 19808 19993 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 19981 19805 19993 19808
rect 20027 19805 20039 19839
rect 20806 19836 20812 19848
rect 20767 19808 20812 19836
rect 19981 19799 20039 19805
rect 20806 19796 20812 19808
rect 20864 19796 20870 19848
rect 21542 19796 21548 19848
rect 21600 19836 21606 19848
rect 22558 19839 22616 19845
rect 22558 19836 22570 19839
rect 21600 19808 22570 19836
rect 21600 19796 21606 19808
rect 22558 19805 22570 19808
rect 22604 19836 22616 19839
rect 22738 19836 22744 19848
rect 22604 19808 22744 19836
rect 22604 19805 22616 19808
rect 22558 19799 22616 19805
rect 22738 19796 22744 19808
rect 22796 19796 22802 19848
rect 23017 19839 23075 19845
rect 23017 19805 23029 19839
rect 23063 19805 23075 19839
rect 23290 19836 23296 19848
rect 23251 19808 23296 19836
rect 23017 19799 23075 19805
rect 14746 19771 14804 19777
rect 14746 19768 14758 19771
rect 13280 19740 14758 19768
rect 12400 19728 12406 19740
rect 14746 19737 14758 19740
rect 14792 19768 14804 19771
rect 15286 19768 15292 19780
rect 14792 19740 15292 19768
rect 14792 19737 14804 19740
rect 14746 19731 14804 19737
rect 15286 19728 15292 19740
rect 15344 19728 15350 19780
rect 15473 19771 15531 19777
rect 15473 19737 15485 19771
rect 15519 19768 15531 19771
rect 16850 19768 16856 19780
rect 15519 19740 16856 19768
rect 15519 19737 15531 19740
rect 15473 19731 15531 19737
rect 16850 19728 16856 19740
rect 16908 19728 16914 19780
rect 18046 19768 18052 19780
rect 18007 19740 18052 19768
rect 18046 19728 18052 19740
rect 18104 19768 18110 19780
rect 19245 19771 19303 19777
rect 19245 19768 19257 19771
rect 18104 19740 19257 19768
rect 18104 19728 18110 19740
rect 19245 19737 19257 19740
rect 19291 19737 19303 19771
rect 19245 19731 19303 19737
rect 21076 19771 21134 19777
rect 21076 19737 21088 19771
rect 21122 19768 21134 19771
rect 21450 19768 21456 19780
rect 21122 19740 21456 19768
rect 21122 19737 21134 19740
rect 21076 19731 21134 19737
rect 21450 19728 21456 19740
rect 21508 19728 21514 19780
rect 22373 19771 22431 19777
rect 22373 19768 22385 19771
rect 22066 19740 22385 19768
rect 11756 19672 12112 19700
rect 11756 19660 11762 19672
rect 12158 19660 12164 19712
rect 12216 19700 12222 19712
rect 12360 19700 12388 19728
rect 12618 19700 12624 19712
rect 12216 19672 12388 19700
rect 12579 19672 12624 19700
rect 12216 19660 12222 19672
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 16574 19700 16580 19712
rect 16535 19672 16580 19700
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 16945 19703 17003 19709
rect 16945 19669 16957 19703
rect 16991 19700 17003 19703
rect 17402 19700 17408 19712
rect 16991 19672 17408 19700
rect 16991 19669 17003 19672
rect 16945 19663 17003 19669
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 18426 19703 18484 19709
rect 18426 19669 18438 19703
rect 18472 19700 18484 19703
rect 19518 19700 19524 19712
rect 18472 19672 19524 19700
rect 18472 19669 18484 19672
rect 18426 19663 18484 19669
rect 19518 19660 19524 19672
rect 19576 19700 19582 19712
rect 19622 19703 19680 19709
rect 19622 19700 19634 19703
rect 19576 19672 19634 19700
rect 19576 19660 19582 19672
rect 19622 19669 19634 19672
rect 19668 19669 19680 19703
rect 20530 19700 20536 19712
rect 20491 19672 20536 19700
rect 19622 19663 19680 19669
rect 20530 19660 20536 19672
rect 20588 19660 20594 19712
rect 21174 19660 21180 19712
rect 21232 19700 21238 19712
rect 22066 19700 22094 19740
rect 22373 19737 22385 19740
rect 22419 19737 22431 19771
rect 22373 19731 22431 19737
rect 22462 19728 22468 19780
rect 22520 19768 22526 19780
rect 23032 19768 23060 19799
rect 23290 19796 23296 19808
rect 23348 19796 23354 19848
rect 23842 19845 23848 19848
rect 23477 19839 23535 19845
rect 23477 19805 23489 19839
rect 23523 19836 23535 19839
rect 23811 19839 23848 19845
rect 23811 19836 23823 19839
rect 23523 19808 23823 19836
rect 23523 19805 23535 19808
rect 23477 19799 23535 19805
rect 23811 19805 23823 19808
rect 23811 19799 23848 19805
rect 23842 19796 23848 19799
rect 23900 19796 23906 19848
rect 24213 19839 24271 19845
rect 24213 19805 24225 19839
rect 24259 19836 24271 19839
rect 24486 19836 24492 19848
rect 24259 19808 24492 19836
rect 24259 19805 24271 19808
rect 24213 19799 24271 19805
rect 24486 19796 24492 19808
rect 24544 19836 24550 19848
rect 24688 19845 24716 19876
rect 25501 19873 25513 19876
rect 25547 19873 25559 19907
rect 25501 19867 25559 19873
rect 24639 19839 24716 19845
rect 24639 19836 24651 19839
rect 24544 19808 24651 19836
rect 24544 19796 24550 19808
rect 24639 19805 24651 19808
rect 24685 19808 24716 19839
rect 24946 19836 24952 19848
rect 24907 19808 24952 19836
rect 24685 19805 24697 19808
rect 24639 19799 24697 19805
rect 24946 19796 24952 19808
rect 25004 19796 25010 19848
rect 25038 19796 25044 19848
rect 25096 19836 25102 19848
rect 25133 19839 25191 19845
rect 25133 19836 25145 19839
rect 25096 19808 25145 19836
rect 25096 19796 25102 19808
rect 25133 19805 25145 19808
rect 25179 19805 25191 19839
rect 25133 19799 25191 19805
rect 23109 19771 23167 19777
rect 23109 19768 23121 19771
rect 22520 19740 23121 19768
rect 22520 19728 22526 19740
rect 23109 19737 23121 19740
rect 23155 19737 23167 19771
rect 23109 19731 23167 19737
rect 23934 19728 23940 19780
rect 23992 19768 23998 19780
rect 24397 19771 24455 19777
rect 24397 19768 24409 19771
rect 23992 19740 24409 19768
rect 23992 19728 23998 19740
rect 24397 19737 24409 19740
rect 24443 19737 24455 19771
rect 24964 19768 24992 19796
rect 25317 19771 25375 19777
rect 25317 19768 25329 19771
rect 24964 19740 25329 19768
rect 24397 19731 24455 19737
rect 25317 19737 25329 19740
rect 25363 19737 25375 19771
rect 25317 19731 25375 19737
rect 21232 19672 22094 19700
rect 23661 19703 23719 19709
rect 21232 19660 21238 19672
rect 23661 19669 23673 19703
rect 23707 19700 23719 19703
rect 24210 19700 24216 19712
rect 23707 19672 24216 19700
rect 23707 19669 23719 19672
rect 23661 19663 23719 19669
rect 24210 19660 24216 19672
rect 24268 19660 24274 19712
rect 1104 19610 26128 19632
rect 1104 19558 9291 19610
rect 9343 19558 9355 19610
rect 9407 19558 9419 19610
rect 9471 19558 9483 19610
rect 9535 19558 9547 19610
rect 9599 19558 17632 19610
rect 17684 19558 17696 19610
rect 17748 19558 17760 19610
rect 17812 19558 17824 19610
rect 17876 19558 17888 19610
rect 17940 19558 26128 19610
rect 1104 19536 26128 19558
rect 3513 19499 3571 19505
rect 3513 19465 3525 19499
rect 3559 19465 3571 19499
rect 3513 19459 3571 19465
rect 3528 19428 3556 19459
rect 3878 19456 3884 19508
rect 3936 19496 3942 19508
rect 4338 19496 4344 19508
rect 3936 19468 4344 19496
rect 3936 19456 3942 19468
rect 4338 19456 4344 19468
rect 4396 19496 4402 19508
rect 4433 19499 4491 19505
rect 4433 19496 4445 19499
rect 4396 19468 4445 19496
rect 4396 19456 4402 19468
rect 4433 19465 4445 19468
rect 4479 19465 4491 19499
rect 4433 19459 4491 19465
rect 5626 19456 5632 19508
rect 5684 19496 5690 19508
rect 6270 19496 6276 19508
rect 5684 19468 6276 19496
rect 5684 19456 5690 19468
rect 6270 19456 6276 19468
rect 6328 19496 6334 19508
rect 8202 19496 8208 19508
rect 6328 19468 8208 19496
rect 6328 19456 6334 19468
rect 8202 19456 8208 19468
rect 8260 19456 8266 19508
rect 8757 19499 8815 19505
rect 8757 19465 8769 19499
rect 8803 19496 8815 19499
rect 10229 19499 10287 19505
rect 8803 19468 8984 19496
rect 8803 19465 8815 19468
rect 8757 19459 8815 19465
rect 5994 19428 6000 19440
rect 3528 19400 6000 19428
rect 1486 19320 1492 19372
rect 1544 19360 1550 19372
rect 3988 19369 4016 19400
rect 5994 19388 6000 19400
rect 6052 19388 6058 19440
rect 6362 19388 6368 19440
rect 6420 19428 6426 19440
rect 8956 19428 8984 19468
rect 10229 19465 10241 19499
rect 10275 19465 10287 19499
rect 10229 19459 10287 19465
rect 10873 19499 10931 19505
rect 10873 19465 10885 19499
rect 10919 19496 10931 19499
rect 11146 19496 11152 19508
rect 10919 19468 11152 19496
rect 10919 19465 10931 19468
rect 10873 19459 10931 19465
rect 9094 19431 9152 19437
rect 9094 19428 9106 19431
rect 6420 19400 8892 19428
rect 8956 19400 9106 19428
rect 6420 19388 6426 19400
rect 2133 19363 2191 19369
rect 2133 19360 2145 19363
rect 1544 19332 2145 19360
rect 1544 19320 1550 19332
rect 2133 19329 2145 19332
rect 2179 19329 2191 19363
rect 2133 19323 2191 19329
rect 2400 19363 2458 19369
rect 2400 19329 2412 19363
rect 2446 19360 2458 19363
rect 3789 19363 3847 19369
rect 3789 19360 3801 19363
rect 2446 19332 3801 19360
rect 2446 19329 2458 19332
rect 2400 19323 2458 19329
rect 3789 19329 3801 19332
rect 3835 19329 3847 19363
rect 3789 19323 3847 19329
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19329 4031 19363
rect 3973 19323 4031 19329
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19360 4123 19363
rect 4154 19360 4160 19372
rect 4111 19332 4160 19360
rect 4111 19329 4123 19332
rect 4065 19323 4123 19329
rect 4154 19320 4160 19332
rect 4212 19320 4218 19372
rect 4338 19360 4344 19372
rect 4299 19332 4344 19360
rect 4338 19320 4344 19332
rect 4396 19320 4402 19372
rect 4617 19363 4675 19369
rect 4617 19329 4629 19363
rect 4663 19360 4675 19363
rect 5534 19360 5540 19372
rect 4663 19332 5540 19360
rect 4663 19329 4675 19332
rect 4617 19323 4675 19329
rect 5534 19320 5540 19332
rect 5592 19320 5598 19372
rect 6549 19363 6607 19369
rect 6549 19329 6561 19363
rect 6595 19360 6607 19363
rect 6638 19360 6644 19372
rect 6595 19332 6644 19360
rect 6595 19329 6607 19332
rect 6549 19323 6607 19329
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 6918 19363 6976 19369
rect 6918 19329 6930 19363
rect 6964 19360 6976 19363
rect 7006 19360 7012 19372
rect 6964 19332 7012 19360
rect 6964 19329 6976 19332
rect 6918 19323 6976 19329
rect 7006 19320 7012 19332
rect 7064 19320 7070 19372
rect 7101 19363 7159 19369
rect 7101 19329 7113 19363
rect 7147 19329 7159 19363
rect 7101 19323 7159 19329
rect 7193 19363 7251 19369
rect 7193 19329 7205 19363
rect 7239 19329 7251 19363
rect 7193 19323 7251 19329
rect 7377 19363 7435 19369
rect 7377 19329 7389 19363
rect 7423 19329 7435 19363
rect 7377 19323 7435 19329
rect 7837 19363 7895 19369
rect 7837 19329 7849 19363
rect 7883 19360 7895 19363
rect 8202 19360 8208 19372
rect 7883 19332 8208 19360
rect 7883 19329 7895 19332
rect 7837 19323 7895 19329
rect 4246 19292 4252 19304
rect 4207 19264 4252 19292
rect 4246 19252 4252 19264
rect 4304 19252 4310 19304
rect 5810 19252 5816 19304
rect 5868 19292 5874 19304
rect 6733 19295 6791 19301
rect 6733 19292 6745 19295
rect 5868 19264 6745 19292
rect 5868 19252 5874 19264
rect 6733 19261 6745 19264
rect 6779 19261 6791 19295
rect 6733 19255 6791 19261
rect 6822 19252 6828 19304
rect 6880 19292 6886 19304
rect 6880 19264 6925 19292
rect 6880 19252 6886 19264
rect 7116 19236 7144 19323
rect 7208 19292 7236 19323
rect 7282 19292 7288 19304
rect 7208 19264 7288 19292
rect 7282 19252 7288 19264
rect 7340 19252 7346 19304
rect 7392 19292 7420 19323
rect 8202 19320 8208 19332
rect 8260 19320 8266 19372
rect 8570 19360 8576 19372
rect 8531 19332 8576 19360
rect 8570 19320 8576 19332
rect 8628 19320 8634 19372
rect 8864 19369 8892 19400
rect 9094 19397 9106 19400
rect 9140 19397 9152 19431
rect 10244 19428 10272 19459
rect 11146 19456 11152 19468
rect 11204 19456 11210 19508
rect 11716 19468 11928 19496
rect 11716 19428 11744 19468
rect 10244 19400 11744 19428
rect 9094 19391 9152 19397
rect 8849 19363 8907 19369
rect 8849 19329 8861 19363
rect 8895 19329 8907 19363
rect 11054 19360 11060 19372
rect 11015 19332 11060 19360
rect 8849 19323 8907 19329
rect 11054 19320 11060 19332
rect 11112 19320 11118 19372
rect 11330 19360 11336 19372
rect 11291 19332 11336 19360
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19329 11575 19363
rect 11698 19360 11704 19372
rect 11659 19332 11704 19360
rect 11517 19323 11575 19329
rect 7392 19264 7604 19292
rect 5442 19184 5448 19236
rect 5500 19224 5506 19236
rect 7098 19224 7104 19236
rect 5500 19196 7104 19224
rect 5500 19184 5506 19196
rect 7098 19184 7104 19196
rect 7156 19184 7162 19236
rect 7466 19224 7472 19236
rect 7427 19196 7472 19224
rect 7466 19184 7472 19196
rect 7524 19184 7530 19236
rect 6454 19156 6460 19168
rect 6415 19128 6460 19156
rect 6454 19116 6460 19128
rect 6512 19116 6518 19168
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 7576 19156 7604 19264
rect 11149 19227 11207 19233
rect 11149 19193 11161 19227
rect 11195 19224 11207 19227
rect 11238 19224 11244 19236
rect 11195 19196 11244 19224
rect 11195 19193 11207 19196
rect 11149 19187 11207 19193
rect 11238 19184 11244 19196
rect 11296 19184 11302 19236
rect 11532 19224 11560 19323
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 11900 19369 11928 19468
rect 12250 19456 12256 19508
rect 12308 19496 12314 19508
rect 14090 19496 14096 19508
rect 12308 19468 14096 19496
rect 12308 19456 12314 19468
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 15286 19456 15292 19508
rect 15344 19496 15350 19508
rect 15758 19499 15816 19505
rect 15758 19496 15770 19499
rect 15344 19468 15770 19496
rect 15344 19456 15350 19468
rect 15758 19465 15770 19468
rect 15804 19465 15816 19499
rect 18690 19496 18696 19508
rect 18651 19468 18696 19496
rect 15758 19459 15816 19465
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 19518 19496 19524 19508
rect 19479 19468 19524 19496
rect 19518 19456 19524 19468
rect 19576 19496 19582 19508
rect 20266 19499 20324 19505
rect 20266 19496 20278 19499
rect 19576 19468 20278 19496
rect 19576 19456 19582 19468
rect 20266 19465 20278 19468
rect 20312 19496 20324 19499
rect 20438 19496 20444 19508
rect 20312 19468 20444 19496
rect 20312 19465 20324 19468
rect 20266 19459 20324 19465
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 21085 19499 21143 19505
rect 21085 19465 21097 19499
rect 21131 19496 21143 19499
rect 21174 19496 21180 19508
rect 21131 19468 21180 19496
rect 21131 19465 21143 19468
rect 21085 19459 21143 19465
rect 21174 19456 21180 19468
rect 21232 19456 21238 19508
rect 21450 19496 21456 19508
rect 21411 19468 21456 19496
rect 21450 19456 21456 19468
rect 21508 19456 21514 19508
rect 22738 19496 22744 19508
rect 22699 19468 22744 19496
rect 22738 19456 22744 19468
rect 22796 19456 22802 19508
rect 23842 19496 23848 19508
rect 22848 19468 23848 19496
rect 11992 19400 12434 19428
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19329 11851 19363
rect 11793 19323 11851 19329
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 11808 19292 11836 19323
rect 11992 19292 12020 19400
rect 12069 19363 12127 19369
rect 12069 19329 12081 19363
rect 12115 19360 12127 19363
rect 12158 19360 12164 19372
rect 12115 19332 12164 19360
rect 12115 19329 12127 19332
rect 12069 19323 12127 19329
rect 12158 19320 12164 19332
rect 12216 19320 12222 19372
rect 11808 19264 12020 19292
rect 11606 19224 11612 19236
rect 11532 19196 11612 19224
rect 11606 19184 11612 19196
rect 11664 19184 11670 19236
rect 11882 19184 11888 19236
rect 11940 19224 11946 19236
rect 12176 19224 12204 19320
rect 12406 19292 12434 19400
rect 12618 19388 12624 19440
rect 12676 19428 12682 19440
rect 12958 19431 13016 19437
rect 12958 19428 12970 19431
rect 12676 19400 12970 19428
rect 12676 19388 12682 19400
rect 12958 19397 12970 19400
rect 13004 19397 13016 19431
rect 12958 19391 13016 19397
rect 14366 19388 14372 19440
rect 14424 19428 14430 19440
rect 15381 19431 15439 19437
rect 15381 19428 15393 19431
rect 14424 19400 15393 19428
rect 14424 19388 14430 19400
rect 15381 19397 15393 19400
rect 15427 19428 15439 19431
rect 18046 19428 18052 19440
rect 15427 19400 18052 19428
rect 15427 19397 15439 19400
rect 15381 19391 15439 19397
rect 18046 19388 18052 19400
rect 18104 19388 18110 19440
rect 18874 19428 18880 19440
rect 18248 19400 18880 19428
rect 16022 19360 16028 19372
rect 15983 19332 16028 19360
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 18248 19369 18276 19400
rect 18874 19388 18880 19400
rect 18932 19388 18938 19440
rect 19610 19388 19616 19440
rect 19668 19428 19674 19440
rect 19889 19431 19947 19437
rect 19889 19428 19901 19431
rect 19668 19400 19901 19428
rect 19668 19388 19674 19400
rect 19889 19397 19901 19400
rect 19935 19397 19947 19431
rect 19889 19391 19947 19397
rect 20548 19400 21680 19428
rect 18233 19363 18291 19369
rect 18233 19329 18245 19363
rect 18279 19329 18291 19363
rect 18233 19323 18291 19329
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 18543 19363 18601 19369
rect 18543 19360 18555 19363
rect 18380 19332 18555 19360
rect 18380 19320 18386 19332
rect 18543 19329 18555 19332
rect 18589 19329 18601 19363
rect 19058 19360 19064 19372
rect 18543 19323 18601 19329
rect 18708 19332 19064 19360
rect 12526 19292 12532 19304
rect 12406 19264 12532 19292
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 12618 19252 12624 19304
rect 12676 19292 12682 19304
rect 12713 19295 12771 19301
rect 12713 19292 12725 19295
rect 12676 19264 12725 19292
rect 12676 19252 12682 19264
rect 12713 19261 12725 19264
rect 12759 19261 12771 19295
rect 12713 19255 12771 19261
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15654 19292 15660 19304
rect 15059 19264 15660 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15654 19252 15660 19264
rect 15712 19252 15718 19304
rect 18141 19295 18199 19301
rect 18141 19261 18153 19295
rect 18187 19292 18199 19295
rect 18708 19292 18736 19332
rect 19058 19320 19064 19332
rect 19116 19320 19122 19372
rect 19702 19360 19708 19372
rect 19663 19332 19708 19360
rect 19702 19320 19708 19332
rect 19760 19360 19766 19372
rect 20548 19369 20576 19400
rect 20533 19363 20591 19369
rect 19760 19332 20484 19360
rect 19760 19320 19766 19332
rect 18187 19264 18736 19292
rect 20456 19292 20484 19332
rect 20533 19329 20545 19363
rect 20579 19329 20591 19363
rect 20990 19360 20996 19372
rect 20951 19332 20996 19360
rect 20533 19323 20591 19329
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 21652 19369 21680 19400
rect 22462 19388 22468 19440
rect 22520 19388 22526 19440
rect 22848 19428 22876 19468
rect 22572 19400 22876 19428
rect 21637 19363 21695 19369
rect 21637 19329 21649 19363
rect 21683 19329 21695 19363
rect 21637 19323 21695 19329
rect 22155 19363 22213 19369
rect 22155 19329 22167 19363
rect 22201 19360 22213 19363
rect 22480 19360 22508 19388
rect 22201 19332 22508 19360
rect 22201 19329 22213 19332
rect 22155 19323 22213 19329
rect 20898 19292 20904 19304
rect 20456 19264 20904 19292
rect 18187 19261 18199 19264
rect 18141 19255 18199 19261
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 21266 19292 21272 19304
rect 21227 19264 21272 19292
rect 21266 19252 21272 19264
rect 21324 19252 21330 19304
rect 22572 19301 22600 19400
rect 23124 19369 23152 19468
rect 23842 19456 23848 19468
rect 23900 19456 23906 19508
rect 24946 19456 24952 19508
rect 25004 19496 25010 19508
rect 25501 19499 25559 19505
rect 25501 19496 25513 19499
rect 25004 19468 25513 19496
rect 25004 19456 25010 19468
rect 25501 19465 25513 19468
rect 25547 19465 25559 19499
rect 25501 19459 25559 19465
rect 23566 19388 23572 19440
rect 23624 19437 23630 19440
rect 23624 19428 23636 19437
rect 25406 19428 25412 19440
rect 23624 19400 23669 19428
rect 23860 19400 25412 19428
rect 23624 19391 23636 19400
rect 23624 19388 23630 19391
rect 23109 19363 23167 19369
rect 23109 19329 23121 19363
rect 23155 19329 23167 19363
rect 23109 19323 23167 19329
rect 23198 19320 23204 19372
rect 23256 19360 23262 19372
rect 23860 19369 23888 19400
rect 25406 19388 25412 19400
rect 25464 19388 25470 19440
rect 23845 19363 23903 19369
rect 23256 19332 23301 19360
rect 23256 19320 23262 19332
rect 23845 19329 23857 19363
rect 23891 19329 23903 19363
rect 23845 19323 23903 19329
rect 24388 19363 24446 19369
rect 24388 19329 24400 19363
rect 24434 19360 24446 19363
rect 25222 19360 25228 19372
rect 24434 19332 25228 19360
rect 24434 19329 24446 19332
rect 24388 19323 24446 19329
rect 25222 19320 25228 19332
rect 25280 19320 25286 19372
rect 22465 19295 22523 19301
rect 22465 19261 22477 19295
rect 22511 19261 22523 19295
rect 22465 19255 22523 19261
rect 22557 19295 22615 19301
rect 22557 19261 22569 19295
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 12345 19227 12403 19233
rect 12345 19224 12357 19227
rect 11940 19196 12357 19224
rect 11940 19184 11946 19196
rect 12345 19193 12357 19196
rect 12391 19193 12403 19227
rect 12345 19187 12403 19193
rect 14734 19184 14740 19236
rect 14792 19224 14798 19236
rect 17954 19224 17960 19236
rect 14792 19196 17960 19224
rect 14792 19184 14798 19196
rect 17954 19184 17960 19196
rect 18012 19184 18018 19236
rect 20625 19227 20683 19233
rect 20625 19224 20637 19227
rect 20272 19196 20637 19224
rect 6880 19128 7604 19156
rect 7745 19159 7803 19165
rect 6880 19116 6886 19128
rect 7745 19125 7757 19159
rect 7791 19156 7803 19159
rect 8294 19156 8300 19168
rect 7791 19128 8300 19156
rect 7791 19125 7803 19128
rect 7745 19119 7803 19125
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 10781 19159 10839 19165
rect 10781 19125 10793 19159
rect 10827 19156 10839 19159
rect 11900 19156 11928 19184
rect 12158 19156 12164 19168
rect 10827 19128 11928 19156
rect 12119 19128 12164 19156
rect 10827 19125 10839 19128
rect 10781 19119 10839 19125
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 15749 19159 15807 19165
rect 15749 19125 15761 19159
rect 15795 19156 15807 19159
rect 16574 19156 16580 19168
rect 15795 19128 16580 19156
rect 15795 19125 15807 19128
rect 15749 19119 15807 19125
rect 16574 19116 16580 19128
rect 16632 19116 16638 19168
rect 20272 19165 20300 19196
rect 20625 19193 20637 19196
rect 20671 19193 20683 19227
rect 20625 19187 20683 19193
rect 22186 19184 22192 19236
rect 22244 19224 22250 19236
rect 22480 19224 22508 19255
rect 22830 19252 22836 19304
rect 22888 19292 22894 19304
rect 23017 19295 23075 19301
rect 23017 19292 23029 19295
rect 22888 19264 23029 19292
rect 22888 19252 22894 19264
rect 23017 19261 23029 19264
rect 23063 19261 23075 19295
rect 23017 19255 23075 19261
rect 24026 19252 24032 19304
rect 24084 19292 24090 19304
rect 24121 19295 24179 19301
rect 24121 19292 24133 19295
rect 24084 19264 24133 19292
rect 24084 19252 24090 19264
rect 24121 19261 24133 19264
rect 24167 19261 24179 19295
rect 24121 19255 24179 19261
rect 22244 19196 23152 19224
rect 22244 19184 22250 19196
rect 20257 19159 20315 19165
rect 20257 19125 20269 19159
rect 20303 19125 20315 19159
rect 20257 19119 20315 19125
rect 20530 19116 20536 19168
rect 20588 19156 20594 19168
rect 21266 19156 21272 19168
rect 20588 19128 21272 19156
rect 20588 19116 20594 19128
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 22005 19159 22063 19165
rect 22005 19125 22017 19159
rect 22051 19156 22063 19159
rect 22278 19156 22284 19168
rect 22051 19128 22284 19156
rect 22051 19125 22063 19128
rect 22005 19119 22063 19125
rect 22278 19116 22284 19128
rect 22336 19116 22342 19168
rect 23124 19165 23152 19196
rect 23109 19159 23167 19165
rect 23109 19125 23121 19159
rect 23155 19156 23167 19159
rect 23290 19156 23296 19168
rect 23155 19128 23296 19156
rect 23155 19125 23167 19128
rect 23109 19119 23167 19125
rect 23290 19116 23296 19128
rect 23348 19116 23354 19168
rect 23474 19116 23480 19168
rect 23532 19156 23538 19168
rect 23569 19159 23627 19165
rect 23569 19156 23581 19159
rect 23532 19128 23581 19156
rect 23532 19116 23538 19128
rect 23569 19125 23581 19128
rect 23615 19125 23627 19159
rect 23569 19119 23627 19125
rect 1104 19066 26128 19088
rect 1104 19014 5120 19066
rect 5172 19014 5184 19066
rect 5236 19014 5248 19066
rect 5300 19014 5312 19066
rect 5364 19014 5376 19066
rect 5428 19014 13462 19066
rect 13514 19014 13526 19066
rect 13578 19014 13590 19066
rect 13642 19014 13654 19066
rect 13706 19014 13718 19066
rect 13770 19014 21803 19066
rect 21855 19014 21867 19066
rect 21919 19014 21931 19066
rect 21983 19014 21995 19066
rect 22047 19014 22059 19066
rect 22111 19014 26128 19066
rect 1104 18992 26128 19014
rect 4890 18912 4896 18964
rect 4948 18952 4954 18964
rect 5537 18955 5595 18961
rect 5537 18952 5549 18955
rect 4948 18924 5549 18952
rect 4948 18912 4954 18924
rect 5537 18921 5549 18924
rect 5583 18952 5595 18955
rect 5902 18952 5908 18964
rect 5583 18924 5908 18952
rect 5583 18921 5595 18924
rect 5537 18915 5595 18921
rect 5902 18912 5908 18924
rect 5960 18952 5966 18964
rect 6822 18952 6828 18964
rect 5960 18924 6828 18952
rect 5960 18912 5966 18924
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 8478 18912 8484 18964
rect 8536 18952 8542 18964
rect 9033 18955 9091 18961
rect 9033 18952 9045 18955
rect 8536 18924 9045 18952
rect 8536 18912 8542 18924
rect 9033 18921 9045 18924
rect 9079 18952 9091 18955
rect 10686 18952 10692 18964
rect 9079 18924 10692 18952
rect 9079 18921 9091 18924
rect 9033 18915 9091 18921
rect 10686 18912 10692 18924
rect 10744 18912 10750 18964
rect 15657 18955 15715 18961
rect 15657 18921 15669 18955
rect 15703 18952 15715 18955
rect 16574 18952 16580 18964
rect 15703 18924 16580 18952
rect 15703 18921 15715 18924
rect 15657 18915 15715 18921
rect 16574 18912 16580 18924
rect 16632 18952 16638 18964
rect 17218 18952 17224 18964
rect 16632 18924 17224 18952
rect 16632 18912 16638 18924
rect 17218 18912 17224 18924
rect 17276 18912 17282 18964
rect 20441 18955 20499 18961
rect 20441 18921 20453 18955
rect 20487 18952 20499 18955
rect 21726 18952 21732 18964
rect 20487 18924 21732 18952
rect 20487 18921 20499 18924
rect 20441 18915 20499 18921
rect 21726 18912 21732 18924
rect 21784 18912 21790 18964
rect 22186 18952 22192 18964
rect 22147 18924 22192 18952
rect 22186 18912 22192 18924
rect 22244 18912 22250 18964
rect 23109 18955 23167 18961
rect 23109 18921 23121 18955
rect 23155 18921 23167 18955
rect 23109 18915 23167 18921
rect 23293 18955 23351 18961
rect 23293 18921 23305 18955
rect 23339 18952 23351 18955
rect 23658 18952 23664 18964
rect 23339 18924 23664 18952
rect 23339 18921 23351 18924
rect 23293 18915 23351 18921
rect 5626 18844 5632 18896
rect 5684 18844 5690 18896
rect 11241 18887 11299 18893
rect 11241 18853 11253 18887
rect 11287 18884 11299 18887
rect 11606 18884 11612 18896
rect 11287 18856 11612 18884
rect 11287 18853 11299 18856
rect 11241 18847 11299 18853
rect 11606 18844 11612 18856
rect 11664 18844 11670 18896
rect 17126 18884 17132 18896
rect 17087 18856 17132 18884
rect 17126 18844 17132 18856
rect 17184 18884 17190 18896
rect 20622 18884 20628 18896
rect 17184 18856 17908 18884
rect 20583 18856 20628 18884
rect 17184 18844 17190 18856
rect 5644 18816 5672 18844
rect 17880 18825 17908 18856
rect 20622 18844 20628 18856
rect 20680 18844 20686 18896
rect 23124 18884 23152 18915
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 25222 18952 25228 18964
rect 25183 18924 25228 18952
rect 25222 18912 25228 18924
rect 25280 18912 25286 18964
rect 24397 18887 24455 18893
rect 24397 18884 24409 18887
rect 23124 18856 24409 18884
rect 24397 18853 24409 18856
rect 24443 18853 24455 18887
rect 24397 18847 24455 18853
rect 5368 18788 5672 18816
rect 17865 18819 17923 18825
rect 4246 18708 4252 18760
rect 4304 18748 4310 18760
rect 5368 18757 5396 18788
rect 17865 18785 17877 18819
rect 17911 18785 17923 18819
rect 17865 18779 17923 18785
rect 20088 18788 20944 18816
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 4304 18720 5365 18748
rect 4304 18708 4310 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5626 18748 5632 18760
rect 5587 18720 5632 18748
rect 5353 18711 5411 18717
rect 5626 18708 5632 18720
rect 5684 18708 5690 18760
rect 5896 18751 5954 18757
rect 5896 18717 5908 18751
rect 5942 18748 5954 18751
rect 6454 18748 6460 18760
rect 5942 18720 6460 18748
rect 5942 18717 5954 18720
rect 5896 18711 5954 18717
rect 6454 18708 6460 18720
rect 6512 18708 6518 18760
rect 7190 18748 7196 18760
rect 7151 18720 7196 18748
rect 7190 18708 7196 18720
rect 7248 18748 7254 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 7248 18720 10425 18748
rect 7248 18708 7254 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11146 18748 11152 18760
rect 11103 18720 11152 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 11146 18708 11152 18720
rect 11204 18708 11210 18760
rect 11514 18748 11520 18760
rect 11475 18720 11520 18748
rect 11514 18708 11520 18720
rect 11572 18708 11578 18760
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18748 11851 18751
rect 12618 18748 12624 18760
rect 11839 18720 12624 18748
rect 11839 18717 11851 18720
rect 11793 18711 11851 18717
rect 12618 18708 12624 18720
rect 12676 18748 12682 18760
rect 13354 18748 13360 18760
rect 12676 18720 13360 18748
rect 12676 18708 12682 18720
rect 13354 18708 13360 18720
rect 13412 18748 13418 18760
rect 14277 18751 14335 18757
rect 14277 18748 14289 18751
rect 13412 18720 14289 18748
rect 13412 18708 13418 18720
rect 14277 18717 14289 18720
rect 14323 18748 14335 18751
rect 15102 18748 15108 18760
rect 14323 18720 15108 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 19610 18708 19616 18760
rect 19668 18748 19674 18760
rect 20088 18757 20116 18788
rect 20073 18751 20131 18757
rect 20073 18748 20085 18751
rect 19668 18720 20085 18748
rect 19668 18708 19674 18720
rect 20073 18717 20085 18720
rect 20119 18717 20131 18751
rect 20806 18748 20812 18760
rect 20767 18720 20812 18748
rect 20073 18711 20131 18717
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 20916 18748 20944 18788
rect 23198 18776 23204 18828
rect 23256 18776 23262 18828
rect 23934 18816 23940 18828
rect 23895 18788 23940 18816
rect 23934 18776 23940 18788
rect 23992 18776 23998 18828
rect 24121 18819 24179 18825
rect 24121 18785 24133 18819
rect 24167 18785 24179 18819
rect 24121 18779 24179 18785
rect 22741 18751 22799 18757
rect 22741 18748 22753 18751
rect 20916 18720 22753 18748
rect 22741 18717 22753 18720
rect 22787 18748 22799 18751
rect 23216 18748 23244 18776
rect 22787 18720 23244 18748
rect 22787 18717 22799 18720
rect 22741 18711 22799 18717
rect 5166 18640 5172 18692
rect 5224 18680 5230 18692
rect 7098 18680 7104 18692
rect 5224 18652 7104 18680
rect 5224 18640 5230 18652
rect 7098 18640 7104 18652
rect 7156 18640 7162 18692
rect 7466 18689 7472 18692
rect 7460 18680 7472 18689
rect 7427 18652 7472 18680
rect 7460 18643 7472 18652
rect 7466 18640 7472 18643
rect 7524 18640 7530 18692
rect 10168 18683 10226 18689
rect 10168 18649 10180 18683
rect 10214 18680 10226 18683
rect 10502 18680 10508 18692
rect 10214 18652 10508 18680
rect 10214 18649 10226 18652
rect 10168 18643 10226 18649
rect 10502 18640 10508 18652
rect 10560 18640 10566 18692
rect 12060 18683 12118 18689
rect 12060 18649 12072 18683
rect 12106 18680 12118 18683
rect 12158 18680 12164 18692
rect 12106 18652 12164 18680
rect 12106 18649 12118 18652
rect 12060 18643 12118 18649
rect 12158 18640 12164 18652
rect 12216 18640 12222 18692
rect 14544 18683 14602 18689
rect 14544 18649 14556 18683
rect 14590 18680 14602 18683
rect 15562 18680 15568 18692
rect 14590 18652 15568 18680
rect 14590 18649 14602 18652
rect 14544 18643 14602 18649
rect 15562 18640 15568 18652
rect 15620 18640 15626 18692
rect 16485 18683 16543 18689
rect 16485 18680 16497 18683
rect 16132 18652 16497 18680
rect 16132 18624 16160 18652
rect 16485 18649 16497 18652
rect 16531 18680 16543 18683
rect 17034 18680 17040 18692
rect 16531 18652 17040 18680
rect 16531 18649 16543 18652
rect 16485 18643 16543 18649
rect 17034 18640 17040 18652
rect 17092 18640 17098 18692
rect 20438 18640 20444 18692
rect 20496 18689 20502 18692
rect 21082 18689 21088 18692
rect 20496 18680 20508 18689
rect 20496 18652 20541 18680
rect 20496 18643 20508 18652
rect 21076 18643 21088 18689
rect 21140 18680 21146 18692
rect 23155 18683 23213 18689
rect 23155 18680 23167 18683
rect 21140 18652 21176 18680
rect 22066 18652 23167 18680
rect 20496 18640 20502 18643
rect 21082 18640 21088 18643
rect 21140 18640 21146 18652
rect 3786 18572 3792 18624
rect 3844 18612 3850 18624
rect 4157 18615 4215 18621
rect 4157 18612 4169 18615
rect 3844 18584 4169 18612
rect 3844 18572 3850 18584
rect 4157 18581 4169 18584
rect 4203 18612 4215 18615
rect 6822 18612 6828 18624
rect 4203 18584 6828 18612
rect 4203 18581 4215 18584
rect 4157 18575 4215 18581
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 6914 18572 6920 18624
rect 6972 18612 6978 18624
rect 7009 18615 7067 18621
rect 7009 18612 7021 18615
rect 6972 18584 7021 18612
rect 6972 18572 6978 18584
rect 7009 18581 7021 18584
rect 7055 18612 7067 18615
rect 7650 18612 7656 18624
rect 7055 18584 7656 18612
rect 7055 18581 7067 18584
rect 7009 18575 7067 18581
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 8386 18572 8392 18624
rect 8444 18612 8450 18624
rect 8573 18615 8631 18621
rect 8573 18612 8585 18615
rect 8444 18584 8585 18612
rect 8444 18572 8450 18584
rect 8573 18581 8585 18584
rect 8619 18581 8631 18615
rect 11330 18612 11336 18624
rect 11243 18584 11336 18612
rect 8573 18575 8631 18581
rect 11330 18572 11336 18584
rect 11388 18612 11394 18624
rect 11974 18612 11980 18624
rect 11388 18584 11980 18612
rect 11388 18572 11394 18584
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12526 18572 12532 18624
rect 12584 18612 12590 18624
rect 13173 18615 13231 18621
rect 13173 18612 13185 18615
rect 12584 18584 13185 18612
rect 12584 18572 12590 18584
rect 13173 18581 13185 18584
rect 13219 18612 13231 18615
rect 14826 18612 14832 18624
rect 13219 18584 14832 18612
rect 13219 18581 13231 18584
rect 13173 18575 13231 18581
rect 14826 18572 14832 18584
rect 14884 18572 14890 18624
rect 16114 18612 16120 18624
rect 16075 18584 16120 18612
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16390 18612 16396 18624
rect 16351 18584 16396 18612
rect 16390 18572 16396 18584
rect 16448 18572 16454 18624
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 16942 18612 16948 18624
rect 16724 18584 16948 18612
rect 16724 18572 16730 18584
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 17218 18572 17224 18624
rect 17276 18612 17282 18624
rect 17313 18615 17371 18621
rect 17313 18612 17325 18615
rect 17276 18584 17325 18612
rect 17276 18572 17282 18584
rect 17313 18581 17325 18584
rect 17359 18581 17371 18615
rect 17313 18575 17371 18581
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 17681 18615 17739 18621
rect 17681 18612 17693 18615
rect 17552 18584 17693 18612
rect 17552 18572 17558 18584
rect 17681 18581 17693 18584
rect 17727 18581 17739 18615
rect 17681 18575 17739 18581
rect 17773 18615 17831 18621
rect 17773 18581 17785 18615
rect 17819 18612 17831 18615
rect 18230 18612 18236 18624
rect 17819 18584 18236 18612
rect 17819 18581 17831 18584
rect 17773 18575 17831 18581
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 21358 18572 21364 18624
rect 21416 18612 21422 18624
rect 22066 18612 22094 18652
rect 23155 18649 23167 18652
rect 23201 18680 23213 18683
rect 23566 18680 23572 18692
rect 23201 18652 23572 18680
rect 23201 18649 23213 18652
rect 23155 18643 23213 18649
rect 23566 18640 23572 18652
rect 23624 18640 23630 18692
rect 24136 18680 24164 18779
rect 24210 18776 24216 18828
rect 24268 18816 24274 18828
rect 24857 18819 24915 18825
rect 24857 18816 24869 18819
rect 24268 18788 24869 18816
rect 24268 18776 24274 18788
rect 24857 18785 24869 18788
rect 24903 18785 24915 18819
rect 24857 18779 24915 18785
rect 25041 18819 25099 18825
rect 25041 18785 25053 18819
rect 25087 18816 25099 18819
rect 25501 18819 25559 18825
rect 25501 18816 25513 18819
rect 25087 18788 25513 18816
rect 25087 18785 25099 18788
rect 25041 18779 25099 18785
rect 24765 18683 24823 18689
rect 24136 18652 24256 18680
rect 24228 18624 24256 18652
rect 24765 18649 24777 18683
rect 24811 18680 24823 18683
rect 25130 18680 25136 18692
rect 24811 18652 25136 18680
rect 24811 18649 24823 18652
rect 24765 18643 24823 18649
rect 25130 18640 25136 18652
rect 25188 18640 25194 18692
rect 23474 18612 23480 18624
rect 21416 18584 22094 18612
rect 23435 18584 23480 18612
rect 21416 18572 21422 18584
rect 23474 18572 23480 18584
rect 23532 18572 23538 18624
rect 23842 18612 23848 18624
rect 23803 18584 23848 18612
rect 23842 18572 23848 18584
rect 23900 18572 23906 18624
rect 24210 18612 24216 18624
rect 24123 18584 24216 18612
rect 24210 18572 24216 18584
rect 24268 18612 24274 18624
rect 25240 18612 25268 18788
rect 25501 18785 25513 18788
rect 25547 18785 25559 18819
rect 25501 18779 25559 18785
rect 25406 18748 25412 18760
rect 25367 18720 25412 18748
rect 25406 18708 25412 18720
rect 25464 18708 25470 18760
rect 24268 18584 25268 18612
rect 24268 18572 24274 18584
rect 1104 18522 26128 18544
rect 1104 18470 9291 18522
rect 9343 18470 9355 18522
rect 9407 18470 9419 18522
rect 9471 18470 9483 18522
rect 9535 18470 9547 18522
rect 9599 18470 17632 18522
rect 17684 18470 17696 18522
rect 17748 18470 17760 18522
rect 17812 18470 17824 18522
rect 17876 18470 17888 18522
rect 17940 18470 26128 18522
rect 1104 18448 26128 18470
rect 3694 18408 3700 18420
rect 3160 18380 3700 18408
rect 3160 18340 3188 18380
rect 3694 18368 3700 18380
rect 3752 18368 3758 18420
rect 4341 18411 4399 18417
rect 4341 18377 4353 18411
rect 4387 18377 4399 18411
rect 5534 18408 5540 18420
rect 4341 18371 4399 18377
rect 4540 18380 5540 18408
rect 3068 18312 3188 18340
rect 3068 18281 3096 18312
rect 3234 18300 3240 18352
rect 3292 18340 3298 18352
rect 4356 18340 4384 18371
rect 3292 18312 4384 18340
rect 3292 18300 3298 18312
rect 3053 18275 3111 18281
rect 3053 18241 3065 18275
rect 3099 18241 3111 18275
rect 3053 18235 3111 18241
rect 3142 18232 3148 18284
rect 3200 18272 3206 18284
rect 3422 18275 3480 18281
rect 3422 18272 3434 18275
rect 3200 18244 3434 18272
rect 3200 18232 3206 18244
rect 3422 18241 3434 18244
rect 3468 18241 3480 18275
rect 3422 18235 3480 18241
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 3786 18272 3792 18284
rect 3747 18244 3792 18272
rect 3605 18235 3663 18241
rect 3234 18204 3240 18216
rect 3195 18176 3240 18204
rect 3234 18164 3240 18176
rect 3292 18164 3298 18216
rect 3329 18207 3387 18213
rect 3329 18173 3341 18207
rect 3375 18173 3387 18207
rect 3620 18204 3648 18235
rect 3786 18232 3792 18244
rect 3844 18232 3850 18284
rect 4246 18272 4252 18284
rect 4207 18244 4252 18272
rect 4246 18232 4252 18244
rect 4304 18232 4310 18284
rect 4540 18281 4568 18380
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 5718 18408 5724 18420
rect 5635 18380 5724 18408
rect 4632 18312 5304 18340
rect 4632 18281 4660 18312
rect 4525 18275 4583 18281
rect 4525 18241 4537 18275
rect 4571 18241 4583 18275
rect 4525 18235 4583 18241
rect 4617 18275 4675 18281
rect 4617 18241 4629 18275
rect 4663 18241 4675 18275
rect 4798 18272 4804 18284
rect 4759 18244 4804 18272
rect 4617 18235 4675 18241
rect 3620 18176 4016 18204
rect 3329 18167 3387 18173
rect 2866 18136 2872 18148
rect 2827 18108 2872 18136
rect 2866 18096 2872 18108
rect 2924 18096 2930 18148
rect 3344 18136 3372 18167
rect 3988 18145 4016 18176
rect 4338 18164 4344 18216
rect 4396 18204 4402 18216
rect 4632 18204 4660 18235
rect 4798 18232 4804 18244
rect 4856 18232 4862 18284
rect 4890 18232 4896 18284
rect 4948 18272 4954 18284
rect 5166 18272 5172 18284
rect 4948 18244 4993 18272
rect 5127 18244 5172 18272
rect 4948 18232 4954 18244
rect 5166 18232 5172 18244
rect 5224 18232 5230 18284
rect 5276 18272 5304 18312
rect 5635 18287 5663 18380
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 7742 18408 7748 18420
rect 6288 18380 7748 18408
rect 5442 18272 5448 18284
rect 5500 18281 5506 18284
rect 5610 18281 5668 18287
rect 5276 18244 5448 18272
rect 5442 18232 5448 18244
rect 5500 18235 5509 18281
rect 5610 18247 5622 18281
rect 5656 18247 5668 18281
rect 5610 18241 5668 18247
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18272 5779 18275
rect 5902 18272 5908 18284
rect 5767 18244 5908 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 5500 18232 5506 18235
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 6288 18272 6316 18380
rect 7742 18368 7748 18380
rect 7800 18368 7806 18420
rect 8481 18411 8539 18417
rect 8481 18377 8493 18411
rect 8527 18408 8539 18411
rect 8570 18408 8576 18420
rect 8527 18380 8576 18408
rect 8527 18377 8539 18380
rect 8481 18371 8539 18377
rect 8570 18368 8576 18380
rect 8628 18368 8634 18420
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 14734 18408 14740 18420
rect 13872 18380 14740 18408
rect 13872 18368 13878 18380
rect 14734 18368 14740 18380
rect 14792 18368 14798 18420
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 15562 18408 15568 18420
rect 14884 18380 15147 18408
rect 15523 18380 15568 18408
rect 14884 18368 14890 18380
rect 7190 18340 7196 18352
rect 6380 18312 7196 18340
rect 6380 18281 6408 18312
rect 7190 18300 7196 18312
rect 7248 18340 7254 18352
rect 7834 18340 7840 18352
rect 7248 18312 7840 18340
rect 7248 18300 7254 18312
rect 7834 18300 7840 18312
rect 7892 18300 7898 18352
rect 8110 18340 8116 18352
rect 8071 18312 8116 18340
rect 8110 18300 8116 18312
rect 8168 18300 8174 18352
rect 8297 18343 8355 18349
rect 8297 18309 8309 18343
rect 8343 18340 8355 18343
rect 8386 18340 8392 18352
rect 8343 18312 8392 18340
rect 8343 18309 8355 18312
rect 8297 18303 8355 18309
rect 8386 18300 8392 18312
rect 8444 18300 8450 18352
rect 9674 18340 9680 18352
rect 9587 18312 9680 18340
rect 9674 18300 9680 18312
rect 9732 18340 9738 18352
rect 11238 18340 11244 18352
rect 9732 18312 11244 18340
rect 9732 18300 9738 18312
rect 11238 18300 11244 18312
rect 11296 18340 11302 18352
rect 11333 18343 11391 18349
rect 11333 18340 11345 18343
rect 11296 18312 11345 18340
rect 11296 18300 11302 18312
rect 11333 18309 11345 18312
rect 11379 18340 11391 18343
rect 11379 18312 11928 18340
rect 11379 18309 11391 18312
rect 11333 18303 11391 18309
rect 11900 18284 11928 18312
rect 15119 18287 15147 18380
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 16666 18368 16672 18420
rect 16724 18408 16730 18420
rect 18969 18411 19027 18417
rect 18969 18408 18981 18411
rect 16724 18380 18981 18408
rect 16724 18368 16730 18380
rect 18969 18377 18981 18380
rect 19015 18408 19027 18411
rect 20806 18408 20812 18420
rect 19015 18380 20812 18408
rect 19015 18377 19027 18380
rect 18969 18371 19027 18377
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 20993 18411 21051 18417
rect 20993 18377 21005 18411
rect 21039 18408 21051 18411
rect 21082 18408 21088 18420
rect 21039 18380 21088 18408
rect 21039 18377 21051 18380
rect 20993 18371 21051 18377
rect 21082 18368 21088 18380
rect 21140 18368 21146 18420
rect 21358 18408 21364 18420
rect 21319 18380 21364 18408
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 21726 18368 21732 18420
rect 21784 18408 21790 18420
rect 21821 18411 21879 18417
rect 21821 18408 21833 18411
rect 21784 18380 21833 18408
rect 21784 18368 21790 18380
rect 21821 18377 21833 18380
rect 21867 18377 21879 18411
rect 22278 18408 22284 18420
rect 22239 18380 22284 18408
rect 21821 18371 21879 18377
rect 22278 18368 22284 18380
rect 22336 18368 22342 18420
rect 23385 18411 23443 18417
rect 23385 18377 23397 18411
rect 23431 18408 23443 18411
rect 24210 18408 24216 18420
rect 23431 18380 24216 18408
rect 23431 18377 23443 18380
rect 23385 18371 23443 18377
rect 15933 18343 15991 18349
rect 15933 18309 15945 18343
rect 15979 18340 15991 18343
rect 16390 18340 16396 18352
rect 15979 18312 16396 18340
rect 15979 18309 15991 18312
rect 15933 18303 15991 18309
rect 16390 18300 16396 18312
rect 16448 18340 16454 18352
rect 18877 18343 18935 18349
rect 18877 18340 18889 18343
rect 16448 18312 18889 18340
rect 16448 18300 16454 18312
rect 18877 18309 18889 18312
rect 18923 18309 18935 18343
rect 18877 18303 18935 18309
rect 21266 18300 21272 18352
rect 21324 18340 21330 18352
rect 21637 18343 21695 18349
rect 21637 18340 21649 18343
rect 21324 18312 21649 18340
rect 21324 18300 21330 18312
rect 21637 18309 21649 18312
rect 21683 18340 21695 18343
rect 21683 18312 22094 18340
rect 21683 18309 21695 18312
rect 21637 18303 21695 18309
rect 6043 18244 6316 18272
rect 6365 18275 6423 18281
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 6365 18241 6377 18275
rect 6411 18241 6423 18275
rect 6621 18275 6679 18281
rect 6621 18272 6633 18275
rect 6365 18235 6423 18241
rect 6472 18244 6633 18272
rect 4396 18176 4660 18204
rect 4985 18207 5043 18213
rect 4396 18164 4402 18176
rect 4985 18173 4997 18207
rect 5031 18204 5043 18207
rect 5810 18204 5816 18216
rect 5031 18176 5816 18204
rect 5031 18173 5043 18176
rect 4985 18167 5043 18173
rect 5460 18148 5488 18176
rect 5810 18164 5816 18176
rect 5868 18164 5874 18216
rect 6181 18207 6239 18213
rect 6181 18173 6193 18207
rect 6227 18204 6239 18207
rect 6472 18204 6500 18244
rect 6621 18241 6633 18244
rect 6667 18241 6679 18275
rect 6621 18235 6679 18241
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 11606 18272 11612 18284
rect 11563 18244 11612 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 11606 18232 11612 18244
rect 11664 18232 11670 18284
rect 11700 18275 11758 18281
rect 11700 18241 11712 18275
rect 11746 18241 11758 18275
rect 11882 18272 11888 18284
rect 11843 18244 11888 18272
rect 11700 18235 11758 18241
rect 6227 18176 6500 18204
rect 6227 18173 6239 18176
rect 6181 18167 6239 18173
rect 10778 18164 10784 18216
rect 10836 18204 10842 18216
rect 11716 18204 11744 18235
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 12066 18272 12072 18284
rect 12027 18244 12072 18272
rect 12066 18232 12072 18244
rect 12124 18232 12130 18284
rect 13354 18272 13360 18284
rect 13315 18244 13360 18272
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 13446 18232 13452 18284
rect 13504 18272 13510 18284
rect 15104 18281 15162 18287
rect 13613 18275 13671 18281
rect 13613 18272 13625 18275
rect 13504 18244 13625 18272
rect 13504 18232 13510 18244
rect 13613 18241 13625 18244
rect 13659 18241 13671 18275
rect 13613 18235 13671 18241
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18241 14979 18275
rect 15104 18247 15116 18281
rect 15150 18247 15162 18281
rect 15104 18241 15162 18247
rect 15197 18275 15255 18281
rect 15197 18241 15209 18275
rect 15243 18272 15255 18275
rect 15473 18275 15531 18281
rect 15243 18244 15424 18272
rect 15243 18241 15255 18244
rect 14921 18235 14979 18241
rect 15197 18235 15255 18241
rect 10836 18176 11744 18204
rect 11793 18207 11851 18213
rect 10836 18164 10842 18176
rect 11793 18173 11805 18207
rect 11839 18173 11851 18207
rect 11793 18167 11851 18173
rect 3973 18139 4031 18145
rect 3344 18108 3832 18136
rect 3804 18080 3832 18108
rect 3973 18105 3985 18139
rect 4019 18136 4031 18139
rect 4522 18136 4528 18148
rect 4019 18108 4528 18136
rect 4019 18105 4031 18108
rect 3973 18099 4031 18105
rect 4522 18096 4528 18108
rect 4580 18096 4586 18148
rect 5442 18096 5448 18148
rect 5500 18096 5506 18148
rect 5534 18096 5540 18148
rect 5592 18136 5598 18148
rect 11808 18136 11836 18167
rect 12894 18136 12900 18148
rect 5592 18108 5948 18136
rect 5592 18096 5598 18108
rect 3786 18028 3792 18080
rect 3844 18068 3850 18080
rect 4065 18071 4123 18077
rect 4065 18068 4077 18071
rect 3844 18040 4077 18068
rect 3844 18028 3850 18040
rect 4065 18037 4077 18040
rect 4111 18037 4123 18071
rect 4065 18031 4123 18037
rect 5261 18071 5319 18077
rect 5261 18037 5273 18071
rect 5307 18068 5319 18071
rect 5810 18068 5816 18080
rect 5307 18040 5816 18068
rect 5307 18037 5319 18040
rect 5261 18031 5319 18037
rect 5810 18028 5816 18040
rect 5868 18028 5874 18080
rect 5920 18068 5948 18108
rect 7300 18108 8340 18136
rect 11808 18108 12900 18136
rect 7300 18068 7328 18108
rect 8312 18080 8340 18108
rect 12894 18096 12900 18108
rect 12952 18096 12958 18148
rect 7742 18068 7748 18080
rect 5920 18040 7328 18068
rect 7703 18040 7748 18068
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 8294 18068 8300 18080
rect 8255 18040 8300 18068
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 12158 18068 12164 18080
rect 12119 18040 12164 18068
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 13078 18028 13084 18080
rect 13136 18068 13142 18080
rect 14936 18068 14964 18235
rect 15286 18204 15292 18216
rect 15247 18176 15292 18204
rect 15286 18164 15292 18176
rect 15344 18164 15350 18216
rect 15396 18204 15424 18244
rect 15473 18241 15485 18275
rect 15519 18272 15531 18275
rect 16574 18272 16580 18284
rect 15519 18244 16580 18272
rect 15519 18241 15531 18244
rect 15473 18235 15531 18241
rect 16574 18232 16580 18244
rect 16632 18232 16638 18284
rect 16761 18275 16819 18281
rect 16761 18241 16773 18275
rect 16807 18272 16819 18275
rect 16942 18272 16948 18284
rect 16807 18244 16948 18272
rect 16807 18241 16819 18244
rect 16761 18235 16819 18241
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 17310 18272 17316 18284
rect 17271 18244 17316 18272
rect 17310 18232 17316 18244
rect 17368 18232 17374 18284
rect 17773 18275 17831 18281
rect 17773 18241 17785 18275
rect 17819 18272 17831 18275
rect 18046 18272 18052 18284
rect 17819 18244 18052 18272
rect 17819 18241 17831 18244
rect 17773 18235 17831 18241
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 18196 18244 18245 18272
rect 18196 18232 18202 18244
rect 18233 18241 18245 18244
rect 18279 18241 18291 18275
rect 18414 18272 18420 18284
rect 18375 18244 18420 18272
rect 18233 18235 18291 18241
rect 18414 18232 18420 18244
rect 18472 18232 18478 18284
rect 20622 18232 20628 18284
rect 20680 18272 20686 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20680 18244 20821 18272
rect 20680 18232 20686 18244
rect 20809 18241 20821 18244
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 21177 18275 21235 18281
rect 21177 18272 21189 18275
rect 20956 18244 21189 18272
rect 20956 18232 20962 18244
rect 21177 18241 21189 18244
rect 21223 18241 21235 18275
rect 21177 18235 21235 18241
rect 16390 18204 16396 18216
rect 15396 18176 16396 18204
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 17221 18207 17279 18213
rect 17221 18173 17233 18207
rect 17267 18204 17279 18207
rect 17494 18204 17500 18216
rect 17267 18176 17500 18204
rect 17267 18173 17279 18176
rect 17221 18167 17279 18173
rect 17494 18164 17500 18176
rect 17552 18204 17558 18216
rect 17865 18207 17923 18213
rect 17865 18204 17877 18207
rect 17552 18176 17877 18204
rect 17552 18164 17558 18176
rect 17865 18173 17877 18176
rect 17911 18173 17923 18207
rect 17865 18167 17923 18173
rect 17957 18207 18015 18213
rect 17957 18173 17969 18207
rect 18003 18173 18015 18207
rect 22066 18204 22094 18312
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18272 22247 18275
rect 22554 18272 22560 18284
rect 22235 18244 22560 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 22465 18207 22523 18213
rect 22465 18204 22477 18207
rect 22066 18176 22477 18204
rect 17957 18167 18015 18173
rect 22465 18173 22477 18176
rect 22511 18204 22523 18207
rect 23400 18204 23428 18371
rect 24210 18368 24216 18380
rect 24268 18368 24274 18420
rect 25314 18368 25320 18420
rect 25372 18408 25378 18420
rect 25409 18411 25467 18417
rect 25409 18408 25421 18411
rect 25372 18380 25421 18408
rect 25372 18368 25378 18380
rect 25409 18377 25421 18380
rect 25455 18377 25467 18411
rect 25409 18371 25467 18377
rect 24296 18343 24354 18349
rect 24296 18309 24308 18343
rect 24342 18340 24354 18343
rect 24578 18340 24584 18352
rect 24342 18312 24584 18340
rect 24342 18309 24354 18312
rect 24296 18303 24354 18309
rect 24578 18300 24584 18312
rect 24636 18300 24642 18352
rect 24026 18204 24032 18216
rect 22511 18176 23428 18204
rect 23939 18176 24032 18204
rect 22511 18173 22523 18176
rect 22465 18167 22523 18173
rect 15102 18096 15108 18148
rect 15160 18136 15166 18148
rect 15749 18139 15807 18145
rect 15749 18136 15761 18139
rect 15160 18108 15761 18136
rect 15160 18096 15166 18108
rect 15749 18105 15761 18108
rect 15795 18105 15807 18139
rect 17402 18136 17408 18148
rect 17363 18108 17408 18136
rect 15749 18099 15807 18105
rect 17402 18096 17408 18108
rect 17460 18096 17466 18148
rect 17972 18136 18000 18167
rect 24026 18164 24032 18176
rect 24084 18164 24090 18216
rect 19153 18139 19211 18145
rect 19153 18136 19165 18139
rect 17972 18108 19165 18136
rect 13136 18040 14964 18068
rect 13136 18028 13142 18040
rect 16942 18028 16948 18080
rect 17000 18068 17006 18080
rect 17972 18068 18000 18108
rect 19153 18105 19165 18108
rect 19199 18136 19211 18139
rect 19242 18136 19248 18148
rect 19199 18108 19248 18136
rect 19199 18105 19211 18108
rect 19153 18099 19211 18105
rect 19242 18096 19248 18108
rect 19300 18096 19306 18148
rect 20806 18096 20812 18148
rect 20864 18136 20870 18148
rect 24044 18136 24072 18164
rect 20864 18108 24072 18136
rect 20864 18096 20870 18108
rect 17000 18040 18000 18068
rect 18601 18071 18659 18077
rect 17000 18028 17006 18040
rect 18601 18037 18613 18071
rect 18647 18068 18659 18071
rect 19058 18068 19064 18080
rect 18647 18040 19064 18068
rect 18647 18037 18659 18040
rect 18601 18031 18659 18037
rect 19058 18028 19064 18040
rect 19116 18028 19122 18080
rect 1104 17978 26128 18000
rect 1104 17926 5120 17978
rect 5172 17926 5184 17978
rect 5236 17926 5248 17978
rect 5300 17926 5312 17978
rect 5364 17926 5376 17978
rect 5428 17926 13462 17978
rect 13514 17926 13526 17978
rect 13578 17926 13590 17978
rect 13642 17926 13654 17978
rect 13706 17926 13718 17978
rect 13770 17926 21803 17978
rect 21855 17926 21867 17978
rect 21919 17926 21931 17978
rect 21983 17926 21995 17978
rect 22047 17926 22059 17978
rect 22111 17926 26128 17978
rect 1104 17904 26128 17926
rect 5353 17867 5411 17873
rect 5353 17833 5365 17867
rect 5399 17864 5411 17867
rect 5442 17864 5448 17876
rect 5399 17836 5448 17864
rect 5399 17833 5411 17836
rect 5353 17827 5411 17833
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 12526 17864 12532 17876
rect 5552 17836 12532 17864
rect 4062 17756 4068 17808
rect 4120 17796 4126 17808
rect 5552 17796 5580 17836
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12894 17864 12900 17876
rect 12855 17836 12900 17864
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 13354 17824 13360 17876
rect 13412 17864 13418 17876
rect 13725 17867 13783 17873
rect 13725 17864 13737 17867
rect 13412 17836 13737 17864
rect 13412 17824 13418 17836
rect 13725 17833 13737 17836
rect 13771 17833 13783 17867
rect 15930 17864 15936 17876
rect 13725 17827 13783 17833
rect 14384 17836 15936 17864
rect 10502 17796 10508 17808
rect 4120 17768 5580 17796
rect 10463 17768 10508 17796
rect 4120 17756 4126 17768
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 11330 17796 11336 17808
rect 10612 17768 11336 17796
rect 3786 17688 3792 17740
rect 3844 17728 3850 17740
rect 4617 17731 4675 17737
rect 4617 17728 4629 17731
rect 3844 17700 4629 17728
rect 3844 17688 3850 17700
rect 4617 17697 4629 17700
rect 4663 17697 4675 17731
rect 4617 17691 4675 17697
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17728 4767 17731
rect 5442 17728 5448 17740
rect 4755 17700 5448 17728
rect 4755 17697 4767 17700
rect 4709 17691 4767 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 2038 17660 2044 17672
rect 1999 17632 2044 17660
rect 2038 17620 2044 17632
rect 2096 17620 2102 17672
rect 4341 17663 4399 17669
rect 4341 17629 4353 17663
rect 4387 17629 4399 17663
rect 4341 17623 4399 17629
rect 4524 17663 4582 17669
rect 4524 17629 4536 17663
rect 4570 17660 4582 17663
rect 4893 17663 4951 17669
rect 4570 17632 4660 17660
rect 4570 17629 4582 17632
rect 4524 17623 4582 17629
rect 2308 17595 2366 17601
rect 2308 17561 2320 17595
rect 2354 17592 2366 17595
rect 2774 17592 2780 17604
rect 2354 17564 2780 17592
rect 2354 17561 2366 17564
rect 2308 17555 2366 17561
rect 2774 17552 2780 17564
rect 2832 17552 2838 17604
rect 2958 17552 2964 17604
rect 3016 17592 3022 17604
rect 3973 17595 4031 17601
rect 3973 17592 3985 17595
rect 3016 17564 3985 17592
rect 3016 17552 3022 17564
rect 3973 17561 3985 17564
rect 4019 17561 4031 17595
rect 4154 17592 4160 17604
rect 4115 17564 4160 17592
rect 3973 17555 4031 17561
rect 4154 17552 4160 17564
rect 4212 17552 4218 17604
rect 4356 17592 4384 17623
rect 4632 17604 4660 17632
rect 4893 17629 4905 17663
rect 4939 17629 4951 17663
rect 5534 17660 5540 17672
rect 5495 17632 5540 17660
rect 4893 17623 4951 17629
rect 4356 17564 4568 17592
rect 4540 17536 4568 17564
rect 4614 17552 4620 17604
rect 4672 17552 4678 17604
rect 4908 17592 4936 17623
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 5626 17620 5632 17672
rect 5684 17660 5690 17672
rect 5721 17663 5779 17669
rect 5721 17660 5733 17663
rect 5684 17632 5733 17660
rect 5684 17620 5690 17632
rect 5721 17629 5733 17632
rect 5767 17629 5779 17663
rect 5721 17623 5779 17629
rect 5810 17620 5816 17672
rect 5868 17660 5874 17672
rect 5977 17663 6035 17669
rect 5977 17660 5989 17663
rect 5868 17632 5989 17660
rect 5868 17620 5874 17632
rect 5977 17629 5989 17632
rect 6023 17629 6035 17663
rect 5977 17623 6035 17629
rect 7834 17620 7840 17672
rect 7892 17660 7898 17672
rect 8941 17663 8999 17669
rect 8941 17660 8953 17663
rect 7892 17632 8953 17660
rect 7892 17620 7898 17632
rect 8941 17629 8953 17632
rect 8987 17629 8999 17663
rect 10612 17660 10640 17768
rect 11330 17756 11336 17768
rect 11388 17756 11394 17808
rect 13170 17756 13176 17808
rect 13228 17796 13234 17808
rect 13228 17768 13492 17796
rect 13228 17756 13234 17768
rect 10962 17688 10968 17740
rect 11020 17728 11026 17740
rect 11020 17700 11065 17728
rect 11020 17688 11026 17700
rect 12710 17688 12716 17740
rect 12768 17728 12774 17740
rect 13464 17737 13492 17768
rect 13357 17731 13415 17737
rect 13357 17728 13369 17731
rect 12768 17700 13369 17728
rect 12768 17688 12774 17700
rect 13357 17697 13369 17700
rect 13403 17697 13415 17731
rect 13357 17691 13415 17697
rect 13449 17731 13507 17737
rect 13449 17697 13461 17731
rect 13495 17697 13507 17731
rect 14384 17728 14412 17836
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 16761 17867 16819 17873
rect 16761 17833 16773 17867
rect 16807 17864 16819 17867
rect 16850 17864 16856 17876
rect 16807 17836 16856 17864
rect 16807 17833 16819 17836
rect 16761 17827 16819 17833
rect 16850 17824 16856 17836
rect 16908 17824 16914 17876
rect 18046 17864 18052 17876
rect 18007 17836 18052 17864
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 18598 17824 18604 17876
rect 18656 17864 18662 17876
rect 19245 17867 19303 17873
rect 19245 17864 19257 17867
rect 18656 17836 19257 17864
rect 18656 17824 18662 17836
rect 19245 17833 19257 17836
rect 19291 17833 19303 17867
rect 19245 17827 19303 17833
rect 14458 17756 14464 17808
rect 14516 17796 14522 17808
rect 14516 17768 14688 17796
rect 14516 17756 14522 17768
rect 14660 17737 14688 17768
rect 17126 17756 17132 17808
rect 17184 17796 17190 17808
rect 17184 17768 18644 17796
rect 17184 17756 17190 17768
rect 14645 17731 14703 17737
rect 14384 17700 14504 17728
rect 13449 17691 13507 17697
rect 8941 17623 8999 17629
rect 9048 17632 10640 17660
rect 6086 17592 6092 17604
rect 4908 17564 6092 17592
rect 6086 17552 6092 17564
rect 6144 17552 6150 17604
rect 6822 17552 6828 17604
rect 6880 17592 6886 17604
rect 9048 17592 9076 17632
rect 10686 17620 10692 17672
rect 10744 17660 10750 17672
rect 10873 17663 10931 17669
rect 11241 17663 11299 17669
rect 10744 17632 10789 17660
rect 10744 17620 10750 17632
rect 10873 17629 10885 17663
rect 10919 17629 10931 17663
rect 10873 17623 10931 17629
rect 11058 17657 11116 17663
rect 11058 17623 11070 17657
rect 11104 17623 11116 17657
rect 11241 17629 11253 17663
rect 11287 17629 11299 17663
rect 11514 17660 11520 17672
rect 11475 17632 11520 17660
rect 11241 17623 11299 17629
rect 6880 17564 9076 17592
rect 9208 17595 9266 17601
rect 6880 17552 6886 17564
rect 9208 17561 9220 17595
rect 9254 17592 9266 17595
rect 9858 17592 9864 17604
rect 9254 17564 9864 17592
rect 9254 17561 9266 17564
rect 9208 17555 9266 17561
rect 9858 17552 9864 17564
rect 9916 17552 9922 17604
rect 10502 17552 10508 17604
rect 10560 17592 10566 17604
rect 10888 17592 10916 17623
rect 11058 17617 11116 17623
rect 10560 17564 10916 17592
rect 10560 17552 10566 17564
rect 3421 17527 3479 17533
rect 3421 17493 3433 17527
rect 3467 17524 3479 17527
rect 3878 17524 3884 17536
rect 3467 17496 3884 17524
rect 3467 17493 3479 17496
rect 3421 17487 3479 17493
rect 3878 17484 3884 17496
rect 3936 17484 3942 17536
rect 4522 17484 4528 17536
rect 4580 17484 4586 17536
rect 4890 17484 4896 17536
rect 4948 17524 4954 17536
rect 4985 17527 5043 17533
rect 4985 17524 4997 17527
rect 4948 17496 4997 17524
rect 4948 17484 4954 17496
rect 4985 17493 4997 17496
rect 5031 17493 5043 17527
rect 7098 17524 7104 17536
rect 7059 17496 7104 17524
rect 4985 17487 5043 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 10226 17484 10232 17536
rect 10284 17524 10290 17536
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 10284 17496 10333 17524
rect 10284 17484 10290 17496
rect 10321 17493 10333 17496
rect 10367 17524 10379 17527
rect 11072 17524 11100 17617
rect 11256 17592 11284 17623
rect 11514 17620 11520 17632
rect 11572 17620 11578 17672
rect 11784 17663 11842 17669
rect 11784 17629 11796 17663
rect 11830 17660 11842 17663
rect 12158 17660 12164 17672
rect 11830 17632 12164 17660
rect 11830 17629 11842 17632
rect 11784 17623 11842 17629
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 12618 17660 12624 17672
rect 12406 17632 12624 17660
rect 12406 17592 12434 17632
rect 12618 17620 12624 17632
rect 12676 17660 12682 17672
rect 13078 17660 13084 17672
rect 12676 17632 13084 17660
rect 12676 17620 12682 17632
rect 13078 17620 13084 17632
rect 13136 17620 13142 17672
rect 13262 17660 13268 17672
rect 13223 17632 13268 17660
rect 13262 17620 13268 17632
rect 13320 17620 13326 17672
rect 13633 17663 13691 17669
rect 13633 17629 13645 17663
rect 13679 17660 13691 17663
rect 13814 17660 13820 17672
rect 13679 17632 13820 17660
rect 13679 17629 13691 17632
rect 13633 17623 13691 17629
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 14369 17663 14427 17669
rect 14369 17629 14381 17663
rect 14415 17629 14427 17663
rect 14476 17660 14504 17700
rect 14645 17697 14657 17731
rect 14691 17697 14703 17731
rect 15105 17731 15163 17737
rect 14645 17691 14703 17697
rect 14844 17700 15056 17728
rect 14534 17663 14592 17669
rect 14534 17660 14546 17663
rect 14476 17632 14546 17660
rect 14369 17623 14427 17629
rect 14534 17629 14546 17632
rect 14580 17629 14592 17663
rect 14734 17660 14740 17672
rect 14695 17632 14740 17660
rect 14534 17623 14592 17629
rect 14384 17592 14412 17623
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 14844 17592 14872 17700
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17629 14979 17663
rect 15028 17660 15056 17700
rect 15105 17697 15117 17731
rect 15151 17728 15163 17731
rect 15151 17700 15332 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 15197 17663 15255 17669
rect 15197 17660 15209 17663
rect 15028 17632 15209 17660
rect 14921 17623 14979 17629
rect 11256 17564 12434 17592
rect 13096 17564 14412 17592
rect 14568 17564 14872 17592
rect 10367 17496 11100 17524
rect 10367 17493 10379 17496
rect 10321 17487 10379 17493
rect 11606 17484 11612 17536
rect 11664 17524 11670 17536
rect 13096 17524 13124 17564
rect 14568 17536 14596 17564
rect 11664 17496 13124 17524
rect 11664 17484 11670 17496
rect 14550 17484 14556 17536
rect 14608 17484 14614 17536
rect 14936 17524 14964 17623
rect 15120 17604 15148 17632
rect 15197 17629 15209 17632
rect 15243 17629 15255 17663
rect 15304 17660 15332 17700
rect 16942 17688 16948 17740
rect 17000 17728 17006 17740
rect 18616 17737 18644 17768
rect 17313 17731 17371 17737
rect 17313 17728 17325 17731
rect 17000 17700 17325 17728
rect 17000 17688 17006 17700
rect 17313 17697 17325 17700
rect 17359 17697 17371 17731
rect 17313 17691 17371 17697
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17697 18659 17731
rect 18601 17691 18659 17697
rect 19242 17688 19248 17740
rect 19300 17728 19306 17740
rect 19797 17731 19855 17737
rect 19797 17728 19809 17731
rect 19300 17700 19809 17728
rect 19300 17688 19306 17700
rect 19797 17697 19809 17700
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 15453 17663 15511 17669
rect 15453 17660 15465 17663
rect 15304 17632 15465 17660
rect 15197 17623 15255 17629
rect 15453 17629 15465 17632
rect 15499 17629 15511 17663
rect 15453 17623 15511 17629
rect 17129 17663 17187 17669
rect 17129 17629 17141 17663
rect 17175 17660 17187 17663
rect 17218 17660 17224 17672
rect 17175 17632 17224 17660
rect 17175 17629 17187 17632
rect 17129 17623 17187 17629
rect 17218 17620 17224 17632
rect 17276 17620 17282 17672
rect 17589 17663 17647 17669
rect 17589 17629 17601 17663
rect 17635 17629 17647 17663
rect 17589 17623 17647 17629
rect 17865 17663 17923 17669
rect 17865 17629 17877 17663
rect 17911 17660 17923 17663
rect 17954 17660 17960 17672
rect 17911 17632 17960 17660
rect 17911 17629 17923 17632
rect 17865 17623 17923 17629
rect 15102 17552 15108 17604
rect 15160 17552 15166 17604
rect 17604 17592 17632 17623
rect 17954 17620 17960 17632
rect 18012 17620 18018 17672
rect 19058 17660 19064 17672
rect 19019 17632 19064 17660
rect 19058 17620 19064 17632
rect 19116 17620 19122 17672
rect 19150 17620 19156 17672
rect 19208 17660 19214 17672
rect 23382 17660 23388 17672
rect 19208 17632 23388 17660
rect 19208 17620 19214 17632
rect 23382 17620 23388 17632
rect 23440 17620 23446 17672
rect 19705 17595 19763 17601
rect 19705 17592 19717 17595
rect 17144 17564 17632 17592
rect 18432 17564 19717 17592
rect 17144 17536 17172 17564
rect 18432 17536 18460 17564
rect 19705 17561 19717 17564
rect 19751 17561 19763 17595
rect 19705 17555 19763 17561
rect 16577 17527 16635 17533
rect 16577 17524 16589 17527
rect 14936 17496 16589 17524
rect 16577 17493 16589 17496
rect 16623 17524 16635 17527
rect 17126 17524 17132 17536
rect 16623 17496 17132 17524
rect 16623 17493 16635 17496
rect 16577 17487 16635 17493
rect 17126 17484 17132 17496
rect 17184 17484 17190 17536
rect 17221 17527 17279 17533
rect 17221 17493 17233 17527
rect 17267 17524 17279 17527
rect 17310 17524 17316 17536
rect 17267 17496 17316 17524
rect 17267 17493 17279 17496
rect 17221 17487 17279 17493
rect 17310 17484 17316 17496
rect 17368 17524 17374 17536
rect 17681 17527 17739 17533
rect 17681 17524 17693 17527
rect 17368 17496 17693 17524
rect 17368 17484 17374 17496
rect 17681 17493 17693 17496
rect 17727 17493 17739 17527
rect 18414 17524 18420 17536
rect 18375 17496 18420 17524
rect 17681 17487 17739 17493
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17524 18567 17527
rect 18877 17527 18935 17533
rect 18877 17524 18889 17527
rect 18555 17496 18889 17524
rect 18555 17493 18567 17496
rect 18509 17487 18567 17493
rect 18877 17493 18889 17496
rect 18923 17493 18935 17527
rect 19610 17524 19616 17536
rect 19571 17496 19616 17524
rect 18877 17487 18935 17493
rect 19610 17484 19616 17496
rect 19668 17484 19674 17536
rect 1104 17434 26128 17456
rect 1104 17382 9291 17434
rect 9343 17382 9355 17434
rect 9407 17382 9419 17434
rect 9471 17382 9483 17434
rect 9535 17382 9547 17434
rect 9599 17382 17632 17434
rect 17684 17382 17696 17434
rect 17748 17382 17760 17434
rect 17812 17382 17824 17434
rect 17876 17382 17888 17434
rect 17940 17382 26128 17434
rect 1104 17360 26128 17382
rect 3237 17323 3295 17329
rect 3237 17289 3249 17323
rect 3283 17320 3295 17323
rect 3970 17320 3976 17332
rect 3283 17292 3976 17320
rect 3283 17289 3295 17292
rect 3237 17283 3295 17289
rect 3970 17280 3976 17292
rect 4028 17280 4034 17332
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 4212 17292 6561 17320
rect 4212 17280 4218 17292
rect 6549 17289 6561 17292
rect 6595 17320 6607 17323
rect 6595 17292 8432 17320
rect 6595 17289 6607 17292
rect 6549 17283 6607 17289
rect 2038 17252 2044 17264
rect 1872 17224 2044 17252
rect 1872 17193 1900 17224
rect 2038 17212 2044 17224
rect 2096 17252 2102 17264
rect 2096 17224 3004 17252
rect 2096 17212 2102 17224
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17153 1915 17187
rect 1857 17147 1915 17153
rect 2124 17187 2182 17193
rect 2124 17153 2136 17187
rect 2170 17184 2182 17187
rect 2170 17156 2912 17184
rect 2170 17153 2182 17156
rect 2124 17147 2182 17153
rect 2884 17048 2912 17156
rect 2976 17128 3004 17224
rect 4062 17212 4068 17264
rect 4120 17252 4126 17264
rect 8404 17261 8432 17292
rect 9030 17280 9036 17332
rect 9088 17320 9094 17332
rect 9674 17320 9680 17332
rect 9088 17292 9680 17320
rect 9088 17280 9094 17292
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 9858 17320 9864 17332
rect 9819 17292 9864 17320
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 12897 17323 12955 17329
rect 12897 17320 12909 17323
rect 10888 17292 12909 17320
rect 8389 17255 8447 17261
rect 4120 17224 5488 17252
rect 4120 17212 4126 17224
rect 5460 17193 5488 17224
rect 5920 17224 8340 17252
rect 3780 17187 3838 17193
rect 3780 17153 3792 17187
rect 3826 17184 3838 17187
rect 5077 17187 5135 17193
rect 5077 17184 5089 17187
rect 3826 17156 5089 17184
rect 3826 17153 3838 17156
rect 3780 17147 3838 17153
rect 5077 17153 5089 17156
rect 5123 17153 5135 17187
rect 5077 17147 5135 17153
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17153 5319 17187
rect 5261 17147 5319 17153
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17153 5503 17187
rect 5445 17147 5503 17153
rect 5665 17190 5724 17196
rect 5665 17156 5677 17190
rect 5711 17156 5724 17190
rect 5665 17150 5724 17156
rect 2958 17076 2964 17128
rect 3016 17116 3022 17128
rect 3513 17119 3571 17125
rect 3513 17116 3525 17119
rect 3016 17088 3525 17116
rect 3016 17076 3022 17088
rect 3513 17085 3525 17088
rect 3559 17085 3571 17119
rect 5276 17116 5304 17147
rect 5718 17144 5724 17150
rect 5776 17144 5782 17196
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 5920 17184 5948 17224
rect 5859 17156 5948 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 3513 17079 3571 17085
rect 4908 17088 5304 17116
rect 5537 17119 5595 17125
rect 3418 17048 3424 17060
rect 2884 17020 3424 17048
rect 3418 17008 3424 17020
rect 3476 17008 3482 17060
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 4908 16989 4936 17088
rect 5537 17085 5549 17119
rect 5583 17085 5595 17119
rect 5537 17079 5595 17085
rect 4893 16983 4951 16989
rect 4893 16980 4905 16983
rect 4764 16952 4905 16980
rect 4764 16940 4770 16952
rect 4893 16949 4905 16952
rect 4939 16949 4951 16983
rect 5552 16980 5580 17079
rect 5920 17057 5948 17156
rect 6089 17187 6147 17193
rect 6089 17153 6101 17187
rect 6135 17153 6147 17187
rect 6089 17147 6147 17153
rect 6641 17187 6699 17193
rect 6641 17153 6653 17187
rect 6687 17184 6699 17187
rect 8312 17184 8340 17224
rect 8389 17221 8401 17255
rect 8435 17221 8447 17255
rect 8389 17215 8447 17221
rect 8680 17224 10548 17252
rect 8680 17184 8708 17224
rect 8846 17184 8852 17196
rect 6687 17156 7144 17184
rect 8312 17156 8708 17184
rect 8807 17156 8852 17184
rect 6687 17153 6699 17156
rect 6641 17147 6699 17153
rect 6104 17116 6132 17147
rect 6822 17116 6828 17128
rect 6104 17088 6828 17116
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 5905 17051 5963 17057
rect 5905 17017 5917 17051
rect 5951 17017 5963 17051
rect 5905 17011 5963 17017
rect 6270 16980 6276 16992
rect 5552 16952 6276 16980
rect 4893 16943 4951 16949
rect 6270 16940 6276 16952
rect 6328 16940 6334 16992
rect 7116 16989 7144 17156
rect 8846 17144 8852 17156
rect 8904 17144 8910 17196
rect 9030 17184 9036 17196
rect 8991 17156 9036 17184
rect 9030 17144 9036 17156
rect 9088 17144 9094 17196
rect 9218 17187 9276 17193
rect 9218 17153 9230 17187
rect 9264 17184 9276 17187
rect 9306 17184 9312 17196
rect 9264 17156 9312 17184
rect 9264 17153 9276 17156
rect 9218 17147 9276 17153
rect 9306 17144 9312 17156
rect 9364 17144 9370 17196
rect 9416 17193 9444 17224
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17153 9459 17187
rect 9401 17147 9459 17153
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 9950 17184 9956 17196
rect 9732 17156 9956 17184
rect 9732 17144 9738 17156
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 10042 17144 10048 17196
rect 10100 17193 10106 17196
rect 10100 17187 10149 17193
rect 10100 17153 10103 17187
rect 10137 17153 10149 17187
rect 10226 17184 10232 17196
rect 10187 17156 10232 17184
rect 10100 17147 10149 17153
rect 10100 17144 10106 17147
rect 10226 17144 10232 17156
rect 10284 17144 10290 17196
rect 10520 17193 10548 17224
rect 10339 17187 10397 17193
rect 10339 17153 10351 17187
rect 10385 17184 10397 17187
rect 10505 17187 10563 17193
rect 10385 17156 10456 17184
rect 10385 17153 10397 17156
rect 10339 17147 10397 17153
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 9048 17116 9076 17144
rect 8251 17088 9076 17116
rect 9125 17119 9183 17125
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 9125 17085 9137 17119
rect 9171 17116 9183 17119
rect 10428 17116 10456 17156
rect 10505 17153 10517 17187
rect 10551 17184 10563 17187
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10551 17156 10609 17184
rect 10551 17153 10563 17156
rect 10505 17147 10563 17153
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10778 17184 10784 17196
rect 10597 17147 10655 17153
rect 10704 17156 10784 17184
rect 10704 17116 10732 17156
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 10888 17193 10916 17292
rect 12897 17289 12909 17292
rect 12943 17320 12955 17323
rect 13262 17320 13268 17332
rect 12943 17292 13268 17320
rect 12943 17289 12955 17292
rect 12897 17283 12955 17289
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 15289 17323 15347 17329
rect 15289 17289 15301 17323
rect 15335 17320 15347 17323
rect 15930 17320 15936 17332
rect 15335 17292 15936 17320
rect 15335 17289 15347 17292
rect 15289 17283 15347 17289
rect 15930 17280 15936 17292
rect 15988 17280 15994 17332
rect 18046 17320 18052 17332
rect 17959 17292 18052 17320
rect 18046 17280 18052 17292
rect 18104 17320 18110 17332
rect 19150 17320 19156 17332
rect 18104 17292 19156 17320
rect 18104 17280 18110 17292
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 19610 17280 19616 17332
rect 19668 17320 19674 17332
rect 19981 17323 20039 17329
rect 19981 17320 19993 17323
rect 19668 17292 19993 17320
rect 19668 17280 19674 17292
rect 19981 17289 19993 17292
rect 20027 17289 20039 17323
rect 19981 17283 20039 17289
rect 20257 17323 20315 17329
rect 20257 17289 20269 17323
rect 20303 17320 20315 17323
rect 20898 17320 20904 17332
rect 20303 17292 20904 17320
rect 20303 17289 20315 17292
rect 20257 17283 20315 17289
rect 20898 17280 20904 17292
rect 20956 17280 20962 17332
rect 11333 17255 11391 17261
rect 11333 17221 11345 17255
rect 11379 17252 11391 17255
rect 11762 17255 11820 17261
rect 11762 17252 11774 17255
rect 11379 17224 11774 17252
rect 11379 17221 11391 17224
rect 11333 17215 11391 17221
rect 11762 17221 11774 17224
rect 11808 17221 11820 17255
rect 11762 17215 11820 17221
rect 12526 17212 12532 17264
rect 12584 17252 12590 17264
rect 13998 17252 14004 17264
rect 12584 17224 14004 17252
rect 12584 17212 12590 17224
rect 13998 17212 14004 17224
rect 14056 17212 14062 17264
rect 18230 17252 18236 17264
rect 18191 17224 18236 17252
rect 18230 17212 18236 17224
rect 18288 17212 18294 17264
rect 19426 17212 19432 17264
rect 19484 17252 19490 17264
rect 21085 17255 21143 17261
rect 21085 17252 21097 17255
rect 19484 17224 21097 17252
rect 19484 17212 19490 17224
rect 21085 17221 21097 17224
rect 21131 17252 21143 17255
rect 21542 17252 21548 17264
rect 21131 17224 21548 17252
rect 21131 17221 21143 17224
rect 21085 17215 21143 17221
rect 21542 17212 21548 17224
rect 21600 17252 21606 17264
rect 23937 17255 23995 17261
rect 23937 17252 23949 17255
rect 21600 17224 23949 17252
rect 21600 17212 21606 17224
rect 23937 17221 23949 17224
rect 23983 17221 23995 17255
rect 23937 17215 23995 17221
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 11238 17184 11244 17196
rect 11195 17156 11244 17184
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 16758 17144 16764 17196
rect 16816 17184 16822 17196
rect 16925 17187 16983 17193
rect 16925 17184 16937 17187
rect 16816 17156 16937 17184
rect 16816 17144 16822 17156
rect 16925 17153 16937 17156
rect 16971 17153 16983 17187
rect 16925 17147 16983 17153
rect 17402 17144 17408 17196
rect 17460 17184 17466 17196
rect 18325 17187 18383 17193
rect 18325 17184 18337 17187
rect 17460 17156 18337 17184
rect 17460 17144 17466 17156
rect 18325 17153 18337 17156
rect 18371 17153 18383 17187
rect 18506 17184 18512 17196
rect 18467 17156 18512 17184
rect 18325 17147 18383 17153
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 18877 17187 18935 17193
rect 18877 17153 18889 17187
rect 18923 17184 18935 17187
rect 19613 17187 19671 17193
rect 19613 17184 19625 17187
rect 18923 17156 19625 17184
rect 18923 17153 18935 17156
rect 18877 17147 18935 17153
rect 19613 17153 19625 17156
rect 19659 17184 19671 17187
rect 19702 17184 19708 17196
rect 19659 17156 19708 17184
rect 19659 17153 19671 17156
rect 19613 17147 19671 17153
rect 19702 17144 19708 17156
rect 19760 17144 19766 17196
rect 19794 17144 19800 17196
rect 19852 17184 19858 17196
rect 20073 17187 20131 17193
rect 20073 17184 20085 17187
rect 19852 17156 20085 17184
rect 19852 17144 19858 17156
rect 20073 17153 20085 17156
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17184 20775 17187
rect 22186 17184 22192 17196
rect 20763 17156 22192 17184
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 24210 17184 24216 17196
rect 24171 17156 24216 17184
rect 24210 17144 24216 17156
rect 24268 17144 24274 17196
rect 10962 17116 10968 17128
rect 9171 17088 10732 17116
rect 10923 17088 10968 17116
rect 9171 17085 9183 17088
rect 9125 17079 9183 17085
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 11514 17116 11520 17128
rect 11427 17088 11520 17116
rect 11514 17076 11520 17088
rect 11572 17076 11578 17128
rect 16666 17116 16672 17128
rect 16627 17088 16672 17116
rect 16666 17076 16672 17088
rect 16724 17076 16730 17128
rect 18138 17076 18144 17128
rect 18196 17116 18202 17128
rect 18693 17119 18751 17125
rect 18693 17116 18705 17119
rect 18196 17088 18705 17116
rect 18196 17076 18202 17088
rect 18693 17085 18705 17088
rect 18739 17085 18751 17119
rect 19426 17116 19432 17128
rect 19387 17088 19432 17116
rect 18693 17079 18751 17085
rect 7834 17008 7840 17060
rect 7892 17048 7898 17060
rect 8573 17051 8631 17057
rect 8573 17048 8585 17051
rect 7892 17020 8585 17048
rect 7892 17008 7898 17020
rect 8573 17017 8585 17020
rect 8619 17048 8631 17051
rect 11532 17048 11560 17076
rect 8619 17020 11560 17048
rect 18708 17048 18736 17079
rect 19426 17076 19432 17088
rect 19484 17076 19490 17128
rect 19518 17076 19524 17128
rect 19576 17116 19582 17128
rect 20533 17119 20591 17125
rect 19576 17088 19621 17116
rect 19576 17076 19582 17088
rect 20533 17085 20545 17119
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 20548 17048 20576 17079
rect 18708 17020 20576 17048
rect 24397 17051 24455 17057
rect 8619 17017 8631 17020
rect 8573 17011 8631 17017
rect 24397 17017 24409 17051
rect 24443 17048 24455 17051
rect 25406 17048 25412 17060
rect 24443 17020 25412 17048
rect 24443 17017 24455 17020
rect 24397 17011 24455 17017
rect 25406 17008 25412 17020
rect 25464 17008 25470 17060
rect 7101 16983 7159 16989
rect 7101 16949 7113 16983
rect 7147 16980 7159 16983
rect 7558 16980 7564 16992
rect 7147 16952 7564 16980
rect 7147 16949 7159 16952
rect 7101 16943 7159 16949
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 8757 16983 8815 16989
rect 8757 16949 8769 16983
rect 8803 16980 8815 16983
rect 9030 16980 9036 16992
rect 8803 16952 9036 16980
rect 8803 16949 8815 16952
rect 8757 16943 8815 16949
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 10042 16940 10048 16992
rect 10100 16980 10106 16992
rect 14274 16980 14280 16992
rect 10100 16952 14280 16980
rect 10100 16940 10106 16952
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 19061 16983 19119 16989
rect 19061 16949 19073 16983
rect 19107 16980 19119 16983
rect 19794 16980 19800 16992
rect 19107 16952 19800 16980
rect 19107 16949 19119 16952
rect 19061 16943 19119 16949
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 20714 16940 20720 16992
rect 20772 16980 20778 16992
rect 20901 16983 20959 16989
rect 20901 16980 20913 16983
rect 20772 16952 20913 16980
rect 20772 16940 20778 16952
rect 20901 16949 20913 16952
rect 20947 16949 20959 16983
rect 20901 16943 20959 16949
rect 21726 16940 21732 16992
rect 21784 16980 21790 16992
rect 21821 16983 21879 16989
rect 21821 16980 21833 16983
rect 21784 16952 21833 16980
rect 21784 16940 21790 16952
rect 21821 16949 21833 16952
rect 21867 16980 21879 16983
rect 22465 16983 22523 16989
rect 22465 16980 22477 16983
rect 21867 16952 22477 16980
rect 21867 16949 21879 16952
rect 21821 16943 21879 16949
rect 22465 16949 22477 16952
rect 22511 16980 22523 16983
rect 23109 16983 23167 16989
rect 23109 16980 23121 16983
rect 22511 16952 23121 16980
rect 22511 16949 22523 16952
rect 22465 16943 22523 16949
rect 23109 16949 23121 16952
rect 23155 16980 23167 16983
rect 23198 16980 23204 16992
rect 23155 16952 23204 16980
rect 23155 16949 23167 16952
rect 23109 16943 23167 16949
rect 23198 16940 23204 16952
rect 23256 16980 23262 16992
rect 23293 16983 23351 16989
rect 23293 16980 23305 16983
rect 23256 16952 23305 16980
rect 23256 16940 23262 16952
rect 23293 16949 23305 16952
rect 23339 16949 23351 16983
rect 24486 16980 24492 16992
rect 24447 16952 24492 16980
rect 23293 16943 23351 16949
rect 24486 16940 24492 16952
rect 24544 16940 24550 16992
rect 1104 16890 26128 16912
rect 1104 16838 5120 16890
rect 5172 16838 5184 16890
rect 5236 16838 5248 16890
rect 5300 16838 5312 16890
rect 5364 16838 5376 16890
rect 5428 16838 13462 16890
rect 13514 16838 13526 16890
rect 13578 16838 13590 16890
rect 13642 16838 13654 16890
rect 13706 16838 13718 16890
rect 13770 16838 21803 16890
rect 21855 16838 21867 16890
rect 21919 16838 21931 16890
rect 21983 16838 21995 16890
rect 22047 16838 22059 16890
rect 22111 16838 26128 16890
rect 1104 16816 26128 16838
rect 3418 16736 3424 16788
rect 3476 16776 3482 16788
rect 3881 16779 3939 16785
rect 3881 16776 3893 16779
rect 3476 16748 3893 16776
rect 3476 16736 3482 16748
rect 3881 16745 3893 16748
rect 3927 16745 3939 16779
rect 5626 16776 5632 16788
rect 3881 16739 3939 16745
rect 4632 16748 5632 16776
rect 2038 16600 2044 16652
rect 2096 16640 2102 16652
rect 4632 16649 4660 16748
rect 5626 16736 5632 16748
rect 5684 16736 5690 16788
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 8846 16776 8852 16788
rect 8803 16748 8852 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 8846 16736 8852 16748
rect 8904 16736 8910 16788
rect 9306 16776 9312 16788
rect 8956 16748 9312 16776
rect 8956 16708 8984 16748
rect 9306 16736 9312 16748
rect 9364 16776 9370 16788
rect 10134 16776 10140 16788
rect 9364 16748 10140 16776
rect 9364 16736 9370 16748
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10505 16779 10563 16785
rect 10505 16745 10517 16779
rect 10551 16776 10563 16779
rect 10778 16776 10784 16788
rect 10551 16748 10784 16776
rect 10551 16745 10563 16748
rect 10505 16739 10563 16745
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 14550 16776 14556 16788
rect 12452 16748 14556 16776
rect 8864 16680 8984 16708
rect 2133 16643 2191 16649
rect 2133 16640 2145 16643
rect 2096 16612 2145 16640
rect 2096 16600 2102 16612
rect 2133 16609 2145 16612
rect 2179 16609 2191 16643
rect 4617 16643 4675 16649
rect 4617 16640 4629 16643
rect 2133 16603 2191 16609
rect 3160 16612 4629 16640
rect 2400 16575 2458 16581
rect 2400 16541 2412 16575
rect 2446 16572 2458 16575
rect 2866 16572 2872 16584
rect 2446 16544 2872 16572
rect 2446 16541 2458 16544
rect 2400 16535 2458 16541
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 2958 16532 2964 16584
rect 3016 16572 3022 16584
rect 3160 16572 3188 16612
rect 4617 16609 4629 16612
rect 4663 16609 4675 16643
rect 4617 16603 4675 16609
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16640 8263 16643
rect 8864 16640 8892 16680
rect 12452 16649 12480 16748
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 16758 16776 16764 16788
rect 16719 16748 16764 16776
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 17034 16736 17040 16788
rect 17092 16776 17098 16788
rect 17957 16779 18015 16785
rect 17957 16776 17969 16779
rect 17092 16748 17969 16776
rect 17092 16736 17098 16748
rect 17957 16745 17969 16748
rect 18003 16745 18015 16779
rect 17957 16739 18015 16745
rect 17218 16668 17224 16720
rect 17276 16708 17282 16720
rect 17972 16708 18000 16739
rect 18506 16736 18512 16788
rect 18564 16776 18570 16788
rect 18693 16779 18751 16785
rect 18693 16776 18705 16779
rect 18564 16748 18705 16776
rect 18564 16736 18570 16748
rect 18693 16745 18705 16748
rect 18739 16745 18751 16779
rect 18693 16739 18751 16745
rect 19242 16736 19248 16788
rect 19300 16776 19306 16788
rect 19429 16779 19487 16785
rect 19429 16776 19441 16779
rect 19300 16748 19441 16776
rect 19300 16736 19306 16748
rect 19429 16745 19441 16748
rect 19475 16745 19487 16779
rect 19429 16739 19487 16745
rect 18138 16708 18144 16720
rect 17276 16680 17724 16708
rect 17972 16680 18144 16708
rect 17276 16668 17282 16680
rect 8251 16612 8892 16640
rect 8941 16643 8999 16649
rect 8251 16609 8263 16612
rect 8205 16603 8263 16609
rect 8941 16609 8953 16643
rect 8987 16609 8999 16643
rect 8941 16603 8999 16609
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16609 12495 16643
rect 14550 16640 14556 16652
rect 14511 16612 14556 16640
rect 12437 16603 12495 16609
rect 3970 16572 3976 16584
rect 3016 16544 3188 16572
rect 3931 16544 3976 16572
rect 3016 16532 3022 16544
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4062 16532 4068 16584
rect 4120 16581 4126 16584
rect 4430 16582 4436 16584
rect 4357 16581 4436 16582
rect 4120 16575 4169 16581
rect 4120 16541 4123 16575
rect 4157 16541 4169 16575
rect 4120 16535 4169 16541
rect 4230 16575 4288 16581
rect 4230 16541 4242 16575
rect 4276 16572 4288 16575
rect 4342 16575 4436 16581
rect 4276 16541 4292 16572
rect 4230 16535 4292 16541
rect 4342 16541 4354 16575
rect 4388 16554 4436 16575
rect 4388 16541 4400 16554
rect 4342 16535 4400 16541
rect 4120 16532 4126 16535
rect 3786 16464 3792 16516
rect 3844 16504 3850 16516
rect 4264 16504 4292 16535
rect 4430 16532 4436 16554
rect 4488 16532 4494 16584
rect 4890 16581 4896 16584
rect 4537 16575 4595 16581
rect 4537 16541 4549 16575
rect 4583 16572 4595 16575
rect 4884 16572 4896 16581
rect 4583 16544 4660 16572
rect 4851 16544 4896 16572
rect 4583 16541 4595 16544
rect 4537 16535 4595 16541
rect 3844 16476 4292 16504
rect 3844 16464 3850 16476
rect 4632 16448 4660 16544
rect 4884 16535 4896 16544
rect 4890 16532 4896 16535
rect 4948 16532 4954 16584
rect 7834 16532 7840 16584
rect 7892 16572 7898 16584
rect 8956 16572 8984 16603
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 16224 16612 16497 16640
rect 7892 16544 8984 16572
rect 7892 16532 7898 16544
rect 9030 16532 9036 16584
rect 9088 16572 9094 16584
rect 9197 16575 9255 16581
rect 9197 16572 9209 16575
rect 9088 16544 9209 16572
rect 9088 16532 9094 16544
rect 9197 16541 9209 16544
rect 9243 16541 9255 16575
rect 9197 16535 9255 16541
rect 10410 16532 10416 16584
rect 10468 16572 10474 16584
rect 10689 16575 10747 16581
rect 10689 16572 10701 16575
rect 10468 16544 10701 16572
rect 10468 16532 10474 16544
rect 10689 16541 10701 16544
rect 10735 16572 10747 16575
rect 11698 16572 11704 16584
rect 10735 16544 11704 16572
rect 10735 16541 10747 16544
rect 10689 16535 10747 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 15896 16544 16129 16572
rect 15896 16532 15902 16544
rect 16117 16541 16129 16544
rect 16163 16541 16175 16575
rect 16117 16535 16175 16541
rect 4798 16464 4804 16516
rect 4856 16504 4862 16516
rect 8018 16504 8024 16516
rect 4856 16476 8024 16504
rect 4856 16464 4862 16476
rect 8018 16464 8024 16476
rect 8076 16464 8082 16516
rect 8386 16504 8392 16516
rect 8347 16476 8392 16504
rect 8386 16464 8392 16476
rect 8444 16464 8450 16516
rect 8478 16464 8484 16516
rect 8536 16504 8542 16516
rect 11790 16504 11796 16516
rect 8536 16476 11796 16504
rect 8536 16464 8542 16476
rect 11790 16464 11796 16476
rect 11848 16464 11854 16516
rect 12704 16507 12762 16513
rect 12704 16473 12716 16507
rect 12750 16504 12762 16507
rect 13078 16504 13084 16516
rect 12750 16476 13084 16504
rect 12750 16473 12762 16476
rect 12704 16467 12762 16473
rect 13078 16464 13084 16476
rect 13136 16464 13142 16516
rect 14826 16513 14832 16516
rect 14820 16467 14832 16513
rect 14884 16504 14890 16516
rect 14884 16476 14920 16504
rect 14826 16464 14832 16467
rect 14884 16464 14890 16476
rect 15286 16464 15292 16516
rect 15344 16504 15350 16516
rect 16022 16504 16028 16516
rect 15344 16476 16028 16504
rect 15344 16464 15350 16476
rect 16022 16464 16028 16476
rect 16080 16504 16086 16516
rect 16224 16504 16252 16612
rect 16485 16609 16497 16612
rect 16531 16609 16543 16643
rect 17310 16640 17316 16652
rect 17271 16612 17316 16640
rect 16485 16603 16543 16609
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 16300 16569 16358 16575
rect 16300 16535 16312 16569
rect 16346 16535 16358 16569
rect 16300 16529 16358 16535
rect 16390 16532 16396 16584
rect 16448 16572 16454 16584
rect 16669 16575 16727 16581
rect 16448 16544 16493 16572
rect 16448 16532 16454 16544
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 17402 16572 17408 16584
rect 17363 16544 17408 16572
rect 16669 16535 16727 16541
rect 16080 16476 16252 16504
rect 16080 16464 16086 16476
rect 3513 16439 3571 16445
rect 3513 16405 3525 16439
rect 3559 16436 3571 16439
rect 3694 16436 3700 16448
rect 3559 16408 3700 16436
rect 3559 16405 3571 16408
rect 3513 16399 3571 16405
rect 3694 16396 3700 16408
rect 3752 16396 3758 16448
rect 4614 16396 4620 16448
rect 4672 16396 4678 16448
rect 5997 16439 6055 16445
rect 5997 16405 6009 16439
rect 6043 16436 6055 16439
rect 6086 16436 6092 16448
rect 6043 16408 6092 16436
rect 6043 16405 6055 16408
rect 5997 16399 6055 16405
rect 6086 16396 6092 16408
rect 6144 16436 6150 16448
rect 6822 16436 6828 16448
rect 6144 16408 6828 16436
rect 6144 16396 6150 16408
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 8294 16436 8300 16448
rect 8255 16408 8300 16436
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 10134 16396 10140 16448
rect 10192 16436 10198 16448
rect 10321 16439 10379 16445
rect 10321 16436 10333 16439
rect 10192 16408 10333 16436
rect 10192 16396 10198 16408
rect 10321 16405 10333 16408
rect 10367 16405 10379 16439
rect 10321 16399 10379 16405
rect 13817 16439 13875 16445
rect 13817 16405 13829 16439
rect 13863 16436 13875 16439
rect 14366 16436 14372 16448
rect 13863 16408 14372 16436
rect 13863 16405 13875 16408
rect 13817 16399 13875 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 14734 16396 14740 16448
rect 14792 16436 14798 16448
rect 15933 16439 15991 16445
rect 15933 16436 15945 16439
rect 14792 16408 15945 16436
rect 14792 16396 14798 16408
rect 15933 16405 15945 16408
rect 15979 16436 15991 16439
rect 16316 16436 16344 16529
rect 16684 16504 16712 16535
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 17696 16581 17724 16680
rect 18138 16668 18144 16680
rect 18196 16708 18202 16720
rect 19334 16708 19340 16720
rect 18196 16680 19340 16708
rect 18196 16668 18202 16680
rect 19334 16668 19340 16680
rect 19392 16668 19398 16720
rect 19444 16708 19472 16739
rect 19610 16736 19616 16788
rect 19668 16776 19674 16788
rect 25590 16776 25596 16788
rect 19668 16748 19713 16776
rect 25551 16748 25596 16776
rect 19668 16736 19674 16748
rect 25590 16736 25596 16748
rect 25648 16736 25654 16788
rect 20901 16711 20959 16717
rect 19444 16680 20484 16708
rect 17865 16643 17923 16649
rect 17865 16609 17877 16643
rect 17911 16640 17923 16643
rect 17954 16640 17960 16652
rect 17911 16612 17960 16640
rect 17911 16609 17923 16612
rect 17865 16603 17923 16609
rect 17954 16600 17960 16612
rect 18012 16640 18018 16652
rect 18230 16640 18236 16652
rect 18012 16612 18236 16640
rect 18012 16600 18018 16612
rect 18230 16600 18236 16612
rect 18288 16600 18294 16652
rect 18506 16600 18512 16652
rect 18564 16640 18570 16652
rect 18564 16612 19334 16640
rect 18564 16600 18570 16612
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16541 17739 16575
rect 17681 16535 17739 16541
rect 19306 16566 19334 16612
rect 19702 16600 19708 16652
rect 19760 16640 19766 16652
rect 20456 16649 20484 16680
rect 20901 16677 20913 16711
rect 20947 16708 20959 16711
rect 20947 16680 21496 16708
rect 20947 16677 20959 16680
rect 20901 16671 20959 16677
rect 21468 16649 21496 16680
rect 20349 16643 20407 16649
rect 20349 16640 20361 16643
rect 19760 16612 20361 16640
rect 19760 16600 19766 16612
rect 20349 16609 20361 16612
rect 20395 16609 20407 16643
rect 20349 16603 20407 16609
rect 20441 16643 20499 16649
rect 20441 16609 20453 16643
rect 20487 16640 20499 16643
rect 21453 16643 21511 16649
rect 20487 16612 21404 16640
rect 20487 16609 20499 16612
rect 20441 16603 20499 16609
rect 19518 16572 19524 16584
rect 19444 16566 19524 16572
rect 19306 16544 19524 16566
rect 19306 16538 19472 16544
rect 19518 16532 19524 16544
rect 19576 16532 19582 16584
rect 19794 16572 19800 16584
rect 19755 16544 19800 16572
rect 19794 16532 19800 16544
rect 19852 16532 19858 16584
rect 20714 16572 20720 16584
rect 20675 16544 20720 16572
rect 20714 16532 20720 16544
rect 20772 16532 20778 16584
rect 21376 16572 21404 16612
rect 21453 16609 21465 16643
rect 21499 16609 21511 16643
rect 21453 16603 21511 16609
rect 21542 16600 21548 16652
rect 21600 16640 21606 16652
rect 21913 16643 21971 16649
rect 21600 16612 21645 16640
rect 21600 16600 21606 16612
rect 21913 16609 21925 16643
rect 21959 16609 21971 16643
rect 23198 16640 23204 16652
rect 23159 16612 23204 16640
rect 21913 16603 21971 16609
rect 21726 16572 21732 16584
rect 21376 16544 21732 16572
rect 21726 16532 21732 16544
rect 21784 16572 21790 16584
rect 21928 16572 21956 16603
rect 23198 16600 23204 16612
rect 23256 16640 23262 16652
rect 24029 16643 24087 16649
rect 24029 16640 24041 16643
rect 23256 16612 24041 16640
rect 23256 16600 23262 16612
rect 24029 16609 24041 16612
rect 24075 16640 24087 16643
rect 24486 16640 24492 16652
rect 24075 16612 24492 16640
rect 24075 16609 24087 16612
rect 24029 16603 24087 16609
rect 24486 16600 24492 16612
rect 24544 16600 24550 16652
rect 24670 16640 24676 16652
rect 24631 16612 24676 16640
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 25608 16640 25636 16736
rect 25424 16612 25636 16640
rect 21784 16544 21956 16572
rect 22189 16575 22247 16581
rect 21784 16532 21790 16544
rect 22189 16541 22201 16575
rect 22235 16572 22247 16575
rect 22235 16544 22784 16572
rect 22235 16541 22247 16544
rect 22189 16535 22247 16541
rect 18046 16504 18052 16516
rect 16684 16476 18052 16504
rect 18046 16464 18052 16476
rect 18104 16464 18110 16516
rect 21361 16507 21419 16513
rect 21361 16473 21373 16507
rect 21407 16504 21419 16507
rect 22094 16504 22100 16516
rect 21407 16476 22100 16504
rect 21407 16473 21419 16476
rect 21361 16467 21419 16473
rect 22094 16464 22100 16476
rect 22152 16504 22158 16516
rect 22756 16504 22784 16544
rect 22830 16532 22836 16584
rect 22888 16572 22894 16584
rect 25424 16581 25452 16612
rect 25317 16575 25375 16581
rect 25317 16572 25329 16575
rect 22888 16544 25329 16572
rect 22888 16532 22894 16544
rect 25317 16541 25329 16544
rect 25363 16541 25375 16575
rect 25317 16535 25375 16541
rect 25409 16575 25467 16581
rect 25409 16541 25421 16575
rect 25455 16541 25467 16575
rect 25409 16535 25467 16541
rect 22922 16504 22928 16516
rect 22152 16476 22245 16504
rect 22756 16476 22928 16504
rect 22152 16464 22158 16476
rect 22922 16464 22928 16476
rect 22980 16464 22986 16516
rect 23109 16507 23167 16513
rect 23109 16473 23121 16507
rect 23155 16504 23167 16507
rect 23658 16504 23664 16516
rect 23155 16476 23664 16504
rect 23155 16473 23167 16476
rect 23109 16467 23167 16473
rect 23658 16464 23664 16476
rect 23716 16464 23722 16516
rect 23845 16507 23903 16513
rect 23845 16473 23857 16507
rect 23891 16504 23903 16507
rect 24946 16504 24952 16516
rect 23891 16476 24952 16504
rect 23891 16473 23903 16476
rect 23845 16467 23903 16473
rect 24946 16464 24952 16476
rect 25004 16464 25010 16516
rect 18322 16436 18328 16448
rect 15979 16408 18328 16436
rect 15979 16405 15991 16408
rect 15933 16399 15991 16405
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 19337 16439 19395 16445
rect 19337 16405 19349 16439
rect 19383 16436 19395 16439
rect 19426 16436 19432 16448
rect 19383 16408 19432 16436
rect 19383 16405 19395 16408
rect 19337 16399 19395 16405
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 19886 16436 19892 16448
rect 19847 16408 19892 16436
rect 19886 16396 19892 16408
rect 19944 16396 19950 16448
rect 20254 16436 20260 16448
rect 20215 16408 20260 16436
rect 20254 16396 20260 16408
rect 20312 16396 20318 16448
rect 20993 16439 21051 16445
rect 20993 16405 21005 16439
rect 21039 16436 21051 16439
rect 21174 16436 21180 16448
rect 21039 16408 21180 16436
rect 21039 16405 21051 16408
rect 20993 16399 21051 16405
rect 21174 16396 21180 16408
rect 21232 16396 21238 16448
rect 22554 16436 22560 16448
rect 22515 16408 22560 16436
rect 22554 16396 22560 16408
rect 22612 16396 22618 16448
rect 22646 16396 22652 16448
rect 22704 16436 22710 16448
rect 23014 16436 23020 16448
rect 22704 16408 22749 16436
rect 22975 16408 23020 16436
rect 22704 16396 22710 16408
rect 23014 16396 23020 16408
rect 23072 16396 23078 16448
rect 23477 16439 23535 16445
rect 23477 16405 23489 16439
rect 23523 16436 23535 16439
rect 23750 16436 23756 16448
rect 23523 16408 23756 16436
rect 23523 16405 23535 16408
rect 23477 16399 23535 16405
rect 23750 16396 23756 16408
rect 23808 16396 23814 16448
rect 23937 16439 23995 16445
rect 23937 16405 23949 16439
rect 23983 16436 23995 16439
rect 24578 16436 24584 16448
rect 23983 16408 24584 16436
rect 23983 16405 23995 16408
rect 23937 16399 23995 16405
rect 24578 16396 24584 16408
rect 24636 16396 24642 16448
rect 24765 16439 24823 16445
rect 24765 16405 24777 16439
rect 24811 16436 24823 16439
rect 24854 16436 24860 16448
rect 24811 16408 24860 16436
rect 24811 16405 24823 16408
rect 24765 16399 24823 16405
rect 24854 16396 24860 16408
rect 24912 16396 24918 16448
rect 25130 16436 25136 16448
rect 25091 16408 25136 16436
rect 25130 16396 25136 16408
rect 25188 16396 25194 16448
rect 1104 16346 26128 16368
rect 1104 16294 9291 16346
rect 9343 16294 9355 16346
rect 9407 16294 9419 16346
rect 9471 16294 9483 16346
rect 9535 16294 9547 16346
rect 9599 16294 17632 16346
rect 17684 16294 17696 16346
rect 17748 16294 17760 16346
rect 17812 16294 17824 16346
rect 17876 16294 17888 16346
rect 17940 16294 26128 16346
rect 1104 16272 26128 16294
rect 3234 16232 3240 16244
rect 3147 16204 3240 16232
rect 3234 16192 3240 16204
rect 3292 16232 3298 16244
rect 4062 16232 4068 16244
rect 3292 16204 4068 16232
rect 3292 16192 3298 16204
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 9769 16235 9827 16241
rect 9769 16232 9781 16235
rect 8352 16204 9781 16232
rect 8352 16192 8358 16204
rect 2774 16124 2780 16176
rect 2832 16164 2838 16176
rect 2869 16167 2927 16173
rect 2869 16164 2881 16167
rect 2832 16136 2881 16164
rect 2832 16124 2838 16136
rect 2869 16133 2881 16136
rect 2915 16133 2927 16167
rect 2869 16127 2927 16133
rect 3252 16105 3280 16192
rect 9416 16176 9444 16204
rect 9769 16201 9781 16204
rect 9815 16201 9827 16235
rect 9950 16232 9956 16244
rect 9911 16204 9956 16232
rect 9769 16195 9827 16201
rect 9950 16192 9956 16204
rect 10008 16192 10014 16244
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 10244 16204 10609 16232
rect 3326 16124 3332 16176
rect 3384 16124 3390 16176
rect 8018 16124 8024 16176
rect 8076 16164 8082 16176
rect 9306 16164 9312 16176
rect 8076 16136 9312 16164
rect 8076 16124 8082 16136
rect 9306 16124 9312 16136
rect 9364 16124 9370 16176
rect 9398 16124 9404 16176
rect 9456 16124 9462 16176
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16065 3111 16099
rect 3053 16059 3111 16065
rect 3237 16099 3295 16105
rect 3237 16065 3249 16099
rect 3283 16065 3295 16099
rect 3344 16096 3372 16124
rect 10244 16108 10272 16204
rect 10597 16201 10609 16204
rect 10643 16201 10655 16235
rect 13078 16232 13084 16244
rect 13039 16204 13084 16232
rect 10597 16195 10655 16201
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 13998 16232 14004 16244
rect 13959 16204 14004 16232
rect 13998 16192 14004 16204
rect 14056 16192 14062 16244
rect 14826 16232 14832 16244
rect 14787 16204 14832 16232
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 19242 16192 19248 16244
rect 19300 16232 19306 16244
rect 20717 16235 20775 16241
rect 19300 16204 19748 16232
rect 19300 16192 19306 16204
rect 12342 16164 12348 16176
rect 10796 16136 12348 16164
rect 3422 16099 3480 16105
rect 3422 16096 3434 16099
rect 3344 16068 3434 16096
rect 3237 16059 3295 16065
rect 3422 16065 3434 16068
rect 3468 16065 3480 16099
rect 3422 16059 3480 16065
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 4614 16096 4620 16108
rect 3651 16068 4620 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 3073 15960 3101 16059
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 8110 16105 8116 16108
rect 8104 16096 8116 16105
rect 8071 16068 8116 16096
rect 8104 16059 8116 16068
rect 8110 16056 8116 16059
rect 8168 16056 8174 16108
rect 9582 16096 9588 16108
rect 9543 16068 9588 16096
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16065 9735 16099
rect 10226 16096 10232 16108
rect 10187 16068 10232 16096
rect 9677 16059 9735 16065
rect 3329 16031 3387 16037
rect 3329 15997 3341 16031
rect 3375 16028 3387 16031
rect 3786 16028 3792 16040
rect 3375 16000 3792 16028
rect 3375 15997 3387 16000
rect 3329 15991 3387 15997
rect 3786 15988 3792 16000
rect 3844 15988 3850 16040
rect 7834 16028 7840 16040
rect 7795 16000 7840 16028
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 9692 16028 9720 16059
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 10796 16105 10824 16136
rect 12342 16124 12348 16136
rect 12400 16164 12406 16176
rect 13814 16164 13820 16176
rect 12400 16136 13820 16164
rect 12400 16124 12406 16136
rect 13814 16124 13820 16136
rect 13872 16124 13878 16176
rect 14090 16124 14096 16176
rect 14148 16164 14154 16176
rect 16393 16167 16451 16173
rect 14148 16136 15801 16164
rect 14148 16124 14154 16136
rect 15773 16122 15801 16136
rect 16393 16133 16405 16167
rect 16439 16164 16451 16167
rect 16914 16167 16972 16173
rect 16914 16164 16926 16167
rect 16439 16136 16926 16164
rect 16439 16133 16451 16136
rect 16393 16127 16451 16133
rect 16914 16133 16926 16136
rect 16960 16133 16972 16167
rect 16914 16127 16972 16133
rect 15773 16111 15848 16122
rect 10781 16099 10839 16105
rect 10781 16065 10793 16099
rect 10827 16065 10839 16099
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 10781 16059 10839 16065
rect 12360 16068 12449 16096
rect 12360 16028 12388 16068
rect 12437 16065 12449 16068
rect 12483 16096 12495 16099
rect 12526 16096 12532 16108
rect 12483 16068 12532 16096
rect 12483 16065 12495 16068
rect 12437 16059 12495 16065
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 12620 16099 12678 16105
rect 12620 16065 12632 16099
rect 12666 16096 12678 16099
rect 12894 16096 12900 16108
rect 12666 16068 12900 16096
rect 12666 16065 12678 16068
rect 12620 16059 12678 16065
rect 12894 16056 12900 16068
rect 12952 16056 12958 16108
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16096 13047 16099
rect 14182 16096 14188 16108
rect 13035 16068 13400 16096
rect 14143 16068 14188 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 12710 16028 12716 16040
rect 9232 16000 9720 16028
rect 10428 16000 12388 16028
rect 12671 16000 12716 16028
rect 3878 15960 3884 15972
rect 3073 15932 3884 15960
rect 3878 15920 3884 15932
rect 3936 15920 3942 15972
rect 9232 15969 9260 16000
rect 9217 15963 9275 15969
rect 9217 15929 9229 15963
rect 9263 15929 9275 15963
rect 9217 15923 9275 15929
rect 9306 15920 9312 15972
rect 9364 15960 9370 15972
rect 10428 15969 10456 16000
rect 12710 15988 12716 16000
rect 12768 15988 12774 16040
rect 12805 16031 12863 16037
rect 12805 15997 12817 16031
rect 12851 16028 12863 16031
rect 13170 16028 13176 16040
rect 12851 16000 13176 16028
rect 12851 15997 12863 16000
rect 12805 15991 12863 15997
rect 10413 15963 10471 15969
rect 9364 15932 9628 15960
rect 9364 15920 9370 15932
rect 3510 15852 3516 15904
rect 3568 15892 3574 15904
rect 7374 15892 7380 15904
rect 3568 15864 7380 15892
rect 3568 15852 3574 15864
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 8754 15852 8760 15904
rect 8812 15892 8818 15904
rect 9493 15895 9551 15901
rect 9493 15892 9505 15895
rect 8812 15864 9505 15892
rect 8812 15852 8818 15864
rect 9493 15861 9505 15864
rect 9539 15861 9551 15895
rect 9600 15892 9628 15932
rect 10413 15929 10425 15963
rect 10459 15929 10471 15963
rect 12434 15960 12440 15972
rect 10413 15923 10471 15929
rect 10520 15932 12440 15960
rect 10520 15892 10548 15932
rect 12434 15920 12440 15932
rect 12492 15920 12498 15972
rect 12820 15960 12848 15991
rect 13170 15988 13176 16000
rect 13228 15988 13234 16040
rect 12636 15932 12848 15960
rect 12636 15904 12664 15932
rect 9600 15864 10548 15892
rect 9493 15855 9551 15861
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 12342 15892 12348 15904
rect 10928 15864 12348 15892
rect 10928 15852 10934 15864
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 12618 15852 12624 15904
rect 12676 15852 12682 15904
rect 13372 15901 13400 16068
rect 14182 16056 14188 16068
rect 14240 16056 14246 16108
rect 14368 16099 14426 16105
rect 14368 16065 14380 16099
rect 14414 16065 14426 16099
rect 14368 16059 14426 16065
rect 13998 15988 14004 16040
rect 14056 16028 14062 16040
rect 14384 16028 14412 16059
rect 14458 16056 14464 16108
rect 14516 16096 14522 16108
rect 14516 16068 14561 16096
rect 14516 16056 14522 16068
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 15773 16105 15863 16111
rect 15657 16099 15715 16105
rect 14792 16068 14837 16096
rect 14792 16056 14798 16068
rect 15657 16065 15669 16099
rect 15703 16065 15715 16099
rect 15773 16094 15817 16105
rect 15805 16071 15817 16094
rect 15851 16071 15863 16105
rect 15805 16065 15863 16071
rect 15657 16059 15715 16065
rect 14056 16000 14412 16028
rect 14553 16031 14611 16037
rect 14056 15988 14062 16000
rect 14553 15997 14565 16031
rect 14599 16028 14611 16031
rect 14642 16028 14648 16040
rect 14599 16000 14648 16028
rect 14599 15997 14611 16000
rect 14553 15991 14611 15997
rect 14642 15988 14648 16000
rect 14700 15988 14706 16040
rect 15672 16028 15700 16059
rect 15930 16056 15936 16108
rect 15988 16096 15994 16108
rect 16209 16099 16267 16105
rect 15988 16068 16160 16096
rect 15988 16056 15994 16068
rect 16022 16028 16028 16040
rect 15672 16000 15884 16028
rect 15983 16000 16028 16028
rect 15856 15972 15884 16000
rect 16022 15988 16028 16000
rect 16080 15988 16086 16040
rect 16132 16028 16160 16068
rect 16209 16065 16221 16099
rect 16255 16096 16267 16099
rect 16255 16068 18092 16096
rect 16255 16065 16267 16068
rect 16209 16059 16267 16065
rect 16390 16028 16396 16040
rect 16132 16000 16396 16028
rect 16390 15988 16396 16000
rect 16448 15988 16454 16040
rect 16666 16028 16672 16040
rect 16627 16000 16672 16028
rect 16666 15988 16672 16000
rect 16724 15988 16730 16040
rect 15838 15920 15844 15972
rect 15896 15920 15902 15972
rect 13357 15895 13415 15901
rect 13357 15861 13369 15895
rect 13403 15892 13415 15895
rect 14366 15892 14372 15904
rect 13403 15864 14372 15892
rect 13403 15861 13415 15864
rect 13357 15855 13415 15861
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 18064 15901 18092 16068
rect 19720 16037 19748 16204
rect 20717 16201 20729 16235
rect 20763 16232 20775 16235
rect 20806 16232 20812 16244
rect 20763 16204 20812 16232
rect 20763 16201 20775 16204
rect 20717 16195 20775 16201
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 21174 16232 21180 16244
rect 21135 16204 21180 16232
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 21266 16192 21272 16244
rect 21324 16232 21330 16244
rect 21324 16204 21369 16232
rect 21324 16192 21330 16204
rect 21450 16192 21456 16244
rect 21508 16232 21514 16244
rect 22830 16232 22836 16244
rect 21508 16204 22836 16232
rect 21508 16192 21514 16204
rect 22830 16192 22836 16204
rect 22888 16192 22894 16244
rect 23014 16192 23020 16244
rect 23072 16232 23078 16244
rect 23201 16235 23259 16241
rect 23201 16232 23213 16235
rect 23072 16204 23213 16232
rect 23072 16192 23078 16204
rect 23201 16201 23213 16204
rect 23247 16201 23259 16235
rect 23201 16195 23259 16201
rect 23842 16192 23848 16244
rect 23900 16232 23906 16244
rect 24029 16235 24087 16241
rect 24029 16232 24041 16235
rect 23900 16204 24041 16232
rect 23900 16192 23906 16204
rect 24029 16201 24041 16204
rect 24075 16201 24087 16235
rect 24854 16232 24860 16244
rect 24815 16204 24860 16232
rect 24029 16195 24087 16201
rect 24854 16192 24860 16204
rect 24912 16192 24918 16244
rect 24946 16192 24952 16244
rect 25004 16232 25010 16244
rect 25406 16232 25412 16244
rect 25004 16204 25049 16232
rect 25367 16204 25412 16232
rect 25004 16192 25010 16204
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 20898 16124 20904 16176
rect 20956 16164 20962 16176
rect 21821 16167 21879 16173
rect 21821 16164 21833 16167
rect 20956 16136 21833 16164
rect 20956 16124 20962 16136
rect 21821 16133 21833 16136
rect 21867 16133 21879 16167
rect 21821 16127 21879 16133
rect 23569 16167 23627 16173
rect 23569 16133 23581 16167
rect 23615 16164 23627 16167
rect 24118 16164 24124 16176
rect 23615 16136 24124 16164
rect 23615 16133 23627 16136
rect 23569 16127 23627 16133
rect 24118 16124 24124 16136
rect 24176 16164 24182 16176
rect 24489 16167 24547 16173
rect 24489 16164 24501 16167
rect 24176 16136 24501 16164
rect 24176 16124 24182 16136
rect 24489 16133 24501 16136
rect 24535 16133 24547 16167
rect 24489 16127 24547 16133
rect 20349 16099 20407 16105
rect 20349 16065 20361 16099
rect 20395 16096 20407 16099
rect 21082 16096 21088 16108
rect 20395 16068 21088 16096
rect 20395 16065 20407 16068
rect 20349 16059 20407 16065
rect 21082 16056 21088 16068
rect 21140 16056 21146 16108
rect 21634 16096 21640 16108
rect 21192 16068 21640 16096
rect 19705 16031 19763 16037
rect 19705 15997 19717 16031
rect 19751 16028 19763 16031
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 19751 16000 19901 16028
rect 19751 15997 19763 16000
rect 19705 15991 19763 15997
rect 19889 15997 19901 16000
rect 19935 16028 19947 16031
rect 20165 16031 20223 16037
rect 20165 16028 20177 16031
rect 19935 16000 20177 16028
rect 19935 15997 19947 16000
rect 19889 15991 19947 15997
rect 20165 15997 20177 16000
rect 20211 15997 20223 16031
rect 20165 15991 20223 15997
rect 20257 16031 20315 16037
rect 20257 15997 20269 16031
rect 20303 16028 20315 16031
rect 21192 16028 21220 16068
rect 21634 16056 21640 16068
rect 21692 16096 21698 16108
rect 22097 16099 22155 16105
rect 22097 16096 22109 16099
rect 21692 16068 22109 16096
rect 21692 16056 21698 16068
rect 22097 16065 22109 16068
rect 22143 16096 22155 16099
rect 22833 16099 22891 16105
rect 22833 16096 22845 16099
rect 22143 16068 22845 16096
rect 22143 16065 22155 16068
rect 22097 16059 22155 16065
rect 22833 16065 22845 16068
rect 22879 16065 22891 16099
rect 22833 16059 22891 16065
rect 23661 16099 23719 16105
rect 23661 16065 23673 16099
rect 23707 16096 23719 16099
rect 24302 16096 24308 16108
rect 23707 16068 24308 16096
rect 23707 16065 23719 16068
rect 23661 16059 23719 16065
rect 24302 16056 24308 16068
rect 24360 16056 24366 16108
rect 25317 16099 25375 16105
rect 25317 16065 25329 16099
rect 25363 16065 25375 16099
rect 25317 16059 25375 16065
rect 20303 16000 21220 16028
rect 21361 16031 21419 16037
rect 20303 15997 20315 16000
rect 20257 15991 20315 15997
rect 21361 15997 21373 16031
rect 21407 15997 21419 16031
rect 21361 15991 21419 15997
rect 21821 16031 21879 16037
rect 21821 15997 21833 16031
rect 21867 16028 21879 16031
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 21867 16000 21925 16028
rect 21867 15997 21879 16000
rect 21821 15991 21879 15997
rect 21913 15997 21925 16000
rect 21959 16028 21971 16031
rect 22554 16028 22560 16040
rect 21959 16000 22094 16028
rect 22515 16000 22560 16028
rect 21959 15997 21971 16000
rect 21913 15991 21971 15997
rect 20180 15960 20208 15991
rect 20809 15963 20867 15969
rect 20180 15932 20300 15960
rect 18049 15895 18107 15901
rect 18049 15861 18061 15895
rect 18095 15892 18107 15895
rect 18966 15892 18972 15904
rect 18095 15864 18972 15892
rect 18095 15861 18107 15864
rect 18049 15855 18107 15861
rect 18966 15852 18972 15864
rect 19024 15852 19030 15904
rect 20272 15892 20300 15932
rect 20809 15929 20821 15963
rect 20855 15960 20867 15963
rect 20990 15960 20996 15972
rect 20855 15932 20996 15960
rect 20855 15929 20867 15932
rect 20809 15923 20867 15929
rect 20990 15920 20996 15932
rect 21048 15920 21054 15972
rect 21376 15892 21404 15991
rect 22066 15960 22094 16000
rect 22554 15988 22560 16000
rect 22612 15988 22618 16040
rect 22738 16028 22744 16040
rect 22699 16000 22744 16028
rect 22738 15988 22744 16000
rect 22796 15988 22802 16040
rect 23198 15988 23204 16040
rect 23256 16028 23262 16040
rect 23385 16031 23443 16037
rect 23385 16028 23397 16031
rect 23256 16000 23397 16028
rect 23256 15988 23262 16000
rect 23385 15997 23397 16000
rect 23431 15997 23443 16031
rect 23385 15991 23443 15997
rect 23474 15988 23480 16040
rect 23532 16028 23538 16040
rect 24213 16031 24271 16037
rect 24213 16028 24225 16031
rect 23532 16000 24225 16028
rect 23532 15988 23538 16000
rect 24213 15997 24225 16000
rect 24259 15997 24271 16031
rect 24213 15991 24271 15997
rect 24397 16031 24455 16037
rect 24397 15997 24409 16031
rect 24443 16028 24455 16031
rect 25222 16028 25228 16040
rect 24443 16000 25228 16028
rect 24443 15997 24455 16000
rect 24397 15991 24455 15997
rect 25222 15988 25228 16000
rect 25280 15988 25286 16040
rect 23750 15960 23756 15972
rect 22066 15932 23756 15960
rect 23750 15920 23756 15932
rect 23808 15920 23814 15972
rect 25332 15960 25360 16059
rect 25498 16028 25504 16040
rect 25459 16000 25504 16028
rect 25498 15988 25504 16000
rect 25556 15988 25562 16040
rect 25240 15932 25360 15960
rect 20272 15864 21404 15892
rect 22281 15895 22339 15901
rect 22281 15861 22293 15895
rect 22327 15892 22339 15895
rect 22646 15892 22652 15904
rect 22327 15864 22652 15892
rect 22327 15861 22339 15864
rect 22281 15855 22339 15861
rect 22646 15852 22652 15864
rect 22704 15852 22710 15904
rect 23658 15852 23664 15904
rect 23716 15892 23722 15904
rect 25240 15892 25268 15932
rect 23716 15864 25268 15892
rect 23716 15852 23722 15864
rect 1104 15802 26128 15824
rect 1104 15750 5120 15802
rect 5172 15750 5184 15802
rect 5236 15750 5248 15802
rect 5300 15750 5312 15802
rect 5364 15750 5376 15802
rect 5428 15750 13462 15802
rect 13514 15750 13526 15802
rect 13578 15750 13590 15802
rect 13642 15750 13654 15802
rect 13706 15750 13718 15802
rect 13770 15750 21803 15802
rect 21855 15750 21867 15802
rect 21919 15750 21931 15802
rect 21983 15750 21995 15802
rect 22047 15750 22059 15802
rect 22111 15750 26128 15802
rect 1104 15728 26128 15750
rect 3881 15691 3939 15697
rect 3881 15657 3893 15691
rect 3927 15688 3939 15691
rect 4798 15688 4804 15700
rect 3927 15660 4804 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 3145 15555 3203 15561
rect 3145 15521 3157 15555
rect 3191 15552 3203 15555
rect 3786 15552 3792 15564
rect 3191 15524 3792 15552
rect 3191 15521 3203 15524
rect 3145 15515 3203 15521
rect 3786 15512 3792 15524
rect 3844 15512 3850 15564
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3050 15484 3056 15496
rect 3007 15456 3056 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 3234 15484 3240 15496
rect 3195 15456 3240 15484
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 3330 15487 3388 15493
rect 3330 15453 3342 15487
rect 3376 15484 3388 15487
rect 3376 15456 3464 15484
rect 3376 15453 3388 15456
rect 3330 15447 3388 15453
rect 2774 15376 2780 15428
rect 2832 15416 2838 15428
rect 3436 15416 3464 15456
rect 3510 15444 3516 15496
rect 3568 15484 3574 15496
rect 3896 15484 3924 15651
rect 4798 15648 4804 15660
rect 4856 15648 4862 15700
rect 6546 15648 6552 15700
rect 6604 15688 6610 15700
rect 7009 15691 7067 15697
rect 7009 15688 7021 15691
rect 6604 15660 7021 15688
rect 6604 15648 6610 15660
rect 7009 15657 7021 15660
rect 7055 15688 7067 15691
rect 8478 15688 8484 15700
rect 7055 15660 8484 15688
rect 7055 15657 7067 15660
rect 7009 15651 7067 15657
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9493 15691 9551 15697
rect 9493 15688 9505 15691
rect 9088 15660 9505 15688
rect 9088 15648 9094 15660
rect 9493 15657 9505 15660
rect 9539 15657 9551 15691
rect 9493 15651 9551 15657
rect 10318 15648 10324 15700
rect 10376 15688 10382 15700
rect 10502 15688 10508 15700
rect 10376 15660 10508 15688
rect 10376 15648 10382 15660
rect 10502 15648 10508 15660
rect 10560 15688 10566 15700
rect 12069 15691 12127 15697
rect 12069 15688 12081 15691
rect 10560 15660 12081 15688
rect 10560 15648 10566 15660
rect 12069 15657 12081 15660
rect 12115 15657 12127 15691
rect 12342 15688 12348 15700
rect 12303 15660 12348 15688
rect 12069 15651 12127 15657
rect 7834 15580 7840 15632
rect 7892 15620 7898 15632
rect 7892 15592 10180 15620
rect 7892 15580 7898 15592
rect 5626 15552 5632 15564
rect 5587 15524 5632 15552
rect 5626 15512 5632 15524
rect 5684 15512 5690 15564
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 10152 15561 10180 15592
rect 11606 15580 11612 15632
rect 11664 15620 11670 15632
rect 11885 15623 11943 15629
rect 11885 15620 11897 15623
rect 11664 15592 11897 15620
rect 11664 15580 11670 15592
rect 11885 15589 11897 15592
rect 11931 15589 11943 15623
rect 11885 15583 11943 15589
rect 8205 15555 8263 15561
rect 8205 15552 8217 15555
rect 8168 15524 8217 15552
rect 8168 15512 8174 15524
rect 8205 15521 8217 15524
rect 8251 15521 8263 15555
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 8205 15515 8263 15521
rect 8404 15524 9045 15552
rect 3568 15456 3924 15484
rect 3568 15444 3574 15456
rect 4062 15444 4068 15496
rect 4120 15484 4126 15496
rect 7377 15487 7435 15493
rect 4120 15456 7328 15484
rect 4120 15444 4126 15456
rect 4246 15416 4252 15428
rect 2832 15388 2877 15416
rect 3436 15388 4252 15416
rect 2832 15376 2838 15388
rect 4246 15376 4252 15388
rect 4304 15376 4310 15428
rect 5896 15419 5954 15425
rect 5896 15385 5908 15419
rect 5942 15416 5954 15419
rect 6270 15416 6276 15428
rect 5942 15388 6276 15416
rect 5942 15385 5954 15388
rect 5896 15379 5954 15385
rect 6270 15376 6276 15388
rect 6328 15376 6334 15428
rect 7300 15416 7328 15456
rect 7377 15453 7389 15487
rect 7423 15484 7435 15487
rect 8018 15484 8024 15496
rect 7423 15456 8024 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 8018 15444 8024 15456
rect 8076 15444 8082 15496
rect 8404 15493 8432 15524
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 10137 15555 10195 15561
rect 9033 15515 9091 15521
rect 9140 15524 10088 15552
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15453 8447 15487
rect 8389 15447 8447 15453
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 8536 15456 8581 15484
rect 8536 15444 8542 15456
rect 9140 15416 9168 15524
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15453 9275 15487
rect 9217 15447 9275 15453
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15453 9367 15487
rect 9309 15447 9367 15453
rect 7300 15388 9168 15416
rect 7282 15308 7288 15360
rect 7340 15348 7346 15360
rect 7926 15348 7932 15360
rect 7340 15320 7932 15348
rect 7340 15308 7346 15320
rect 7926 15308 7932 15320
rect 7984 15348 7990 15360
rect 8021 15351 8079 15357
rect 8021 15348 8033 15351
rect 7984 15320 8033 15348
rect 7984 15308 7990 15320
rect 8021 15317 8033 15320
rect 8067 15348 8079 15351
rect 8478 15348 8484 15360
rect 8067 15320 8484 15348
rect 8067 15317 8079 15320
rect 8021 15311 8079 15317
rect 8478 15308 8484 15320
rect 8536 15308 8542 15360
rect 9232 15348 9260 15447
rect 9324 15416 9352 15447
rect 9398 15444 9404 15496
rect 9456 15484 9462 15496
rect 9585 15487 9643 15493
rect 9585 15484 9597 15487
rect 9456 15456 9597 15484
rect 9456 15444 9462 15456
rect 9585 15453 9597 15456
rect 9631 15453 9643 15487
rect 10060 15484 10088 15524
rect 10137 15521 10149 15555
rect 10183 15521 10195 15555
rect 12084 15552 12112 15651
rect 12342 15648 12348 15660
rect 12400 15648 12406 15700
rect 13541 15691 13599 15697
rect 13541 15657 13553 15691
rect 13587 15688 13599 15691
rect 14458 15688 14464 15700
rect 13587 15660 14464 15688
rect 13587 15657 13599 15660
rect 13541 15651 13599 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 16022 15688 16028 15700
rect 14783 15660 16028 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 16022 15648 16028 15660
rect 16080 15648 16086 15700
rect 19061 15691 19119 15697
rect 19061 15657 19073 15691
rect 19107 15688 19119 15691
rect 19242 15688 19248 15700
rect 19107 15660 19248 15688
rect 19107 15657 19119 15660
rect 19061 15651 19119 15657
rect 19242 15648 19248 15660
rect 19300 15648 19306 15700
rect 19978 15688 19984 15700
rect 19939 15660 19984 15688
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 20254 15648 20260 15700
rect 20312 15688 20318 15700
rect 20441 15691 20499 15697
rect 20441 15688 20453 15691
rect 20312 15660 20453 15688
rect 20312 15648 20318 15660
rect 20441 15657 20453 15660
rect 20487 15657 20499 15691
rect 20441 15651 20499 15657
rect 21082 15648 21088 15700
rect 21140 15688 21146 15700
rect 21269 15691 21327 15697
rect 21269 15688 21281 15691
rect 21140 15660 21281 15688
rect 21140 15648 21146 15660
rect 21269 15657 21281 15660
rect 21315 15657 21327 15691
rect 21269 15651 21327 15657
rect 22738 15648 22744 15700
rect 22796 15688 22802 15700
rect 22833 15691 22891 15697
rect 22833 15688 22845 15691
rect 22796 15660 22845 15688
rect 22796 15648 22802 15660
rect 22833 15657 22845 15660
rect 22879 15657 22891 15691
rect 22833 15651 22891 15657
rect 22922 15648 22928 15700
rect 22980 15688 22986 15700
rect 24121 15691 24179 15697
rect 22980 15660 23025 15688
rect 22980 15648 22986 15660
rect 24121 15657 24133 15691
rect 24167 15688 24179 15691
rect 24210 15688 24216 15700
rect 24167 15660 24216 15688
rect 24167 15657 24179 15660
rect 24121 15651 24179 15657
rect 24210 15648 24216 15660
rect 24268 15648 24274 15700
rect 24302 15648 24308 15700
rect 24360 15688 24366 15700
rect 24397 15691 24455 15697
rect 24397 15688 24409 15691
rect 24360 15660 24409 15688
rect 24360 15648 24366 15660
rect 24397 15657 24409 15660
rect 24443 15657 24455 15691
rect 25222 15688 25228 15700
rect 25183 15660 25228 15688
rect 24397 15651 24455 15657
rect 25222 15648 25228 15660
rect 25280 15648 25286 15700
rect 14277 15623 14335 15629
rect 14277 15589 14289 15623
rect 14323 15620 14335 15623
rect 15930 15620 15936 15632
rect 14323 15592 15936 15620
rect 14323 15589 14335 15592
rect 14277 15583 14335 15589
rect 15930 15580 15936 15592
rect 15988 15580 15994 15632
rect 21450 15620 21456 15632
rect 17236 15592 21456 15620
rect 12434 15552 12440 15564
rect 12084 15524 12440 15552
rect 10137 15515 10195 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 13262 15552 13268 15564
rect 12544 15524 13268 15552
rect 10060 15456 11100 15484
rect 9585 15447 9643 15453
rect 11072 15428 11100 15456
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11698 15484 11704 15496
rect 11204 15456 11704 15484
rect 11204 15444 11210 15456
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 12250 15484 12256 15496
rect 12211 15456 12256 15484
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 12544 15493 12572 15524
rect 13262 15512 13268 15524
rect 13320 15552 13326 15564
rect 13320 15524 14136 15552
rect 13320 15512 13326 15524
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15453 12587 15487
rect 13357 15487 13415 15493
rect 13357 15484 13369 15487
rect 12529 15447 12587 15453
rect 12635 15456 13369 15484
rect 9766 15416 9772 15428
rect 9324 15388 9772 15416
rect 9766 15376 9772 15388
rect 9824 15376 9830 15428
rect 10404 15419 10462 15425
rect 10404 15385 10416 15419
rect 10450 15416 10462 15419
rect 10594 15416 10600 15428
rect 10450 15388 10600 15416
rect 10450 15385 10462 15388
rect 10404 15379 10462 15385
rect 10594 15376 10600 15388
rect 10652 15376 10658 15428
rect 11054 15376 11060 15428
rect 11112 15376 11118 15428
rect 11440 15388 11744 15416
rect 11440 15348 11468 15388
rect 9232 15320 11468 15348
rect 11514 15308 11520 15360
rect 11572 15348 11578 15360
rect 11716 15348 11744 15388
rect 12434 15376 12440 15428
rect 12492 15416 12498 15428
rect 12635 15416 12663 15456
rect 13357 15453 13369 15456
rect 13403 15453 13415 15487
rect 13630 15484 13636 15496
rect 13591 15456 13636 15484
rect 13357 15447 13415 15453
rect 13630 15444 13636 15456
rect 13688 15444 13694 15496
rect 14108 15493 14136 15524
rect 14093 15487 14151 15493
rect 14093 15453 14105 15487
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 17236 15416 17264 15592
rect 21450 15580 21456 15592
rect 21508 15580 21514 15632
rect 24762 15620 24768 15632
rect 23492 15592 24768 15620
rect 23492 15564 23520 15592
rect 24762 15580 24768 15592
rect 24820 15620 24826 15632
rect 25498 15620 25504 15632
rect 24820 15592 25504 15620
rect 24820 15580 24826 15592
rect 19242 15512 19248 15564
rect 19300 15552 19306 15564
rect 19337 15555 19395 15561
rect 19337 15552 19349 15555
rect 19300 15524 19349 15552
rect 19300 15512 19306 15524
rect 19337 15521 19349 15524
rect 19383 15521 19395 15555
rect 19337 15515 19395 15521
rect 19521 15555 19579 15561
rect 19521 15521 19533 15555
rect 19567 15552 19579 15555
rect 20530 15552 20536 15564
rect 19567 15524 20536 15552
rect 19567 15521 19579 15524
rect 19521 15515 19579 15521
rect 20530 15512 20536 15524
rect 20588 15512 20594 15564
rect 20714 15512 20720 15564
rect 20772 15552 20778 15564
rect 20901 15555 20959 15561
rect 20901 15552 20913 15555
rect 20772 15524 20913 15552
rect 20772 15512 20778 15524
rect 20901 15521 20913 15524
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 21085 15555 21143 15561
rect 21085 15521 21097 15555
rect 21131 15552 21143 15555
rect 21542 15552 21548 15564
rect 21131 15524 21548 15552
rect 21131 15521 21143 15524
rect 21085 15515 21143 15521
rect 21542 15512 21548 15524
rect 21600 15552 21606 15564
rect 21821 15555 21879 15561
rect 21821 15552 21833 15555
rect 21600 15524 21833 15552
rect 21600 15512 21606 15524
rect 21821 15521 21833 15524
rect 21867 15552 21879 15555
rect 22097 15555 22155 15561
rect 22097 15552 22109 15555
rect 21867 15524 22109 15552
rect 21867 15521 21879 15524
rect 21821 15515 21879 15521
rect 22097 15521 22109 15524
rect 22143 15552 22155 15555
rect 22281 15555 22339 15561
rect 22281 15552 22293 15555
rect 22143 15524 22293 15552
rect 22143 15521 22155 15524
rect 22097 15515 22155 15521
rect 22281 15521 22293 15524
rect 22327 15552 22339 15555
rect 22465 15555 22523 15561
rect 22465 15552 22477 15555
rect 22327 15524 22477 15552
rect 22327 15521 22339 15524
rect 22281 15515 22339 15521
rect 22465 15521 22477 15524
rect 22511 15552 22523 15555
rect 22554 15552 22560 15564
rect 22511 15524 22560 15552
rect 22511 15521 22523 15524
rect 22465 15515 22523 15521
rect 22554 15512 22560 15524
rect 22612 15552 22618 15564
rect 23474 15552 23480 15564
rect 22612 15524 23480 15552
rect 22612 15512 22618 15524
rect 23474 15512 23480 15524
rect 23532 15512 23538 15564
rect 23750 15552 23756 15564
rect 23711 15524 23756 15552
rect 23750 15512 23756 15524
rect 23808 15512 23814 15564
rect 24964 15561 24992 15592
rect 25498 15580 25504 15592
rect 25556 15580 25562 15632
rect 24949 15555 25007 15561
rect 24949 15521 24961 15555
rect 24995 15521 25007 15555
rect 24949 15515 25007 15521
rect 18690 15484 18696 15496
rect 18651 15456 18696 15484
rect 18690 15444 18696 15456
rect 18748 15444 18754 15496
rect 20162 15484 20168 15496
rect 20123 15456 20168 15484
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 20809 15487 20867 15493
rect 20809 15453 20821 15487
rect 20855 15484 20867 15487
rect 20990 15484 20996 15496
rect 20855 15456 20996 15484
rect 20855 15453 20867 15456
rect 20809 15447 20867 15453
rect 20990 15444 20996 15456
rect 21048 15444 21054 15496
rect 22646 15484 22652 15496
rect 22607 15456 22652 15484
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 23658 15444 23664 15496
rect 23716 15484 23722 15496
rect 23937 15487 23995 15493
rect 23937 15484 23949 15487
rect 23716 15456 23949 15484
rect 23716 15444 23722 15456
rect 23937 15453 23949 15456
rect 23983 15484 23995 15487
rect 24026 15484 24032 15496
rect 23983 15456 24032 15484
rect 23983 15453 23995 15456
rect 23937 15447 23995 15453
rect 24026 15444 24032 15456
rect 24084 15444 24090 15496
rect 24578 15444 24584 15496
rect 24636 15484 24642 15496
rect 24765 15487 24823 15493
rect 24765 15484 24777 15487
rect 24636 15456 24777 15484
rect 24636 15444 24642 15456
rect 24765 15453 24777 15456
rect 24811 15453 24823 15487
rect 25406 15484 25412 15496
rect 25367 15456 25412 15484
rect 24765 15447 24823 15453
rect 25406 15444 25412 15456
rect 25464 15444 25470 15496
rect 18230 15416 18236 15428
rect 12492 15388 12663 15416
rect 13280 15388 17264 15416
rect 18191 15388 18236 15416
rect 12492 15376 12498 15388
rect 13280 15348 13308 15388
rect 18230 15376 18236 15388
rect 18288 15376 18294 15428
rect 18322 15376 18328 15428
rect 18380 15416 18386 15428
rect 18417 15419 18475 15425
rect 18417 15416 18429 15419
rect 18380 15388 18429 15416
rect 18380 15376 18386 15388
rect 18417 15385 18429 15388
rect 18463 15385 18475 15419
rect 18598 15416 18604 15428
rect 18559 15388 18604 15416
rect 18417 15379 18475 15385
rect 18598 15376 18604 15388
rect 18656 15376 18662 15428
rect 21729 15419 21787 15425
rect 21729 15416 21741 15419
rect 20364 15388 21741 15416
rect 11572 15320 11617 15348
rect 11716 15320 13308 15348
rect 13817 15351 13875 15357
rect 11572 15308 11578 15320
rect 13817 15317 13829 15351
rect 13863 15348 13875 15351
rect 14737 15351 14795 15357
rect 14737 15348 14749 15351
rect 13863 15320 14749 15348
rect 13863 15317 13875 15320
rect 13817 15311 13875 15317
rect 14737 15317 14749 15320
rect 14783 15317 14795 15351
rect 14737 15311 14795 15317
rect 14921 15351 14979 15357
rect 14921 15317 14933 15351
rect 14967 15348 14979 15351
rect 15194 15348 15200 15360
rect 14967 15320 15200 15348
rect 14967 15317 14979 15320
rect 14921 15311 14979 15317
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 18506 15308 18512 15360
rect 18564 15348 18570 15360
rect 18877 15351 18935 15357
rect 18877 15348 18889 15351
rect 18564 15320 18889 15348
rect 18564 15308 18570 15320
rect 18877 15317 18889 15320
rect 18923 15317 18935 15351
rect 18877 15311 18935 15317
rect 19610 15308 19616 15360
rect 19668 15348 19674 15360
rect 20364 15357 20392 15388
rect 21729 15385 21741 15388
rect 21775 15385 21787 15419
rect 21729 15379 21787 15385
rect 23293 15419 23351 15425
rect 23293 15385 23305 15419
rect 23339 15416 23351 15419
rect 23339 15388 24164 15416
rect 23339 15385 23351 15388
rect 23293 15379 23351 15385
rect 20349 15351 20407 15357
rect 19668 15320 19713 15348
rect 19668 15308 19674 15320
rect 20349 15317 20361 15351
rect 20395 15317 20407 15351
rect 20349 15311 20407 15317
rect 20530 15308 20536 15360
rect 20588 15348 20594 15360
rect 21637 15351 21695 15357
rect 21637 15348 21649 15351
rect 20588 15320 21649 15348
rect 20588 15308 20594 15320
rect 21637 15317 21649 15320
rect 21683 15317 21695 15351
rect 21637 15311 21695 15317
rect 23382 15308 23388 15360
rect 23440 15348 23446 15360
rect 24136 15348 24164 15388
rect 24210 15376 24216 15428
rect 24268 15416 24274 15428
rect 24857 15419 24915 15425
rect 24857 15416 24869 15419
rect 24268 15388 24869 15416
rect 24268 15376 24274 15388
rect 24857 15385 24869 15388
rect 24903 15385 24915 15419
rect 24857 15379 24915 15385
rect 24670 15348 24676 15360
rect 23440 15320 23485 15348
rect 24136 15320 24676 15348
rect 23440 15308 23446 15320
rect 24670 15308 24676 15320
rect 24728 15308 24734 15360
rect 1104 15258 26128 15280
rect 1104 15206 9291 15258
rect 9343 15206 9355 15258
rect 9407 15206 9419 15258
rect 9471 15206 9483 15258
rect 9535 15206 9547 15258
rect 9599 15206 17632 15258
rect 17684 15206 17696 15258
rect 17748 15206 17760 15258
rect 17812 15206 17824 15258
rect 17876 15206 17888 15258
rect 17940 15206 26128 15258
rect 1104 15184 26128 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 3050 15144 3056 15156
rect 1627 15116 3056 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 4246 15144 4252 15156
rect 4207 15116 4252 15144
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 4706 15144 4712 15156
rect 4667 15116 4712 15144
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 8662 15144 8668 15156
rect 6564 15116 8668 15144
rect 2774 15076 2780 15088
rect 2746 15036 2780 15076
rect 2832 15036 2838 15088
rect 6564 15076 6592 15116
rect 8662 15104 8668 15116
rect 8720 15144 8726 15156
rect 8757 15147 8815 15153
rect 8757 15144 8769 15147
rect 8720 15116 8769 15144
rect 8720 15104 8726 15116
rect 8757 15113 8769 15116
rect 8803 15113 8815 15147
rect 10594 15144 10600 15156
rect 10555 15116 10600 15144
rect 8757 15107 8815 15113
rect 10594 15104 10600 15116
rect 10652 15104 10658 15156
rect 14182 15104 14188 15156
rect 14240 15144 14246 15156
rect 16114 15144 16120 15156
rect 14240 15116 16120 15144
rect 14240 15104 14246 15116
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 18138 15104 18144 15156
rect 18196 15144 18202 15156
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 18196 15116 18245 15144
rect 18196 15104 18202 15116
rect 18233 15113 18245 15116
rect 18279 15113 18291 15147
rect 18782 15144 18788 15156
rect 18743 15116 18788 15144
rect 18233 15107 18291 15113
rect 18782 15104 18788 15116
rect 18840 15104 18846 15156
rect 19153 15147 19211 15153
rect 19153 15113 19165 15147
rect 19199 15144 19211 15147
rect 19610 15144 19616 15156
rect 19199 15116 19616 15144
rect 19199 15113 19211 15116
rect 19153 15107 19211 15113
rect 19610 15104 19616 15116
rect 19668 15104 19674 15156
rect 20162 15104 20168 15156
rect 20220 15144 20226 15156
rect 20257 15147 20315 15153
rect 20257 15144 20269 15147
rect 20220 15116 20269 15144
rect 20220 15104 20226 15116
rect 20257 15113 20269 15116
rect 20303 15113 20315 15147
rect 20257 15107 20315 15113
rect 20622 15104 20628 15156
rect 20680 15144 20686 15156
rect 20809 15147 20867 15153
rect 20809 15144 20821 15147
rect 20680 15116 20821 15144
rect 20680 15104 20686 15116
rect 20809 15113 20821 15116
rect 20855 15113 20867 15147
rect 21266 15144 21272 15156
rect 21227 15116 21272 15144
rect 20809 15107 20867 15113
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 23293 15147 23351 15153
rect 23293 15113 23305 15147
rect 23339 15144 23351 15147
rect 23382 15144 23388 15156
rect 23339 15116 23388 15144
rect 23339 15113 23351 15116
rect 23293 15107 23351 15113
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 24305 15147 24363 15153
rect 24305 15113 24317 15147
rect 24351 15144 24363 15147
rect 25406 15144 25412 15156
rect 24351 15116 25412 15144
rect 24351 15113 24363 15116
rect 24305 15107 24363 15113
rect 25406 15104 25412 15116
rect 25464 15104 25470 15156
rect 7834 15076 7840 15088
rect 3160 15048 6592 15076
rect 6656 15048 7840 15076
rect 2746 15017 2774 15036
rect 2705 15011 2774 15017
rect 2705 14977 2717 15011
rect 2751 14980 2774 15011
rect 2958 15008 2964 15020
rect 2919 14980 2964 15008
rect 2751 14977 2763 14980
rect 2705 14971 2763 14977
rect 2958 14968 2964 14980
rect 3016 14968 3022 15020
rect 2682 14764 2688 14816
rect 2740 14804 2746 14816
rect 3160 14804 3188 15048
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 3510 15008 3516 15020
rect 3467 14980 3516 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 3602 14968 3608 15020
rect 3660 15008 3666 15020
rect 3973 15011 4031 15017
rect 3660 14980 3704 15008
rect 3660 14968 3666 14980
rect 3973 14977 3985 15011
rect 4019 15008 4031 15011
rect 4614 15008 4620 15020
rect 4019 14980 4476 15008
rect 4575 14980 4620 15008
rect 4019 14977 4031 14980
rect 3973 14971 4031 14977
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 3697 14943 3755 14949
rect 3697 14940 3709 14943
rect 3292 14912 3709 14940
rect 3292 14900 3298 14912
rect 3697 14909 3709 14912
rect 3743 14909 3755 14943
rect 3697 14903 3755 14909
rect 3786 14900 3792 14952
rect 3844 14940 3850 14952
rect 3844 14912 3889 14940
rect 3844 14900 3850 14912
rect 4448 14872 4476 14980
rect 4614 14968 4620 14980
rect 4672 15008 4678 15020
rect 5077 15011 5135 15017
rect 5077 15008 5089 15011
rect 4672 14980 5089 15008
rect 4672 14968 4678 14980
rect 5077 14977 5089 14980
rect 5123 14977 5135 15011
rect 6546 15008 6552 15020
rect 6507 14980 6552 15008
rect 5077 14971 5135 14977
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 6656 15017 6684 15048
rect 7834 15036 7840 15048
rect 7892 15036 7898 15088
rect 10226 15076 10232 15088
rect 8956 15048 10232 15076
rect 6914 15017 6920 15020
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 6908 14971 6920 15017
rect 6972 15008 6978 15020
rect 6972 14980 7008 15008
rect 6914 14968 6920 14971
rect 6972 14968 6978 14980
rect 8570 14968 8576 15020
rect 8628 15008 8634 15020
rect 8956 15017 8984 15048
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 12986 15036 12992 15088
rect 13044 15076 13050 15088
rect 19978 15076 19984 15088
rect 13044 15048 19984 15076
rect 13044 15036 13050 15048
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 24762 15076 24768 15088
rect 24723 15048 24768 15076
rect 24762 15036 24768 15048
rect 24820 15036 24826 15088
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8628 14980 8953 15008
rect 8628 14968 8634 14980
rect 8941 14977 8953 14980
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 9122 14968 9128 15020
rect 9180 15008 9186 15020
rect 9953 15011 10011 15017
rect 9953 15008 9965 15011
rect 9180 14980 9965 15008
rect 9180 14968 9186 14980
rect 9953 14977 9965 14980
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 10134 14968 10140 15020
rect 10192 15008 10198 15020
rect 10192 14980 10236 15008
rect 10192 14968 10198 14980
rect 10318 14968 10324 15020
rect 10376 15008 10382 15020
rect 10505 15011 10563 15017
rect 10376 14980 10421 15008
rect 10376 14968 10382 14980
rect 10505 14977 10517 15011
rect 10551 15008 10563 15011
rect 11514 15008 11520 15020
rect 10551 14980 11520 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 12894 15008 12900 15020
rect 12855 14980 12900 15008
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 14921 15011 14979 15017
rect 14921 15008 14933 15011
rect 13872 14980 14933 15008
rect 13872 14968 13878 14980
rect 14921 14977 14933 14980
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 15102 14968 15108 15020
rect 15160 15008 15166 15020
rect 15269 15011 15327 15017
rect 15269 15008 15281 15011
rect 15160 14980 15281 15008
rect 15160 14968 15166 14980
rect 15269 14977 15281 14980
rect 15315 14977 15327 15011
rect 16666 15008 16672 15020
rect 16627 14980 16672 15008
rect 15269 14971 15327 14977
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 16925 15011 16983 15017
rect 16925 15008 16937 15011
rect 16816 14980 16937 15008
rect 16816 14968 16822 14980
rect 16925 14977 16937 14980
rect 16971 14977 16983 15011
rect 16925 14971 16983 14977
rect 18524 14980 19334 15008
rect 4522 14900 4528 14952
rect 4580 14940 4586 14952
rect 4801 14943 4859 14949
rect 4801 14940 4813 14943
rect 4580 14912 4813 14940
rect 4580 14900 4586 14912
rect 4801 14909 4813 14912
rect 4847 14909 4859 14943
rect 4801 14903 4859 14909
rect 10229 14943 10287 14949
rect 10229 14909 10241 14943
rect 10275 14940 10287 14943
rect 10870 14940 10876 14952
rect 10275 14912 10876 14940
rect 10275 14909 10287 14912
rect 10229 14903 10287 14909
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 14550 14900 14556 14952
rect 14608 14940 14614 14952
rect 15013 14943 15071 14949
rect 15013 14940 15025 14943
rect 14608 14912 15025 14940
rect 14608 14900 14614 14912
rect 15013 14909 15025 14912
rect 15059 14909 15071 14943
rect 15013 14903 15071 14909
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 18524 14949 18552 14980
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18196 14912 18521 14940
rect 18196 14900 18202 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14940 18751 14943
rect 19058 14940 19064 14952
rect 18739 14912 19064 14940
rect 18739 14909 18751 14912
rect 18693 14903 18751 14909
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 19306 14940 19334 14980
rect 19518 14968 19524 15020
rect 19576 15008 19582 15020
rect 20441 15011 20499 15017
rect 19576 14980 19621 15008
rect 19576 14968 19582 14980
rect 20441 14977 20453 15011
rect 20487 15008 20499 15011
rect 20530 15008 20536 15020
rect 20487 14980 20536 15008
rect 20487 14977 20499 14980
rect 20441 14971 20499 14977
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 20806 15008 20812 15020
rect 20767 14980 20812 15008
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 21082 15008 21088 15020
rect 21043 14980 21088 15008
rect 21082 14968 21088 14980
rect 21140 14968 21146 15020
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 14977 21235 15011
rect 23290 15008 23296 15020
rect 23251 14980 23296 15008
rect 21177 14971 21235 14977
rect 19981 14943 20039 14949
rect 19981 14940 19993 14943
rect 19306 14912 19993 14940
rect 19981 14909 19993 14912
rect 20027 14909 20039 14943
rect 19981 14903 20039 14909
rect 20625 14943 20683 14949
rect 20625 14909 20637 14943
rect 20671 14940 20683 14943
rect 20714 14940 20720 14952
rect 20671 14912 20720 14940
rect 20671 14909 20683 14912
rect 20625 14903 20683 14909
rect 20714 14900 20720 14912
rect 20772 14900 20778 14952
rect 20824 14940 20852 14968
rect 21192 14940 21220 14971
rect 23290 14968 23296 14980
rect 23348 14968 23354 15020
rect 23569 15011 23627 15017
rect 23569 14977 23581 15011
rect 23615 15008 23627 15011
rect 23658 15008 23664 15020
rect 23615 14980 23664 15008
rect 23615 14977 23627 14980
rect 23569 14971 23627 14977
rect 23658 14968 23664 14980
rect 23716 14968 23722 15020
rect 23750 14968 23756 15020
rect 23808 15008 23814 15020
rect 23937 15011 23995 15017
rect 23937 15008 23949 15011
rect 23808 14980 23949 15008
rect 23808 14968 23814 14980
rect 23937 14977 23949 14980
rect 23983 14977 23995 15011
rect 24118 15008 24124 15020
rect 24079 14980 24124 15008
rect 23937 14971 23995 14977
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 20824 14912 21220 14940
rect 5534 14872 5540 14884
rect 4448 14844 5540 14872
rect 5534 14832 5540 14844
rect 5592 14832 5598 14884
rect 14734 14872 14740 14884
rect 7576 14844 14740 14872
rect 4062 14804 4068 14816
rect 2740 14776 3188 14804
rect 4023 14776 4068 14804
rect 2740 14764 2746 14776
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 6546 14764 6552 14816
rect 6604 14804 6610 14816
rect 7576 14804 7604 14844
rect 14734 14832 14740 14844
rect 14792 14832 14798 14884
rect 19518 14872 19524 14884
rect 17972 14844 19524 14872
rect 8018 14804 8024 14816
rect 6604 14776 7604 14804
rect 7979 14776 8024 14804
rect 6604 14764 6610 14776
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 9122 14804 9128 14816
rect 9083 14776 9128 14804
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 10873 14807 10931 14813
rect 10873 14773 10885 14807
rect 10919 14804 10931 14807
rect 11514 14804 11520 14816
rect 10919 14776 11520 14804
rect 10919 14773 10931 14776
rect 10873 14767 10931 14773
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 12805 14807 12863 14813
rect 12805 14773 12817 14807
rect 12851 14804 12863 14807
rect 12894 14804 12900 14816
rect 12851 14776 12900 14804
rect 12851 14773 12863 14776
rect 12805 14767 12863 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 14182 14804 14188 14816
rect 14143 14776 14188 14804
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 14918 14764 14924 14816
rect 14976 14804 14982 14816
rect 16390 14804 16396 14816
rect 14976 14776 16396 14804
rect 14976 14764 14982 14776
rect 16390 14764 16396 14776
rect 16448 14804 16454 14816
rect 17972 14804 18000 14844
rect 19518 14832 19524 14844
rect 19576 14832 19582 14884
rect 16448 14776 18000 14804
rect 18049 14807 18107 14813
rect 16448 14764 16454 14776
rect 18049 14773 18061 14807
rect 18095 14804 18107 14807
rect 18138 14804 18144 14816
rect 18095 14776 18144 14804
rect 18095 14773 18107 14776
rect 18049 14767 18107 14773
rect 18138 14764 18144 14776
rect 18196 14764 18202 14816
rect 19610 14804 19616 14816
rect 19571 14776 19616 14804
rect 19610 14764 19616 14776
rect 19668 14764 19674 14816
rect 21082 14764 21088 14816
rect 21140 14804 21146 14816
rect 21545 14807 21603 14813
rect 21545 14804 21557 14807
rect 21140 14776 21557 14804
rect 21140 14764 21146 14776
rect 21545 14773 21557 14776
rect 21591 14804 21603 14807
rect 23658 14804 23664 14816
rect 21591 14776 23664 14804
rect 21591 14773 21603 14776
rect 21545 14767 21603 14773
rect 23658 14764 23664 14776
rect 23716 14804 23722 14816
rect 24489 14807 24547 14813
rect 24489 14804 24501 14807
rect 23716 14776 24501 14804
rect 23716 14764 23722 14776
rect 24489 14773 24501 14776
rect 24535 14773 24547 14807
rect 24489 14767 24547 14773
rect 1104 14714 26128 14736
rect 1104 14662 5120 14714
rect 5172 14662 5184 14714
rect 5236 14662 5248 14714
rect 5300 14662 5312 14714
rect 5364 14662 5376 14714
rect 5428 14662 13462 14714
rect 13514 14662 13526 14714
rect 13578 14662 13590 14714
rect 13642 14662 13654 14714
rect 13706 14662 13718 14714
rect 13770 14662 21803 14714
rect 21855 14662 21867 14714
rect 21919 14662 21931 14714
rect 21983 14662 21995 14714
rect 22047 14662 22059 14714
rect 22111 14662 26128 14714
rect 1104 14640 26128 14662
rect 2406 14560 2412 14612
rect 2464 14600 2470 14612
rect 5169 14603 5227 14609
rect 2464 14572 3832 14600
rect 2464 14560 2470 14572
rect 3050 14424 3056 14476
rect 3108 14473 3114 14476
rect 3804 14473 3832 14572
rect 5169 14569 5181 14603
rect 5215 14600 5227 14603
rect 5534 14600 5540 14612
rect 5215 14572 5540 14600
rect 5215 14569 5227 14572
rect 5169 14563 5227 14569
rect 5534 14560 5540 14572
rect 5592 14600 5598 14612
rect 6086 14600 6092 14612
rect 5592 14572 6092 14600
rect 5592 14560 5598 14572
rect 6086 14560 6092 14572
rect 6144 14560 6150 14612
rect 6270 14600 6276 14612
rect 6231 14572 6276 14600
rect 6270 14560 6276 14572
rect 6328 14560 6334 14612
rect 6380 14572 6961 14600
rect 3108 14464 3116 14473
rect 3789 14467 3847 14473
rect 3108 14436 3153 14464
rect 3108 14427 3116 14436
rect 3789 14433 3801 14467
rect 3835 14433 3847 14467
rect 5902 14464 5908 14476
rect 5863 14436 5908 14464
rect 3789 14427 3847 14433
rect 3108 14424 3114 14427
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 2777 14399 2835 14405
rect 2777 14365 2789 14399
rect 2823 14396 2835 14399
rect 2866 14396 2872 14408
rect 2823 14368 2872 14396
rect 2823 14365 2835 14368
rect 2777 14359 2835 14365
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 2958 14356 2964 14408
rect 3016 14396 3022 14408
rect 3016 14368 3061 14396
rect 3016 14356 3022 14368
rect 3142 14356 3148 14408
rect 3200 14396 3206 14408
rect 4062 14405 4068 14408
rect 3329 14399 3387 14405
rect 3200 14368 3245 14396
rect 3200 14356 3206 14368
rect 3329 14365 3341 14399
rect 3375 14365 3387 14399
rect 4056 14396 4068 14405
rect 4023 14368 4068 14396
rect 3329 14359 3387 14365
rect 4056 14359 4068 14368
rect 3344 14328 3372 14359
rect 4062 14356 4068 14359
rect 4120 14356 4126 14408
rect 5626 14396 5632 14408
rect 5587 14368 5632 14396
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 5812 14399 5870 14405
rect 5812 14365 5824 14399
rect 5858 14396 5870 14399
rect 5997 14399 6055 14405
rect 5858 14368 5948 14396
rect 5858 14365 5870 14368
rect 5812 14359 5870 14365
rect 3510 14328 3516 14340
rect 3344 14300 3516 14328
rect 3510 14288 3516 14300
rect 3568 14328 3574 14340
rect 5644 14328 5672 14356
rect 5920 14340 5948 14368
rect 5997 14365 6009 14399
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 3568 14300 5672 14328
rect 3568 14288 3574 14300
rect 5902 14288 5908 14340
rect 5960 14288 5966 14340
rect 6012 14328 6040 14359
rect 6178 14356 6184 14408
rect 6236 14396 6242 14408
rect 6380 14396 6408 14572
rect 6638 14532 6644 14544
rect 6564 14504 6644 14532
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6236 14368 6281 14396
rect 6380 14368 6469 14396
rect 6236 14356 6242 14368
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 6564 14328 6592 14504
rect 6638 14492 6644 14504
rect 6696 14532 6702 14544
rect 6933 14532 6961 14572
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 7101 14603 7159 14609
rect 7101 14600 7113 14603
rect 7064 14572 7113 14600
rect 7064 14560 7070 14572
rect 7101 14569 7113 14572
rect 7147 14569 7159 14603
rect 7282 14600 7288 14612
rect 7243 14572 7288 14600
rect 7101 14563 7159 14569
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 8110 14600 8116 14612
rect 7432 14572 8116 14600
rect 7432 14560 7438 14572
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 8386 14560 8392 14612
rect 8444 14600 8450 14612
rect 8662 14600 8668 14612
rect 8444 14572 8668 14600
rect 8444 14560 8450 14572
rect 8662 14560 8668 14572
rect 8720 14600 8726 14612
rect 8720 14572 9260 14600
rect 8720 14560 8726 14572
rect 7190 14532 7196 14544
rect 6696 14504 6868 14532
rect 6933 14504 7196 14532
rect 6696 14492 6702 14504
rect 6730 14464 6736 14476
rect 6691 14436 6736 14464
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 6840 14473 6868 14504
rect 7190 14492 7196 14504
rect 7248 14492 7254 14544
rect 8588 14504 8984 14532
rect 6825 14467 6883 14473
rect 6825 14433 6837 14467
rect 6871 14433 6883 14467
rect 6825 14427 6883 14433
rect 7098 14424 7104 14476
rect 7156 14464 7162 14476
rect 7745 14467 7803 14473
rect 7745 14464 7757 14467
rect 7156 14436 7757 14464
rect 7156 14424 7162 14436
rect 7745 14433 7757 14436
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 7834 14424 7840 14476
rect 7892 14464 7898 14476
rect 7892 14436 7937 14464
rect 7892 14424 7898 14436
rect 6640 14399 6698 14405
rect 6640 14365 6652 14399
rect 6686 14396 6698 14399
rect 7009 14399 7067 14405
rect 6686 14368 6961 14396
rect 6686 14365 6698 14368
rect 6640 14359 6698 14365
rect 6012 14300 6592 14328
rect 6933 14328 6961 14368
rect 7009 14365 7021 14399
rect 7055 14396 7067 14399
rect 8018 14396 8024 14408
rect 7055 14368 8024 14396
rect 7055 14365 7067 14368
rect 7009 14359 7067 14365
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 8588 14405 8616 14504
rect 8754 14405 8760 14408
rect 8573 14399 8631 14405
rect 8573 14396 8585 14399
rect 8168 14368 8585 14396
rect 8168 14356 8174 14368
rect 8573 14365 8585 14368
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 8751 14359 8760 14405
rect 8812 14396 8818 14408
rect 8956 14405 8984 14504
rect 9232 14405 9260 14572
rect 11054 14560 11060 14612
rect 11112 14600 11118 14612
rect 11425 14603 11483 14609
rect 11425 14600 11437 14603
rect 11112 14572 11437 14600
rect 11112 14560 11118 14572
rect 11425 14569 11437 14572
rect 11471 14569 11483 14603
rect 11425 14563 11483 14569
rect 12176 14572 13768 14600
rect 11146 14464 11152 14476
rect 9324 14436 11152 14464
rect 8941 14399 8999 14405
rect 8812 14368 8851 14396
rect 8754 14356 8760 14359
rect 8812 14356 8818 14368
rect 8941 14365 8953 14399
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 7282 14328 7288 14340
rect 6933 14300 7288 14328
rect 7282 14288 7288 14300
rect 7340 14288 7346 14340
rect 7653 14331 7711 14337
rect 7653 14297 7665 14331
rect 7699 14328 7711 14331
rect 8202 14328 8208 14340
rect 7699 14300 8208 14328
rect 7699 14297 7711 14300
rect 7653 14291 7711 14297
rect 8202 14288 8208 14300
rect 8260 14288 8266 14340
rect 9324 14328 9352 14436
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 11440 14464 11468 14563
rect 11974 14464 11980 14476
rect 11440 14436 11744 14464
rect 11935 14436 11980 14464
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14365 9459 14399
rect 11606 14396 11612 14408
rect 11567 14368 11612 14396
rect 9401 14359 9459 14365
rect 8312 14300 9352 14328
rect 2682 14260 2688 14272
rect 2643 14232 2688 14260
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 3418 14220 3424 14272
rect 3476 14260 3482 14272
rect 8312 14260 8340 14300
rect 3476 14232 8340 14260
rect 8389 14263 8447 14269
rect 3476 14220 3482 14232
rect 8389 14229 8401 14263
rect 8435 14260 8447 14263
rect 8662 14260 8668 14272
rect 8435 14232 8668 14260
rect 8435 14229 8447 14232
rect 8389 14223 8447 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 8846 14220 8852 14272
rect 8904 14260 8910 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8904 14232 9045 14260
rect 8904 14220 8910 14232
rect 9033 14229 9045 14232
rect 9079 14229 9091 14263
rect 9416 14260 9444 14359
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 11716 14396 11744 14436
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 11774 14399 11832 14405
rect 11774 14396 11786 14399
rect 11716 14368 11786 14396
rect 11774 14365 11786 14368
rect 11820 14365 11832 14399
rect 11774 14359 11832 14365
rect 11882 14356 11888 14408
rect 11940 14396 11946 14408
rect 12176 14405 12204 14572
rect 13740 14532 13768 14572
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14274 14600 14280 14612
rect 13872 14572 14280 14600
rect 13872 14560 13878 14572
rect 14274 14560 14280 14572
rect 14332 14560 14338 14612
rect 14829 14603 14887 14609
rect 14829 14569 14841 14603
rect 14875 14600 14887 14603
rect 15102 14600 15108 14612
rect 14875 14572 15108 14600
rect 14875 14569 14887 14572
rect 14829 14563 14887 14569
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 16022 14560 16028 14612
rect 16080 14600 16086 14612
rect 16485 14603 16543 14609
rect 16080 14572 16252 14600
rect 16080 14560 16086 14572
rect 14093 14535 14151 14541
rect 14093 14532 14105 14535
rect 13740 14504 14105 14532
rect 14093 14501 14105 14504
rect 14139 14501 14151 14535
rect 14093 14495 14151 14501
rect 14476 14504 15332 14532
rect 14476 14476 14504 14504
rect 14458 14464 14464 14476
rect 14419 14436 14464 14464
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 14642 14464 14648 14476
rect 14599 14436 14648 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 15304 14473 15332 14504
rect 15930 14492 15936 14544
rect 15988 14532 15994 14544
rect 15988 14504 16160 14532
rect 15988 14492 15994 14504
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 15436 14436 15481 14464
rect 15436 14424 15442 14436
rect 15654 14424 15660 14476
rect 15712 14464 15718 14476
rect 16132 14473 16160 14504
rect 16224 14473 16252 14572
rect 16485 14569 16497 14603
rect 16531 14600 16543 14603
rect 16758 14600 16764 14612
rect 16531 14572 16764 14600
rect 16531 14569 16543 14572
rect 16485 14563 16543 14569
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 19426 14560 19432 14612
rect 19484 14600 19490 14612
rect 21082 14600 21088 14612
rect 19484 14572 21088 14600
rect 19484 14560 19490 14572
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 18690 14532 18696 14544
rect 18651 14504 18696 14532
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 20165 14535 20223 14541
rect 20165 14501 20177 14535
rect 20211 14532 20223 14535
rect 20806 14532 20812 14544
rect 20211 14504 20812 14532
rect 20211 14501 20223 14504
rect 20165 14495 20223 14501
rect 20806 14492 20812 14504
rect 20864 14492 20870 14544
rect 23290 14492 23296 14544
rect 23348 14532 23354 14544
rect 23348 14504 24440 14532
rect 23348 14492 23354 14504
rect 15749 14467 15807 14473
rect 15749 14464 15761 14467
rect 15712 14436 15761 14464
rect 15712 14424 15718 14436
rect 15749 14433 15761 14436
rect 15795 14433 15807 14467
rect 15749 14427 15807 14433
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 16209 14467 16267 14473
rect 16209 14433 16221 14467
rect 16255 14433 16267 14467
rect 16209 14427 16267 14433
rect 18141 14467 18199 14473
rect 18141 14433 18153 14467
rect 18187 14464 18199 14467
rect 18322 14464 18328 14476
rect 18187 14436 18328 14464
rect 18187 14433 18199 14436
rect 18141 14427 18199 14433
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 19610 14464 19616 14476
rect 19571 14436 19616 14464
rect 19610 14424 19616 14436
rect 19668 14424 19674 14476
rect 20254 14424 20260 14476
rect 20312 14464 20318 14476
rect 20625 14467 20683 14473
rect 20625 14464 20637 14467
rect 20312 14436 20637 14464
rect 20312 14424 20318 14436
rect 20625 14433 20637 14436
rect 20671 14433 20683 14467
rect 20625 14427 20683 14433
rect 23014 14424 23020 14476
rect 23072 14464 23078 14476
rect 23658 14464 23664 14476
rect 23072 14436 23664 14464
rect 23072 14424 23078 14436
rect 23658 14424 23664 14436
rect 23716 14464 23722 14476
rect 24210 14464 24216 14476
rect 23716 14436 23888 14464
rect 24171 14436 24216 14464
rect 23716 14424 23722 14436
rect 12161 14399 12219 14405
rect 11940 14368 11985 14396
rect 11940 14356 11946 14368
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 12437 14399 12495 14405
rect 12437 14365 12449 14399
rect 12483 14396 12495 14399
rect 13078 14396 13084 14408
rect 12483 14368 13084 14396
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 14090 14396 14096 14408
rect 13372 14368 14096 14396
rect 9769 14263 9827 14269
rect 9769 14260 9781 14263
rect 9416 14232 9781 14260
rect 9033 14223 9091 14229
rect 9769 14229 9781 14232
rect 9815 14260 9827 14263
rect 10778 14260 10784 14272
rect 9815 14232 10784 14260
rect 9815 14229 9827 14232
rect 9769 14223 9827 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 11624 14260 11652 14356
rect 12345 14331 12403 14337
rect 12345 14297 12357 14331
rect 12391 14328 12403 14331
rect 12682 14331 12740 14337
rect 12682 14328 12694 14331
rect 12391 14300 12694 14328
rect 12391 14297 12403 14300
rect 12345 14291 12403 14297
rect 12682 14297 12694 14300
rect 12728 14297 12740 14331
rect 12682 14291 12740 14297
rect 13372 14260 13400 14368
rect 14090 14356 14096 14368
rect 14148 14396 14154 14408
rect 14185 14399 14243 14405
rect 14185 14396 14197 14399
rect 14148 14368 14197 14396
rect 14148 14356 14154 14368
rect 14185 14365 14197 14368
rect 14231 14365 14243 14399
rect 14185 14359 14243 14365
rect 14200 14328 14228 14359
rect 14274 14356 14280 14408
rect 14332 14396 14338 14408
rect 14368 14399 14426 14405
rect 14368 14396 14380 14399
rect 14332 14368 14380 14396
rect 14332 14356 14338 14368
rect 14368 14365 14380 14368
rect 14414 14365 14426 14399
rect 14368 14359 14426 14365
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14396 14795 14399
rect 14918 14396 14924 14408
rect 14783 14368 14924 14396
rect 14783 14365 14795 14368
rect 14737 14359 14795 14365
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 15028 14328 15056 14359
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 15562 14396 15568 14408
rect 15252 14368 15424 14396
rect 15523 14368 15568 14396
rect 15252 14356 15258 14368
rect 14200 14300 15056 14328
rect 15396 14328 15424 14368
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 15838 14396 15844 14408
rect 15799 14368 15844 14396
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 16024 14399 16082 14405
rect 16024 14365 16036 14399
rect 16070 14396 16082 14399
rect 16393 14399 16451 14405
rect 16070 14368 16344 14396
rect 16070 14365 16082 14368
rect 16024 14359 16082 14365
rect 15930 14328 15936 14340
rect 15396 14300 15936 14328
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 16316 14328 16344 14368
rect 16393 14365 16405 14399
rect 16439 14396 16451 14399
rect 17954 14396 17960 14408
rect 16439 14368 17960 14396
rect 16439 14365 16451 14368
rect 16393 14359 16451 14365
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14365 18107 14399
rect 18049 14359 18107 14365
rect 16482 14328 16488 14340
rect 16316 14300 16488 14328
rect 16482 14288 16488 14300
rect 16540 14288 16546 14340
rect 18064 14328 18092 14359
rect 18230 14356 18236 14408
rect 18288 14396 18294 14408
rect 18451 14399 18509 14405
rect 18451 14396 18463 14399
rect 18288 14368 18463 14396
rect 18288 14356 18294 14368
rect 18451 14365 18463 14368
rect 18497 14365 18509 14399
rect 18451 14359 18509 14365
rect 19797 14399 19855 14405
rect 19797 14365 19809 14399
rect 19843 14396 19855 14399
rect 20070 14396 20076 14408
rect 19843 14368 20076 14396
rect 19843 14365 19855 14368
rect 19797 14359 19855 14365
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20438 14396 20444 14408
rect 20399 14368 20444 14396
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 23477 14399 23535 14405
rect 23477 14365 23489 14399
rect 23523 14365 23535 14399
rect 23477 14359 23535 14365
rect 18598 14328 18604 14340
rect 18064 14300 18604 14328
rect 18598 14288 18604 14300
rect 18656 14328 18662 14340
rect 19242 14328 19248 14340
rect 18656 14300 19248 14328
rect 18656 14288 18662 14300
rect 19242 14288 19248 14300
rect 19300 14328 19306 14340
rect 19429 14331 19487 14337
rect 19429 14328 19441 14331
rect 19300 14300 19441 14328
rect 19300 14288 19306 14300
rect 19429 14297 19441 14300
rect 19475 14297 19487 14331
rect 19429 14291 19487 14297
rect 19521 14331 19579 14337
rect 19521 14297 19533 14331
rect 19567 14328 19579 14331
rect 19702 14328 19708 14340
rect 19567 14300 19708 14328
rect 19567 14297 19579 14300
rect 19521 14291 19579 14297
rect 19702 14288 19708 14300
rect 19760 14288 19766 14340
rect 23492 14328 23520 14359
rect 23566 14356 23572 14408
rect 23624 14396 23630 14408
rect 23860 14405 23888 14436
rect 24210 14424 24216 14436
rect 24268 14424 24274 14476
rect 23845 14399 23903 14405
rect 23624 14368 23669 14396
rect 23624 14356 23630 14368
rect 23845 14365 23857 14399
rect 23891 14365 23903 14399
rect 23845 14359 23903 14365
rect 24121 14399 24179 14405
rect 24121 14365 24133 14399
rect 24167 14396 24179 14399
rect 24302 14396 24308 14408
rect 24167 14368 24308 14396
rect 24167 14365 24179 14368
rect 24121 14359 24179 14365
rect 24302 14356 24308 14368
rect 24360 14356 24366 14408
rect 24412 14405 24440 14504
rect 24397 14399 24455 14405
rect 24397 14365 24409 14399
rect 24443 14365 24455 14399
rect 24397 14359 24455 14365
rect 23750 14328 23756 14340
rect 23492 14300 23756 14328
rect 23750 14288 23756 14300
rect 23808 14288 23814 14340
rect 11624 14232 13400 14260
rect 13817 14263 13875 14269
rect 13817 14229 13829 14263
rect 13863 14260 13875 14263
rect 13998 14260 14004 14272
rect 13863 14232 14004 14260
rect 13863 14229 13875 14232
rect 13817 14223 13875 14229
rect 13998 14220 14004 14232
rect 14056 14260 14062 14272
rect 14093 14263 14151 14269
rect 14093 14260 14105 14263
rect 14056 14232 14105 14260
rect 14056 14220 14062 14232
rect 14093 14229 14105 14232
rect 14139 14229 14151 14263
rect 14093 14223 14151 14229
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 15010 14260 15016 14272
rect 14332 14232 15016 14260
rect 14332 14220 14338 14232
rect 15010 14220 15016 14232
rect 15068 14260 15074 14272
rect 16669 14263 16727 14269
rect 16669 14260 16681 14263
rect 15068 14232 16681 14260
rect 15068 14220 15074 14232
rect 16669 14229 16681 14232
rect 16715 14229 16727 14263
rect 16669 14223 16727 14229
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 20806 14260 20812 14272
rect 17460 14232 20812 14260
rect 17460 14220 17466 14232
rect 20806 14220 20812 14232
rect 20864 14260 20870 14272
rect 21174 14260 21180 14272
rect 20864 14232 21180 14260
rect 20864 14220 20870 14232
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 23198 14220 23204 14272
rect 23256 14260 23262 14272
rect 23385 14263 23443 14269
rect 23385 14260 23397 14263
rect 23256 14232 23397 14260
rect 23256 14220 23262 14232
rect 23385 14229 23397 14232
rect 23431 14229 23443 14263
rect 23385 14223 23443 14229
rect 24489 14263 24547 14269
rect 24489 14229 24501 14263
rect 24535 14260 24547 14263
rect 24670 14260 24676 14272
rect 24535 14232 24676 14260
rect 24535 14229 24547 14232
rect 24489 14223 24547 14229
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 1104 14170 26128 14192
rect 1104 14118 9291 14170
rect 9343 14118 9355 14170
rect 9407 14118 9419 14170
rect 9471 14118 9483 14170
rect 9535 14118 9547 14170
rect 9599 14118 17632 14170
rect 17684 14118 17696 14170
rect 17748 14118 17760 14170
rect 17812 14118 17824 14170
rect 17876 14118 17888 14170
rect 17940 14118 26128 14170
rect 1104 14096 26128 14118
rect 2958 14016 2964 14068
rect 3016 14056 3022 14068
rect 3016 14028 3188 14056
rect 3016 14016 3022 14028
rect 3160 13988 3188 14028
rect 3602 14016 3608 14068
rect 3660 14056 3666 14068
rect 3697 14059 3755 14065
rect 3697 14056 3709 14059
rect 3660 14028 3709 14056
rect 3660 14016 3666 14028
rect 3697 14025 3709 14028
rect 3743 14025 3755 14059
rect 3697 14019 3755 14025
rect 3786 14016 3792 14068
rect 3844 14056 3850 14068
rect 4801 14059 4859 14065
rect 4801 14056 4813 14059
rect 3844 14028 4813 14056
rect 3844 14016 3850 14028
rect 4801 14025 4813 14028
rect 4847 14025 4859 14059
rect 4801 14019 4859 14025
rect 5445 14059 5503 14065
rect 5445 14025 5457 14059
rect 5491 14056 5503 14059
rect 5626 14056 5632 14068
rect 5491 14028 5632 14056
rect 5491 14025 5503 14028
rect 5445 14019 5503 14025
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 5902 14056 5908 14068
rect 5863 14028 5908 14056
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 5994 14016 6000 14068
rect 6052 14056 6058 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 6052 14028 6377 14056
rect 6052 14016 6058 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 6822 14056 6828 14068
rect 6783 14028 6828 14056
rect 6365 14019 6423 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 7650 14056 7656 14068
rect 7611 14028 7656 14056
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 8110 14056 8116 14068
rect 8071 14028 8116 14056
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 11146 14056 11152 14068
rect 11107 14028 11152 14056
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 11882 14056 11888 14068
rect 11664 14028 11888 14056
rect 11664 14016 11670 14028
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 12250 14016 12256 14068
rect 12308 14056 12314 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12308 14028 12909 14056
rect 12308 14016 12314 14028
rect 12897 14025 12909 14028
rect 12943 14056 12955 14059
rect 12986 14056 12992 14068
rect 12943 14028 12992 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 14829 14059 14887 14065
rect 14829 14025 14841 14059
rect 14875 14056 14887 14059
rect 15194 14056 15200 14068
rect 14875 14028 15200 14056
rect 14875 14025 14887 14028
rect 14829 14019 14887 14025
rect 15194 14016 15200 14028
rect 15252 14056 15258 14068
rect 15838 14056 15844 14068
rect 15252 14028 15844 14056
rect 15252 14016 15258 14028
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 16393 14059 16451 14065
rect 16393 14056 16405 14059
rect 16316 14028 16405 14056
rect 3804 13988 3832 14016
rect 3160 13960 3832 13988
rect 4065 13991 4123 13997
rect 2958 13920 2964 13932
rect 2919 13892 2964 13920
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3160 13929 3188 13960
rect 4065 13957 4077 13991
rect 4111 13988 4123 13991
rect 4890 13988 4896 14000
rect 4111 13960 4896 13988
rect 4111 13957 4123 13960
rect 4065 13951 4123 13957
rect 4890 13948 4896 13960
rect 4948 13948 4954 14000
rect 8205 13991 8263 13997
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13889 3203 13923
rect 3326 13920 3332 13932
rect 3288 13892 3332 13920
rect 3145 13883 3203 13889
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 3510 13920 3516 13932
rect 3471 13892 3516 13920
rect 3510 13880 3516 13892
rect 3568 13880 3574 13932
rect 3694 13880 3700 13932
rect 3752 13920 3758 13932
rect 4157 13923 4215 13929
rect 4157 13920 4169 13923
rect 3752 13892 4169 13920
rect 3752 13880 3758 13892
rect 4157 13889 4169 13892
rect 4203 13889 4215 13923
rect 4706 13920 4712 13932
rect 4667 13892 4712 13920
rect 4157 13883 4215 13889
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 5718 13929 5724 13958
rect 4985 13923 5043 13929
rect 4985 13889 4997 13923
rect 5031 13920 5043 13923
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 5031 13892 5089 13920
rect 5031 13889 5043 13892
rect 4985 13883 5043 13889
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5620 13923 5678 13929
rect 5620 13889 5632 13923
rect 5666 13889 5678 13923
rect 5620 13883 5678 13889
rect 5713 13906 5724 13929
rect 5776 13906 5782 13958
rect 8205 13957 8217 13991
rect 8251 13988 8263 13991
rect 8386 13988 8392 14000
rect 8251 13960 8392 13988
rect 8251 13957 8263 13960
rect 8205 13951 8263 13957
rect 8386 13948 8392 13960
rect 8444 13948 8450 14000
rect 9214 13948 9220 14000
rect 9272 13988 9278 14000
rect 9272 13960 9444 13988
rect 9272 13948 9278 13960
rect 5997 13923 6055 13929
rect 5997 13920 6009 13923
rect 5713 13889 5725 13906
rect 5759 13889 5771 13906
rect 5911 13904 6009 13920
rect 5713 13883 5771 13889
rect 5828 13892 6009 13904
rect 3050 13812 3056 13864
rect 3108 13852 3114 13864
rect 3237 13855 3295 13861
rect 3237 13852 3249 13855
rect 3108 13824 3249 13852
rect 3108 13812 3114 13824
rect 3237 13821 3249 13824
rect 3283 13852 3295 13855
rect 4338 13852 4344 13864
rect 3283 13824 4200 13852
rect 4299 13824 4344 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 4172 13796 4200 13824
rect 4338 13812 4344 13824
rect 4396 13852 4402 13864
rect 4522 13852 4528 13864
rect 4396 13824 4528 13852
rect 4396 13812 4402 13824
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 5000 13852 5028 13883
rect 4663 13824 5028 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 2774 13744 2780 13796
rect 2832 13784 2838 13796
rect 2832 13756 2877 13784
rect 2832 13744 2838 13756
rect 4154 13744 4160 13796
rect 4212 13744 4218 13796
rect 5261 13787 5319 13793
rect 5261 13753 5273 13787
rect 5307 13784 5319 13787
rect 5442 13784 5448 13796
rect 5307 13756 5448 13784
rect 5307 13753 5319 13756
rect 5261 13747 5319 13753
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 5635 13716 5663 13883
rect 5828 13876 5939 13892
rect 5997 13889 6009 13892
rect 6043 13920 6055 13923
rect 6546 13920 6552 13932
rect 6043 13892 6552 13920
rect 6043 13889 6055 13892
rect 5997 13883 6055 13889
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 7282 13920 7288 13932
rect 6779 13892 7288 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 7282 13880 7288 13892
rect 7340 13880 7346 13932
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 8294 13920 8300 13932
rect 7607 13892 8300 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 8662 13920 8668 13932
rect 8623 13892 8668 13920
rect 8662 13880 8668 13892
rect 8720 13880 8726 13932
rect 8846 13920 8852 13932
rect 8772 13892 8852 13920
rect 5828 13716 5856 13876
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 7650 13852 7656 13864
rect 6972 13824 7656 13852
rect 6972 13812 6978 13824
rect 7650 13812 7656 13824
rect 7708 13852 7714 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7708 13824 7757 13852
rect 7708 13812 7714 13824
rect 7745 13821 7757 13824
rect 7791 13852 7803 13855
rect 7834 13852 7840 13864
rect 7791 13824 7840 13852
rect 7791 13821 7803 13824
rect 7745 13815 7803 13821
rect 7834 13812 7840 13824
rect 7892 13852 7898 13864
rect 8772 13852 8800 13892
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9125 13923 9183 13929
rect 9125 13889 9137 13923
rect 9171 13889 9183 13923
rect 9125 13883 9183 13889
rect 9309 13923 9367 13929
rect 9309 13889 9321 13923
rect 9355 13918 9367 13923
rect 9416 13918 9444 13960
rect 9674 13948 9680 14000
rect 9732 13988 9738 14000
rect 9769 13991 9827 13997
rect 9769 13988 9781 13991
rect 9732 13960 9781 13988
rect 9732 13948 9738 13960
rect 9769 13957 9781 13960
rect 9815 13957 9827 13991
rect 14090 13988 14096 14000
rect 9769 13951 9827 13957
rect 13096 13960 14096 13988
rect 13096 13932 13124 13960
rect 14090 13948 14096 13960
rect 14148 13988 14154 14000
rect 15280 13991 15338 13997
rect 14148 13960 15056 13988
rect 14148 13948 14154 13960
rect 9355 13890 9444 13918
rect 9585 13923 9643 13929
rect 9355 13889 9367 13890
rect 9309 13883 9367 13889
rect 9585 13889 9597 13923
rect 9631 13920 9643 13923
rect 9950 13920 9956 13932
rect 9631 13892 9956 13920
rect 9631 13889 9643 13892
rect 9585 13883 9643 13889
rect 8938 13852 8944 13864
rect 7892 13824 8800 13852
rect 8899 13824 8944 13852
rect 7892 13812 7898 13824
rect 8938 13812 8944 13824
rect 8996 13812 9002 13864
rect 9140 13852 9168 13883
rect 9600 13852 9628 13883
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 11790 13929 11796 13932
rect 11784 13883 11796 13929
rect 11848 13920 11854 13932
rect 13078 13920 13084 13932
rect 11848 13892 11884 13920
rect 13039 13892 13084 13920
rect 11790 13880 11796 13883
rect 11848 13880 11854 13892
rect 13078 13880 13084 13892
rect 13136 13880 13142 13932
rect 13170 13880 13176 13932
rect 13228 13920 13234 13932
rect 13337 13923 13395 13929
rect 13337 13920 13349 13923
rect 13228 13892 13349 13920
rect 13228 13880 13234 13892
rect 13337 13889 13349 13892
rect 13383 13889 13395 13923
rect 13337 13883 13395 13889
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13920 14703 13923
rect 14734 13920 14740 13932
rect 14691 13892 14740 13920
rect 14691 13889 14703 13892
rect 14645 13883 14703 13889
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 15028 13929 15056 13960
rect 15280 13957 15292 13991
rect 15326 13988 15338 13991
rect 15654 13988 15660 14000
rect 15326 13960 15660 13988
rect 15326 13957 15338 13960
rect 15280 13951 15338 13957
rect 15654 13948 15660 13960
rect 15712 13948 15718 14000
rect 16316 13988 16344 14028
rect 16393 14025 16405 14028
rect 16439 14025 16451 14059
rect 16393 14019 16451 14025
rect 16482 14016 16488 14068
rect 16540 14056 16546 14068
rect 17218 14056 17224 14068
rect 16540 14028 17224 14056
rect 16540 14016 16546 14028
rect 17218 14016 17224 14028
rect 17276 14056 17282 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17276 14028 17785 14056
rect 17276 14016 17282 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 18322 14016 18328 14068
rect 18380 14056 18386 14068
rect 18601 14059 18659 14065
rect 18601 14056 18613 14059
rect 18380 14028 18613 14056
rect 18380 14016 18386 14028
rect 18601 14025 18613 14028
rect 18647 14025 18659 14059
rect 19058 14056 19064 14068
rect 19019 14028 19064 14056
rect 18601 14019 18659 14025
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 19705 14059 19763 14065
rect 19705 14056 19717 14059
rect 19300 14028 19717 14056
rect 19300 14016 19306 14028
rect 19705 14025 19717 14028
rect 19751 14025 19763 14059
rect 19705 14019 19763 14025
rect 20070 14016 20076 14068
rect 20128 14056 20134 14068
rect 20257 14059 20315 14065
rect 20257 14056 20269 14059
rect 20128 14028 20269 14056
rect 20128 14016 20134 14028
rect 20257 14025 20269 14028
rect 20303 14025 20315 14059
rect 23290 14056 23296 14068
rect 23251 14028 23296 14056
rect 20257 14019 20315 14025
rect 23290 14016 23296 14028
rect 23348 14016 23354 14068
rect 24397 14059 24455 14065
rect 24397 14025 24409 14059
rect 24443 14056 24455 14059
rect 24578 14056 24584 14068
rect 24443 14028 24584 14056
rect 24443 14025 24455 14028
rect 24397 14019 24455 14025
rect 24578 14016 24584 14028
rect 24636 14016 24642 14068
rect 16316 13960 19564 13988
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 15562 13880 15568 13932
rect 15620 13920 15626 13932
rect 16316 13920 16344 13960
rect 15620 13892 16344 13920
rect 15620 13880 15626 13892
rect 17586 13880 17592 13932
rect 17644 13920 17650 13932
rect 17681 13923 17739 13929
rect 17681 13920 17693 13923
rect 17644 13892 17693 13920
rect 17644 13880 17650 13892
rect 17681 13889 17693 13892
rect 17727 13889 17739 13923
rect 17681 13883 17739 13889
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18509 13923 18567 13929
rect 18509 13920 18521 13923
rect 18472 13892 18521 13920
rect 18472 13880 18478 13892
rect 18509 13889 18521 13892
rect 18555 13889 18567 13923
rect 19058 13920 19064 13932
rect 19019 13892 19064 13920
rect 18509 13883 18567 13889
rect 19058 13880 19064 13892
rect 19116 13880 19122 13932
rect 19337 13923 19395 13929
rect 19337 13889 19349 13923
rect 19383 13920 19395 13923
rect 19426 13920 19432 13932
rect 19383 13892 19432 13920
rect 19383 13889 19395 13892
rect 19337 13883 19395 13889
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 11514 13852 11520 13864
rect 9140 13824 9628 13852
rect 11475 13824 11520 13852
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 17402 13852 17408 13864
rect 14108 13824 15056 13852
rect 8757 13787 8815 13793
rect 8757 13753 8769 13787
rect 8803 13784 8815 13787
rect 9306 13784 9312 13796
rect 8803 13756 9312 13784
rect 8803 13753 8815 13756
rect 8757 13747 8815 13753
rect 9306 13744 9312 13756
rect 9364 13744 9370 13796
rect 9401 13787 9459 13793
rect 9401 13753 9413 13787
rect 9447 13784 9459 13787
rect 9582 13784 9588 13796
rect 9447 13756 9588 13784
rect 9447 13753 9459 13756
rect 9401 13747 9459 13753
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 14108 13784 14136 13824
rect 14016 13756 14136 13784
rect 14016 13728 14044 13756
rect 6178 13716 6184 13728
rect 5635 13688 5856 13716
rect 6139 13688 6184 13716
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 6972 13688 7205 13716
rect 6972 13676 6978 13688
rect 7193 13685 7205 13688
rect 7239 13685 7251 13719
rect 9950 13716 9956 13728
rect 9911 13688 9956 13716
rect 7193 13679 7251 13685
rect 9950 13676 9956 13688
rect 10008 13716 10014 13728
rect 10045 13719 10103 13725
rect 10045 13716 10057 13719
rect 10008 13688 10057 13716
rect 10008 13676 10014 13688
rect 10045 13685 10057 13688
rect 10091 13716 10103 13719
rect 10229 13719 10287 13725
rect 10229 13716 10241 13719
rect 10091 13688 10241 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 10229 13685 10241 13688
rect 10275 13685 10287 13719
rect 10229 13679 10287 13685
rect 13998 13676 14004 13728
rect 14056 13676 14062 13728
rect 14461 13719 14519 13725
rect 14461 13685 14473 13719
rect 14507 13716 14519 13719
rect 14550 13716 14556 13728
rect 14507 13688 14556 13716
rect 14507 13685 14519 13688
rect 14461 13679 14519 13685
rect 14550 13676 14556 13688
rect 14608 13676 14614 13728
rect 15028 13716 15056 13824
rect 16040 13824 17408 13852
rect 16040 13784 16068 13824
rect 17402 13812 17408 13824
rect 17460 13812 17466 13864
rect 17865 13855 17923 13861
rect 17865 13821 17877 13855
rect 17911 13821 17923 13855
rect 17865 13815 17923 13821
rect 18693 13855 18751 13861
rect 18693 13821 18705 13855
rect 18739 13821 18751 13855
rect 18693 13815 18751 13821
rect 19536 13852 19564 13960
rect 19978 13948 19984 14000
rect 20036 13988 20042 14000
rect 20036 13960 23336 13988
rect 20036 13948 20042 13960
rect 19610 13880 19616 13932
rect 19668 13920 19674 13932
rect 19889 13923 19947 13929
rect 19889 13920 19901 13923
rect 19668 13892 19901 13920
rect 19668 13880 19674 13892
rect 19889 13889 19901 13892
rect 19935 13889 19947 13923
rect 19889 13883 19947 13889
rect 20073 13923 20131 13929
rect 20073 13889 20085 13923
rect 20119 13920 20131 13923
rect 20346 13920 20352 13932
rect 20119 13892 20352 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 20438 13880 20444 13932
rect 20496 13920 20502 13932
rect 20806 13920 20812 13932
rect 20496 13892 20589 13920
rect 20767 13892 20812 13920
rect 20496 13880 20502 13892
rect 20806 13880 20812 13892
rect 20864 13880 20870 13932
rect 21091 13929 21119 13960
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 21174 13880 21180 13932
rect 21232 13920 21238 13932
rect 21269 13923 21327 13929
rect 21269 13920 21281 13923
rect 21232 13892 21281 13920
rect 21232 13880 21238 13892
rect 21269 13889 21281 13892
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 21358 13880 21364 13932
rect 21416 13920 21422 13932
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 21416 13892 21833 13920
rect 21416 13880 21422 13892
rect 21821 13889 21833 13892
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 22189 13923 22247 13929
rect 22189 13889 22201 13923
rect 22235 13920 22247 13923
rect 23198 13920 23204 13932
rect 22235 13892 23204 13920
rect 22235 13889 22247 13892
rect 22189 13883 22247 13889
rect 23198 13880 23204 13892
rect 23256 13880 23262 13932
rect 23308 13920 23336 13960
rect 23658 13948 23664 14000
rect 23716 13988 23722 14000
rect 23716 13960 24164 13988
rect 23716 13948 23722 13960
rect 23566 13920 23572 13932
rect 23308 13892 23572 13920
rect 23566 13880 23572 13892
rect 23624 13880 23630 13932
rect 23842 13880 23848 13932
rect 23900 13920 23906 13932
rect 24136 13929 24164 13960
rect 23937 13923 23995 13929
rect 23937 13920 23949 13923
rect 23900 13892 23949 13920
rect 23900 13880 23906 13892
rect 23937 13889 23949 13892
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 24121 13923 24179 13929
rect 24121 13889 24133 13923
rect 24167 13889 24179 13923
rect 24302 13920 24308 13932
rect 24263 13892 24308 13920
rect 24121 13883 24179 13889
rect 24302 13880 24308 13892
rect 24360 13880 24366 13932
rect 20456 13852 20484 13880
rect 19536 13824 20484 13852
rect 20901 13855 20959 13861
rect 15948 13756 16068 13784
rect 17037 13787 17095 13793
rect 15948 13716 15976 13756
rect 17037 13753 17049 13787
rect 17083 13784 17095 13787
rect 17218 13784 17224 13796
rect 17083 13756 17224 13784
rect 17083 13753 17095 13756
rect 17037 13747 17095 13753
rect 17218 13744 17224 13756
rect 17276 13784 17282 13796
rect 17880 13784 17908 13815
rect 18708 13784 18736 13815
rect 17276 13756 18736 13784
rect 17276 13744 17282 13756
rect 17310 13716 17316 13728
rect 15028 13688 15976 13716
rect 17271 13688 17316 13716
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 18138 13716 18144 13728
rect 18099 13688 18144 13716
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 19536 13716 19564 13824
rect 20901 13821 20913 13855
rect 20947 13852 20959 13855
rect 22005 13855 22063 13861
rect 22005 13852 22017 13855
rect 20947 13824 22017 13852
rect 20947 13821 20959 13824
rect 20901 13815 20959 13821
rect 22005 13821 22017 13824
rect 22051 13821 22063 13855
rect 23750 13852 23756 13864
rect 23711 13824 23756 13852
rect 22005 13815 22063 13821
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 21450 13784 21456 13796
rect 21411 13756 21456 13784
rect 21450 13744 21456 13756
rect 21508 13744 21514 13796
rect 22186 13784 22192 13796
rect 22147 13756 22192 13784
rect 22186 13744 22192 13756
rect 22244 13744 22250 13796
rect 23934 13784 23940 13796
rect 23895 13756 23940 13784
rect 23934 13744 23940 13756
rect 23992 13744 23998 13796
rect 19889 13719 19947 13725
rect 19889 13716 19901 13719
rect 19536 13688 19901 13716
rect 19889 13685 19901 13688
rect 19935 13685 19947 13719
rect 19889 13679 19947 13685
rect 23566 13676 23572 13728
rect 23624 13716 23630 13728
rect 24026 13716 24032 13728
rect 23624 13688 24032 13716
rect 23624 13676 23630 13688
rect 24026 13676 24032 13688
rect 24084 13676 24090 13728
rect 1104 13626 26128 13648
rect 1104 13574 5120 13626
rect 5172 13574 5184 13626
rect 5236 13574 5248 13626
rect 5300 13574 5312 13626
rect 5364 13574 5376 13626
rect 5428 13574 13462 13626
rect 13514 13574 13526 13626
rect 13578 13574 13590 13626
rect 13642 13574 13654 13626
rect 13706 13574 13718 13626
rect 13770 13574 21803 13626
rect 21855 13574 21867 13626
rect 21919 13574 21931 13626
rect 21983 13574 21995 13626
rect 22047 13574 22059 13626
rect 22111 13574 26128 13626
rect 1104 13552 26128 13574
rect 3142 13472 3148 13524
rect 3200 13512 3206 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3200 13484 3801 13512
rect 3200 13472 3206 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 3789 13475 3847 13481
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4617 13515 4675 13521
rect 4617 13512 4629 13515
rect 4212 13484 4629 13512
rect 4212 13472 4218 13484
rect 4617 13481 4629 13484
rect 4663 13481 4675 13515
rect 4617 13475 4675 13481
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 7098 13512 7104 13524
rect 6236 13484 7104 13512
rect 6236 13472 6242 13484
rect 7098 13472 7104 13484
rect 7156 13472 7162 13524
rect 8662 13472 8668 13524
rect 8720 13512 8726 13524
rect 8846 13512 8852 13524
rect 8720 13484 8852 13512
rect 8720 13472 8726 13484
rect 8846 13472 8852 13484
rect 8904 13512 8910 13524
rect 9769 13515 9827 13521
rect 8904 13484 9339 13512
rect 8904 13472 8910 13484
rect 7006 13444 7012 13456
rect 5460 13416 7012 13444
rect 3970 13336 3976 13388
rect 4028 13376 4034 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 4028 13348 4261 13376
rect 4028 13336 4034 13348
rect 4249 13345 4261 13348
rect 4295 13345 4307 13379
rect 4249 13339 4307 13345
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 4396 13348 4441 13376
rect 4396 13336 4402 13348
rect 1670 13268 1676 13320
rect 1728 13308 1734 13320
rect 2406 13308 2412 13320
rect 1728 13280 2412 13308
rect 1728 13268 1734 13280
rect 2406 13268 2412 13280
rect 2464 13308 2470 13320
rect 2961 13311 3019 13317
rect 2961 13308 2973 13311
rect 2464 13280 2973 13308
rect 2464 13268 2470 13280
rect 2961 13277 2973 13280
rect 3007 13308 3019 13311
rect 4706 13308 4712 13320
rect 3007 13280 4712 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 4798 13268 4804 13320
rect 4856 13308 4862 13320
rect 4856 13280 4901 13308
rect 4856 13268 4862 13280
rect 2682 13200 2688 13252
rect 2740 13249 2746 13252
rect 2740 13240 2752 13249
rect 4157 13243 4215 13249
rect 2740 13212 2785 13240
rect 2740 13203 2752 13212
rect 4157 13209 4169 13243
rect 4203 13240 4215 13243
rect 5460 13240 5488 13416
rect 7006 13404 7012 13416
rect 7064 13404 7070 13456
rect 8941 13447 8999 13453
rect 8941 13413 8953 13447
rect 8987 13444 8999 13447
rect 9030 13444 9036 13456
rect 8987 13416 9036 13444
rect 8987 13413 8999 13416
rect 8941 13407 8999 13413
rect 9030 13404 9036 13416
rect 9088 13444 9094 13456
rect 9214 13444 9220 13456
rect 9088 13416 9220 13444
rect 9088 13404 9094 13416
rect 9214 13404 9220 13416
rect 9272 13404 9278 13456
rect 5902 13376 5908 13388
rect 5863 13348 5908 13376
rect 5902 13336 5908 13348
rect 5960 13336 5966 13388
rect 7374 13376 7380 13388
rect 6472 13348 7380 13376
rect 5626 13308 5632 13320
rect 5587 13280 5632 13308
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 5810 13308 5816 13320
rect 5771 13280 5816 13308
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6015 13311 6073 13317
rect 6015 13277 6027 13311
rect 6061 13308 6073 13311
rect 6061 13280 6132 13308
rect 6061 13277 6073 13280
rect 6015 13271 6073 13277
rect 4203 13212 5488 13240
rect 6104 13240 6132 13280
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6472 13317 6500 13348
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 7650 13376 7656 13388
rect 7611 13348 7656 13376
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 9311 13376 9339 13484
rect 9769 13481 9781 13515
rect 9815 13481 9827 13515
rect 9769 13475 9827 13481
rect 9784 13376 9812 13475
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 11204 13484 11560 13512
rect 11204 13472 11210 13484
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 11112 13416 11468 13444
rect 11112 13404 11118 13416
rect 10870 13376 10876 13388
rect 9311 13348 9812 13376
rect 10831 13348 10876 13376
rect 6457 13311 6515 13317
rect 6236 13280 6281 13308
rect 6236 13268 6242 13280
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6638 13308 6644 13320
rect 6599 13280 6644 13308
rect 6457 13271 6515 13277
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 6914 13317 6920 13320
rect 6861 13311 6920 13317
rect 6788 13280 6833 13308
rect 6788 13268 6794 13280
rect 6861 13277 6873 13311
rect 6907 13277 6920 13311
rect 6861 13271 6920 13277
rect 6914 13268 6920 13271
rect 6972 13268 6978 13320
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 7098 13308 7104 13320
rect 7055 13280 7104 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 7742 13308 7748 13320
rect 7607 13280 7748 13308
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 7742 13268 7748 13280
rect 7800 13268 7806 13320
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 9311 13317 9339 13348
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 9183 13311 9241 13317
rect 9183 13308 9195 13311
rect 9088 13280 9195 13308
rect 9088 13268 9094 13280
rect 9183 13277 9195 13280
rect 9229 13277 9241 13311
rect 9183 13271 9241 13277
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9438 13311 9496 13317
rect 9438 13308 9450 13311
rect 9416 13298 9450 13308
rect 9309 13271 9367 13277
rect 7469 13243 7527 13249
rect 6104 13212 7144 13240
rect 4203 13209 4215 13212
rect 4157 13203 4215 13209
rect 2740 13200 2746 13203
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 2866 13172 2872 13184
rect 1627 13144 2872 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 2866 13132 2872 13144
rect 2924 13172 2930 13184
rect 3970 13172 3976 13184
rect 2924 13144 3976 13172
rect 2924 13132 2930 13144
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 5534 13172 5540 13184
rect 5495 13144 5540 13172
rect 5534 13132 5540 13144
rect 5592 13132 5598 13184
rect 6365 13175 6423 13181
rect 6365 13141 6377 13175
rect 6411 13172 6423 13175
rect 6454 13172 6460 13184
rect 6411 13144 6460 13172
rect 6411 13141 6423 13144
rect 6365 13135 6423 13141
rect 6454 13132 6460 13144
rect 6512 13132 6518 13184
rect 7116 13181 7144 13212
rect 7469 13209 7481 13243
rect 7515 13240 7527 13243
rect 8846 13240 8852 13252
rect 7515 13212 8852 13240
rect 7515 13209 7527 13212
rect 7469 13203 7527 13209
rect 8846 13200 8852 13212
rect 8904 13200 8910 13252
rect 9398 13246 9404 13298
rect 9484 13277 9496 13311
rect 9585 13311 9643 13317
rect 9585 13308 9597 13311
rect 9456 13271 9496 13277
rect 9580 13277 9597 13308
rect 9631 13277 9643 13311
rect 9580 13271 9643 13277
rect 9456 13246 9462 13271
rect 7101 13175 7159 13181
rect 7101 13141 7113 13175
rect 7147 13141 7159 13175
rect 7101 13135 7159 13141
rect 9122 13132 9128 13184
rect 9180 13172 9186 13184
rect 9580 13172 9608 13271
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 9861 13311 9919 13317
rect 9732 13280 9777 13308
rect 9732 13268 9738 13280
rect 9861 13277 9873 13311
rect 9907 13308 9919 13311
rect 9950 13308 9956 13320
rect 9907 13280 9956 13308
rect 9907 13277 9919 13280
rect 9861 13271 9919 13277
rect 9950 13268 9956 13280
rect 10008 13308 10014 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 10008 13280 10241 13308
rect 10008 13268 10014 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10686 13308 10692 13320
rect 10647 13280 10692 13308
rect 10229 13271 10287 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 10965 13311 11023 13317
rect 11146 13314 11152 13320
rect 10965 13308 10977 13311
rect 10888 13280 10977 13308
rect 10888 13252 10916 13280
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 11093 13308 11152 13314
rect 11093 13274 11105 13308
rect 11139 13274 11152 13308
rect 11093 13268 11152 13274
rect 11204 13268 11210 13320
rect 11339 13311 11397 13317
rect 11241 13285 11299 13291
rect 10134 13200 10140 13252
rect 10192 13240 10198 13252
rect 10192 13212 10732 13240
rect 10192 13200 10198 13212
rect 10042 13172 10048 13184
rect 9180 13144 9608 13172
rect 10003 13144 10048 13172
rect 9180 13132 9186 13144
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 10594 13172 10600 13184
rect 10555 13144 10600 13172
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 10704 13172 10732 13212
rect 10870 13200 10876 13252
rect 10928 13200 10934 13252
rect 11241 13251 11253 13285
rect 11287 13251 11299 13285
rect 11339 13277 11351 13311
rect 11385 13308 11397 13311
rect 11440 13308 11468 13416
rect 11532 13317 11560 13484
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 11977 13515 12035 13521
rect 11977 13512 11989 13515
rect 11848 13484 11989 13512
rect 11848 13472 11854 13484
rect 11977 13481 11989 13484
rect 12023 13481 12035 13515
rect 14642 13512 14648 13524
rect 11977 13475 12035 13481
rect 12360 13484 13952 13512
rect 14603 13484 14648 13512
rect 12250 13444 12256 13456
rect 11900 13416 12256 13444
rect 11701 13379 11759 13385
rect 11701 13345 11713 13379
rect 11747 13376 11759 13379
rect 11790 13376 11796 13388
rect 11747 13348 11796 13376
rect 11747 13345 11759 13348
rect 11701 13339 11759 13345
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 11385 13280 11468 13308
rect 11385 13277 11397 13280
rect 11339 13271 11397 13277
rect 11241 13245 11299 13251
rect 11256 13172 11284 13245
rect 11440 13240 11468 13280
rect 11516 13311 11574 13317
rect 11516 13277 11528 13311
rect 11562 13277 11574 13311
rect 11516 13271 11574 13277
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 11900 13317 11928 13416
rect 12250 13404 12256 13416
rect 12308 13404 12314 13456
rect 12360 13376 12388 13484
rect 12526 13444 12532 13456
rect 12452 13416 12532 13444
rect 12452 13385 12480 13416
rect 12526 13404 12532 13416
rect 12584 13404 12590 13456
rect 12897 13447 12955 13453
rect 12897 13413 12909 13447
rect 12943 13444 12955 13447
rect 13170 13444 13176 13456
rect 12943 13416 13176 13444
rect 12943 13413 12955 13416
rect 12897 13407 12955 13413
rect 13170 13404 13176 13416
rect 13228 13404 13234 13456
rect 12268 13348 12388 13376
rect 12437 13379 12495 13385
rect 11885 13311 11943 13317
rect 11664 13280 11709 13308
rect 11664 13268 11670 13280
rect 11885 13277 11897 13311
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 12161 13311 12219 13317
rect 12161 13277 12173 13311
rect 12207 13277 12219 13311
rect 12268 13305 12296 13348
rect 12437 13345 12449 13379
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 13924 13385 13952 13484
rect 14642 13472 14648 13484
rect 14700 13472 14706 13524
rect 17037 13515 17095 13521
rect 17037 13481 17049 13515
rect 17083 13512 17095 13515
rect 17494 13512 17500 13524
rect 17083 13484 17500 13512
rect 17083 13481 17095 13484
rect 17037 13475 17095 13481
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 20346 13472 20352 13524
rect 20404 13512 20410 13524
rect 21358 13512 21364 13524
rect 20404 13484 21364 13512
rect 20404 13472 20410 13484
rect 21358 13472 21364 13484
rect 21416 13512 21422 13524
rect 21453 13515 21511 13521
rect 21453 13512 21465 13515
rect 21416 13484 21465 13512
rect 21416 13472 21422 13484
rect 21453 13481 21465 13484
rect 21499 13481 21511 13515
rect 21453 13475 21511 13481
rect 21542 13472 21548 13524
rect 21600 13512 21606 13524
rect 21637 13515 21695 13521
rect 21637 13512 21649 13515
rect 21600 13484 21649 13512
rect 21600 13472 21606 13484
rect 21637 13481 21649 13484
rect 21683 13512 21695 13515
rect 23109 13515 23167 13521
rect 23109 13512 23121 13515
rect 21683 13484 23121 13512
rect 21683 13481 21695 13484
rect 21637 13475 21695 13481
rect 23109 13481 23121 13484
rect 23155 13512 23167 13515
rect 23658 13512 23664 13524
rect 23155 13484 23664 13512
rect 23155 13481 23167 13484
rect 23109 13475 23167 13481
rect 23658 13472 23664 13484
rect 23716 13472 23722 13524
rect 24118 13472 24124 13524
rect 24176 13512 24182 13524
rect 24489 13515 24547 13521
rect 24489 13512 24501 13515
rect 24176 13484 24501 13512
rect 24176 13472 24182 13484
rect 24489 13481 24501 13484
rect 24535 13481 24547 13515
rect 24489 13475 24547 13481
rect 14090 13444 14096 13456
rect 14051 13416 14096 13444
rect 14090 13404 14096 13416
rect 14148 13404 14154 13456
rect 23382 13444 23388 13456
rect 15120 13416 23388 13444
rect 13357 13379 13415 13385
rect 13357 13376 13369 13379
rect 12676 13348 13369 13376
rect 12676 13336 12682 13348
rect 13357 13345 13369 13348
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 13909 13379 13967 13385
rect 13909 13345 13921 13379
rect 13955 13376 13967 13379
rect 15120 13376 15148 13416
rect 23382 13404 23388 13416
rect 23440 13404 23446 13456
rect 17586 13376 17592 13388
rect 13955 13348 15148 13376
rect 17547 13348 17592 13376
rect 13955 13345 13967 13348
rect 13909 13339 13967 13345
rect 17586 13336 17592 13348
rect 17644 13336 17650 13388
rect 17678 13336 17684 13388
rect 17736 13376 17742 13388
rect 18414 13376 18420 13388
rect 17736 13348 17781 13376
rect 18375 13348 18420 13376
rect 17736 13336 17742 13348
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 18601 13379 18659 13385
rect 18601 13345 18613 13379
rect 18647 13376 18659 13379
rect 19334 13376 19340 13388
rect 18647 13348 19340 13376
rect 18647 13345 18659 13348
rect 18601 13339 18659 13345
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 20346 13336 20352 13388
rect 20404 13376 20410 13388
rect 20533 13379 20591 13385
rect 20533 13376 20545 13379
rect 20404 13348 20545 13376
rect 20404 13336 20410 13348
rect 20533 13345 20545 13348
rect 20579 13345 20591 13379
rect 20533 13339 20591 13345
rect 21450 13336 21456 13388
rect 21508 13376 21514 13388
rect 21729 13379 21787 13385
rect 21729 13376 21741 13379
rect 21508 13348 21741 13376
rect 21508 13336 21514 13348
rect 21729 13345 21741 13348
rect 21775 13345 21787 13379
rect 23477 13379 23535 13385
rect 23477 13376 23489 13379
rect 21729 13339 21787 13345
rect 22940 13348 23489 13376
rect 12326 13308 12384 13314
rect 12326 13305 12338 13308
rect 12268 13277 12338 13305
rect 12161 13271 12219 13277
rect 12326 13274 12338 13277
rect 12372 13274 12384 13308
rect 12176 13240 12204 13271
rect 12326 13268 12384 13274
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13277 12587 13311
rect 12529 13271 12587 13277
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13277 12771 13311
rect 12713 13271 12771 13277
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13078 13308 13084 13320
rect 13035 13280 13084 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 12544 13240 12572 13271
rect 11440 13212 12204 13240
rect 12268 13212 12572 13240
rect 12728 13240 12756 13271
rect 13078 13268 13084 13280
rect 13136 13268 13142 13320
rect 13172 13311 13230 13317
rect 13172 13277 13184 13311
rect 13218 13277 13230 13311
rect 13172 13271 13230 13277
rect 13187 13240 13225 13271
rect 13262 13268 13268 13320
rect 13320 13308 13326 13320
rect 13320 13280 13365 13308
rect 13320 13268 13326 13280
rect 13538 13268 13544 13320
rect 13596 13308 13602 13320
rect 14458 13308 14464 13320
rect 13596 13280 13641 13308
rect 14419 13280 14464 13308
rect 13596 13268 13602 13280
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 14734 13308 14740 13320
rect 14695 13280 14740 13308
rect 14734 13268 14740 13280
rect 14792 13268 14798 13320
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 17497 13311 17555 13317
rect 17497 13308 17509 13311
rect 17368 13280 17509 13308
rect 17368 13268 17374 13280
rect 17497 13277 17509 13280
rect 17543 13277 17555 13311
rect 17497 13271 17555 13277
rect 18138 13268 18144 13320
rect 18196 13308 18202 13320
rect 18325 13311 18383 13317
rect 18325 13308 18337 13311
rect 18196 13280 18337 13308
rect 18196 13268 18202 13280
rect 18325 13277 18337 13280
rect 18371 13277 18383 13311
rect 18325 13271 18383 13277
rect 20438 13268 20444 13320
rect 20496 13308 20502 13320
rect 20717 13311 20775 13317
rect 20717 13308 20729 13311
rect 20496 13280 20729 13308
rect 20496 13268 20502 13280
rect 20717 13277 20729 13280
rect 20763 13277 20775 13311
rect 20717 13271 20775 13277
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 21266 13308 21272 13320
rect 20855 13280 21272 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 21637 13311 21695 13317
rect 21637 13277 21649 13311
rect 21683 13308 21695 13311
rect 21910 13308 21916 13320
rect 21683 13280 21772 13308
rect 21871 13280 21916 13308
rect 21683 13277 21695 13280
rect 21637 13271 21695 13277
rect 14274 13240 14280 13252
rect 12728 13212 13768 13240
rect 14235 13212 14280 13240
rect 12268 13184 12296 13212
rect 10704 13144 11284 13172
rect 11330 13132 11336 13184
rect 11388 13172 11394 13184
rect 11606 13172 11612 13184
rect 11388 13144 11612 13172
rect 11388 13132 11394 13144
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 11790 13132 11796 13184
rect 11848 13172 11854 13184
rect 12250 13172 12256 13184
rect 11848 13144 12256 13172
rect 11848 13132 11854 13144
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 13630 13172 13636 13184
rect 13591 13144 13636 13172
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 13740 13172 13768 13212
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 21744 13240 21772 13280
rect 21910 13268 21916 13280
rect 21968 13308 21974 13320
rect 22940 13317 22968 13348
rect 23477 13345 23489 13348
rect 23523 13376 23535 13379
rect 23842 13376 23848 13388
rect 23523 13348 23848 13376
rect 23523 13345 23535 13348
rect 23477 13339 23535 13345
rect 23842 13336 23848 13348
rect 23900 13336 23906 13388
rect 23934 13336 23940 13388
rect 23992 13376 23998 13388
rect 24029 13379 24087 13385
rect 24029 13376 24041 13379
rect 23992 13348 24041 13376
rect 23992 13336 23998 13348
rect 24029 13345 24041 13348
rect 24075 13376 24087 13379
rect 24949 13379 25007 13385
rect 24075 13348 24808 13376
rect 24075 13345 24087 13348
rect 24029 13339 24087 13345
rect 22373 13311 22431 13317
rect 22373 13308 22385 13311
rect 21968 13280 22385 13308
rect 21968 13268 21974 13280
rect 22373 13277 22385 13280
rect 22419 13277 22431 13311
rect 22373 13271 22431 13277
rect 22925 13311 22983 13317
rect 22925 13277 22937 13311
rect 22971 13277 22983 13311
rect 22925 13271 22983 13277
rect 23017 13311 23075 13317
rect 23017 13277 23029 13311
rect 23063 13277 23075 13311
rect 23658 13308 23664 13320
rect 23619 13280 23664 13308
rect 23017 13271 23075 13277
rect 22002 13240 22008 13252
rect 14608 13212 21772 13240
rect 21963 13212 22008 13240
rect 14608 13200 14614 13212
rect 14568 13172 14596 13200
rect 14918 13172 14924 13184
rect 13740 13144 14596 13172
rect 14879 13144 14924 13172
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 17126 13172 17132 13184
rect 17087 13144 17132 13172
rect 17126 13132 17132 13144
rect 17184 13132 17190 13184
rect 17954 13172 17960 13184
rect 17915 13144 17960 13172
rect 17954 13132 17960 13144
rect 18012 13132 18018 13184
rect 20346 13172 20352 13184
rect 20307 13144 20352 13172
rect 20346 13132 20352 13144
rect 20404 13132 20410 13184
rect 20898 13132 20904 13184
rect 20956 13172 20962 13184
rect 21177 13175 21235 13181
rect 21177 13172 21189 13175
rect 20956 13144 21189 13172
rect 20956 13132 20962 13144
rect 21177 13141 21189 13144
rect 21223 13141 21235 13175
rect 21744 13172 21772 13212
rect 22002 13200 22008 13212
rect 22060 13200 22066 13252
rect 22189 13243 22247 13249
rect 22189 13209 22201 13243
rect 22235 13240 22247 13243
rect 22462 13240 22468 13252
rect 22235 13212 22468 13240
rect 22235 13209 22247 13212
rect 22189 13203 22247 13209
rect 22462 13200 22468 13212
rect 22520 13200 22526 13252
rect 23032 13240 23060 13271
rect 23658 13268 23664 13280
rect 23716 13268 23722 13320
rect 24780 13317 24808 13348
rect 24949 13345 24961 13379
rect 24995 13376 25007 13379
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 24995 13348 25145 13376
rect 24995 13345 25007 13348
rect 24949 13339 25007 13345
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 24765 13311 24823 13317
rect 23768 13280 24716 13308
rect 23768 13240 23796 13280
rect 22940 13212 23796 13240
rect 23937 13243 23995 13249
rect 22940 13184 22968 13212
rect 23937 13209 23949 13243
rect 23983 13240 23995 13243
rect 24302 13240 24308 13252
rect 23983 13212 24308 13240
rect 23983 13209 23995 13212
rect 23937 13203 23995 13209
rect 24302 13200 24308 13212
rect 24360 13200 24366 13252
rect 24397 13243 24455 13249
rect 24397 13209 24409 13243
rect 24443 13209 24455 13243
rect 24688 13240 24716 13280
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 25041 13311 25099 13317
rect 25041 13277 25053 13311
rect 25087 13277 25099 13311
rect 25041 13271 25099 13277
rect 25056 13240 25084 13271
rect 24688 13212 25084 13240
rect 24397 13203 24455 13209
rect 22922 13172 22928 13184
rect 21744 13144 22928 13172
rect 21177 13135 21235 13141
rect 22922 13132 22928 13144
rect 22980 13132 22986 13184
rect 23293 13175 23351 13181
rect 23293 13141 23305 13175
rect 23339 13172 23351 13175
rect 23750 13172 23756 13184
rect 23339 13144 23756 13172
rect 23339 13141 23351 13144
rect 23293 13135 23351 13141
rect 23750 13132 23756 13144
rect 23808 13172 23814 13184
rect 24412 13172 24440 13203
rect 23808 13144 24440 13172
rect 23808 13132 23814 13144
rect 1104 13082 26128 13104
rect 1104 13030 9291 13082
rect 9343 13030 9355 13082
rect 9407 13030 9419 13082
rect 9471 13030 9483 13082
rect 9535 13030 9547 13082
rect 9599 13030 17632 13082
rect 17684 13030 17696 13082
rect 17748 13030 17760 13082
rect 17812 13030 17824 13082
rect 17876 13030 17888 13082
rect 17940 13030 26128 13082
rect 1104 13008 26128 13030
rect 2958 12928 2964 12980
rect 3016 12968 3022 12980
rect 3237 12971 3295 12977
rect 3237 12968 3249 12971
rect 3016 12940 3249 12968
rect 3016 12928 3022 12940
rect 3237 12937 3249 12940
rect 3283 12937 3295 12971
rect 3237 12931 3295 12937
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 3421 12971 3479 12977
rect 3421 12968 3433 12971
rect 3384 12940 3433 12968
rect 3384 12928 3390 12940
rect 3421 12937 3433 12940
rect 3467 12937 3479 12971
rect 3421 12931 3479 12937
rect 3789 12971 3847 12977
rect 3789 12937 3801 12971
rect 3835 12968 3847 12971
rect 5442 12968 5448 12980
rect 3835 12940 5448 12968
rect 3835 12937 3847 12940
rect 3789 12931 3847 12937
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 5626 12928 5632 12980
rect 5684 12968 5690 12980
rect 6089 12971 6147 12977
rect 6089 12968 6101 12971
rect 5684 12940 6101 12968
rect 5684 12928 5690 12940
rect 6089 12937 6101 12940
rect 6135 12968 6147 12971
rect 6178 12968 6184 12980
rect 6135 12940 6184 12968
rect 6135 12937 6147 12940
rect 6089 12931 6147 12937
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 7432 12940 7757 12968
rect 7432 12928 7438 12940
rect 7745 12937 7757 12940
rect 7791 12937 7803 12971
rect 7745 12931 7803 12937
rect 9030 12928 9036 12980
rect 9088 12928 9094 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 9953 12971 10011 12977
rect 9732 12940 9777 12968
rect 9732 12928 9738 12940
rect 9953 12937 9965 12971
rect 9999 12968 10011 12971
rect 10134 12968 10140 12980
rect 9999 12940 10140 12968
rect 9999 12937 10011 12940
rect 9953 12931 10011 12937
rect 10134 12928 10140 12940
rect 10192 12968 10198 12980
rect 10686 12968 10692 12980
rect 10192 12940 10692 12968
rect 10192 12928 10198 12940
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 11517 12971 11575 12977
rect 11517 12968 11529 12971
rect 10928 12940 11529 12968
rect 10928 12928 10934 12940
rect 11517 12937 11529 12940
rect 11563 12968 11575 12971
rect 11793 12971 11851 12977
rect 11793 12968 11805 12971
rect 11563 12940 11805 12968
rect 11563 12937 11575 12940
rect 11517 12931 11575 12937
rect 11793 12937 11805 12940
rect 11839 12937 11851 12971
rect 11793 12931 11851 12937
rect 14090 12928 14096 12980
rect 14148 12928 14154 12980
rect 16393 12971 16451 12977
rect 16393 12937 16405 12971
rect 16439 12937 16451 12971
rect 16393 12931 16451 12937
rect 2124 12903 2182 12909
rect 2124 12869 2136 12903
rect 2170 12900 2182 12903
rect 2774 12900 2780 12912
rect 2170 12872 2780 12900
rect 2170 12869 2182 12872
rect 2124 12863 2182 12869
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 3878 12900 3884 12912
rect 3839 12872 3884 12900
rect 3878 12860 3884 12872
rect 3936 12860 3942 12912
rect 4724 12872 6408 12900
rect 4724 12844 4752 12872
rect 4706 12832 4712 12844
rect 4619 12804 4712 12832
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 4976 12835 5034 12841
rect 4976 12801 4988 12835
rect 5022 12832 5034 12835
rect 5534 12832 5540 12844
rect 5022 12804 5540 12832
rect 5022 12801 5034 12804
rect 4976 12795 5034 12801
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 6380 12841 6408 12872
rect 8662 12860 8668 12912
rect 8720 12860 8726 12912
rect 8941 12903 8999 12909
rect 8941 12869 8953 12903
rect 8987 12900 8999 12903
rect 9048 12900 9076 12928
rect 9858 12900 9864 12912
rect 8987 12872 9864 12900
rect 8987 12869 8999 12872
rect 8941 12863 8999 12869
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 6621 12835 6679 12841
rect 6621 12832 6633 12835
rect 6512 12804 6633 12832
rect 6512 12792 6518 12804
rect 6621 12801 6633 12804
rect 6667 12801 6679 12835
rect 8680 12832 8708 12860
rect 9324 12841 9352 12872
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 10594 12860 10600 12912
rect 10652 12900 10658 12912
rect 11066 12903 11124 12909
rect 11066 12900 11078 12903
rect 10652 12872 11078 12900
rect 10652 12860 10658 12872
rect 11066 12869 11078 12872
rect 11112 12869 11124 12903
rect 14108 12900 14136 12928
rect 14108 12872 14412 12900
rect 11066 12863 11124 12869
rect 9033 12835 9091 12841
rect 9033 12832 9045 12835
rect 8680 12804 9045 12832
rect 6621 12795 6679 12801
rect 9033 12801 9045 12804
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9309 12835 9367 12841
rect 9309 12801 9321 12835
rect 9355 12801 9367 12835
rect 9309 12795 9367 12801
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 1670 12724 1676 12776
rect 1728 12764 1734 12776
rect 1857 12767 1915 12773
rect 1857 12764 1869 12767
rect 1728 12736 1869 12764
rect 1728 12724 1734 12736
rect 1857 12733 1869 12736
rect 1903 12733 1915 12767
rect 1857 12727 1915 12733
rect 4065 12767 4123 12773
rect 4065 12733 4077 12767
rect 4111 12764 4123 12767
rect 4338 12764 4344 12776
rect 4111 12736 4344 12764
rect 4111 12733 4123 12736
rect 4065 12727 4123 12733
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 8938 12764 8944 12776
rect 8720 12736 8944 12764
rect 8720 12724 8726 12736
rect 8938 12724 8944 12736
rect 8996 12764 9002 12776
rect 9508 12764 9536 12795
rect 10042 12792 10048 12844
rect 10100 12832 10106 12844
rect 11333 12835 11391 12841
rect 10100 12804 11284 12832
rect 10100 12792 10106 12804
rect 8996 12736 9536 12764
rect 11256 12764 11284 12804
rect 11333 12801 11345 12835
rect 11379 12832 11391 12835
rect 11514 12832 11520 12844
rect 11379 12804 11520 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 11606 12764 11612 12776
rect 11256 12736 11612 12764
rect 8996 12724 9002 12736
rect 11606 12724 11612 12736
rect 11664 12764 11670 12776
rect 11716 12764 11744 12795
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 12161 12835 12219 12841
rect 11940 12804 11985 12832
rect 11940 12792 11946 12804
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 12434 12832 12440 12844
rect 12207 12804 12440 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 12621 12835 12679 12841
rect 12621 12801 12633 12835
rect 12667 12832 12679 12835
rect 12986 12832 12992 12844
rect 12667 12804 12992 12832
rect 12667 12801 12679 12804
rect 12621 12795 12679 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 14384 12841 14412 12872
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 16408 12900 16436 12931
rect 18138 12928 18144 12980
rect 18196 12968 18202 12980
rect 18325 12971 18383 12977
rect 18325 12968 18337 12971
rect 18196 12940 18337 12968
rect 18196 12928 18202 12940
rect 18325 12937 18337 12940
rect 18371 12968 18383 12971
rect 18782 12968 18788 12980
rect 18371 12940 18788 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 20993 12971 21051 12977
rect 20993 12937 21005 12971
rect 21039 12968 21051 12971
rect 21266 12968 21272 12980
rect 21039 12940 21272 12968
rect 21039 12937 21051 12940
rect 20993 12931 21051 12937
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 21545 12971 21603 12977
rect 21545 12937 21557 12971
rect 21591 12968 21603 12971
rect 21634 12968 21640 12980
rect 21591 12940 21640 12968
rect 21591 12937 21603 12940
rect 21545 12931 21603 12937
rect 21634 12928 21640 12940
rect 21692 12928 21698 12980
rect 22005 12971 22063 12977
rect 22005 12937 22017 12971
rect 22051 12968 22063 12971
rect 23385 12971 23443 12977
rect 22051 12940 22508 12968
rect 22051 12937 22063 12940
rect 22005 12931 22063 12937
rect 22370 12900 22376 12912
rect 15988 12872 22376 12900
rect 15988 12860 15994 12872
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 14102 12835 14160 12841
rect 14102 12832 14114 12835
rect 13688 12804 14114 12832
rect 13688 12792 13694 12804
rect 14102 12801 14114 12804
rect 14148 12801 14160 12835
rect 14102 12795 14160 12801
rect 14369 12835 14427 12841
rect 14369 12801 14381 12835
rect 14415 12832 14427 12835
rect 15010 12832 15016 12844
rect 14415 12804 15016 12832
rect 14415 12801 14427 12804
rect 14369 12795 14427 12801
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 15280 12835 15338 12841
rect 15280 12801 15292 12835
rect 15326 12832 15338 12835
rect 15562 12832 15568 12844
rect 15326 12804 15568 12832
rect 15326 12801 15338 12804
rect 15280 12795 15338 12801
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 18414 12832 18420 12844
rect 18327 12804 18420 12832
rect 18414 12792 18420 12804
rect 18472 12832 18478 12844
rect 19058 12832 19064 12844
rect 18472 12804 19064 12832
rect 18472 12792 18478 12804
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 20806 12792 20812 12844
rect 20864 12832 20870 12844
rect 21361 12835 21419 12841
rect 21361 12832 21373 12835
rect 20864 12804 21373 12832
rect 20864 12792 20870 12804
rect 21361 12801 21373 12804
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 21821 12835 21879 12841
rect 21821 12801 21833 12835
rect 21867 12832 21879 12835
rect 21910 12832 21916 12844
rect 21867 12804 21916 12832
rect 21867 12801 21879 12804
rect 21821 12795 21879 12801
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 22480 12832 22508 12940
rect 23385 12937 23397 12971
rect 23431 12968 23443 12971
rect 23845 12971 23903 12977
rect 23845 12968 23857 12971
rect 23431 12940 23857 12968
rect 23431 12937 23443 12940
rect 23385 12931 23443 12937
rect 23845 12937 23857 12940
rect 23891 12937 23903 12971
rect 23845 12931 23903 12937
rect 24118 12928 24124 12980
rect 24176 12968 24182 12980
rect 24213 12971 24271 12977
rect 24213 12968 24225 12971
rect 24176 12940 24225 12968
rect 24176 12928 24182 12940
rect 24213 12937 24225 12940
rect 24259 12937 24271 12971
rect 24213 12931 24271 12937
rect 22922 12860 22928 12912
rect 22980 12900 22986 12912
rect 24305 12903 24363 12909
rect 24305 12900 24317 12903
rect 22980 12872 24317 12900
rect 22980 12860 22986 12872
rect 24305 12869 24317 12872
rect 24351 12869 24363 12903
rect 24305 12863 24363 12869
rect 22556 12835 22614 12841
rect 22556 12832 22568 12835
rect 22480 12804 22568 12832
rect 22556 12801 22568 12804
rect 22602 12832 22614 12835
rect 23842 12832 23848 12844
rect 22602 12804 23848 12832
rect 22602 12801 22614 12804
rect 22556 12795 22614 12801
rect 23842 12792 23848 12804
rect 23900 12792 23906 12844
rect 24118 12792 24124 12844
rect 24176 12792 24182 12844
rect 11664 12736 11744 12764
rect 11793 12767 11851 12773
rect 11664 12724 11670 12736
rect 11793 12733 11805 12767
rect 11839 12764 11851 12767
rect 13262 12764 13268 12776
rect 11839 12736 13268 12764
rect 11839 12733 11851 12736
rect 11793 12727 11851 12733
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 17865 12767 17923 12773
rect 17865 12764 17877 12767
rect 17552 12736 17877 12764
rect 17552 12724 17558 12736
rect 17865 12733 17877 12736
rect 17911 12764 17923 12767
rect 19153 12767 19211 12773
rect 19153 12764 19165 12767
rect 17911 12736 19165 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 19153 12733 19165 12736
rect 19199 12764 19211 12767
rect 19334 12764 19340 12776
rect 19199 12736 19340 12764
rect 19199 12733 19211 12736
rect 19153 12727 19211 12733
rect 19334 12724 19340 12736
rect 19392 12764 19398 12776
rect 19794 12764 19800 12776
rect 19392 12736 19800 12764
rect 19392 12724 19398 12736
rect 19794 12724 19800 12736
rect 19852 12764 19858 12776
rect 20349 12767 20407 12773
rect 20349 12764 20361 12767
rect 19852 12736 20361 12764
rect 19852 12724 19858 12736
rect 20349 12733 20361 12736
rect 20395 12764 20407 12767
rect 21085 12767 21143 12773
rect 21085 12764 21097 12767
rect 20395 12736 21097 12764
rect 20395 12733 20407 12736
rect 20349 12727 20407 12733
rect 21085 12733 21097 12736
rect 21131 12764 21143 12767
rect 21450 12764 21456 12776
rect 21131 12736 21456 12764
rect 21131 12733 21143 12736
rect 21085 12727 21143 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 21634 12724 21640 12776
rect 21692 12764 21698 12776
rect 22002 12764 22008 12776
rect 21692 12736 22008 12764
rect 21692 12724 21698 12736
rect 22002 12724 22008 12736
rect 22060 12764 22066 12776
rect 22097 12767 22155 12773
rect 22097 12764 22109 12767
rect 22060 12736 22109 12764
rect 22060 12724 22066 12736
rect 22097 12733 22109 12736
rect 22143 12733 22155 12767
rect 22097 12727 22155 12733
rect 22189 12767 22247 12773
rect 22189 12733 22201 12767
rect 22235 12764 22247 12767
rect 23109 12767 23167 12773
rect 23109 12764 23121 12767
rect 22235 12736 22508 12764
rect 22235 12733 22247 12736
rect 22189 12727 22247 12733
rect 22480 12708 22508 12736
rect 22848 12736 23121 12764
rect 9122 12696 9128 12708
rect 9083 12668 9128 12696
rect 9122 12656 9128 12668
rect 9180 12656 9186 12708
rect 11330 12656 11336 12708
rect 11388 12696 11394 12708
rect 12345 12699 12403 12705
rect 12345 12696 12357 12699
rect 11388 12668 12357 12696
rect 11388 12656 11394 12668
rect 12345 12665 12357 12668
rect 12391 12696 12403 12699
rect 12434 12696 12440 12708
rect 12391 12668 12440 12696
rect 12391 12665 12403 12668
rect 12345 12659 12403 12665
rect 12434 12656 12440 12668
rect 12492 12656 12498 12708
rect 12710 12656 12716 12708
rect 12768 12696 12774 12708
rect 12989 12699 13047 12705
rect 12989 12696 13001 12699
rect 12768 12668 13001 12696
rect 12768 12656 12774 12668
rect 12989 12665 13001 12668
rect 13035 12665 13047 12699
rect 12989 12659 13047 12665
rect 22462 12656 22468 12708
rect 22520 12656 22526 12708
rect 22848 12640 22876 12736
rect 23109 12733 23121 12736
rect 23155 12733 23167 12767
rect 23109 12727 23167 12733
rect 23293 12767 23351 12773
rect 23293 12733 23305 12767
rect 23339 12764 23351 12767
rect 24136 12764 24164 12792
rect 23339 12736 24164 12764
rect 24397 12767 24455 12773
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 24397 12733 24409 12767
rect 24443 12733 24455 12767
rect 24397 12727 24455 12733
rect 24118 12656 24124 12708
rect 24176 12696 24182 12708
rect 24412 12696 24440 12727
rect 24176 12668 24440 12696
rect 24176 12656 24182 12668
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 10318 12628 10324 12640
rect 8536 12600 10324 12628
rect 8536 12588 8542 12600
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 11422 12588 11428 12640
rect 11480 12628 11486 12640
rect 11882 12628 11888 12640
rect 11480 12600 11888 12628
rect 11480 12588 11486 12600
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 12069 12631 12127 12637
rect 12069 12597 12081 12631
rect 12115 12628 12127 12631
rect 12250 12628 12256 12640
rect 12115 12600 12256 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 12526 12628 12532 12640
rect 12487 12600 12532 12628
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 13078 12588 13084 12640
rect 13136 12628 13142 12640
rect 14918 12628 14924 12640
rect 13136 12600 14924 12628
rect 13136 12588 13142 12600
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 20533 12631 20591 12637
rect 20533 12597 20545 12631
rect 20579 12628 20591 12631
rect 21082 12628 21088 12640
rect 20579 12600 21088 12628
rect 20579 12597 20591 12600
rect 20533 12591 20591 12597
rect 21082 12588 21088 12600
rect 21140 12588 21146 12640
rect 22646 12588 22652 12640
rect 22704 12628 22710 12640
rect 22704 12600 22749 12628
rect 22704 12588 22710 12600
rect 22830 12588 22836 12640
rect 22888 12628 22894 12640
rect 23750 12628 23756 12640
rect 22888 12600 22933 12628
rect 23711 12600 23756 12628
rect 22888 12588 22894 12600
rect 23750 12588 23756 12600
rect 23808 12588 23814 12640
rect 1104 12538 26128 12560
rect 1104 12486 5120 12538
rect 5172 12486 5184 12538
rect 5236 12486 5248 12538
rect 5300 12486 5312 12538
rect 5364 12486 5376 12538
rect 5428 12486 13462 12538
rect 13514 12486 13526 12538
rect 13578 12486 13590 12538
rect 13642 12486 13654 12538
rect 13706 12486 13718 12538
rect 13770 12486 21803 12538
rect 21855 12486 21867 12538
rect 21919 12486 21931 12538
rect 21983 12486 21995 12538
rect 22047 12486 22059 12538
rect 22111 12486 26128 12538
rect 1104 12464 26128 12486
rect 7926 12384 7932 12436
rect 7984 12424 7990 12436
rect 9214 12424 9220 12436
rect 7984 12396 9220 12424
rect 7984 12384 7990 12396
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 9582 12384 9588 12436
rect 9640 12424 9646 12436
rect 10413 12427 10471 12433
rect 10413 12424 10425 12427
rect 9640 12396 10425 12424
rect 9640 12384 9646 12396
rect 10413 12393 10425 12396
rect 10459 12424 10471 12427
rect 10459 12396 10548 12424
rect 10459 12393 10471 12396
rect 10413 12387 10471 12393
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 9030 12356 9036 12368
rect 8352 12328 9036 12356
rect 8352 12316 8358 12328
rect 9030 12316 9036 12328
rect 9088 12316 9094 12368
rect 9769 12359 9827 12365
rect 9769 12356 9781 12359
rect 9416 12328 9781 12356
rect 8386 12248 8392 12300
rect 8444 12288 8450 12300
rect 9416 12297 9444 12328
rect 9769 12325 9781 12328
rect 9815 12325 9827 12359
rect 9769 12319 9827 12325
rect 10045 12359 10103 12365
rect 10045 12325 10057 12359
rect 10091 12325 10103 12359
rect 10520 12356 10548 12396
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 11606 12424 11612 12436
rect 11204 12396 11612 12424
rect 11204 12384 11210 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 12345 12427 12403 12433
rect 12345 12393 12357 12427
rect 12391 12424 12403 12427
rect 12618 12424 12624 12436
rect 12391 12396 12624 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 20073 12427 20131 12433
rect 20073 12424 20085 12427
rect 12820 12396 20085 12424
rect 10520 12328 11468 12356
rect 10045 12319 10103 12325
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 8444 12260 9413 12288
rect 8444 12248 8450 12260
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 10060 12288 10088 12319
rect 9401 12251 9459 12257
rect 9692 12260 10824 12288
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 6917 12223 6975 12229
rect 6917 12220 6929 12223
rect 6604 12192 6929 12220
rect 6604 12180 6610 12192
rect 6917 12189 6929 12192
rect 6963 12220 6975 12223
rect 8662 12220 8668 12232
rect 6963 12192 8668 12220
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 8772 12152 8800 12183
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 9088 12192 9137 12220
rect 9088 12180 9094 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 9272 12192 9321 12220
rect 9272 12180 9278 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9494 12223 9552 12229
rect 9494 12189 9506 12223
rect 9540 12220 9552 12223
rect 9582 12220 9588 12232
rect 9540 12192 9588 12220
rect 9540 12189 9552 12192
rect 9494 12183 9552 12189
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 9692 12229 9720 12260
rect 9677 12223 9735 12229
rect 9677 12189 9689 12223
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 9953 12223 10011 12229
rect 9953 12220 9965 12223
rect 9824 12192 9965 12220
rect 9824 12180 9830 12192
rect 9953 12189 9965 12192
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10796 12220 10824 12260
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 11330 12288 11336 12300
rect 10928 12260 11192 12288
rect 11291 12260 11336 12288
rect 10928 12248 10934 12260
rect 11054 12220 11060 12232
rect 10796 12192 11060 12220
rect 10229 12183 10287 12189
rect 10244 12152 10272 12183
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11164 12220 11192 12260
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 11440 12288 11468 12328
rect 11440 12260 12434 12288
rect 11222 12223 11280 12229
rect 11222 12220 11234 12223
rect 11164 12192 11234 12220
rect 11222 12189 11234 12192
rect 11268 12189 11280 12223
rect 11222 12183 11280 12189
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 11440 12152 11468 12183
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 12066 12220 12072 12232
rect 11664 12192 12072 12220
rect 11664 12180 11670 12192
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 12250 12152 12256 12164
rect 8772 12124 11008 12152
rect 11440 12124 12256 12152
rect 6822 12044 6828 12096
rect 6880 12084 6886 12096
rect 7009 12087 7067 12093
rect 7009 12084 7021 12087
rect 6880 12056 7021 12084
rect 6880 12044 6886 12056
rect 7009 12053 7021 12056
rect 7055 12053 7067 12087
rect 7009 12047 7067 12053
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 7800 12056 8585 12084
rect 7800 12044 7806 12056
rect 8573 12053 8585 12056
rect 8619 12053 8631 12087
rect 9030 12084 9036 12096
rect 8991 12056 9036 12084
rect 8573 12047 8631 12053
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 10410 12044 10416 12096
rect 10468 12084 10474 12096
rect 10870 12084 10876 12096
rect 10468 12056 10876 12084
rect 10468 12044 10474 12056
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 10980 12084 11008 12124
rect 12250 12112 12256 12124
rect 12308 12112 12314 12164
rect 12406 12152 12434 12260
rect 12618 12248 12624 12300
rect 12676 12288 12682 12300
rect 12820 12288 12848 12396
rect 20073 12393 20085 12396
rect 20119 12393 20131 12427
rect 20073 12387 20131 12393
rect 22741 12427 22799 12433
rect 22741 12393 22753 12427
rect 22787 12424 22799 12427
rect 23566 12424 23572 12436
rect 22787 12396 23572 12424
rect 22787 12393 22799 12396
rect 22741 12387 22799 12393
rect 23566 12384 23572 12396
rect 23624 12384 23630 12436
rect 12897 12359 12955 12365
rect 12897 12325 12909 12359
rect 12943 12356 12955 12359
rect 15746 12356 15752 12368
rect 12943 12328 15752 12356
rect 12943 12325 12955 12328
rect 12897 12319 12955 12325
rect 15304 12297 15332 12328
rect 15746 12316 15752 12328
rect 15804 12316 15810 12368
rect 16758 12316 16764 12368
rect 16816 12356 16822 12368
rect 17218 12356 17224 12368
rect 16816 12328 17224 12356
rect 16816 12316 16822 12328
rect 17218 12316 17224 12328
rect 17276 12316 17282 12368
rect 17313 12359 17371 12365
rect 17313 12325 17325 12359
rect 17359 12356 17371 12359
rect 17494 12356 17500 12368
rect 17359 12328 17500 12356
rect 17359 12325 17371 12328
rect 17313 12319 17371 12325
rect 17494 12316 17500 12328
rect 17552 12316 17558 12368
rect 18414 12356 18420 12368
rect 18375 12328 18420 12356
rect 18414 12316 18420 12328
rect 18472 12316 18478 12368
rect 20346 12356 20352 12368
rect 18892 12328 20352 12356
rect 12676 12260 12848 12288
rect 15289 12291 15347 12297
rect 12676 12248 12682 12260
rect 15289 12257 15301 12291
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 15562 12248 15568 12300
rect 15620 12288 15626 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15620 12260 15669 12288
rect 15620 12248 15626 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 16117 12291 16175 12297
rect 16117 12257 16129 12291
rect 16163 12288 16175 12291
rect 16574 12288 16580 12300
rect 16163 12260 16580 12288
rect 16163 12257 16175 12260
rect 16117 12251 16175 12257
rect 16574 12248 16580 12260
rect 16632 12288 16638 12300
rect 17236 12288 17264 12316
rect 18892 12297 18920 12328
rect 20346 12316 20352 12328
rect 20404 12316 20410 12368
rect 20806 12356 20812 12368
rect 20767 12328 20812 12356
rect 20806 12316 20812 12328
rect 20864 12316 20870 12368
rect 21284 12328 21588 12356
rect 17589 12291 17647 12297
rect 17589 12288 17601 12291
rect 16632 12260 16988 12288
rect 17236 12260 17601 12288
rect 16632 12248 16638 12260
rect 12526 12220 12532 12232
rect 12487 12192 12532 12220
rect 12526 12180 12532 12192
rect 12584 12220 12590 12232
rect 12713 12223 12771 12229
rect 12713 12220 12725 12223
rect 12584 12192 12725 12220
rect 12584 12180 12590 12192
rect 12713 12189 12725 12192
rect 12759 12189 12771 12223
rect 12986 12220 12992 12232
rect 12947 12192 12992 12220
rect 12713 12183 12771 12189
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 14918 12220 14924 12232
rect 14879 12192 14924 12220
rect 14918 12180 14924 12192
rect 14976 12180 14982 12232
rect 15102 12220 15108 12232
rect 15063 12192 15108 12220
rect 15102 12180 15108 12192
rect 15160 12180 15166 12232
rect 15197 12223 15255 12229
rect 15197 12189 15209 12223
rect 15243 12189 15255 12223
rect 15197 12183 15255 12189
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12220 15531 12223
rect 15930 12220 15936 12232
rect 15519 12192 15936 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 12802 12152 12808 12164
rect 12406 12124 12808 12152
rect 12802 12112 12808 12124
rect 12860 12112 12866 12164
rect 15212 12152 15240 12183
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 16960 12229 16988 12260
rect 17589 12257 17601 12260
rect 17635 12288 17647 12291
rect 18877 12291 18935 12297
rect 18877 12288 18889 12291
rect 17635 12260 18889 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 18877 12257 18889 12260
rect 18923 12257 18935 12291
rect 19702 12288 19708 12300
rect 19663 12260 19708 12288
rect 18877 12251 18935 12257
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 19794 12248 19800 12300
rect 19852 12288 19858 12300
rect 20073 12291 20131 12297
rect 19852 12260 19897 12288
rect 19852 12248 19858 12260
rect 20073 12257 20085 12291
rect 20119 12288 20131 12291
rect 20257 12291 20315 12297
rect 20257 12288 20269 12291
rect 20119 12260 20269 12288
rect 20119 12257 20131 12260
rect 20073 12251 20131 12257
rect 20257 12257 20269 12260
rect 20303 12288 20315 12291
rect 21284 12288 21312 12328
rect 21450 12288 21456 12300
rect 20303 12260 21312 12288
rect 21411 12260 21456 12288
rect 20303 12257 20315 12260
rect 20257 12251 20315 12257
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 21560 12288 21588 12328
rect 24118 12316 24124 12368
rect 24176 12356 24182 12368
rect 24176 12328 24992 12356
rect 24176 12316 24182 12328
rect 21910 12288 21916 12300
rect 21560 12260 21916 12288
rect 21910 12248 21916 12260
rect 21968 12248 21974 12300
rect 23658 12248 23664 12300
rect 23716 12288 23722 12300
rect 24964 12297 24992 12328
rect 24857 12291 24915 12297
rect 24857 12288 24869 12291
rect 23716 12260 24869 12288
rect 23716 12248 23722 12260
rect 24857 12257 24869 12260
rect 24903 12257 24915 12291
rect 24857 12251 24915 12257
rect 24949 12291 25007 12297
rect 24949 12257 24961 12291
rect 24995 12257 25007 12291
rect 24949 12251 25007 12257
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 16484 12223 16542 12229
rect 16484 12189 16496 12223
rect 16530 12220 16542 12223
rect 16945 12223 17003 12229
rect 16530 12192 16896 12220
rect 16530 12189 16542 12192
rect 16484 12183 16542 12189
rect 15378 12152 15384 12164
rect 15212 12124 15384 12152
rect 11606 12084 11612 12096
rect 10980 12056 11612 12084
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 11701 12087 11759 12093
rect 11701 12053 11713 12087
rect 11747 12084 11759 12087
rect 11790 12084 11796 12096
rect 11747 12056 11796 12084
rect 11747 12053 11759 12056
rect 11701 12047 11759 12053
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 13173 12087 13231 12093
rect 13173 12053 13185 12087
rect 13219 12084 13231 12087
rect 13262 12084 13268 12096
rect 13219 12056 13268 12084
rect 13219 12053 13231 12056
rect 13173 12047 13231 12053
rect 13262 12044 13268 12056
rect 13320 12084 13326 12096
rect 15212 12084 15240 12124
rect 15378 12112 15384 12124
rect 15436 12112 15442 12164
rect 16040 12152 16068 12183
rect 16761 12155 16819 12161
rect 16761 12152 16773 12155
rect 15488 12124 16773 12152
rect 15488 12096 15516 12124
rect 16761 12121 16773 12124
rect 16807 12121 16819 12155
rect 16761 12115 16819 12121
rect 13320 12056 15240 12084
rect 13320 12044 13326 12056
rect 15470 12044 15476 12096
rect 15528 12044 15534 12096
rect 16577 12087 16635 12093
rect 16577 12053 16589 12087
rect 16623 12084 16635 12087
rect 16666 12084 16672 12096
rect 16623 12056 16672 12084
rect 16623 12053 16635 12056
rect 16577 12047 16635 12053
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 16868 12084 16896 12192
rect 16945 12189 16957 12223
rect 16991 12189 17003 12223
rect 16945 12183 17003 12189
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12220 18199 12223
rect 18322 12220 18328 12232
rect 18187 12192 18328 12220
rect 18187 12189 18199 12192
rect 18141 12183 18199 12189
rect 17129 12155 17187 12161
rect 17129 12121 17141 12155
rect 17175 12152 17187 12155
rect 17972 12152 18000 12183
rect 18322 12180 18328 12192
rect 18380 12180 18386 12232
rect 18506 12220 18512 12232
rect 18467 12192 18512 12220
rect 18506 12180 18512 12192
rect 18564 12180 18570 12232
rect 18598 12180 18604 12232
rect 18656 12220 18662 12232
rect 20165 12223 20223 12229
rect 18656 12192 18701 12220
rect 18656 12180 18662 12192
rect 20165 12189 20177 12223
rect 20211 12189 20223 12223
rect 20165 12183 20223 12189
rect 20624 12223 20682 12229
rect 20624 12189 20636 12223
rect 20670 12220 20682 12223
rect 21634 12220 21640 12232
rect 20670 12192 21640 12220
rect 20670 12189 20682 12192
rect 20624 12183 20682 12189
rect 18782 12152 18788 12164
rect 17175 12124 18788 12152
rect 17175 12121 17187 12124
rect 17129 12115 17187 12121
rect 17144 12084 17172 12115
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 19334 12152 19340 12164
rect 18984 12124 19340 12152
rect 16868 12056 17172 12084
rect 18693 12087 18751 12093
rect 18693 12053 18705 12087
rect 18739 12084 18751 12087
rect 18984 12084 19012 12124
rect 19334 12112 19340 12124
rect 19392 12112 19398 12164
rect 20180 12152 20208 12183
rect 21634 12180 21640 12192
rect 21692 12220 21698 12232
rect 22097 12223 22155 12229
rect 22097 12220 22109 12223
rect 21692 12192 22109 12220
rect 21692 12180 21698 12192
rect 22097 12189 22109 12192
rect 22143 12189 22155 12223
rect 22554 12220 22560 12232
rect 22515 12192 22560 12220
rect 22097 12183 22155 12189
rect 22554 12180 22560 12192
rect 22612 12180 22618 12232
rect 24578 12180 24584 12232
rect 24636 12220 24642 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 24636 12192 24777 12220
rect 24636 12180 24642 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 20438 12152 20444 12164
rect 20180 12124 20444 12152
rect 20438 12112 20444 12124
rect 20496 12152 20502 12164
rect 21729 12155 21787 12161
rect 21729 12152 21741 12155
rect 20496 12124 21741 12152
rect 20496 12112 20502 12124
rect 21729 12121 21741 12124
rect 21775 12121 21787 12155
rect 21910 12152 21916 12164
rect 21871 12124 21916 12152
rect 21729 12115 21787 12121
rect 21910 12112 21916 12124
rect 21968 12112 21974 12164
rect 18739 12056 19012 12084
rect 18739 12053 18751 12056
rect 18693 12047 18751 12053
rect 19058 12044 19064 12096
rect 19116 12084 19122 12096
rect 19245 12087 19303 12093
rect 19245 12084 19257 12087
rect 19116 12056 19257 12084
rect 19116 12044 19122 12056
rect 19245 12053 19257 12056
rect 19291 12053 19303 12087
rect 19610 12084 19616 12096
rect 19571 12056 19616 12084
rect 19245 12047 19303 12053
rect 19610 12044 19616 12056
rect 19668 12044 19674 12096
rect 20898 12084 20904 12096
rect 20859 12056 20904 12084
rect 20898 12044 20904 12056
rect 20956 12044 20962 12096
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 21269 12087 21327 12093
rect 21269 12084 21281 12087
rect 21048 12056 21281 12084
rect 21048 12044 21054 12056
rect 21269 12053 21281 12056
rect 21315 12053 21327 12087
rect 21269 12047 21327 12053
rect 21358 12044 21364 12096
rect 21416 12084 21422 12096
rect 22094 12084 22100 12096
rect 21416 12056 22100 12084
rect 21416 12044 21422 12056
rect 22094 12044 22100 12056
rect 22152 12044 22158 12096
rect 22186 12044 22192 12096
rect 22244 12084 22250 12096
rect 22830 12084 22836 12096
rect 22244 12056 22836 12084
rect 22244 12044 22250 12056
rect 22830 12044 22836 12056
rect 22888 12044 22894 12096
rect 23658 12084 23664 12096
rect 23619 12056 23664 12084
rect 23658 12044 23664 12056
rect 23716 12084 23722 12096
rect 24118 12084 24124 12096
rect 23716 12056 24124 12084
rect 23716 12044 23722 12056
rect 24118 12044 24124 12056
rect 24176 12044 24182 12096
rect 24394 12084 24400 12096
rect 24355 12056 24400 12084
rect 24394 12044 24400 12056
rect 24452 12044 24458 12096
rect 1104 11994 26128 12016
rect 1104 11942 9291 11994
rect 9343 11942 9355 11994
rect 9407 11942 9419 11994
rect 9471 11942 9483 11994
rect 9535 11942 9547 11994
rect 9599 11942 17632 11994
rect 17684 11942 17696 11994
rect 17748 11942 17760 11994
rect 17812 11942 17824 11994
rect 17876 11942 17888 11994
rect 17940 11942 26128 11994
rect 1104 11920 26128 11942
rect 3234 11880 3240 11892
rect 3195 11852 3240 11880
rect 3234 11840 3240 11852
rect 3292 11840 3298 11892
rect 8938 11840 8944 11892
rect 8996 11880 9002 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 8996 11852 10701 11880
rect 8996 11840 9002 11852
rect 10689 11849 10701 11852
rect 10735 11880 10747 11883
rect 16850 11880 16856 11892
rect 10735 11852 16528 11880
rect 16811 11852 16856 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 3252 11812 3280 11840
rect 2976 11784 3280 11812
rect 1762 11704 1768 11756
rect 1820 11744 1826 11756
rect 2590 11744 2596 11756
rect 1820 11716 2596 11744
rect 1820 11704 1826 11716
rect 2590 11704 2596 11716
rect 2648 11744 2654 11756
rect 2976 11753 3004 11784
rect 4706 11772 4712 11824
rect 4764 11812 4770 11824
rect 5169 11815 5227 11821
rect 5169 11812 5181 11815
rect 4764 11784 5181 11812
rect 4764 11772 4770 11784
rect 5169 11781 5181 11784
rect 5215 11781 5227 11815
rect 5169 11775 5227 11781
rect 5353 11815 5411 11821
rect 5353 11781 5365 11815
rect 5399 11812 5411 11815
rect 7190 11812 7196 11824
rect 5399 11784 7196 11812
rect 5399 11781 5411 11784
rect 5353 11775 5411 11781
rect 7190 11772 7196 11784
rect 7248 11812 7254 11824
rect 9033 11815 9091 11821
rect 9033 11812 9045 11815
rect 7248 11784 9045 11812
rect 7248 11772 7254 11784
rect 9033 11781 9045 11784
rect 9079 11781 9091 11815
rect 9033 11775 9091 11781
rect 9324 11784 11008 11812
rect 2685 11747 2743 11753
rect 2685 11744 2697 11747
rect 2648 11716 2697 11744
rect 2648 11704 2654 11716
rect 2685 11713 2697 11716
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11713 3019 11747
rect 3142 11744 3148 11756
rect 3103 11716 3148 11744
rect 2961 11707 3019 11713
rect 3142 11704 3148 11716
rect 3200 11704 3206 11756
rect 6546 11744 6552 11756
rect 6507 11716 6552 11744
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 7800 11716 7941 11744
rect 7800 11704 7806 11716
rect 7929 11713 7941 11716
rect 7975 11713 7987 11747
rect 8094 11747 8152 11753
rect 8094 11744 8106 11747
rect 7929 11707 7987 11713
rect 8036 11716 8106 11744
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 3786 11676 3792 11688
rect 2832 11648 3792 11676
rect 2832 11636 2838 11648
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 8036 11676 8064 11716
rect 8094 11713 8106 11716
rect 8140 11713 8152 11747
rect 8094 11707 8152 11713
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11744 8263 11747
rect 8386 11744 8392 11756
rect 8251 11716 8392 11744
rect 8251 11713 8263 11716
rect 8205 11707 8263 11713
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11744 8539 11747
rect 8662 11744 8668 11756
rect 8527 11716 8668 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 8662 11704 8668 11716
rect 8720 11744 8726 11756
rect 8846 11744 8852 11756
rect 8720 11716 8852 11744
rect 8720 11704 8726 11716
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 9324 11753 9352 11784
rect 9217 11747 9275 11753
rect 9217 11744 9229 11747
rect 8996 11716 9229 11744
rect 8996 11704 9002 11716
rect 9217 11713 9229 11716
rect 9263 11744 9275 11747
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 9263 11716 9321 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9565 11747 9623 11753
rect 9565 11744 9577 11747
rect 9309 11707 9367 11713
rect 9416 11716 9577 11744
rect 7760 11648 8064 11676
rect 8297 11679 8355 11685
rect 2869 11611 2927 11617
rect 2869 11577 2881 11611
rect 2915 11608 2927 11611
rect 3418 11608 3424 11620
rect 2915 11580 3424 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 2498 11540 2504 11552
rect 2459 11512 2504 11540
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 5994 11500 6000 11552
rect 6052 11540 6058 11552
rect 6365 11543 6423 11549
rect 6365 11540 6377 11543
rect 6052 11512 6377 11540
rect 6052 11500 6058 11512
rect 6365 11509 6377 11512
rect 6411 11509 6423 11543
rect 6365 11503 6423 11509
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 7760 11549 7788 11648
rect 8297 11645 8309 11679
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 8312 11608 8340 11639
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 9416 11676 9444 11716
rect 9565 11713 9577 11716
rect 9611 11713 9623 11747
rect 9565 11707 9623 11713
rect 9088 11648 9444 11676
rect 10980 11676 11008 11784
rect 15194 11772 15200 11824
rect 15252 11812 15258 11824
rect 16390 11812 16396 11824
rect 15252 11784 16396 11812
rect 15252 11772 15258 11784
rect 16390 11772 16396 11784
rect 16448 11772 16454 11824
rect 16500 11812 16528 11852
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 17313 11883 17371 11889
rect 17313 11849 17325 11883
rect 17359 11880 17371 11883
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 17359 11852 17785 11880
rect 17359 11849 17371 11852
rect 17313 11843 17371 11849
rect 17773 11849 17785 11852
rect 17819 11849 17831 11883
rect 18138 11880 18144 11892
rect 18099 11852 18144 11880
rect 17773 11843 17831 11849
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 18506 11840 18512 11892
rect 18564 11880 18570 11892
rect 18877 11883 18935 11889
rect 18877 11880 18889 11883
rect 18564 11852 18889 11880
rect 18564 11840 18570 11852
rect 18877 11849 18889 11852
rect 18923 11880 18935 11883
rect 19337 11883 19395 11889
rect 18923 11852 19288 11880
rect 18923 11849 18935 11852
rect 18877 11843 18935 11849
rect 17405 11815 17463 11821
rect 16500 11784 17264 11812
rect 11790 11753 11796 11756
rect 11784 11744 11796 11753
rect 11751 11716 11796 11744
rect 11784 11707 11796 11716
rect 11790 11704 11796 11707
rect 11848 11704 11854 11756
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 15280 11747 15338 11753
rect 12124 11716 12940 11744
rect 12124 11704 12130 11716
rect 11514 11676 11520 11688
rect 10980 11648 11520 11676
rect 9088 11636 9094 11648
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 9214 11608 9220 11620
rect 8312 11580 9220 11608
rect 9214 11568 9220 11580
rect 9272 11568 9278 11620
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 6972 11512 7757 11540
rect 6972 11500 6978 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 8573 11543 8631 11549
rect 8573 11509 8585 11543
rect 8619 11540 8631 11543
rect 9030 11540 9036 11552
rect 8619 11512 9036 11540
rect 8619 11509 8631 11512
rect 8573 11503 8631 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 12618 11540 12624 11552
rect 10652 11512 12624 11540
rect 10652 11500 10658 11512
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 12912 11549 12940 11716
rect 15280 11713 15292 11747
rect 15326 11744 15338 11747
rect 15654 11744 15660 11756
rect 15326 11716 15660 11744
rect 15326 11713 15338 11716
rect 15280 11707 15338 11713
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 16666 11744 16672 11756
rect 16627 11716 16672 11744
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 13998 11676 14004 11688
rect 13228 11648 14004 11676
rect 13228 11636 13234 11648
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 14458 11636 14464 11688
rect 14516 11676 14522 11688
rect 15010 11676 15016 11688
rect 14516 11648 15016 11676
rect 14516 11636 14522 11648
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 17236 11608 17264 11784
rect 17405 11781 17417 11815
rect 17451 11812 17463 11815
rect 18156 11812 18184 11840
rect 17451 11784 18184 11812
rect 18233 11815 18291 11821
rect 17451 11781 17463 11784
rect 17405 11775 17463 11781
rect 18233 11781 18245 11815
rect 18279 11812 18291 11815
rect 18322 11812 18328 11824
rect 18279 11784 18328 11812
rect 18279 11781 18291 11784
rect 18233 11775 18291 11781
rect 18322 11772 18328 11784
rect 18380 11812 18386 11824
rect 18380 11784 18644 11812
rect 18380 11772 18386 11784
rect 17310 11704 17316 11756
rect 17368 11744 17374 11756
rect 18616 11753 18644 11784
rect 18601 11747 18659 11753
rect 17368 11716 18368 11744
rect 17368 11704 17374 11716
rect 17494 11676 17500 11688
rect 17455 11648 17500 11676
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 18340 11685 18368 11716
rect 18601 11713 18613 11747
rect 18647 11713 18659 11747
rect 18782 11744 18788 11756
rect 18743 11716 18788 11744
rect 18601 11707 18659 11713
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 18325 11679 18383 11685
rect 18325 11645 18337 11679
rect 18371 11676 18383 11679
rect 18874 11676 18880 11688
rect 18371 11648 18880 11676
rect 18371 11645 18383 11648
rect 18325 11639 18383 11645
rect 18874 11636 18880 11648
rect 18932 11676 18938 11688
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 18932 11648 19165 11676
rect 18932 11636 18938 11648
rect 19153 11645 19165 11648
rect 19199 11645 19211 11679
rect 19260 11676 19288 11852
rect 19337 11849 19349 11883
rect 19383 11880 19395 11883
rect 19518 11880 19524 11892
rect 19383 11852 19524 11880
rect 19383 11849 19395 11852
rect 19337 11843 19395 11849
rect 19518 11840 19524 11852
rect 19576 11840 19582 11892
rect 19610 11840 19616 11892
rect 19668 11880 19674 11892
rect 19797 11883 19855 11889
rect 19797 11880 19809 11883
rect 19668 11852 19809 11880
rect 19668 11840 19674 11852
rect 19797 11849 19809 11852
rect 19843 11849 19855 11883
rect 19797 11843 19855 11849
rect 19886 11840 19892 11892
rect 19944 11880 19950 11892
rect 20625 11883 20683 11889
rect 20625 11880 20637 11883
rect 19944 11852 20637 11880
rect 19944 11840 19950 11852
rect 20625 11849 20637 11852
rect 20671 11849 20683 11883
rect 20625 11843 20683 11849
rect 21177 11883 21235 11889
rect 21177 11849 21189 11883
rect 21223 11880 21235 11883
rect 21821 11883 21879 11889
rect 21821 11880 21833 11883
rect 21223 11852 21833 11880
rect 21223 11849 21235 11852
rect 21177 11843 21235 11849
rect 21821 11849 21833 11852
rect 21867 11849 21879 11883
rect 21821 11843 21879 11849
rect 21910 11840 21916 11892
rect 21968 11880 21974 11892
rect 22281 11883 22339 11889
rect 22281 11880 22293 11883
rect 21968 11852 22293 11880
rect 21968 11840 21974 11852
rect 22281 11849 22293 11852
rect 22327 11849 22339 11883
rect 22281 11843 22339 11849
rect 23293 11883 23351 11889
rect 23293 11849 23305 11883
rect 23339 11880 23351 11883
rect 23566 11880 23572 11892
rect 23339 11852 23572 11880
rect 23339 11849 23351 11852
rect 23293 11843 23351 11849
rect 23566 11840 23572 11852
rect 23624 11840 23630 11892
rect 24121 11883 24179 11889
rect 24121 11849 24133 11883
rect 24167 11880 24179 11883
rect 24394 11880 24400 11892
rect 24167 11852 24400 11880
rect 24167 11849 24179 11852
rect 24121 11843 24179 11849
rect 24394 11840 24400 11852
rect 24452 11840 24458 11892
rect 19429 11815 19487 11821
rect 19429 11781 19441 11815
rect 19475 11812 19487 11815
rect 19702 11812 19708 11824
rect 19475 11784 19708 11812
rect 19475 11781 19487 11784
rect 19429 11775 19487 11781
rect 19702 11772 19708 11784
rect 19760 11772 19766 11824
rect 20349 11815 20407 11821
rect 20349 11781 20361 11815
rect 20395 11812 20407 11815
rect 20530 11812 20536 11824
rect 20395 11784 20536 11812
rect 20395 11781 20407 11784
rect 20349 11775 20407 11781
rect 20530 11772 20536 11784
rect 20588 11772 20594 11824
rect 21269 11815 21327 11821
rect 21269 11781 21281 11815
rect 21315 11812 21327 11815
rect 21726 11812 21732 11824
rect 21315 11784 21732 11812
rect 21315 11781 21327 11784
rect 21269 11775 21327 11781
rect 21726 11772 21732 11784
rect 21784 11812 21790 11824
rect 22189 11815 22247 11821
rect 22189 11812 22201 11815
rect 21784 11784 22201 11812
rect 21784 11772 21790 11784
rect 22189 11781 22201 11784
rect 22235 11781 22247 11815
rect 22189 11775 22247 11781
rect 24213 11815 24271 11821
rect 24213 11781 24225 11815
rect 24259 11812 24271 11815
rect 24578 11812 24584 11824
rect 24259 11784 24584 11812
rect 24259 11781 24271 11784
rect 24213 11775 24271 11781
rect 24578 11772 24584 11784
rect 24636 11772 24642 11824
rect 19334 11704 19340 11756
rect 19392 11744 19398 11756
rect 19889 11747 19947 11753
rect 19889 11744 19901 11747
rect 19392 11716 19901 11744
rect 19392 11704 19398 11716
rect 19889 11713 19901 11716
rect 19935 11713 19947 11747
rect 19889 11707 19947 11713
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11713 20131 11747
rect 20438 11744 20444 11756
rect 20399 11716 20444 11744
rect 20073 11707 20131 11713
rect 20088 11676 20116 11707
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 21542 11744 21548 11756
rect 20772 11716 21548 11744
rect 20772 11704 20778 11716
rect 21542 11704 21548 11716
rect 21600 11704 21606 11756
rect 22756 11716 23520 11744
rect 21450 11676 21456 11688
rect 19260 11648 20116 11676
rect 21411 11648 21456 11676
rect 19153 11639 19211 11645
rect 21450 11636 21456 11648
rect 21508 11676 21514 11688
rect 22186 11676 22192 11688
rect 21508 11648 22192 11676
rect 21508 11636 21514 11648
rect 22186 11636 22192 11648
rect 22244 11636 22250 11688
rect 22370 11676 22376 11688
rect 22331 11648 22376 11676
rect 22370 11636 22376 11648
rect 22428 11676 22434 11688
rect 22756 11685 22784 11716
rect 23492 11685 23520 11716
rect 22741 11679 22799 11685
rect 22741 11676 22753 11679
rect 22428 11648 22753 11676
rect 22428 11636 22434 11648
rect 22741 11645 22753 11648
rect 22787 11645 22799 11679
rect 22741 11639 22799 11645
rect 23385 11679 23443 11685
rect 23385 11645 23397 11679
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 23477 11679 23535 11685
rect 23477 11645 23489 11679
rect 23523 11676 23535 11679
rect 23658 11676 23664 11688
rect 23523 11648 23664 11676
rect 23523 11645 23535 11648
rect 23477 11639 23535 11645
rect 22462 11608 22468 11620
rect 17236 11580 22468 11608
rect 22462 11568 22468 11580
rect 22520 11608 22526 11620
rect 23400 11608 23428 11639
rect 23658 11636 23664 11648
rect 23716 11636 23722 11688
rect 24302 11676 24308 11688
rect 24263 11648 24308 11676
rect 24302 11636 24308 11648
rect 24360 11636 24366 11688
rect 22520 11580 23428 11608
rect 22520 11568 22526 11580
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 13998 11540 14004 11552
rect 12943 11512 14004 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 14182 11500 14188 11552
rect 14240 11540 14246 11552
rect 14461 11543 14519 11549
rect 14461 11540 14473 11543
rect 14240 11512 14473 11540
rect 14240 11500 14246 11512
rect 14461 11509 14473 11512
rect 14507 11540 14519 11543
rect 14642 11540 14648 11552
rect 14507 11512 14648 11540
rect 14507 11509 14519 11512
rect 14461 11503 14519 11509
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 16172 11512 16405 11540
rect 16172 11500 16178 11512
rect 16393 11509 16405 11512
rect 16439 11509 16451 11543
rect 16393 11503 16451 11509
rect 16942 11500 16948 11552
rect 17000 11540 17006 11552
rect 17000 11512 17045 11540
rect 17000 11500 17006 11512
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 20714 11540 20720 11552
rect 17276 11512 20720 11540
rect 17276 11500 17282 11512
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 20809 11543 20867 11549
rect 20809 11509 20821 11543
rect 20855 11540 20867 11543
rect 21266 11540 21272 11552
rect 20855 11512 21272 11540
rect 20855 11509 20867 11512
rect 20809 11503 20867 11509
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 22925 11543 22983 11549
rect 22925 11509 22937 11543
rect 22971 11540 22983 11543
rect 23198 11540 23204 11552
rect 22971 11512 23204 11540
rect 22971 11509 22983 11512
rect 22925 11503 22983 11509
rect 23198 11500 23204 11512
rect 23256 11500 23262 11552
rect 23753 11543 23811 11549
rect 23753 11509 23765 11543
rect 23799 11540 23811 11543
rect 23842 11540 23848 11552
rect 23799 11512 23848 11540
rect 23799 11509 23811 11512
rect 23753 11503 23811 11509
rect 23842 11500 23848 11512
rect 23900 11500 23906 11552
rect 1104 11450 26128 11472
rect 1104 11398 5120 11450
rect 5172 11398 5184 11450
rect 5236 11398 5248 11450
rect 5300 11398 5312 11450
rect 5364 11398 5376 11450
rect 5428 11398 13462 11450
rect 13514 11398 13526 11450
rect 13578 11398 13590 11450
rect 13642 11398 13654 11450
rect 13706 11398 13718 11450
rect 13770 11398 21803 11450
rect 21855 11398 21867 11450
rect 21919 11398 21931 11450
rect 21983 11398 21995 11450
rect 22047 11398 22059 11450
rect 22111 11398 26128 11450
rect 1104 11376 26128 11398
rect 1762 11336 1768 11348
rect 1723 11308 1768 11336
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 8478 11336 8484 11348
rect 6880 11308 8484 11336
rect 6880 11296 6886 11308
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 8754 11336 8760 11348
rect 8667 11308 8760 11336
rect 8754 11296 8760 11308
rect 8812 11336 8818 11348
rect 9214 11336 9220 11348
rect 8812 11308 9220 11336
rect 8812 11296 8818 11308
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 10321 11339 10379 11345
rect 10321 11305 10333 11339
rect 10367 11336 10379 11339
rect 10594 11336 10600 11348
rect 10367 11308 10600 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 6730 11268 6736 11280
rect 6691 11240 6736 11268
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 8294 11268 8300 11280
rect 8255 11240 8300 11268
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 4764 11172 5365 11200
rect 4764 11160 4770 11172
rect 5353 11169 5365 11172
rect 5399 11169 5411 11203
rect 8938 11200 8944 11212
rect 5353 11163 5411 11169
rect 8404 11172 8944 11200
rect 3145 11135 3203 11141
rect 3145 11132 3157 11135
rect 2746 11104 3157 11132
rect 1670 10956 1676 11008
rect 1728 10996 1734 11008
rect 2746 10996 2774 11104
rect 3145 11101 3157 11104
rect 3191 11101 3203 11135
rect 3326 11132 3332 11144
rect 3287 11104 3332 11132
rect 3145 11095 3203 11101
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11132 3571 11135
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3559 11104 3801 11132
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 2900 11067 2958 11073
rect 2900 11033 2912 11067
rect 2946 11064 2958 11067
rect 3237 11067 3295 11073
rect 3237 11064 3249 11067
rect 2946 11036 3249 11064
rect 2946 11033 2958 11036
rect 2900 11027 2958 11033
rect 3237 11033 3249 11036
rect 3283 11033 3295 11067
rect 3237 11027 3295 11033
rect 1728 10968 2774 10996
rect 1728 10956 1734 10968
rect 3050 10956 3056 11008
rect 3108 10996 3114 11008
rect 3528 10996 3556 11095
rect 4890 11092 4896 11144
rect 4948 11132 4954 11144
rect 6730 11132 6736 11144
rect 4948 11104 6736 11132
rect 4948 11092 4954 11104
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 8404 11132 8432 11172
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 6963 11104 8432 11132
rect 8481 11135 8539 11141
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 8481 11101 8493 11135
rect 8527 11132 8539 11135
rect 8573 11135 8631 11141
rect 8573 11132 8585 11135
rect 8527 11104 8585 11132
rect 8527 11101 8539 11104
rect 8481 11095 8539 11101
rect 8573 11101 8585 11104
rect 8619 11101 8631 11135
rect 8573 11095 8631 11101
rect 9030 11092 9036 11144
rect 9088 11132 9094 11144
rect 9197 11135 9255 11141
rect 9197 11132 9209 11135
rect 9088 11104 9209 11132
rect 9088 11092 9094 11104
rect 9197 11101 9209 11104
rect 9243 11101 9255 11135
rect 9197 11095 9255 11101
rect 5626 11073 5632 11076
rect 5077 11067 5135 11073
rect 5077 11033 5089 11067
rect 5123 11064 5135 11067
rect 5123 11036 5580 11064
rect 5123 11033 5135 11036
rect 5077 11027 5135 11033
rect 3108 10968 3556 10996
rect 5552 10996 5580 11036
rect 5620 11027 5632 11073
rect 5684 11064 5690 11076
rect 5684 11036 5720 11064
rect 5626 11024 5632 11027
rect 5684 11024 5690 11036
rect 5810 11024 5816 11076
rect 5868 11064 5874 11076
rect 7162 11067 7220 11073
rect 5868 11036 6776 11064
rect 5868 11024 5874 11036
rect 5718 10996 5724 11008
rect 5552 10968 5724 10996
rect 3108 10956 3114 10968
rect 5718 10956 5724 10968
rect 5776 10956 5782 11008
rect 6748 10996 6776 11036
rect 7162 11033 7174 11067
rect 7208 11033 7220 11067
rect 7162 11027 7220 11033
rect 7177 10996 7205 11027
rect 8662 11024 8668 11076
rect 8720 11064 8726 11076
rect 10336 11064 10364 11299
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 15654 11336 15660 11348
rect 12544 11308 15424 11336
rect 15615 11308 15660 11336
rect 12544 11209 12572 11308
rect 13262 11268 13268 11280
rect 12636 11240 13268 11268
rect 12636 11209 12664 11240
rect 13262 11228 13268 11240
rect 13320 11228 13326 11280
rect 13372 11209 13400 11308
rect 13446 11228 13452 11280
rect 13504 11268 13510 11280
rect 13817 11271 13875 11277
rect 13817 11268 13829 11271
rect 13504 11240 13829 11268
rect 13504 11228 13510 11240
rect 13817 11237 13829 11240
rect 13863 11268 13875 11271
rect 14090 11268 14096 11280
rect 13863 11240 14096 11268
rect 13863 11237 13875 11240
rect 13817 11231 13875 11237
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 14461 11271 14519 11277
rect 14461 11237 14473 11271
rect 14507 11268 14519 11271
rect 15102 11268 15108 11280
rect 14507 11240 15108 11268
rect 14507 11237 14519 11240
rect 14461 11231 14519 11237
rect 15102 11228 15108 11240
rect 15160 11228 15166 11280
rect 15286 11228 15292 11280
rect 15344 11228 15350 11280
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11169 12587 11203
rect 12529 11163 12587 11169
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11169 12679 11203
rect 12621 11163 12679 11169
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11169 13415 11203
rect 13357 11163 13415 11169
rect 14274 11160 14280 11212
rect 14332 11200 14338 11212
rect 15304 11200 15332 11228
rect 15396 11209 15424 11308
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 18322 11336 18328 11348
rect 18283 11308 18328 11336
rect 18322 11296 18328 11308
rect 18380 11296 18386 11348
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 20438 11336 20444 11348
rect 18739 11308 20444 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 20990 11336 20996 11348
rect 20951 11308 20996 11336
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 22186 11296 22192 11348
rect 22244 11336 22250 11348
rect 22649 11339 22707 11345
rect 22649 11336 22661 11339
rect 22244 11308 22661 11336
rect 22244 11296 22250 11308
rect 22649 11305 22661 11308
rect 22695 11305 22707 11339
rect 22649 11299 22707 11305
rect 16574 11228 16580 11280
rect 16632 11228 16638 11280
rect 17037 11271 17095 11277
rect 17037 11237 17049 11271
rect 17083 11237 17095 11271
rect 17037 11231 17095 11237
rect 14332 11172 14872 11200
rect 14332 11160 14338 11172
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 12032 11104 12357 11132
rect 12032 11092 12038 11104
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12714 11135 12772 11141
rect 12714 11132 12726 11135
rect 12492 11104 12726 11132
rect 12492 11092 12498 11104
rect 12714 11101 12726 11104
rect 12760 11101 12772 11135
rect 12714 11095 12772 11101
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11132 12955 11135
rect 12986 11132 12992 11144
rect 12943 11104 12992 11132
rect 12943 11101 12955 11104
rect 12897 11095 12955 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13170 11132 13176 11144
rect 13131 11104 13176 11132
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 13320 11104 13365 11132
rect 13320 11092 13326 11104
rect 13446 11092 13452 11144
rect 13504 11141 13510 11144
rect 13504 11135 13553 11141
rect 13504 11101 13507 11135
rect 13541 11101 13553 11135
rect 14182 11132 14188 11144
rect 13504 11095 13553 11101
rect 13648 11104 14188 11132
rect 13504 11092 13510 11095
rect 8720 11036 10364 11064
rect 12161 11067 12219 11073
rect 8720 11024 8726 11036
rect 12161 11033 12173 11067
rect 12207 11064 12219 11067
rect 12802 11064 12808 11076
rect 12207 11036 12808 11064
rect 12207 11033 12219 11036
rect 12161 11027 12219 11033
rect 12802 11024 12808 11036
rect 12860 11024 12866 11076
rect 6748 10968 7205 10996
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 10226 10996 10232 11008
rect 8352 10968 10232 10996
rect 8352 10956 8358 10968
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 13648 10996 13676 11104
rect 14182 11092 14188 11104
rect 14240 11132 14246 11144
rect 14240 11104 14320 11132
rect 14240 11092 14246 11104
rect 13725 11067 13783 11073
rect 13725 11033 13737 11067
rect 13771 11064 13783 11067
rect 13998 11064 14004 11076
rect 13771 11036 14004 11064
rect 13771 11033 13783 11036
rect 13725 11027 13783 11033
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 14090 11024 14096 11076
rect 14148 11064 14154 11076
rect 14292 11073 14320 11104
rect 14844 11076 14872 11172
rect 15028 11172 15332 11200
rect 15381 11203 15439 11209
rect 15028 11141 15056 11172
rect 15381 11169 15393 11203
rect 15427 11200 15439 11203
rect 15746 11200 15752 11212
rect 15427 11172 15752 11200
rect 15427 11169 15439 11172
rect 15381 11163 15439 11169
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 16393 11203 16451 11209
rect 16393 11169 16405 11203
rect 16439 11200 16451 11203
rect 16439 11172 16473 11200
rect 16439 11169 16451 11172
rect 16393 11163 16451 11169
rect 15013 11135 15071 11141
rect 15013 11101 15025 11135
rect 15059 11101 15071 11135
rect 15194 11132 15200 11144
rect 15155 11104 15200 11132
rect 15013 11095 15071 11101
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 15565 11135 15623 11141
rect 15344 11104 15389 11132
rect 15344 11092 15350 11104
rect 15565 11101 15577 11135
rect 15611 11132 15623 11135
rect 15930 11132 15936 11144
rect 15611 11104 15936 11132
rect 15611 11101 15623 11104
rect 15565 11095 15623 11101
rect 15930 11092 15936 11104
rect 15988 11132 15994 11144
rect 16114 11132 16120 11144
rect 15988 11104 16120 11132
rect 15988 11092 15994 11104
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 16209 11135 16267 11141
rect 16209 11101 16221 11135
rect 16255 11132 16267 11135
rect 16408 11132 16436 11163
rect 16482 11132 16488 11144
rect 16255 11104 16488 11132
rect 16255 11101 16267 11104
rect 16209 11095 16267 11101
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 16592 11141 16620 11228
rect 16850 11200 16856 11212
rect 16684 11172 16856 11200
rect 16684 11141 16712 11172
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 16577 11135 16635 11141
rect 16577 11101 16589 11135
rect 16623 11101 16635 11135
rect 16577 11095 16635 11101
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 17052 11132 17080 11231
rect 17494 11228 17500 11280
rect 17552 11268 17558 11280
rect 17552 11240 17724 11268
rect 17552 11228 17558 11240
rect 17696 11209 17724 11240
rect 18874 11228 18880 11280
rect 18932 11268 18938 11280
rect 18969 11271 19027 11277
rect 18969 11268 18981 11271
rect 18932 11240 18981 11268
rect 18932 11228 18938 11240
rect 18969 11237 18981 11240
rect 19015 11237 19027 11271
rect 18969 11231 19027 11237
rect 19245 11271 19303 11277
rect 19245 11237 19257 11271
rect 19291 11268 19303 11271
rect 19334 11268 19340 11280
rect 19291 11240 19340 11268
rect 19291 11237 19303 11240
rect 19245 11231 19303 11237
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11169 17739 11203
rect 18782 11200 18788 11212
rect 17681 11163 17739 11169
rect 18340 11172 18788 11200
rect 18340 11141 18368 11172
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 18984 11200 19012 11231
rect 19334 11228 19340 11240
rect 19392 11228 19398 11280
rect 22370 11268 22376 11280
rect 20824 11240 21588 11268
rect 20824 11209 20852 11240
rect 19797 11203 19855 11209
rect 19797 11200 19809 11203
rect 18984 11172 19809 11200
rect 19797 11169 19809 11172
rect 19843 11200 19855 11203
rect 20809 11203 20867 11209
rect 20809 11200 20821 11203
rect 19843 11172 20821 11200
rect 19843 11169 19855 11172
rect 19797 11163 19855 11169
rect 20809 11169 20821 11172
rect 20855 11169 20867 11203
rect 20809 11163 20867 11169
rect 21174 11160 21180 11212
rect 21232 11200 21238 11212
rect 21560 11209 21588 11240
rect 22066 11240 22376 11268
rect 21453 11203 21511 11209
rect 21453 11200 21465 11203
rect 21232 11172 21465 11200
rect 21232 11160 21238 11172
rect 21453 11169 21465 11172
rect 21499 11169 21511 11203
rect 21453 11163 21511 11169
rect 21545 11203 21603 11209
rect 21545 11169 21557 11203
rect 21591 11200 21603 11203
rect 21821 11203 21879 11209
rect 21821 11200 21833 11203
rect 21591 11172 21833 11200
rect 21591 11169 21603 11172
rect 21545 11163 21603 11169
rect 21821 11169 21833 11172
rect 21867 11200 21879 11203
rect 22066 11200 22094 11240
rect 22370 11228 22376 11240
rect 22428 11228 22434 11280
rect 21867 11172 22094 11200
rect 22664 11200 22692 11299
rect 23290 11228 23296 11280
rect 23348 11268 23354 11280
rect 24397 11271 24455 11277
rect 24397 11268 24409 11271
rect 23348 11240 24409 11268
rect 23348 11228 23354 11240
rect 24397 11237 24409 11240
rect 24443 11237 24455 11271
rect 24397 11231 24455 11237
rect 23385 11203 23443 11209
rect 23385 11200 23397 11203
rect 22664 11172 23397 11200
rect 21867 11169 21879 11172
rect 21821 11163 21879 11169
rect 23385 11169 23397 11172
rect 23431 11200 23443 11203
rect 23661 11203 23719 11209
rect 23661 11200 23673 11203
rect 23431 11172 23673 11200
rect 23431 11169 23443 11172
rect 23385 11163 23443 11169
rect 23661 11169 23673 11172
rect 23707 11200 23719 11203
rect 24121 11203 24179 11209
rect 24121 11200 24133 11203
rect 23707 11172 24133 11200
rect 23707 11169 23719 11172
rect 23661 11163 23719 11169
rect 24121 11169 24133 11172
rect 24167 11200 24179 11203
rect 24302 11200 24308 11212
rect 24167 11172 24308 11200
rect 24167 11169 24179 11172
rect 24121 11163 24179 11169
rect 24302 11160 24308 11172
rect 24360 11160 24366 11212
rect 24670 11160 24676 11212
rect 24728 11200 24734 11212
rect 24857 11203 24915 11209
rect 24857 11200 24869 11203
rect 24728 11172 24869 11200
rect 24728 11160 24734 11172
rect 24857 11169 24869 11172
rect 24903 11169 24915 11203
rect 24857 11163 24915 11169
rect 24949 11203 25007 11209
rect 24949 11169 24961 11203
rect 24995 11169 25007 11203
rect 24949 11163 25007 11169
rect 17497 11135 17555 11141
rect 17497 11132 17509 11135
rect 16715 11104 16988 11132
rect 17052 11104 17509 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 14277 11067 14335 11073
rect 14148 11036 14193 11064
rect 14148 11024 14154 11036
rect 14277 11033 14289 11067
rect 14323 11033 14335 11067
rect 14642 11064 14648 11076
rect 14555 11036 14648 11064
rect 14277 11027 14335 11033
rect 14642 11024 14648 11036
rect 14700 11024 14706 11076
rect 14826 11064 14832 11076
rect 14787 11036 14832 11064
rect 14826 11024 14832 11036
rect 14884 11024 14890 11076
rect 16850 11064 16856 11076
rect 14936 11036 16856 11064
rect 10652 10968 13676 10996
rect 14660 10996 14688 11024
rect 14936 10996 14964 11036
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 16960 11064 16988 11104
rect 17497 11101 17509 11104
rect 17543 11101 17555 11135
rect 17497 11095 17555 11101
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11101 18383 11135
rect 18325 11095 18383 11101
rect 18414 11092 18420 11144
rect 18472 11132 18478 11144
rect 19610 11132 19616 11144
rect 18472 11104 18517 11132
rect 19523 11104 19616 11132
rect 18472 11092 18478 11104
rect 19610 11092 19616 11104
rect 19668 11132 19674 11144
rect 20530 11132 20536 11144
rect 19668 11104 20536 11132
rect 19668 11092 19674 11104
rect 20530 11092 20536 11104
rect 20588 11092 20594 11144
rect 21358 11132 21364 11144
rect 21319 11104 21364 11132
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 23198 11132 23204 11144
rect 23159 11104 23204 11132
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 23293 11135 23351 11141
rect 23293 11101 23305 11135
rect 23339 11132 23351 11135
rect 23566 11132 23572 11144
rect 23339 11104 23572 11132
rect 23339 11101 23351 11104
rect 23293 11095 23351 11101
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 24320 11132 24348 11160
rect 24964 11132 24992 11163
rect 24320 11104 24992 11132
rect 17589 11067 17647 11073
rect 17589 11064 17601 11067
rect 16960 11036 17601 11064
rect 17589 11033 17601 11036
rect 17635 11033 17647 11067
rect 18432 11064 18460 11092
rect 19705 11067 19763 11073
rect 19705 11064 19717 11067
rect 18432 11036 19717 11064
rect 17589 11027 17647 11033
rect 19705 11033 19717 11036
rect 19751 11033 19763 11067
rect 19705 11027 19763 11033
rect 14660 10968 14964 10996
rect 10652 10956 10658 10968
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 17129 10999 17187 11005
rect 17129 10996 17141 10999
rect 16632 10968 17141 10996
rect 16632 10956 16638 10968
rect 17129 10965 17141 10968
rect 17175 10965 17187 10999
rect 22830 10996 22836 11008
rect 22791 10968 22836 10996
rect 17129 10959 17187 10965
rect 22830 10956 22836 10968
rect 22888 10956 22894 11008
rect 24762 10996 24768 11008
rect 24723 10968 24768 10996
rect 24762 10956 24768 10968
rect 24820 10956 24826 11008
rect 1104 10906 26128 10928
rect 1104 10854 9291 10906
rect 9343 10854 9355 10906
rect 9407 10854 9419 10906
rect 9471 10854 9483 10906
rect 9535 10854 9547 10906
rect 9599 10854 17632 10906
rect 17684 10854 17696 10906
rect 17748 10854 17760 10906
rect 17812 10854 17824 10906
rect 17876 10854 17888 10906
rect 17940 10854 26128 10906
rect 1104 10832 26128 10854
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5810 10792 5816 10804
rect 5307 10764 5816 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 7190 10792 7196 10804
rect 7151 10764 7196 10792
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 8662 10792 8668 10804
rect 7760 10764 8668 10792
rect 7760 10736 7788 10764
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 10781 10795 10839 10801
rect 10781 10792 10793 10795
rect 9508 10764 10793 10792
rect 9508 10736 9536 10764
rect 10781 10761 10793 10764
rect 10827 10792 10839 10795
rect 10827 10764 15516 10792
rect 10827 10761 10839 10764
rect 10781 10755 10839 10761
rect 2124 10727 2182 10733
rect 2124 10693 2136 10727
rect 2170 10724 2182 10727
rect 2498 10724 2504 10736
rect 2170 10696 2504 10724
rect 2170 10693 2182 10696
rect 2124 10687 2182 10693
rect 2498 10684 2504 10696
rect 2556 10684 2562 10736
rect 3142 10684 3148 10736
rect 3200 10724 3206 10736
rect 3513 10727 3571 10733
rect 3513 10724 3525 10727
rect 3200 10696 3525 10724
rect 3200 10684 3206 10696
rect 3513 10693 3525 10696
rect 3559 10693 3571 10727
rect 3513 10687 3571 10693
rect 4246 10684 4252 10736
rect 4304 10724 4310 10736
rect 4982 10724 4988 10736
rect 4304 10696 4988 10724
rect 4304 10684 4310 10696
rect 3418 10656 3424 10668
rect 3379 10628 3424 10656
rect 3418 10616 3424 10628
rect 3476 10616 3482 10668
rect 3786 10656 3792 10668
rect 3747 10628 3792 10656
rect 3786 10616 3792 10628
rect 3844 10656 3850 10668
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3844 10628 4077 10656
rect 3844 10616 3850 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4341 10659 4399 10665
rect 4341 10656 4353 10659
rect 4212 10628 4353 10656
rect 4212 10616 4218 10628
rect 4341 10625 4353 10628
rect 4387 10625 4399 10659
rect 4522 10656 4528 10668
rect 4483 10628 4528 10656
rect 4341 10619 4399 10625
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 4632 10665 4660 10696
rect 4982 10684 4988 10696
rect 5040 10684 5046 10736
rect 5077 10727 5135 10733
rect 5077 10693 5089 10727
rect 5123 10724 5135 10727
rect 5626 10724 5632 10736
rect 5123 10696 5632 10724
rect 5123 10693 5135 10696
rect 5077 10687 5135 10693
rect 5626 10684 5632 10696
rect 5684 10684 5690 10736
rect 7742 10724 7748 10736
rect 5920 10696 7748 10724
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10625 4675 10659
rect 4890 10656 4896 10668
rect 4851 10628 4896 10656
rect 4617 10619 4675 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 5442 10656 5448 10668
rect 5399 10628 5448 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 5920 10665 5948 10696
rect 7742 10684 7748 10696
rect 7800 10684 7806 10736
rect 8294 10724 8300 10736
rect 7852 10696 8300 10724
rect 5905 10659 5963 10665
rect 5776 10628 5821 10656
rect 5776 10616 5782 10628
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 6822 10656 6828 10668
rect 6595 10628 6828 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10656 7343 10659
rect 7558 10656 7564 10668
rect 7331 10628 7564 10656
rect 7331 10625 7343 10628
rect 7285 10619 7343 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 7852 10665 7880 10696
rect 8294 10684 8300 10696
rect 8352 10724 8358 10736
rect 8352 10696 8984 10724
rect 8352 10684 8358 10696
rect 8956 10668 8984 10696
rect 9490 10684 9496 10736
rect 9548 10684 9554 10736
rect 12802 10684 12808 10736
rect 12860 10724 12866 10736
rect 13182 10727 13240 10733
rect 13182 10724 13194 10727
rect 12860 10696 13194 10724
rect 12860 10684 12866 10696
rect 13182 10693 13194 10696
rect 13228 10693 13240 10727
rect 13182 10687 13240 10693
rect 13998 10684 14004 10736
rect 14056 10724 14062 10736
rect 14746 10727 14804 10733
rect 14746 10724 14758 10727
rect 14056 10696 14758 10724
rect 14056 10684 14062 10696
rect 14746 10693 14758 10696
rect 14792 10693 14804 10727
rect 15488 10724 15516 10764
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 15841 10795 15899 10801
rect 15841 10792 15853 10795
rect 15620 10764 15853 10792
rect 15620 10752 15626 10764
rect 15841 10761 15853 10764
rect 15887 10761 15899 10795
rect 17034 10792 17040 10804
rect 16947 10764 17040 10792
rect 15841 10755 15899 10761
rect 17034 10752 17040 10764
rect 17092 10792 17098 10804
rect 17494 10792 17500 10804
rect 17092 10764 17500 10792
rect 17092 10752 17098 10764
rect 17494 10752 17500 10764
rect 17552 10792 17558 10804
rect 18785 10795 18843 10801
rect 18785 10792 18797 10795
rect 17552 10764 18797 10792
rect 17552 10752 17558 10764
rect 18785 10761 18797 10764
rect 18831 10761 18843 10795
rect 19334 10792 19340 10804
rect 19295 10764 19340 10792
rect 18785 10755 18843 10761
rect 18322 10724 18328 10736
rect 15488 10696 18328 10724
rect 14746 10687 14804 10693
rect 18322 10684 18328 10696
rect 18380 10684 18386 10736
rect 8110 10665 8116 10668
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 8104 10619 8116 10665
rect 8168 10656 8174 10668
rect 8168 10628 8204 10656
rect 8110 10616 8116 10619
rect 8168 10616 8174 10628
rect 8938 10616 8944 10668
rect 8996 10656 9002 10668
rect 9674 10665 9680 10668
rect 9401 10659 9459 10665
rect 9401 10656 9413 10659
rect 8996 10628 9413 10656
rect 8996 10616 9002 10628
rect 9401 10625 9413 10628
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 9668 10619 9680 10665
rect 9732 10656 9738 10668
rect 13449 10659 13507 10665
rect 9732 10628 9768 10656
rect 10428 10628 13400 10656
rect 9674 10616 9680 10619
rect 9732 10616 9738 10628
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 1857 10591 1915 10597
rect 1857 10588 1869 10591
rect 1728 10560 1869 10588
rect 1728 10548 1734 10560
rect 1857 10557 1869 10560
rect 1903 10557 1915 10591
rect 3602 10588 3608 10600
rect 3563 10560 3608 10588
rect 1857 10551 1915 10557
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 4709 10591 4767 10597
rect 4709 10557 4721 10591
rect 4755 10557 4767 10591
rect 4709 10551 4767 10557
rect 5537 10591 5595 10597
rect 5537 10557 5549 10591
rect 5583 10557 5595 10591
rect 5537 10551 5595 10557
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10588 5687 10591
rect 5994 10588 6000 10600
rect 5675 10560 6000 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 2866 10480 2872 10532
rect 2924 10520 2930 10532
rect 4157 10523 4215 10529
rect 4157 10520 4169 10523
rect 2924 10492 4169 10520
rect 2924 10480 2930 10492
rect 4157 10489 4169 10492
rect 4203 10489 4215 10523
rect 4157 10483 4215 10489
rect 4338 10480 4344 10532
rect 4396 10520 4402 10532
rect 4724 10520 4752 10551
rect 5552 10520 5580 10551
rect 5994 10548 6000 10560
rect 6052 10548 6058 10600
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6181 10591 6239 10597
rect 6181 10588 6193 10591
rect 6135 10560 6193 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 6181 10557 6193 10560
rect 6227 10588 6239 10591
rect 7466 10588 7472 10600
rect 6227 10560 7472 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 6365 10523 6423 10529
rect 6365 10520 6377 10523
rect 4396 10492 6377 10520
rect 4396 10480 4402 10492
rect 6365 10489 6377 10492
rect 6411 10489 6423 10523
rect 6365 10483 6423 10489
rect 3234 10452 3240 10464
rect 3195 10424 3240 10452
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 6086 10452 6092 10464
rect 4580 10424 6092 10452
rect 4580 10412 4586 10424
rect 6086 10412 6092 10424
rect 6144 10452 6150 10464
rect 6181 10455 6239 10461
rect 6181 10452 6193 10455
rect 6144 10424 6193 10452
rect 6144 10412 6150 10424
rect 6181 10421 6193 10424
rect 6227 10421 6239 10455
rect 6181 10415 6239 10421
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 9217 10455 9275 10461
rect 9217 10452 9229 10455
rect 8260 10424 9229 10452
rect 8260 10412 8266 10424
rect 9217 10421 9229 10424
rect 9263 10452 9275 10455
rect 10428 10452 10456 10628
rect 13372 10588 13400 10628
rect 13449 10625 13461 10659
rect 13495 10656 13507 10659
rect 14458 10656 14464 10668
rect 13495 10628 14464 10656
rect 13495 10625 13507 10628
rect 13449 10619 13507 10625
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 15102 10656 15108 10668
rect 15063 10628 15108 10656
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 15470 10616 15476 10668
rect 15528 10665 15534 10668
rect 15528 10659 15565 10665
rect 15553 10625 15565 10659
rect 15528 10619 15565 10625
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 16025 10659 16083 10665
rect 16025 10656 16037 10659
rect 15795 10628 16037 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 16025 10625 16037 10628
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 15528 10616 15534 10619
rect 15010 10588 15016 10600
rect 13372 10560 14044 10588
rect 14971 10560 15016 10588
rect 13446 10480 13452 10532
rect 13504 10480 13510 10532
rect 9263 10424 10456 10452
rect 9263 10421 9275 10424
rect 9217 10415 9275 10421
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12069 10455 12127 10461
rect 12069 10452 12081 10455
rect 12032 10424 12081 10452
rect 12032 10412 12038 10424
rect 12069 10421 12081 10424
rect 12115 10421 12127 10455
rect 12069 10415 12127 10421
rect 13078 10412 13084 10464
rect 13136 10452 13142 10464
rect 13464 10452 13492 10480
rect 13633 10455 13691 10461
rect 13633 10452 13645 10455
rect 13136 10424 13645 10452
rect 13136 10412 13142 10424
rect 13633 10421 13645 10424
rect 13679 10421 13691 10455
rect 14016 10452 14044 10560
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 15194 10588 15200 10600
rect 15155 10560 15200 10588
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 18800 10588 18828 10755
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 23474 10752 23480 10804
rect 23532 10792 23538 10804
rect 23753 10795 23811 10801
rect 23753 10792 23765 10795
rect 23532 10764 23765 10792
rect 23532 10752 23538 10764
rect 23753 10761 23765 10764
rect 23799 10761 23811 10795
rect 23753 10755 23811 10761
rect 24213 10795 24271 10801
rect 24213 10761 24225 10795
rect 24259 10792 24271 10795
rect 24762 10792 24768 10804
rect 24259 10764 24768 10792
rect 24259 10761 24271 10764
rect 24213 10755 24271 10761
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 19245 10727 19303 10733
rect 19245 10693 19257 10727
rect 19291 10724 19303 10727
rect 19610 10724 19616 10736
rect 19291 10696 19616 10724
rect 19291 10693 19303 10696
rect 19245 10687 19303 10693
rect 19610 10684 19616 10696
rect 19668 10684 19674 10736
rect 23385 10727 23443 10733
rect 23385 10693 23397 10727
rect 23431 10724 23443 10727
rect 23658 10724 23664 10736
rect 23431 10696 23664 10724
rect 23431 10693 23443 10696
rect 23385 10687 23443 10693
rect 23584 10597 23612 10696
rect 23658 10684 23664 10696
rect 23716 10684 23722 10736
rect 23845 10727 23903 10733
rect 23845 10693 23857 10727
rect 23891 10724 23903 10727
rect 24670 10724 24676 10736
rect 23891 10696 24676 10724
rect 23891 10693 23903 10696
rect 23845 10687 23903 10693
rect 24670 10684 24676 10696
rect 24728 10684 24734 10736
rect 19061 10591 19119 10597
rect 19061 10588 19073 10591
rect 18800 10560 19073 10588
rect 19061 10557 19073 10560
rect 19107 10557 19119 10591
rect 19061 10551 19119 10557
rect 23569 10591 23627 10597
rect 23569 10557 23581 10591
rect 23615 10557 23627 10591
rect 23569 10551 23627 10557
rect 18414 10520 18420 10532
rect 16868 10492 18420 10520
rect 16868 10452 16896 10492
rect 18414 10480 18420 10492
rect 18472 10480 18478 10532
rect 19702 10452 19708 10464
rect 14016 10424 16896 10452
rect 19663 10424 19708 10452
rect 13633 10415 13691 10421
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 1104 10362 26128 10384
rect 1104 10310 5120 10362
rect 5172 10310 5184 10362
rect 5236 10310 5248 10362
rect 5300 10310 5312 10362
rect 5364 10310 5376 10362
rect 5428 10310 13462 10362
rect 13514 10310 13526 10362
rect 13578 10310 13590 10362
rect 13642 10310 13654 10362
rect 13706 10310 13718 10362
rect 13770 10310 21803 10362
rect 21855 10310 21867 10362
rect 21919 10310 21931 10362
rect 21983 10310 21995 10362
rect 22047 10310 22059 10362
rect 22111 10310 26128 10362
rect 1104 10288 26128 10310
rect 2409 10251 2467 10257
rect 2409 10217 2421 10251
rect 2455 10248 2467 10251
rect 3326 10248 3332 10260
rect 2455 10220 3332 10248
rect 2455 10217 2467 10220
rect 2409 10211 2467 10217
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 7282 10208 7288 10260
rect 7340 10208 7346 10260
rect 8021 10251 8079 10257
rect 8021 10217 8033 10251
rect 8067 10248 8079 10251
rect 8110 10248 8116 10260
rect 8067 10220 8116 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 8757 10251 8815 10257
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 9585 10251 9643 10257
rect 8803 10220 9536 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 3237 10183 3295 10189
rect 3237 10180 3249 10183
rect 2792 10152 3249 10180
rect 2682 10112 2688 10124
rect 2643 10084 2688 10112
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 2792 10121 2820 10152
rect 3237 10149 3249 10152
rect 3283 10180 3295 10183
rect 3418 10180 3424 10192
rect 3283 10152 3424 10180
rect 3283 10149 3295 10152
rect 3237 10143 3295 10149
rect 3418 10140 3424 10152
rect 3476 10140 3482 10192
rect 7300 10180 7328 10208
rect 9508 10180 9536 10220
rect 9585 10217 9597 10251
rect 9631 10248 9643 10251
rect 9674 10248 9680 10260
rect 9631 10220 9680 10248
rect 9631 10217 9643 10220
rect 9585 10211 9643 10217
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 13354 10208 13360 10260
rect 13412 10248 13418 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 13412 10220 13553 10248
rect 13412 10208 13418 10220
rect 13541 10217 13553 10220
rect 13587 10217 13599 10251
rect 13906 10248 13912 10260
rect 13867 10220 13912 10248
rect 13541 10211 13599 10217
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 15197 10251 15255 10257
rect 15197 10217 15209 10251
rect 15243 10248 15255 10251
rect 15470 10248 15476 10260
rect 15243 10220 15476 10248
rect 15243 10217 15255 10220
rect 15197 10211 15255 10217
rect 15470 10208 15476 10220
rect 15528 10208 15534 10260
rect 10594 10180 10600 10192
rect 7300 10152 9444 10180
rect 9508 10152 10600 10180
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10081 2835 10115
rect 2777 10075 2835 10081
rect 2866 10072 2872 10124
rect 2924 10112 2930 10124
rect 3513 10115 3571 10121
rect 3513 10112 3525 10115
rect 2924 10084 2969 10112
rect 3068 10084 3525 10112
rect 2924 10072 2930 10084
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 3068 10053 3096 10084
rect 3513 10081 3525 10084
rect 3559 10081 3571 10115
rect 3513 10075 3571 10081
rect 3786 10072 3792 10124
rect 3844 10112 3850 10124
rect 4338 10112 4344 10124
rect 3844 10084 4108 10112
rect 4299 10084 4344 10112
rect 3844 10072 3850 10084
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 3234 10004 3240 10056
rect 3292 10044 3298 10056
rect 3329 10047 3387 10053
rect 3329 10044 3341 10047
rect 3292 10016 3341 10044
rect 3292 10004 3298 10016
rect 3329 10013 3341 10016
rect 3375 10013 3387 10047
rect 3602 10044 3608 10056
rect 3563 10016 3608 10044
rect 3329 10007 3387 10013
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 4080 10044 4108 10084
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 4706 10072 4712 10124
rect 4764 10112 4770 10124
rect 4801 10115 4859 10121
rect 4801 10112 4813 10115
rect 4764 10084 4813 10112
rect 4764 10072 4770 10084
rect 4801 10081 4813 10084
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10112 8355 10115
rect 8754 10112 8760 10124
rect 8343 10084 8760 10112
rect 8343 10081 8355 10084
rect 8297 10075 8355 10081
rect 4138 10047 4196 10053
rect 4138 10044 4150 10047
rect 4080 10016 4150 10044
rect 3973 10007 4031 10013
rect 4138 10013 4150 10016
rect 4184 10013 4196 10047
rect 4138 10007 4196 10013
rect 2608 9976 2636 10004
rect 3620 9976 3648 10004
rect 2608 9948 3648 9976
rect 3988 9976 4016 10007
rect 4246 10004 4252 10056
rect 4304 10044 4310 10056
rect 4522 10044 4528 10056
rect 4304 10016 4349 10044
rect 4483 10016 4528 10044
rect 4304 10004 4310 10016
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 4816 10044 4844 10075
rect 8754 10072 8760 10084
rect 8812 10112 8818 10124
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 8812 10084 9321 10112
rect 8812 10072 8818 10084
rect 9309 10081 9321 10084
rect 9355 10081 9367 10115
rect 9309 10075 9367 10081
rect 6365 10047 6423 10053
rect 6365 10044 6377 10047
rect 4816 10016 6377 10044
rect 6365 10013 6377 10016
rect 6411 10013 6423 10047
rect 6365 10007 6423 10013
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10044 8171 10047
rect 8202 10044 8208 10056
rect 8159 10016 8208 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8386 10044 8392 10056
rect 8347 10016 8392 10044
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 8478 10004 8484 10056
rect 8536 10044 8542 10056
rect 8662 10044 8668 10056
rect 8536 10016 8581 10044
rect 8623 10016 8668 10044
rect 8536 10004 8542 10016
rect 8662 10004 8668 10016
rect 8720 10044 8726 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8720 10016 8953 10044
rect 8720 10004 8726 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 9122 10044 9128 10056
rect 9083 10016 9128 10044
rect 8941 10007 8999 10013
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9416 10044 9444 10152
rect 10594 10140 10600 10152
rect 10652 10140 10658 10192
rect 23106 10180 23112 10192
rect 12176 10152 22094 10180
rect 23067 10152 23112 10180
rect 9858 10112 9864 10124
rect 9771 10084 9864 10112
rect 9858 10072 9864 10084
rect 9916 10112 9922 10124
rect 12176 10112 12204 10152
rect 14182 10112 14188 10124
rect 9916 10084 12204 10112
rect 14143 10084 14188 10112
rect 9916 10072 9922 10084
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 15102 10072 15108 10124
rect 15160 10072 15166 10124
rect 21450 10112 21456 10124
rect 21411 10084 21456 10112
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 9490 10044 9496 10056
rect 9403 10016 9496 10044
rect 9217 10007 9275 10013
rect 4614 9976 4620 9988
rect 3988 9948 4620 9976
rect 4172 9920 4200 9948
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 4709 9979 4767 9985
rect 4709 9945 4721 9979
rect 4755 9976 4767 9979
rect 5046 9979 5104 9985
rect 5046 9976 5058 9979
rect 4755 9948 5058 9976
rect 4755 9945 4767 9948
rect 4709 9939 4767 9945
rect 5046 9945 5058 9948
rect 5092 9945 5104 9979
rect 5046 9939 5104 9945
rect 5534 9936 5540 9988
rect 5592 9976 5598 9988
rect 6610 9979 6668 9985
rect 6610 9976 6622 9979
rect 5592 9948 6622 9976
rect 5592 9936 5598 9948
rect 6610 9945 6622 9948
rect 6656 9945 6668 9979
rect 8018 9976 8024 9988
rect 6610 9939 6668 9945
rect 6748 9948 8024 9976
rect 3786 9908 3792 9920
rect 3747 9880 3792 9908
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 4154 9868 4160 9920
rect 4212 9868 4218 9920
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 5626 9908 5632 9920
rect 4580 9880 5632 9908
rect 4580 9868 4586 9880
rect 5626 9868 5632 9880
rect 5684 9908 5690 9920
rect 6181 9911 6239 9917
rect 6181 9908 6193 9911
rect 5684 9880 6193 9908
rect 5684 9868 5690 9880
rect 6181 9877 6193 9880
rect 6227 9908 6239 9911
rect 6748 9908 6776 9948
rect 8018 9936 8024 9948
rect 8076 9936 8082 9988
rect 8404 9976 8432 10004
rect 9232 9976 9260 10007
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10013 13783 10047
rect 14090 10044 14096 10056
rect 14051 10016 14096 10044
rect 13725 10007 13783 10013
rect 8404 9948 9260 9976
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 13740 9976 13768 10007
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 14552 10047 14610 10053
rect 14552 10013 14564 10047
rect 14598 10044 14610 10047
rect 14921 10047 14979 10053
rect 14921 10044 14933 10047
rect 14598 10016 14933 10044
rect 14598 10013 14610 10016
rect 14552 10007 14610 10013
rect 14921 10013 14933 10016
rect 14967 10044 14979 10047
rect 15120 10044 15148 10072
rect 20714 10044 20720 10056
rect 14967 10016 15148 10044
rect 20675 10016 20720 10044
rect 14967 10013 14979 10016
rect 14921 10007 14979 10013
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 20898 10004 20904 10056
rect 20956 10044 20962 10056
rect 21177 10047 21235 10053
rect 21177 10044 21189 10047
rect 20956 10016 21189 10044
rect 20956 10004 20962 10016
rect 21177 10013 21189 10016
rect 21223 10013 21235 10047
rect 21177 10007 21235 10013
rect 22066 9988 22094 10152
rect 23106 10140 23112 10152
rect 23164 10140 23170 10192
rect 24578 10004 24584 10056
rect 24636 10044 24642 10056
rect 24946 10044 24952 10056
rect 24636 10016 24681 10044
rect 24907 10016 24952 10044
rect 24636 10004 24642 10016
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10044 25099 10047
rect 25590 10044 25596 10056
rect 25087 10016 25596 10044
rect 25087 10013 25099 10016
rect 25041 10007 25099 10013
rect 25590 10004 25596 10016
rect 25648 10004 25654 10056
rect 14737 9979 14795 9985
rect 14737 9976 14749 9979
rect 9732 9948 13676 9976
rect 13740 9948 14749 9976
rect 9732 9936 9738 9948
rect 6227 9880 6776 9908
rect 6227 9877 6239 9880
rect 6181 9871 6239 9877
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7745 9911 7803 9917
rect 7745 9908 7757 9911
rect 7064 9880 7757 9908
rect 7064 9868 7070 9880
rect 7745 9877 7757 9880
rect 7791 9908 7803 9911
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 7791 9880 8769 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 9858 9908 9864 9920
rect 9180 9880 9864 9908
rect 9180 9868 9186 9880
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 13648 9908 13676 9948
rect 14737 9945 14749 9948
rect 14783 9945 14795 9979
rect 14737 9939 14795 9945
rect 15105 9979 15163 9985
rect 15105 9945 15117 9979
rect 15151 9945 15163 9979
rect 22066 9948 22100 9988
rect 15105 9939 15163 9945
rect 15120 9908 15148 9939
rect 22094 9936 22100 9948
rect 22152 9936 22158 9988
rect 22646 9936 22652 9988
rect 22704 9976 22710 9988
rect 22833 9979 22891 9985
rect 22833 9976 22845 9979
rect 22704 9948 22845 9976
rect 22704 9936 22710 9948
rect 22833 9945 22845 9948
rect 22879 9945 22891 9979
rect 24394 9976 24400 9988
rect 24355 9948 24400 9976
rect 22833 9939 22891 9945
rect 24394 9936 24400 9948
rect 24452 9936 24458 9988
rect 15194 9908 15200 9920
rect 13648 9880 15200 9908
rect 15194 9868 15200 9880
rect 15252 9908 15258 9920
rect 15470 9908 15476 9920
rect 15252 9880 15476 9908
rect 15252 9868 15258 9880
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 20530 9908 20536 9920
rect 20491 9880 20536 9908
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 20806 9908 20812 9920
rect 20767 9880 20812 9908
rect 20806 9868 20812 9880
rect 20864 9868 20870 9920
rect 21269 9911 21327 9917
rect 21269 9877 21281 9911
rect 21315 9908 21327 9911
rect 22278 9908 22284 9920
rect 21315 9880 22284 9908
rect 21315 9877 21327 9880
rect 21269 9871 21327 9877
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 23198 9868 23204 9920
rect 23256 9908 23262 9920
rect 23293 9911 23351 9917
rect 23293 9908 23305 9911
rect 23256 9880 23305 9908
rect 23256 9868 23262 9880
rect 23293 9877 23305 9880
rect 23339 9877 23351 9911
rect 23293 9871 23351 9877
rect 1104 9818 26128 9840
rect 1104 9766 9291 9818
rect 9343 9766 9355 9818
rect 9407 9766 9419 9818
rect 9471 9766 9483 9818
rect 9535 9766 9547 9818
rect 9599 9766 17632 9818
rect 17684 9766 17696 9818
rect 17748 9766 17760 9818
rect 17812 9766 17824 9818
rect 17876 9766 17888 9818
rect 17940 9766 26128 9818
rect 1104 9744 26128 9766
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 3329 9707 3387 9713
rect 3329 9704 3341 9707
rect 2832 9676 3341 9704
rect 2832 9664 2838 9676
rect 3329 9673 3341 9676
rect 3375 9673 3387 9707
rect 5626 9704 5632 9716
rect 3329 9667 3387 9673
rect 4264 9676 5212 9704
rect 5587 9676 5632 9704
rect 2314 9596 2320 9648
rect 2372 9636 2378 9648
rect 3050 9636 3056 9648
rect 2372 9608 3056 9636
rect 2372 9596 2378 9608
rect 3050 9596 3056 9608
rect 3108 9596 3114 9648
rect 4062 9636 4068 9648
rect 3712 9608 4068 9636
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2547 9540 2697 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2866 9568 2872 9580
rect 2827 9540 2872 9568
rect 2685 9531 2743 9537
rect 2866 9528 2872 9540
rect 2924 9528 2930 9580
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9568 3203 9571
rect 3234 9568 3240 9580
rect 3191 9540 3240 9568
rect 3191 9537 3203 9540
rect 3145 9531 3203 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3712 9577 3740 9608
rect 4062 9596 4068 9608
rect 4120 9636 4126 9648
rect 4264 9636 4292 9676
rect 4120 9608 4292 9636
rect 4120 9596 4126 9608
rect 4338 9596 4344 9648
rect 4396 9636 4402 9648
rect 5184 9636 5212 9676
rect 5626 9664 5632 9676
rect 5684 9664 5690 9716
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 9674 9704 9680 9716
rect 6788 9676 9680 9704
rect 6788 9664 6794 9676
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 13173 9707 13231 9713
rect 13173 9704 13185 9707
rect 9824 9676 13185 9704
rect 9824 9664 9830 9676
rect 13173 9673 13185 9676
rect 13219 9704 13231 9707
rect 13354 9704 13360 9716
rect 13219 9676 13360 9704
rect 13219 9673 13231 9676
rect 13173 9667 13231 9673
rect 13354 9664 13360 9676
rect 13412 9664 13418 9716
rect 13906 9664 13912 9716
rect 13964 9704 13970 9716
rect 14366 9704 14372 9716
rect 13964 9676 14372 9704
rect 13964 9664 13970 9676
rect 14366 9664 14372 9676
rect 14424 9704 14430 9716
rect 14553 9707 14611 9713
rect 14553 9704 14565 9707
rect 14424 9676 14565 9704
rect 14424 9664 14430 9676
rect 14553 9673 14565 9676
rect 14599 9673 14611 9707
rect 14553 9667 14611 9673
rect 15381 9707 15439 9713
rect 15381 9673 15393 9707
rect 15427 9704 15439 9707
rect 15562 9704 15568 9716
rect 15427 9676 15568 9704
rect 15427 9673 15439 9676
rect 15381 9667 15439 9673
rect 15562 9664 15568 9676
rect 15620 9664 15626 9716
rect 22833 9707 22891 9713
rect 20732 9676 21864 9704
rect 5445 9639 5503 9645
rect 4396 9608 5120 9636
rect 5184 9608 5396 9636
rect 4396 9596 4402 9608
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9537 3755 9571
rect 4706 9568 4712 9580
rect 4667 9540 4712 9568
rect 3697 9531 3755 9537
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 5092 9577 5120 9608
rect 4892 9571 4950 9577
rect 4892 9568 4904 9571
rect 4856 9540 4904 9568
rect 4856 9528 4862 9540
rect 4892 9537 4904 9540
rect 4938 9537 4950 9571
rect 4892 9531 4950 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5368 9568 5396 9608
rect 5445 9605 5457 9639
rect 5491 9636 5503 9639
rect 5534 9636 5540 9648
rect 5491 9608 5540 9636
rect 5491 9605 5503 9608
rect 5445 9599 5503 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 5644 9608 10548 9636
rect 5644 9568 5672 9608
rect 5368 9540 5672 9568
rect 8021 9571 8079 9577
rect 5261 9531 5319 9537
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8297 9571 8355 9577
rect 8297 9568 8309 9571
rect 8067 9540 8309 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8297 9537 8309 9540
rect 8343 9568 8355 9571
rect 8570 9568 8576 9580
rect 8343 9540 8576 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 3605 9503 3663 9509
rect 2271 9472 2728 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9432 2467 9435
rect 2590 9432 2596 9444
rect 2455 9404 2596 9432
rect 2455 9401 2467 9404
rect 2409 9395 2467 9401
rect 2590 9392 2596 9404
rect 2648 9392 2654 9444
rect 2700 9432 2728 9472
rect 2976 9472 3280 9500
rect 2976 9432 3004 9472
rect 2700 9404 3004 9432
rect 3053 9435 3111 9441
rect 3053 9401 3065 9435
rect 3099 9432 3111 9435
rect 3142 9432 3148 9444
rect 3099 9404 3148 9432
rect 3099 9401 3111 9404
rect 3053 9395 3111 9401
rect 1946 9324 1952 9376
rect 2004 9364 2010 9376
rect 2041 9367 2099 9373
rect 2041 9364 2053 9367
rect 2004 9336 2053 9364
rect 2004 9324 2010 9336
rect 2041 9333 2053 9336
rect 2087 9333 2099 9367
rect 2041 9327 2099 9333
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 3068 9364 3096 9395
rect 3142 9392 3148 9404
rect 3200 9392 3206 9444
rect 3252 9432 3280 9472
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 3878 9500 3884 9512
rect 3651 9472 3884 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 3878 9460 3884 9472
rect 3936 9460 3942 9512
rect 4246 9460 4252 9512
rect 4304 9500 4310 9512
rect 4985 9503 5043 9509
rect 4985 9500 4997 9503
rect 4304 9472 4997 9500
rect 4304 9460 4310 9472
rect 4985 9469 4997 9472
rect 5031 9469 5043 9503
rect 5276 9500 5304 9531
rect 8570 9528 8576 9540
rect 8628 9528 8634 9580
rect 8846 9528 8852 9580
rect 8904 9568 8910 9580
rect 9677 9571 9735 9577
rect 9677 9568 9689 9571
rect 8904 9540 9689 9568
rect 8904 9528 8910 9540
rect 9677 9537 9689 9540
rect 9723 9537 9735 9571
rect 10318 9568 10324 9580
rect 10279 9540 10324 9568
rect 9677 9531 9735 9537
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10520 9568 10548 9608
rect 10778 9596 10784 9648
rect 10836 9636 10842 9648
rect 17954 9636 17960 9648
rect 10836 9608 17448 9636
rect 17915 9608 17960 9636
rect 10836 9596 10842 9608
rect 12158 9568 12164 9580
rect 10520 9540 12164 9568
rect 10413 9531 10471 9537
rect 7006 9500 7012 9512
rect 5276 9472 7012 9500
rect 4985 9463 5043 9469
rect 7006 9460 7012 9472
rect 7064 9460 7070 9512
rect 7098 9460 7104 9512
rect 7156 9500 7162 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 7156 9472 8401 9500
rect 7156 9460 7162 9472
rect 8389 9469 8401 9472
rect 8435 9500 8447 9503
rect 8478 9500 8484 9512
rect 8435 9472 8484 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 10336 9500 10364 9528
rect 9876 9472 10364 9500
rect 4430 9432 4436 9444
rect 3252 9404 4436 9432
rect 4430 9392 4436 9404
rect 4488 9392 4494 9444
rect 4706 9392 4712 9444
rect 4764 9432 4770 9444
rect 7837 9435 7895 9441
rect 7837 9432 7849 9435
rect 4764 9404 7849 9432
rect 4764 9392 4770 9404
rect 7837 9401 7849 9404
rect 7883 9432 7895 9435
rect 8662 9432 8668 9444
rect 7883 9404 8668 9432
rect 7883 9401 7895 9404
rect 7837 9395 7895 9401
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 9876 9441 9904 9472
rect 9861 9435 9919 9441
rect 9861 9401 9873 9435
rect 9907 9401 9919 9435
rect 10226 9432 10232 9444
rect 10187 9404 10232 9432
rect 9861 9395 9919 9401
rect 10226 9392 10232 9404
rect 10284 9392 10290 9444
rect 3694 9364 3700 9376
rect 2832 9336 3096 9364
rect 3655 9336 3700 9364
rect 2832 9324 2838 9336
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4522 9364 4528 9376
rect 4483 9336 4528 9364
rect 4522 9324 4528 9336
rect 4580 9364 4586 9376
rect 4798 9364 4804 9376
rect 4580 9336 4804 9364
rect 4580 9324 4586 9336
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 7926 9364 7932 9376
rect 5500 9336 7932 9364
rect 5500 9324 5506 9336
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 8110 9364 8116 9376
rect 8071 9336 8116 9364
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 8202 9324 8208 9376
rect 8260 9364 8266 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 8260 9336 9965 9364
rect 8260 9324 8266 9336
rect 9953 9333 9965 9336
rect 9999 9364 10011 9367
rect 10428 9364 10456 9531
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9568 13323 9571
rect 13354 9568 13360 9580
rect 13311 9540 13360 9568
rect 13311 9537 13323 9540
rect 13265 9531 13323 9537
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 14182 9528 14188 9580
rect 14240 9568 14246 9580
rect 14645 9571 14703 9577
rect 14645 9568 14657 9571
rect 14240 9540 14657 9568
rect 14240 9528 14246 9540
rect 14645 9537 14657 9540
rect 14691 9537 14703 9571
rect 15470 9568 15476 9580
rect 15431 9540 15476 9568
rect 14645 9531 14703 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 17310 9568 17316 9580
rect 17271 9540 17316 9568
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 17420 9568 17448 9608
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 20732 9636 20760 9676
rect 18064 9608 20760 9636
rect 20809 9639 20867 9645
rect 18064 9568 18092 9608
rect 20809 9605 20821 9639
rect 20855 9636 20867 9639
rect 21082 9636 21088 9648
rect 20855 9608 21088 9636
rect 20855 9605 20867 9608
rect 20809 9599 20867 9605
rect 21082 9596 21088 9608
rect 21140 9596 21146 9648
rect 21637 9639 21695 9645
rect 21637 9636 21649 9639
rect 21376 9608 21649 9636
rect 17420 9540 18092 9568
rect 20622 9528 20628 9580
rect 20680 9568 20686 9580
rect 21376 9568 21404 9608
rect 21637 9605 21649 9608
rect 21683 9636 21695 9639
rect 21726 9636 21732 9648
rect 21683 9608 21732 9636
rect 21683 9605 21695 9608
rect 21637 9599 21695 9605
rect 21726 9596 21732 9608
rect 21784 9596 21790 9648
rect 21836 9636 21864 9676
rect 22833 9673 22845 9707
rect 22879 9704 22891 9707
rect 23106 9704 23112 9716
rect 22879 9676 23112 9704
rect 22879 9673 22891 9676
rect 22833 9667 22891 9673
rect 23106 9664 23112 9676
rect 23164 9664 23170 9716
rect 24946 9664 24952 9716
rect 25004 9704 25010 9716
rect 25041 9707 25099 9713
rect 25041 9704 25053 9707
rect 25004 9676 25053 9704
rect 25004 9664 25010 9676
rect 25041 9673 25053 9676
rect 25087 9673 25099 9707
rect 25041 9667 25099 9673
rect 22186 9636 22192 9648
rect 21836 9608 22192 9636
rect 22186 9596 22192 9608
rect 22244 9596 22250 9648
rect 23293 9639 23351 9645
rect 23293 9605 23305 9639
rect 23339 9636 23351 9639
rect 24394 9636 24400 9648
rect 23339 9608 24400 9636
rect 23339 9605 23351 9608
rect 23293 9599 23351 9605
rect 24394 9596 24400 9608
rect 24452 9596 24458 9648
rect 25056 9636 25084 9667
rect 25409 9639 25467 9645
rect 25409 9636 25421 9639
rect 25056 9608 25421 9636
rect 25409 9605 25421 9608
rect 25455 9605 25467 9639
rect 25409 9599 25467 9605
rect 20680 9540 21404 9568
rect 21453 9571 21511 9577
rect 20680 9528 20686 9540
rect 21453 9537 21465 9571
rect 21499 9568 21511 9571
rect 21542 9568 21548 9580
rect 21499 9540 21548 9568
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 21542 9528 21548 9540
rect 21600 9528 21606 9580
rect 23201 9571 23259 9577
rect 23201 9537 23213 9571
rect 23247 9537 23259 9571
rect 23201 9531 23259 9537
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 13998 9500 14004 9512
rect 13863 9472 14004 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 13998 9460 14004 9472
rect 14056 9500 14062 9512
rect 14093 9503 14151 9509
rect 14093 9500 14105 9503
rect 14056 9472 14105 9500
rect 14056 9460 14062 9472
rect 14093 9469 14105 9472
rect 14139 9500 14151 9503
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14139 9472 14841 9500
rect 14139 9469 14151 9472
rect 14093 9463 14151 9469
rect 14829 9469 14841 9472
rect 14875 9500 14887 9503
rect 15657 9503 15715 9509
rect 15657 9500 15669 9503
rect 14875 9472 15669 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 15657 9469 15669 9472
rect 15703 9500 15715 9503
rect 16666 9500 16672 9512
rect 15703 9472 16672 9500
rect 15703 9469 15715 9472
rect 15657 9463 15715 9469
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 18046 9460 18052 9472
rect 18104 9460 18110 9512
rect 18141 9503 18199 9509
rect 18141 9469 18153 9503
rect 18187 9469 18199 9503
rect 19794 9500 19800 9512
rect 19755 9472 19800 9500
rect 18141 9463 18199 9469
rect 13357 9435 13415 9441
rect 13357 9401 13369 9435
rect 13403 9432 13415 9435
rect 13906 9432 13912 9444
rect 13403 9404 13912 9432
rect 13403 9401 13415 9404
rect 13357 9395 13415 9401
rect 13906 9392 13912 9404
rect 13964 9432 13970 9444
rect 14918 9432 14924 9444
rect 13964 9404 14924 9432
rect 13964 9392 13970 9404
rect 14918 9392 14924 9404
rect 14976 9392 14982 9444
rect 17218 9392 17224 9444
rect 17276 9432 17282 9444
rect 17589 9435 17647 9441
rect 17589 9432 17601 9435
rect 17276 9404 17601 9432
rect 17276 9392 17282 9404
rect 17589 9401 17601 9404
rect 17635 9401 17647 9435
rect 17589 9395 17647 9401
rect 17954 9392 17960 9444
rect 18012 9432 18018 9444
rect 18156 9432 18184 9463
rect 19794 9460 19800 9472
rect 19852 9460 19858 9512
rect 20898 9500 20904 9512
rect 20859 9472 20904 9500
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 21085 9503 21143 9509
rect 21085 9469 21097 9503
rect 21131 9469 21143 9503
rect 23216 9500 23244 9531
rect 23474 9528 23480 9580
rect 23532 9568 23538 9580
rect 23917 9571 23975 9577
rect 23917 9568 23929 9571
rect 23532 9540 23929 9568
rect 23532 9528 23538 9540
rect 23917 9537 23929 9540
rect 23963 9537 23975 9571
rect 25590 9568 25596 9580
rect 25551 9540 25596 9568
rect 23917 9531 23975 9537
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 23290 9500 23296 9512
rect 23216 9472 23296 9500
rect 21085 9463 21143 9469
rect 18012 9404 18184 9432
rect 20165 9435 20223 9441
rect 18012 9392 18018 9404
rect 20165 9401 20177 9435
rect 20211 9432 20223 9435
rect 20441 9435 20499 9441
rect 20441 9432 20453 9435
rect 20211 9404 20453 9432
rect 20211 9401 20223 9404
rect 20165 9395 20223 9401
rect 20441 9401 20453 9404
rect 20487 9401 20499 9435
rect 21100 9432 21128 9463
rect 23290 9460 23296 9472
rect 23348 9460 23354 9512
rect 23382 9460 23388 9512
rect 23440 9500 23446 9512
rect 23658 9500 23664 9512
rect 23440 9472 23485 9500
rect 23619 9472 23664 9500
rect 23440 9460 23446 9472
rect 23658 9460 23664 9472
rect 23716 9460 23722 9512
rect 21450 9432 21456 9444
rect 21100 9404 21456 9432
rect 20441 9395 20499 9401
rect 21450 9392 21456 9404
rect 21508 9432 21514 9444
rect 23400 9432 23428 9460
rect 21508 9404 23428 9432
rect 25225 9435 25283 9441
rect 21508 9392 21514 9404
rect 25225 9401 25237 9435
rect 25271 9401 25283 9435
rect 25225 9395 25283 9401
rect 10686 9364 10692 9376
rect 9999 9336 10692 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 11609 9367 11667 9373
rect 11609 9333 11621 9367
rect 11655 9364 11667 9367
rect 11882 9364 11888 9376
rect 11655 9336 11888 9364
rect 11655 9333 11667 9336
rect 11609 9327 11667 9333
rect 11882 9324 11888 9336
rect 11940 9364 11946 9376
rect 12250 9364 12256 9376
rect 11940 9336 12256 9364
rect 11940 9324 11946 9336
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 14185 9367 14243 9373
rect 14185 9333 14197 9367
rect 14231 9364 14243 9367
rect 14458 9364 14464 9376
rect 14231 9336 14464 9364
rect 14231 9333 14243 9336
rect 14185 9327 14243 9333
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 15013 9367 15071 9373
rect 15013 9333 15025 9367
rect 15059 9364 15071 9367
rect 15286 9364 15292 9376
rect 15059 9336 15292 9364
rect 15059 9333 15071 9336
rect 15013 9327 15071 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 20257 9367 20315 9373
rect 20257 9333 20269 9367
rect 20303 9364 20315 9367
rect 20714 9364 20720 9376
rect 20303 9336 20720 9364
rect 20303 9333 20315 9336
rect 20257 9327 20315 9333
rect 20714 9324 20720 9336
rect 20772 9324 20778 9376
rect 21358 9364 21364 9376
rect 21319 9336 21364 9364
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 22922 9324 22928 9376
rect 22980 9364 22986 9376
rect 24578 9364 24584 9376
rect 22980 9336 24584 9364
rect 22980 9324 22986 9336
rect 24578 9324 24584 9336
rect 24636 9364 24642 9376
rect 25240 9364 25268 9395
rect 24636 9336 25268 9364
rect 24636 9324 24642 9336
rect 1104 9274 26128 9296
rect 1104 9222 5120 9274
rect 5172 9222 5184 9274
rect 5236 9222 5248 9274
rect 5300 9222 5312 9274
rect 5364 9222 5376 9274
rect 5428 9222 13462 9274
rect 13514 9222 13526 9274
rect 13578 9222 13590 9274
rect 13642 9222 13654 9274
rect 13706 9222 13718 9274
rect 13770 9222 21803 9274
rect 21855 9222 21867 9274
rect 21919 9222 21931 9274
rect 21983 9222 21995 9274
rect 22047 9222 22059 9274
rect 22111 9222 26128 9274
rect 1104 9200 26128 9222
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 3789 9163 3847 9169
rect 3789 9160 3801 9163
rect 3660 9132 3801 9160
rect 3660 9120 3666 9132
rect 3789 9129 3801 9132
rect 3835 9129 3847 9163
rect 3789 9123 3847 9129
rect 4249 9163 4307 9169
rect 4249 9129 4261 9163
rect 4295 9160 4307 9163
rect 11054 9160 11060 9172
rect 4295 9132 11060 9160
rect 4295 9129 4307 9132
rect 4249 9123 4307 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 12713 9163 12771 9169
rect 12713 9129 12725 9163
rect 12759 9160 12771 9163
rect 13354 9160 13360 9172
rect 12759 9132 13360 9160
rect 12759 9129 12771 9132
rect 12713 9123 12771 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13633 9163 13691 9169
rect 13633 9129 13645 9163
rect 13679 9160 13691 9163
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 13679 9132 13737 9160
rect 13679 9129 13691 9132
rect 13633 9123 13691 9129
rect 13725 9129 13737 9132
rect 13771 9160 13783 9163
rect 13998 9160 14004 9172
rect 13771 9132 14004 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 17034 9160 17040 9172
rect 15295 9132 17040 9160
rect 3053 9095 3111 9101
rect 3053 9061 3065 9095
rect 3099 9061 3111 9095
rect 3053 9055 3111 9061
rect 10597 9095 10655 9101
rect 10597 9061 10609 9095
rect 10643 9092 10655 9095
rect 10962 9092 10968 9104
rect 10643 9064 10968 9092
rect 10643 9061 10655 9064
rect 10597 9055 10655 9061
rect 1670 9024 1676 9036
rect 1631 8996 1676 9024
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 3068 9024 3096 9055
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 13906 9092 13912 9104
rect 12820 9064 13912 9092
rect 3878 9024 3884 9036
rect 3068 8996 3884 9024
rect 3878 8984 3884 8996
rect 3936 8984 3942 9036
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 7098 9024 7104 9036
rect 4028 8996 7104 9024
rect 4028 8984 4034 8996
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 9030 9024 9036 9036
rect 8536 8996 9036 9024
rect 8536 8984 8542 8996
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 12820 9033 12848 9064
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 14829 9095 14887 9101
rect 14200 9064 14504 9092
rect 12805 9027 12863 9033
rect 12805 8993 12817 9027
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 12897 9027 12955 9033
rect 12897 8993 12909 9027
rect 12943 9024 12955 9027
rect 13725 9027 13783 9033
rect 13725 9024 13737 9027
rect 12943 8996 13737 9024
rect 12943 8993 12955 8996
rect 12897 8987 12955 8993
rect 13725 8993 13737 8996
rect 13771 8993 13783 9027
rect 13725 8987 13783 8993
rect 13817 9027 13875 9033
rect 13817 8993 13829 9027
rect 13863 9024 13875 9027
rect 13998 9024 14004 9036
rect 13863 8996 14004 9024
rect 13863 8993 13875 8996
rect 13817 8987 13875 8993
rect 1946 8965 1952 8968
rect 1940 8956 1952 8965
rect 1907 8928 1952 8956
rect 1940 8919 1952 8928
rect 1946 8916 1952 8919
rect 2004 8916 2010 8968
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3694 8956 3700 8968
rect 3108 8928 3700 8956
rect 3108 8916 3114 8928
rect 3694 8916 3700 8928
rect 3752 8956 3758 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3752 8928 3801 8956
rect 3752 8916 3758 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8956 7343 8959
rect 8294 8956 8300 8968
rect 7331 8928 8300 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 3234 8848 3240 8900
rect 3292 8888 3298 8900
rect 4080 8888 4108 8919
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 8904 8928 9137 8956
rect 8904 8916 8910 8928
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8956 9367 8959
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 9355 8928 10241 8956
rect 9355 8925 9367 8928
rect 9309 8919 9367 8925
rect 10229 8925 10241 8928
rect 10275 8956 10287 8959
rect 10870 8956 10876 8968
rect 10275 8928 10876 8956
rect 10275 8925 10287 8928
rect 10229 8919 10287 8925
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8925 12035 8959
rect 12250 8956 12256 8968
rect 12211 8928 12256 8956
rect 11977 8919 12035 8925
rect 3292 8860 4108 8888
rect 7552 8891 7610 8897
rect 3292 8848 3298 8860
rect 7552 8857 7564 8891
rect 7598 8888 7610 8891
rect 8018 8888 8024 8900
rect 7598 8860 8024 8888
rect 7598 8857 7610 8860
rect 7552 8851 7610 8857
rect 8018 8848 8024 8860
rect 8076 8848 8082 8900
rect 8938 8888 8944 8900
rect 8128 8860 8944 8888
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 8128 8820 8156 8860
rect 8938 8848 8944 8860
rect 8996 8848 9002 8900
rect 9214 8848 9220 8900
rect 9272 8888 9278 8900
rect 9861 8891 9919 8897
rect 9861 8888 9873 8891
rect 9272 8860 9873 8888
rect 9272 8848 9278 8860
rect 9861 8857 9873 8860
rect 9907 8857 9919 8891
rect 9861 8851 9919 8857
rect 10045 8891 10103 8897
rect 10045 8857 10057 8891
rect 10091 8888 10103 8891
rect 11146 8888 11152 8900
rect 10091 8860 11152 8888
rect 10091 8857 10103 8860
rect 10045 8851 10103 8857
rect 11146 8848 11152 8860
rect 11204 8848 11210 8900
rect 11606 8848 11612 8900
rect 11664 8888 11670 8900
rect 11710 8891 11768 8897
rect 11710 8888 11722 8891
rect 11664 8860 11722 8888
rect 11664 8848 11670 8860
rect 11710 8857 11722 8860
rect 11756 8857 11768 8891
rect 11992 8888 12020 8919
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 12618 8916 12624 8968
rect 12676 8956 12682 8968
rect 12912 8956 12940 8987
rect 13998 8984 14004 8996
rect 14056 9024 14062 9036
rect 14200 9033 14228 9064
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 14056 8996 14197 9024
rect 14056 8984 14062 8996
rect 14185 8993 14197 8996
rect 14231 8993 14243 9027
rect 14366 9024 14372 9036
rect 14327 8996 14372 9024
rect 14185 8987 14243 8993
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 14476 9024 14504 9064
rect 14829 9061 14841 9095
rect 14875 9092 14887 9095
rect 15194 9092 15200 9104
rect 14875 9064 15200 9092
rect 14875 9061 14887 9064
rect 14829 9055 14887 9061
rect 15194 9052 15200 9064
rect 15252 9052 15258 9104
rect 15105 9027 15163 9033
rect 15105 9024 15117 9027
rect 14476 8996 15117 9024
rect 15105 8993 15117 8996
rect 15151 9024 15163 9027
rect 15295 9024 15323 9132
rect 17034 9120 17040 9132
rect 17092 9120 17098 9172
rect 20070 9160 20076 9172
rect 20031 9132 20076 9160
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 21450 9160 21456 9172
rect 20732 9132 21456 9160
rect 15151 8996 15323 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 17954 8984 17960 9036
rect 18012 9024 18018 9036
rect 18693 9027 18751 9033
rect 18693 9024 18705 9027
rect 18012 8996 18705 9024
rect 18012 8984 18018 8996
rect 18693 8993 18705 8996
rect 18739 8993 18751 9027
rect 18693 8987 18751 8993
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19797 9027 19855 9033
rect 19797 9024 19809 9027
rect 19392 8996 19809 9024
rect 19392 8984 19398 8996
rect 19797 8993 19809 8996
rect 19843 8993 19855 9027
rect 19797 8987 19855 8993
rect 20533 9027 20591 9033
rect 20533 8993 20545 9027
rect 20579 9024 20591 9027
rect 20732 9024 20760 9132
rect 21450 9120 21456 9132
rect 21508 9120 21514 9172
rect 23385 9163 23443 9169
rect 23385 9129 23397 9163
rect 23431 9160 23443 9163
rect 23474 9160 23480 9172
rect 23431 9132 23480 9160
rect 23431 9129 23443 9132
rect 23385 9123 23443 9129
rect 23474 9120 23480 9132
rect 23532 9120 23538 9172
rect 22097 9095 22155 9101
rect 22097 9061 22109 9095
rect 22143 9061 22155 9095
rect 22278 9092 22284 9104
rect 22239 9064 22284 9092
rect 22097 9055 22155 9061
rect 20579 8996 20760 9024
rect 20579 8993 20591 8996
rect 20533 8987 20591 8993
rect 22002 8984 22008 9036
rect 22060 9024 22066 9036
rect 22112 9024 22140 9055
rect 22278 9052 22284 9064
rect 22336 9052 22342 9104
rect 22833 9027 22891 9033
rect 22833 9024 22845 9027
rect 22060 8996 22845 9024
rect 22060 8984 22066 8996
rect 22833 8993 22845 8996
rect 22879 8993 22891 9027
rect 22833 8987 22891 8993
rect 23382 8984 23388 9036
rect 23440 9024 23446 9036
rect 24029 9027 24087 9033
rect 24029 9024 24041 9027
rect 23440 8996 24041 9024
rect 23440 8984 23446 8996
rect 24029 8993 24041 8996
rect 24075 8993 24087 9027
rect 24029 8987 24087 8993
rect 24949 9027 25007 9033
rect 24949 8993 24961 9027
rect 24995 9024 25007 9027
rect 24995 8996 25360 9024
rect 24995 8993 25007 8996
rect 24949 8987 25007 8993
rect 13078 8956 13084 8968
rect 12676 8928 12940 8956
rect 13039 8928 13084 8956
rect 12676 8916 12682 8928
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8956 13231 8959
rect 13354 8956 13360 8968
rect 13219 8928 13360 8956
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 14458 8956 14464 8968
rect 14419 8928 14464 8956
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 16393 8959 16451 8965
rect 16393 8956 16405 8959
rect 15028 8928 16405 8956
rect 15028 8900 15056 8928
rect 16393 8925 16405 8928
rect 16439 8925 16451 8959
rect 16393 8919 16451 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8956 18567 8959
rect 19058 8956 19064 8968
rect 18555 8928 19064 8956
rect 18555 8925 18567 8928
rect 18509 8919 18567 8925
rect 19058 8916 19064 8928
rect 19116 8916 19122 8968
rect 20254 8965 20260 8968
rect 19487 8959 19545 8965
rect 19487 8925 19499 8959
rect 19533 8956 19545 8959
rect 19889 8959 19947 8965
rect 19533 8928 19840 8956
rect 19533 8925 19545 8928
rect 19487 8919 19545 8925
rect 15010 8888 15016 8900
rect 11992 8860 15016 8888
rect 11710 8851 11768 8857
rect 15010 8848 15016 8860
rect 15068 8848 15074 8900
rect 15286 8888 15292 8900
rect 15247 8860 15292 8888
rect 15286 8848 15292 8860
rect 15344 8848 15350 8900
rect 15562 8888 15568 8900
rect 15488 8860 15568 8888
rect 6972 8792 8156 8820
rect 6972 8780 6978 8792
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 8665 8823 8723 8829
rect 8665 8820 8677 8823
rect 8628 8792 8677 8820
rect 8628 8780 8634 8792
rect 8665 8789 8677 8792
rect 8711 8789 8723 8823
rect 8665 8783 8723 8789
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 12069 8823 12127 8829
rect 12069 8820 12081 8823
rect 11848 8792 12081 8820
rect 11848 8780 11854 8792
rect 12069 8789 12081 8792
rect 12115 8789 12127 8823
rect 12069 8783 12127 8789
rect 12529 8823 12587 8829
rect 12529 8789 12541 8823
rect 12575 8820 12587 8823
rect 13170 8820 13176 8832
rect 12575 8792 13176 8820
rect 12575 8789 12587 8792
rect 12529 8783 12587 8789
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13354 8820 13360 8832
rect 13315 8792 13360 8820
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 15197 8823 15255 8829
rect 15197 8789 15209 8823
rect 15243 8820 15255 8823
rect 15488 8820 15516 8860
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 15838 8848 15844 8900
rect 15896 8888 15902 8900
rect 16638 8891 16696 8897
rect 16638 8888 16650 8891
rect 15896 8860 16650 8888
rect 15896 8848 15902 8860
rect 16638 8857 16650 8860
rect 16684 8857 16696 8891
rect 16638 8851 16696 8857
rect 18601 8891 18659 8897
rect 18601 8857 18613 8891
rect 18647 8888 18659 8891
rect 19245 8891 19303 8897
rect 19245 8888 19257 8891
rect 18647 8860 19257 8888
rect 18647 8857 18659 8860
rect 18601 8851 18659 8857
rect 19245 8857 19257 8860
rect 19291 8857 19303 8891
rect 19812 8888 19840 8928
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 20223 8959 20260 8965
rect 20223 8956 20235 8959
rect 19935 8928 20235 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 20223 8925 20235 8928
rect 20223 8919 20260 8925
rect 20254 8916 20260 8919
rect 20312 8916 20318 8968
rect 20622 8956 20628 8968
rect 20583 8928 20628 8956
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 20717 8959 20775 8965
rect 20717 8925 20729 8959
rect 20763 8956 20775 8959
rect 20763 8928 21404 8956
rect 20763 8925 20775 8928
rect 20717 8919 20775 8925
rect 19978 8888 19984 8900
rect 19812 8860 19984 8888
rect 19245 8851 19303 8857
rect 19978 8848 19984 8860
rect 20036 8848 20042 8900
rect 15654 8820 15660 8832
rect 15243 8792 15516 8820
rect 15615 8792 15660 8820
rect 15243 8789 15255 8792
rect 15197 8783 15255 8789
rect 15654 8780 15660 8792
rect 15712 8780 15718 8832
rect 17402 8780 17408 8832
rect 17460 8820 17466 8832
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 17460 8792 17785 8820
rect 17460 8780 17466 8792
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 18138 8820 18144 8832
rect 18099 8792 18144 8820
rect 17773 8783 17831 8789
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 20162 8780 20168 8832
rect 20220 8820 20226 8832
rect 20732 8820 20760 8919
rect 20990 8897 20996 8900
rect 20984 8888 20996 8897
rect 20951 8860 20996 8888
rect 20984 8851 20996 8860
rect 20990 8848 20996 8851
rect 21048 8848 21054 8900
rect 21376 8888 21404 8928
rect 21726 8916 21732 8968
rect 21784 8956 21790 8968
rect 22466 8959 22524 8965
rect 22466 8956 22478 8959
rect 21784 8928 22478 8956
rect 21784 8916 21790 8928
rect 22466 8925 22478 8928
rect 22512 8925 22524 8959
rect 22922 8956 22928 8968
rect 22883 8928 22928 8956
rect 22466 8919 22524 8925
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 23198 8956 23204 8968
rect 23159 8928 23204 8956
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 23750 8916 23756 8968
rect 23808 8956 23814 8968
rect 23845 8959 23903 8965
rect 23845 8956 23857 8959
rect 23808 8928 23857 8956
rect 23808 8916 23814 8928
rect 23845 8925 23857 8928
rect 23891 8925 23903 8959
rect 23845 8919 23903 8925
rect 24639 8959 24697 8965
rect 24639 8925 24651 8959
rect 24685 8956 24697 8959
rect 24685 8928 24808 8956
rect 24685 8925 24697 8928
rect 24639 8919 24697 8925
rect 22738 8888 22744 8900
rect 21376 8860 22744 8888
rect 22738 8848 22744 8860
rect 22796 8848 22802 8900
rect 23937 8891 23995 8897
rect 23937 8857 23949 8891
rect 23983 8888 23995 8891
rect 24397 8891 24455 8897
rect 24397 8888 24409 8891
rect 23983 8860 24409 8888
rect 23983 8857 23995 8860
rect 23937 8851 23995 8857
rect 24397 8857 24409 8860
rect 24443 8857 24455 8891
rect 24780 8888 24808 8928
rect 24854 8916 24860 8968
rect 24912 8956 24918 8968
rect 25041 8959 25099 8965
rect 25041 8956 25053 8959
rect 24912 8928 25053 8956
rect 24912 8916 24918 8928
rect 25041 8925 25053 8928
rect 25087 8956 25099 8959
rect 25133 8959 25191 8965
rect 25133 8956 25145 8959
rect 25087 8928 25145 8956
rect 25087 8925 25099 8928
rect 25041 8919 25099 8925
rect 25133 8925 25145 8928
rect 25179 8925 25191 8959
rect 25133 8919 25191 8925
rect 25222 8916 25228 8968
rect 25280 8956 25286 8968
rect 25332 8965 25360 8996
rect 25317 8959 25375 8965
rect 25317 8956 25329 8959
rect 25280 8928 25329 8956
rect 25280 8916 25286 8928
rect 25317 8925 25329 8928
rect 25363 8925 25375 8959
rect 25317 8919 25375 8925
rect 25501 8891 25559 8897
rect 25501 8888 25513 8891
rect 24780 8860 25513 8888
rect 24397 8851 24455 8857
rect 25501 8857 25513 8860
rect 25547 8888 25559 8891
rect 25590 8888 25596 8900
rect 25547 8860 25596 8888
rect 25547 8857 25559 8860
rect 25501 8851 25559 8857
rect 25590 8848 25596 8860
rect 25648 8848 25654 8900
rect 20220 8792 20760 8820
rect 20220 8780 20226 8792
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 23532 8792 23577 8820
rect 23532 8780 23538 8792
rect 1104 8730 26128 8752
rect 1104 8678 9291 8730
rect 9343 8678 9355 8730
rect 9407 8678 9419 8730
rect 9471 8678 9483 8730
rect 9535 8678 9547 8730
rect 9599 8678 17632 8730
rect 17684 8678 17696 8730
rect 17748 8678 17760 8730
rect 17812 8678 17824 8730
rect 17876 8678 17888 8730
rect 17940 8678 26128 8730
rect 1104 8656 26128 8678
rect 2590 8616 2596 8628
rect 2551 8588 2596 8616
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 3878 8576 3884 8628
rect 3936 8576 3942 8628
rect 6086 8616 6092 8628
rect 5459 8588 6092 8616
rect 3896 8548 3924 8576
rect 2792 8520 3924 8548
rect 2792 8489 2820 8520
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8449 2835 8483
rect 3050 8480 3056 8492
rect 3011 8452 3056 8480
rect 2777 8443 2835 8449
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 3160 8489 3188 8520
rect 5459 8492 5487 8588
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 7098 8616 7104 8628
rect 7059 8588 7104 8616
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 8018 8616 8024 8628
rect 7979 8588 8024 8616
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8570 8576 8576 8628
rect 8628 8576 8634 8628
rect 9030 8616 9036 8628
rect 8991 8588 9036 8616
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 11146 8616 11152 8628
rect 11107 8588 11152 8616
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11606 8616 11612 8628
rect 11567 8588 11612 8616
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 12342 8576 12348 8628
rect 12400 8616 12406 8628
rect 12805 8619 12863 8625
rect 12400 8576 12434 8616
rect 12805 8585 12817 8619
rect 12851 8585 12863 8619
rect 13354 8616 13360 8628
rect 13315 8588 13360 8616
rect 12805 8579 12863 8585
rect 6914 8548 6920 8560
rect 6840 8520 6920 8548
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 3234 8440 3240 8492
rect 3292 8480 3298 8492
rect 3881 8483 3939 8489
rect 3292 8452 3337 8480
rect 3292 8440 3298 8452
rect 3881 8449 3893 8483
rect 3927 8480 3939 8483
rect 4062 8480 4068 8492
rect 3927 8452 4068 8480
rect 3927 8449 3939 8452
rect 3881 8443 3939 8449
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 5261 8483 5319 8489
rect 5261 8480 5273 8483
rect 4212 8452 5273 8480
rect 4212 8440 4218 8452
rect 5261 8449 5273 8452
rect 5307 8480 5319 8483
rect 5350 8480 5356 8492
rect 5307 8452 5356 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 5444 8486 5502 8492
rect 5444 8452 5456 8486
rect 5490 8452 5502 8486
rect 5444 8446 5502 8452
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5902 8480 5908 8492
rect 5859 8452 5908 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5902 8440 5908 8452
rect 5960 8440 5966 8492
rect 6840 8489 6868 8520
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 7653 8551 7711 8557
rect 7653 8548 7665 8551
rect 7064 8520 7665 8548
rect 7064 8508 7070 8520
rect 7653 8517 7665 8520
rect 7699 8548 7711 8551
rect 7926 8548 7932 8560
rect 7699 8520 7932 8548
rect 7699 8517 7711 8520
rect 7653 8511 7711 8517
rect 7926 8508 7932 8520
rect 7984 8508 7990 8560
rect 8588 8548 8616 8576
rect 8128 8520 8616 8548
rect 8128 8489 8156 8520
rect 10962 8508 10968 8560
rect 11020 8548 11026 8560
rect 11020 8520 11100 8548
rect 11020 8508 11026 8520
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 6825 8443 6883 8449
rect 6932 8452 7297 8480
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 2961 8347 3019 8353
rect 2961 8313 2973 8347
rect 3007 8344 3019 8347
rect 3234 8344 3240 8356
rect 3007 8316 3240 8344
rect 3007 8313 3019 8316
rect 2961 8307 3019 8313
rect 3234 8304 3240 8316
rect 3292 8344 3298 8356
rect 3697 8347 3755 8353
rect 3697 8344 3709 8347
rect 3292 8316 3709 8344
rect 3292 8304 3298 8316
rect 3697 8313 3709 8316
rect 3743 8313 3755 8347
rect 3697 8307 3755 8313
rect 5552 8344 5580 8375
rect 5626 8372 5632 8424
rect 5684 8412 5690 8424
rect 6362 8412 6368 8424
rect 5684 8384 5729 8412
rect 5828 8384 6368 8412
rect 5684 8372 5690 8384
rect 5828 8344 5856 8384
rect 6362 8372 6368 8384
rect 6420 8412 6426 8424
rect 6730 8412 6736 8424
rect 6420 8384 6736 8412
rect 6420 8372 6426 8384
rect 6730 8372 6736 8384
rect 6788 8372 6794 8424
rect 5994 8344 6000 8356
rect 5552 8316 5856 8344
rect 5955 8316 6000 8344
rect 3142 8276 3148 8288
rect 3103 8248 3148 8276
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 3326 8236 3332 8288
rect 3384 8276 3390 8288
rect 3513 8279 3571 8285
rect 3513 8276 3525 8279
rect 3384 8248 3525 8276
rect 3384 8236 3390 8248
rect 3513 8245 3525 8248
rect 3559 8245 3571 8279
rect 3513 8239 3571 8245
rect 4338 8236 4344 8288
rect 4396 8276 4402 8288
rect 5552 8276 5580 8316
rect 5994 8304 6000 8316
rect 6052 8304 6058 8356
rect 6638 8304 6644 8356
rect 6696 8344 6702 8356
rect 6932 8353 6960 8452
rect 7285 8449 7297 8452
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 8662 8480 8668 8492
rect 8536 8452 8581 8480
rect 8623 8452 8668 8480
rect 8536 8440 8542 8452
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8938 8480 8944 8492
rect 8899 8452 8944 8480
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 11072 8489 11100 8520
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 11940 8520 11985 8548
rect 11940 8508 11946 8520
rect 12406 8489 12434 8576
rect 12820 8548 12848 8579
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 13998 8616 14004 8628
rect 13959 8588 14004 8616
rect 13998 8576 14004 8588
rect 14056 8616 14062 8628
rect 14093 8619 14151 8625
rect 14093 8616 14105 8619
rect 14056 8588 14105 8616
rect 14056 8576 14062 8588
rect 14093 8585 14105 8588
rect 14139 8585 14151 8619
rect 15010 8616 15016 8628
rect 14971 8588 15016 8616
rect 14093 8579 14151 8585
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15838 8616 15844 8628
rect 15799 8588 15844 8616
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 16025 8619 16083 8625
rect 16025 8585 16037 8619
rect 16071 8585 16083 8619
rect 16025 8579 16083 8585
rect 17037 8619 17095 8625
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 17126 8616 17132 8628
rect 17083 8588 17132 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 12544 8520 12848 8548
rect 13265 8551 13323 8557
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 11057 8483 11115 8489
rect 10827 8452 11008 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 8202 8412 8208 8424
rect 7484 8384 8208 8412
rect 7484 8353 7512 8384
rect 8202 8372 8208 8384
rect 8260 8412 8266 8424
rect 8297 8415 8355 8421
rect 8297 8412 8309 8415
rect 8260 8384 8309 8412
rect 8260 8372 8266 8384
rect 8297 8381 8309 8384
rect 8343 8381 8355 8415
rect 8297 8375 8355 8381
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 10226 8412 10232 8424
rect 8444 8384 8800 8412
rect 10139 8384 10232 8412
rect 8444 8372 8450 8384
rect 8772 8353 8800 8384
rect 10226 8372 10232 8384
rect 10284 8412 10290 8424
rect 10870 8412 10876 8424
rect 10284 8384 10732 8412
rect 10831 8384 10876 8412
rect 10284 8372 10290 8384
rect 6917 8347 6975 8353
rect 6917 8344 6929 8347
rect 6696 8316 6929 8344
rect 6696 8304 6702 8316
rect 6917 8313 6929 8316
rect 6963 8313 6975 8347
rect 6917 8307 6975 8313
rect 7469 8347 7527 8353
rect 7469 8313 7481 8347
rect 7515 8313 7527 8347
rect 7469 8307 7527 8313
rect 8757 8347 8815 8353
rect 8757 8313 8769 8347
rect 8803 8344 8815 8347
rect 9214 8344 9220 8356
rect 8803 8316 9220 8344
rect 8803 8313 8815 8316
rect 8757 8307 8815 8313
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 10505 8347 10563 8353
rect 10505 8313 10517 8347
rect 10551 8344 10563 8347
rect 10594 8344 10600 8356
rect 10551 8316 10600 8344
rect 10551 8313 10563 8316
rect 10505 8307 10563 8313
rect 10594 8304 10600 8316
rect 10652 8304 10658 8356
rect 10704 8344 10732 8384
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 10980 8412 11008 8452
rect 11057 8449 11069 8483
rect 11103 8480 11115 8483
rect 11716 8480 11827 8486
rect 12299 8483 12357 8489
rect 12299 8480 12311 8483
rect 11103 8458 12311 8480
rect 11103 8452 11744 8458
rect 11799 8452 12311 8458
rect 11103 8449 11115 8452
rect 11057 8443 11115 8449
rect 12299 8449 12311 8452
rect 12345 8449 12357 8483
rect 12406 8483 12483 8489
rect 12406 8452 12437 8483
rect 12299 8443 12357 8449
rect 12425 8449 12437 8452
rect 12471 8449 12483 8483
rect 12425 8443 12483 8449
rect 11606 8412 11612 8424
rect 10980 8384 11612 8412
rect 11606 8372 11612 8384
rect 11664 8372 11670 8424
rect 11790 8372 11796 8424
rect 11848 8412 11854 8424
rect 12069 8415 12127 8421
rect 11848 8384 11941 8412
rect 11848 8372 11854 8384
rect 12069 8381 12081 8415
rect 12115 8412 12127 8415
rect 12544 8412 12572 8520
rect 13265 8517 13277 8551
rect 13311 8548 13323 8551
rect 13906 8548 13912 8560
rect 13311 8520 13912 8548
rect 13311 8517 13323 8520
rect 13265 8511 13323 8517
rect 13906 8508 13912 8520
rect 13964 8508 13970 8560
rect 14826 8508 14832 8560
rect 14884 8548 14890 8560
rect 14921 8551 14979 8557
rect 14921 8548 14933 8551
rect 14884 8520 14933 8548
rect 14884 8508 14890 8520
rect 14921 8517 14933 8520
rect 14967 8517 14979 8551
rect 14921 8511 14979 8517
rect 12621 8483 12679 8489
rect 12621 8449 12633 8483
rect 12667 8478 12679 8483
rect 12710 8478 12716 8492
rect 12667 8450 12716 8478
rect 12667 8449 12679 8450
rect 12621 8443 12679 8449
rect 12710 8440 12716 8450
rect 12768 8440 12774 8492
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8480 15715 8483
rect 16040 8480 16068 8579
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8585 17923 8619
rect 17865 8579 17923 8585
rect 17880 8548 17908 8579
rect 18046 8576 18052 8628
rect 18104 8616 18110 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 18104 8588 19441 8616
rect 18104 8576 18110 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 21542 8616 21548 8628
rect 21503 8588 21548 8616
rect 19429 8579 19487 8585
rect 21542 8576 21548 8588
rect 21600 8576 21606 8628
rect 25222 8616 25228 8628
rect 25183 8588 25228 8616
rect 25222 8576 25228 8588
rect 25280 8576 25286 8628
rect 19334 8548 19340 8560
rect 17880 8520 19340 8548
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 19794 8508 19800 8560
rect 19852 8548 19858 8560
rect 20432 8551 20490 8557
rect 19852 8520 20392 8548
rect 19852 8508 19858 8520
rect 15703 8452 16068 8480
rect 15703 8449 15715 8452
rect 15657 8443 15715 8449
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 17681 8483 17739 8489
rect 16356 8452 17264 8480
rect 16356 8440 16362 8452
rect 13173 8415 13231 8421
rect 13173 8412 13185 8415
rect 12115 8384 12572 8412
rect 12605 8384 13185 8412
rect 12115 8381 12127 8384
rect 12069 8375 12127 8381
rect 10778 8344 10784 8356
rect 10704 8316 10784 8344
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 4396 8248 5580 8276
rect 4396 8236 4402 8248
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 11808 8276 11836 8372
rect 12161 8347 12219 8353
rect 12161 8313 12173 8347
rect 12207 8344 12219 8347
rect 12605 8344 12633 8384
rect 13173 8381 13185 8384
rect 13219 8412 13231 8415
rect 13262 8412 13268 8424
rect 13219 8384 13268 8412
rect 13219 8381 13231 8384
rect 13173 8375 13231 8381
rect 13262 8372 13268 8384
rect 13320 8412 13326 8424
rect 13998 8412 14004 8424
rect 13320 8384 14004 8412
rect 13320 8372 13326 8384
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 16482 8412 16488 8424
rect 16443 8384 16488 8412
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 17126 8412 17132 8424
rect 17087 8384 17132 8412
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17236 8421 17264 8452
rect 17681 8449 17693 8483
rect 17727 8480 17739 8483
rect 17954 8480 17960 8492
rect 17727 8452 17960 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18598 8440 18604 8492
rect 18656 8480 18662 8492
rect 18978 8483 19036 8489
rect 18978 8480 18990 8483
rect 18656 8452 18990 8480
rect 18656 8440 18662 8452
rect 18978 8449 18990 8452
rect 19024 8449 19036 8483
rect 18978 8443 19036 8449
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 20162 8480 20168 8492
rect 19576 8452 19621 8480
rect 20123 8452 20168 8480
rect 19576 8440 19582 8452
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 20364 8480 20392 8520
rect 20432 8517 20444 8551
rect 20478 8548 20490 8551
rect 20530 8548 20536 8560
rect 20478 8520 20536 8548
rect 20478 8517 20490 8520
rect 20432 8511 20490 8517
rect 20530 8508 20536 8520
rect 20588 8508 20594 8560
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 21821 8551 21879 8557
rect 21821 8548 21833 8551
rect 21784 8520 21833 8548
rect 21784 8508 21790 8520
rect 21821 8517 21833 8520
rect 21867 8517 21879 8551
rect 22002 8548 22008 8560
rect 21963 8520 22008 8548
rect 21821 8511 21879 8517
rect 22002 8508 22008 8520
rect 22060 8508 22066 8560
rect 22189 8551 22247 8557
rect 22189 8517 22201 8551
rect 22235 8548 22247 8551
rect 22922 8548 22928 8560
rect 22235 8520 22928 8548
rect 22235 8517 22247 8520
rect 22189 8511 22247 8517
rect 22922 8508 22928 8520
rect 22980 8508 22986 8560
rect 20364 8452 22094 8480
rect 17221 8415 17279 8421
rect 17221 8381 17233 8415
rect 17267 8412 17279 8415
rect 17862 8412 17868 8424
rect 17267 8384 17868 8412
rect 17267 8381 17279 8384
rect 17221 8375 17279 8381
rect 12207 8316 12633 8344
rect 12207 8313 12219 8316
rect 12161 8307 12219 8313
rect 13354 8304 13360 8356
rect 13412 8344 13418 8356
rect 17512 8353 17540 8384
rect 17862 8372 17868 8384
rect 17920 8372 17926 8424
rect 19245 8415 19303 8421
rect 19245 8381 19257 8415
rect 19291 8412 19303 8415
rect 19886 8412 19892 8424
rect 19291 8384 19748 8412
rect 19847 8384 19892 8412
rect 19291 8381 19303 8384
rect 19245 8375 19303 8381
rect 13725 8347 13783 8353
rect 13725 8344 13737 8347
rect 13412 8316 13737 8344
rect 13412 8304 13418 8316
rect 13725 8313 13737 8316
rect 13771 8313 13783 8347
rect 13725 8307 13783 8313
rect 16209 8347 16267 8353
rect 16209 8313 16221 8347
rect 16255 8344 16267 8347
rect 16669 8347 16727 8353
rect 16669 8344 16681 8347
rect 16255 8316 16681 8344
rect 16255 8313 16267 8316
rect 16209 8307 16267 8313
rect 16669 8313 16681 8316
rect 16715 8313 16727 8347
rect 16669 8307 16727 8313
rect 17497 8347 17555 8353
rect 17497 8313 17509 8347
rect 17543 8313 17555 8347
rect 19720 8344 19748 8384
rect 19886 8372 19892 8384
rect 19944 8372 19950 8424
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 20036 8384 20081 8412
rect 20036 8372 20042 8384
rect 20162 8344 20168 8356
rect 19720 8316 20168 8344
rect 17497 8307 17555 8313
rect 20162 8304 20168 8316
rect 20220 8304 20226 8356
rect 22066 8344 22094 8452
rect 22738 8440 22744 8492
rect 22796 8480 22802 8492
rect 23658 8480 23664 8492
rect 22796 8452 23664 8480
rect 22796 8440 22802 8452
rect 23658 8440 23664 8452
rect 23716 8480 23722 8492
rect 23845 8483 23903 8489
rect 23845 8480 23857 8483
rect 23716 8452 23857 8480
rect 23716 8440 23722 8452
rect 23845 8449 23857 8452
rect 23891 8449 23903 8483
rect 23845 8443 23903 8449
rect 23934 8440 23940 8492
rect 23992 8480 23998 8492
rect 24101 8483 24159 8489
rect 24101 8480 24113 8483
rect 23992 8452 24113 8480
rect 23992 8440 23998 8452
rect 24101 8449 24113 8452
rect 24147 8449 24159 8483
rect 24101 8443 24159 8449
rect 22646 8372 22652 8424
rect 22704 8412 22710 8424
rect 23017 8415 23075 8421
rect 23017 8412 23029 8415
rect 22704 8384 23029 8412
rect 22704 8372 22710 8384
rect 23017 8381 23029 8384
rect 23063 8381 23075 8415
rect 23474 8412 23480 8424
rect 23017 8375 23075 8381
rect 23400 8384 23480 8412
rect 22664 8344 22692 8372
rect 23400 8353 23428 8384
rect 23474 8372 23480 8384
rect 23532 8372 23538 8424
rect 22066 8316 22692 8344
rect 23385 8347 23443 8353
rect 23385 8313 23397 8347
rect 23431 8313 23443 8347
rect 23385 8307 23443 8313
rect 12526 8276 12532 8288
rect 11020 8248 11836 8276
rect 12487 8248 12532 8276
rect 11020 8236 11026 8248
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 23477 8279 23535 8285
rect 23477 8245 23489 8279
rect 23523 8276 23535 8279
rect 23658 8276 23664 8288
rect 23523 8248 23664 8276
rect 23523 8245 23535 8248
rect 23477 8239 23535 8245
rect 23658 8236 23664 8248
rect 23716 8236 23722 8288
rect 1104 8186 26128 8208
rect 1104 8134 5120 8186
rect 5172 8134 5184 8186
rect 5236 8134 5248 8186
rect 5300 8134 5312 8186
rect 5364 8134 5376 8186
rect 5428 8134 13462 8186
rect 13514 8134 13526 8186
rect 13578 8134 13590 8186
rect 13642 8134 13654 8186
rect 13706 8134 13718 8186
rect 13770 8134 21803 8186
rect 21855 8134 21867 8186
rect 21919 8134 21931 8186
rect 21983 8134 21995 8186
rect 22047 8134 22059 8186
rect 22111 8134 26128 8186
rect 1104 8112 26128 8134
rect 2961 8075 3019 8081
rect 2961 8041 2973 8075
rect 3007 8072 3019 8075
rect 3050 8072 3056 8084
rect 3007 8044 3056 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 5626 8072 5632 8084
rect 4448 8044 5632 8072
rect 3786 7896 3792 7948
rect 3844 7936 3850 7948
rect 4338 7936 4344 7948
rect 3844 7908 4200 7936
rect 4299 7908 4344 7936
rect 3844 7896 3850 7908
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 1627 7840 2774 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 1848 7803 1906 7809
rect 1848 7769 1860 7803
rect 1894 7800 1906 7803
rect 2130 7800 2136 7812
rect 1894 7772 2136 7800
rect 1894 7769 1906 7772
rect 1848 7763 1906 7769
rect 2130 7760 2136 7772
rect 2188 7760 2194 7812
rect 2746 7800 2774 7840
rect 3050 7828 3056 7880
rect 3108 7868 3114 7880
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 3108 7840 3341 7868
rect 3108 7828 3114 7840
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 3329 7831 3387 7837
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 4172 7868 4200 7908
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 4448 7945 4476 8044
rect 5626 8032 5632 8044
rect 5684 8072 5690 8084
rect 6454 8072 6460 8084
rect 5684 8044 6460 8072
rect 5684 8032 5690 8044
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 6730 8072 6736 8084
rect 6691 8044 6736 8072
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7006 8032 7012 8084
rect 7064 8072 7070 8084
rect 7834 8072 7840 8084
rect 7064 8044 7840 8072
rect 7064 8032 7070 8044
rect 7834 8032 7840 8044
rect 7892 8072 7898 8084
rect 8110 8072 8116 8084
rect 7892 8044 8116 8072
rect 7892 8032 7898 8044
rect 8110 8032 8116 8044
rect 8168 8072 8174 8084
rect 8757 8075 8815 8081
rect 8757 8072 8769 8075
rect 8168 8044 8769 8072
rect 8168 8032 8174 8044
rect 8757 8041 8769 8044
rect 8803 8041 8815 8075
rect 8757 8035 8815 8041
rect 9030 8032 9036 8084
rect 9088 8072 9094 8084
rect 9858 8072 9864 8084
rect 9088 8044 9864 8072
rect 9088 8032 9094 8044
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 10962 8032 10968 8084
rect 11020 8072 11026 8084
rect 16301 8075 16359 8081
rect 11020 8044 15700 8072
rect 11020 8032 11026 8044
rect 8294 8004 8300 8016
rect 7300 7976 8300 8004
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7905 4491 7939
rect 4433 7899 4491 7905
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7300 7945 7328 7976
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 9122 7964 9128 8016
rect 9180 8004 9186 8016
rect 11698 8004 11704 8016
rect 9180 7976 9444 8004
rect 11611 7976 11704 8004
rect 9180 7964 9186 7976
rect 7285 7939 7343 7945
rect 7156 7908 7236 7936
rect 7156 7896 7162 7908
rect 4230 7871 4288 7877
rect 4230 7868 4242 7871
rect 4172 7840 4242 7868
rect 4230 7837 4242 7840
rect 4276 7837 4288 7871
rect 4230 7831 4288 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4798 7868 4804 7880
rect 4663 7840 4804 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 4908 7840 6377 7868
rect 4338 7800 4344 7812
rect 2746 7772 4344 7800
rect 4338 7760 4344 7772
rect 4396 7800 4402 7812
rect 4908 7800 4936 7840
rect 6365 7837 6377 7840
rect 6411 7837 6423 7871
rect 6638 7868 6644 7880
rect 6599 7840 6644 7868
rect 6365 7831 6423 7837
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 6914 7868 6920 7880
rect 6875 7840 6920 7868
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 7208 7877 7236 7908
rect 7285 7905 7297 7939
rect 7331 7905 7343 7939
rect 7285 7899 7343 7905
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7936 7435 7939
rect 8202 7936 8208 7948
rect 7423 7908 8208 7936
rect 7423 7905 7435 7908
rect 7377 7899 7435 7905
rect 8202 7896 8208 7908
rect 8260 7936 8266 7948
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 8260 7908 9321 7936
rect 8260 7896 8266 7908
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 7192 7871 7250 7877
rect 7064 7840 7109 7868
rect 7064 7828 7070 7840
rect 7192 7837 7204 7871
rect 7238 7837 7250 7871
rect 7192 7831 7250 7837
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7868 7619 7871
rect 7834 7868 7840 7880
rect 7607 7840 7696 7868
rect 7795 7840 7840 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 4396 7772 4936 7800
rect 4396 7760 4402 7772
rect 5994 7760 6000 7812
rect 6052 7800 6058 7812
rect 6098 7803 6156 7809
rect 6098 7800 6110 7803
rect 6052 7772 6110 7800
rect 6052 7760 6058 7772
rect 6098 7769 6110 7772
rect 6144 7769 6156 7803
rect 6098 7763 6156 7769
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 3418 7732 3424 7744
rect 3283 7704 3424 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 3786 7692 3792 7744
rect 3844 7732 3850 7744
rect 3881 7735 3939 7741
rect 3881 7732 3893 7735
rect 3844 7704 3893 7732
rect 3844 7692 3850 7704
rect 3881 7701 3893 7704
rect 3927 7701 3939 7735
rect 4706 7732 4712 7744
rect 4667 7704 4712 7732
rect 3881 7695 3939 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 4985 7735 5043 7741
rect 4985 7701 4997 7735
rect 5031 7732 5043 7735
rect 5902 7732 5908 7744
rect 5031 7704 5908 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 7668 7732 7696 7840
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 8020 7871 8078 7877
rect 8020 7868 8032 7871
rect 7984 7840 8032 7868
rect 7984 7828 7990 7840
rect 8020 7837 8032 7840
rect 8066 7837 8078 7871
rect 8020 7831 8078 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7868 8171 7871
rect 8294 7868 8300 7880
rect 8159 7840 8300 7868
rect 8159 7837 8171 7840
rect 8113 7831 8171 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 8757 7871 8815 7877
rect 8444 7840 8489 7868
rect 8444 7828 8450 7840
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8803 7840 8953 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9124 7871 9182 7877
rect 9124 7868 9136 7871
rect 9088 7840 9136 7868
rect 9088 7828 9094 7840
rect 9124 7837 9136 7840
rect 9170 7837 9182 7871
rect 9124 7831 9182 7837
rect 9214 7828 9220 7880
rect 9272 7868 9278 7880
rect 9416 7868 9444 7976
rect 11698 7964 11704 7976
rect 11756 8004 11762 8016
rect 11756 7976 11928 8004
rect 11756 7964 11762 7976
rect 11900 7945 11928 7976
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7905 11943 7939
rect 11885 7899 11943 7905
rect 12158 7896 12164 7948
rect 12216 7936 12222 7948
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 12216 7908 12357 7936
rect 12216 7896 12222 7908
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 13262 7896 13268 7948
rect 13320 7936 13326 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 13320 7908 13369 7936
rect 13320 7896 13326 7908
rect 13357 7905 13369 7908
rect 13403 7936 13415 7939
rect 13446 7936 13452 7948
rect 13403 7908 13452 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9272 7840 9317 7868
rect 9416 7840 9505 7868
rect 9272 7828 9278 7840
rect 9493 7837 9505 7840
rect 9539 7837 9551 7871
rect 10318 7868 10324 7880
rect 10279 7840 10324 7868
rect 9493 7831 9551 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10594 7877 10600 7880
rect 10588 7868 10600 7877
rect 10555 7840 10600 7868
rect 10588 7831 10600 7840
rect 10594 7828 10600 7831
rect 10652 7828 10658 7880
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11112 7840 12081 7868
rect 11112 7828 11118 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 7745 7803 7803 7809
rect 7745 7769 7757 7803
rect 7791 7800 7803 7803
rect 10134 7800 10140 7812
rect 7791 7772 10140 7800
rect 7791 7769 7803 7772
rect 7745 7763 7803 7769
rect 10134 7760 10140 7772
rect 10192 7760 10198 7812
rect 12084 7800 12112 7831
rect 12250 7828 12256 7880
rect 12308 7868 12314 7880
rect 13556 7877 13584 8044
rect 14185 8007 14243 8013
rect 14185 7973 14197 8007
rect 14231 7973 14243 8007
rect 14185 7967 14243 7973
rect 13814 7896 13820 7948
rect 13872 7936 13878 7948
rect 13909 7939 13967 7945
rect 13909 7936 13921 7939
rect 13872 7908 13921 7936
rect 13872 7896 13878 7908
rect 13909 7905 13921 7908
rect 13955 7936 13967 7939
rect 14200 7936 14228 7967
rect 13955 7908 14228 7936
rect 13955 7905 13967 7908
rect 13909 7899 13967 7905
rect 12437 7871 12495 7877
rect 12437 7868 12449 7871
rect 12308 7840 12449 7868
rect 12308 7828 12314 7840
rect 12437 7837 12449 7840
rect 12483 7868 12495 7871
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12483 7840 12909 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 15068 7840 15577 7868
rect 15068 7828 15074 7840
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 15672 7868 15700 8044
rect 16301 8041 16313 8075
rect 16347 8072 16359 8075
rect 17126 8072 17132 8084
rect 16347 8044 17132 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 17310 8072 17316 8084
rect 17271 8044 17316 8072
rect 17310 8032 17316 8044
rect 17368 8032 17374 8084
rect 19334 8032 19340 8084
rect 19392 8072 19398 8084
rect 19521 8075 19579 8081
rect 19521 8072 19533 8075
rect 19392 8044 19533 8072
rect 19392 8032 19398 8044
rect 19521 8041 19533 8044
rect 19567 8041 19579 8075
rect 19521 8035 19579 8041
rect 19889 8075 19947 8081
rect 19889 8041 19901 8075
rect 19935 8072 19947 8075
rect 19978 8072 19984 8084
rect 19935 8044 19984 8072
rect 19935 8041 19947 8044
rect 19889 8035 19947 8041
rect 17218 8004 17224 8016
rect 17179 7976 17224 8004
rect 17218 7964 17224 7976
rect 17276 7964 17282 8016
rect 18877 8007 18935 8013
rect 18877 7973 18889 8007
rect 18923 7973 18935 8007
rect 19536 8004 19564 8035
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20990 8032 20996 8084
rect 21048 8072 21054 8084
rect 21085 8075 21143 8081
rect 21085 8072 21097 8075
rect 21048 8044 21097 8072
rect 21048 8032 21054 8044
rect 21085 8041 21097 8044
rect 21131 8041 21143 8075
rect 21085 8035 21143 8041
rect 23845 8075 23903 8081
rect 23845 8041 23857 8075
rect 23891 8072 23903 8075
rect 23934 8072 23940 8084
rect 23891 8044 23940 8072
rect 23891 8041 23903 8044
rect 23845 8035 23903 8041
rect 23934 8032 23940 8044
rect 23992 8032 23998 8084
rect 20806 8004 20812 8016
rect 19536 7976 20024 8004
rect 20767 7976 20812 8004
rect 18877 7967 18935 7973
rect 16390 7896 16396 7948
rect 16448 7936 16454 7948
rect 17497 7939 17555 7945
rect 17497 7936 17509 7939
rect 16448 7908 17509 7936
rect 16448 7896 16454 7908
rect 17497 7905 17509 7908
rect 17543 7905 17555 7939
rect 18892 7936 18920 7967
rect 19613 7939 19671 7945
rect 19613 7936 19625 7939
rect 18892 7908 19625 7936
rect 17497 7899 17555 7905
rect 19613 7905 19625 7908
rect 19659 7936 19671 7939
rect 19886 7936 19892 7948
rect 19659 7908 19892 7936
rect 19659 7905 19671 7908
rect 19613 7899 19671 7905
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 16485 7871 16543 7877
rect 16485 7868 16497 7871
rect 15672 7840 16497 7868
rect 15565 7831 15623 7837
rect 16485 7837 16497 7840
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 16669 7871 16727 7877
rect 16669 7837 16681 7871
rect 16715 7868 16727 7871
rect 17402 7868 17408 7880
rect 16715 7840 17408 7868
rect 16715 7837 16727 7840
rect 16669 7831 16727 7837
rect 17402 7828 17408 7840
rect 17460 7828 17466 7880
rect 19996 7877 20024 7976
rect 20806 7964 20812 7976
rect 20864 7964 20870 8016
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 19981 7871 20039 7877
rect 19981 7837 19993 7871
rect 20027 7837 20039 7871
rect 19981 7831 20039 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7868 20223 7871
rect 20254 7868 20260 7880
rect 20211 7840 20260 7868
rect 20211 7837 20223 7840
rect 20165 7831 20223 7837
rect 12342 7800 12348 7812
rect 12084 7772 12348 7800
rect 12342 7760 12348 7772
rect 12400 7760 12406 7812
rect 12529 7803 12587 7809
rect 12529 7769 12541 7803
rect 12575 7800 12587 7803
rect 13081 7803 13139 7809
rect 12575 7772 13032 7800
rect 12575 7769 12587 7772
rect 12529 7763 12587 7769
rect 8294 7732 8300 7744
rect 7668 7704 8300 7732
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8478 7732 8484 7744
rect 8439 7704 8484 7732
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 9585 7735 9643 7741
rect 9585 7732 9597 7735
rect 9272 7704 9597 7732
rect 9272 7692 9278 7704
rect 9585 7701 9597 7704
rect 9631 7701 9643 7735
rect 9585 7695 9643 7701
rect 12618 7692 12624 7744
rect 12676 7732 12682 7744
rect 12713 7735 12771 7741
rect 12713 7732 12725 7735
rect 12676 7704 12725 7732
rect 12676 7692 12682 7704
rect 12713 7701 12725 7704
rect 12759 7701 12771 7735
rect 12713 7695 12771 7701
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 13004 7732 13032 7772
rect 13081 7769 13093 7803
rect 13127 7800 13139 7803
rect 13262 7800 13268 7812
rect 13127 7772 13268 7800
rect 13127 7769 13139 7772
rect 13081 7763 13139 7769
rect 13262 7760 13268 7772
rect 13320 7760 13326 7812
rect 13998 7760 14004 7812
rect 14056 7800 14062 7812
rect 15298 7803 15356 7809
rect 15298 7800 15310 7803
rect 14056 7772 15310 7800
rect 14056 7760 14062 7772
rect 15298 7769 15310 7772
rect 15344 7769 15356 7803
rect 15298 7763 15356 7769
rect 16761 7803 16819 7809
rect 16761 7769 16773 7803
rect 16807 7769 16819 7803
rect 16761 7763 16819 7769
rect 16853 7803 16911 7809
rect 16853 7769 16865 7803
rect 16899 7800 16911 7803
rect 17034 7800 17040 7812
rect 16899 7772 17040 7800
rect 16899 7769 16911 7772
rect 16853 7763 16911 7769
rect 13170 7732 13176 7744
rect 12860 7704 12905 7732
rect 13004 7704 13176 7732
rect 12860 7692 12866 7704
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 13817 7735 13875 7741
rect 13817 7701 13829 7735
rect 13863 7732 13875 7735
rect 13906 7732 13912 7744
rect 13863 7704 13912 7732
rect 13863 7701 13875 7704
rect 13817 7695 13875 7701
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 16776 7732 16804 7763
rect 17034 7760 17040 7772
rect 17092 7760 17098 7812
rect 17494 7760 17500 7812
rect 17552 7800 17558 7812
rect 17742 7803 17800 7809
rect 17742 7800 17754 7803
rect 17552 7772 17754 7800
rect 17552 7760 17558 7772
rect 17742 7769 17754 7772
rect 17788 7769 17800 7803
rect 19720 7800 19748 7831
rect 20180 7800 20208 7831
rect 20254 7828 20260 7840
rect 20312 7828 20318 7880
rect 21269 7871 21327 7877
rect 21269 7868 21281 7871
rect 20916 7840 21281 7868
rect 19720 7772 20208 7800
rect 20441 7803 20499 7809
rect 17742 7763 17800 7769
rect 20441 7769 20453 7803
rect 20487 7769 20499 7803
rect 20441 7763 20499 7769
rect 18322 7732 18328 7744
rect 16776 7704 18328 7732
rect 18322 7692 18328 7704
rect 18380 7732 18386 7744
rect 19337 7735 19395 7741
rect 19337 7732 19349 7735
rect 18380 7704 19349 7732
rect 18380 7692 18386 7704
rect 19337 7701 19349 7704
rect 19383 7732 19395 7735
rect 19518 7732 19524 7744
rect 19383 7704 19524 7732
rect 19383 7701 19395 7704
rect 19337 7695 19395 7701
rect 19518 7692 19524 7704
rect 19576 7692 19582 7744
rect 19794 7692 19800 7744
rect 19852 7732 19858 7744
rect 20456 7732 20484 7763
rect 20916 7741 20944 7840
rect 21269 7837 21281 7840
rect 21315 7837 21327 7871
rect 23290 7868 23296 7880
rect 23251 7840 23296 7868
rect 21269 7831 21327 7837
rect 23290 7828 23296 7840
rect 23348 7828 23354 7880
rect 23658 7868 23664 7880
rect 23619 7840 23664 7868
rect 23658 7828 23664 7840
rect 23716 7828 23722 7880
rect 19852 7704 20484 7732
rect 20901 7735 20959 7741
rect 19852 7692 19858 7704
rect 20901 7701 20913 7735
rect 20947 7701 20959 7735
rect 20901 7695 20959 7701
rect 23014 7692 23020 7744
rect 23072 7732 23078 7744
rect 23109 7735 23167 7741
rect 23109 7732 23121 7735
rect 23072 7704 23121 7732
rect 23072 7692 23078 7704
rect 23109 7701 23121 7704
rect 23155 7701 23167 7735
rect 23109 7695 23167 7701
rect 1104 7642 26128 7664
rect 1104 7590 9291 7642
rect 9343 7590 9355 7642
rect 9407 7590 9419 7642
rect 9471 7590 9483 7642
rect 9535 7590 9547 7642
rect 9599 7590 17632 7642
rect 17684 7590 17696 7642
rect 17748 7590 17760 7642
rect 17812 7590 17824 7642
rect 17876 7590 17888 7642
rect 17940 7590 26128 7642
rect 1104 7568 26128 7590
rect 2130 7528 2136 7540
rect 2091 7500 2136 7528
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 4856 7500 5733 7528
rect 4856 7488 4862 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 5721 7491 5779 7497
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 9030 7528 9036 7540
rect 8352 7500 9036 7528
rect 8352 7488 8358 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 11606 7528 11612 7540
rect 11567 7500 11612 7528
rect 11606 7488 11612 7500
rect 11664 7528 11670 7540
rect 12526 7528 12532 7540
rect 11664 7500 12532 7528
rect 11664 7488 11670 7500
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 13449 7531 13507 7537
rect 13449 7497 13461 7531
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 3418 7460 3424 7472
rect 2792 7432 3424 7460
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2240 7324 2268 7355
rect 2314 7352 2320 7404
rect 2372 7392 2378 7404
rect 2792 7401 2820 7432
rect 3418 7420 3424 7432
rect 3476 7420 3482 7472
rect 4608 7463 4666 7469
rect 4608 7429 4620 7463
rect 4654 7460 4666 7463
rect 4706 7460 4712 7472
rect 4654 7432 4712 7460
rect 4654 7429 4666 7432
rect 4608 7423 4666 7429
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 10962 7460 10968 7472
rect 6932 7432 10968 7460
rect 2777 7395 2835 7401
rect 2372 7364 2417 7392
rect 2372 7352 2378 7364
rect 2777 7361 2789 7395
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7361 2927 7395
rect 2869 7355 2927 7361
rect 2593 7327 2651 7333
rect 2593 7324 2605 7327
rect 2240 7296 2605 7324
rect 2593 7293 2605 7296
rect 2639 7293 2651 7327
rect 2884 7324 2912 7355
rect 3050 7352 3056 7404
rect 3108 7392 3114 7404
rect 3145 7395 3203 7401
rect 3145 7392 3157 7395
rect 3108 7364 3157 7392
rect 3108 7352 3114 7364
rect 3145 7361 3157 7364
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 3326 7392 3332 7404
rect 3283 7364 3332 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 4338 7392 4344 7404
rect 4299 7364 4344 7392
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 6932 7392 6960 7432
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 11241 7463 11299 7469
rect 11241 7429 11253 7463
rect 11287 7460 11299 7463
rect 12802 7460 12808 7472
rect 11287 7432 12808 7460
rect 11287 7429 11299 7432
rect 11241 7423 11299 7429
rect 12802 7420 12808 7432
rect 12860 7460 12866 7472
rect 12860 7432 12940 7460
rect 12860 7420 12866 7432
rect 4448 7364 6960 7392
rect 4448 7324 4476 7364
rect 7006 7352 7012 7404
rect 7064 7392 7070 7404
rect 7570 7395 7628 7401
rect 7570 7392 7582 7395
rect 7064 7364 7582 7392
rect 7064 7352 7070 7364
rect 7570 7361 7582 7364
rect 7616 7361 7628 7395
rect 7570 7355 7628 7361
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 9502 7395 9560 7401
rect 9502 7392 9514 7395
rect 9272 7364 9514 7392
rect 9272 7352 9278 7364
rect 9502 7361 9514 7364
rect 9548 7361 9560 7395
rect 9502 7355 9560 7361
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 11112 7364 11161 7392
rect 11112 7352 11118 7364
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11698 7392 11704 7404
rect 11659 7364 11704 7392
rect 11149 7355 11207 7361
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 12434 7392 12440 7404
rect 12395 7364 12440 7392
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 12912 7401 12940 7432
rect 12897 7395 12955 7401
rect 12897 7361 12909 7395
rect 12943 7361 12955 7395
rect 13262 7392 13268 7404
rect 13223 7364 13268 7392
rect 12897 7355 12955 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 13464 7392 13492 7491
rect 13538 7488 13544 7540
rect 13596 7528 13602 7540
rect 13998 7528 14004 7540
rect 13596 7500 13641 7528
rect 13959 7500 14004 7528
rect 13596 7488 13602 7500
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 17402 7488 17408 7540
rect 17460 7528 17466 7540
rect 18598 7528 18604 7540
rect 17460 7500 18184 7528
rect 18559 7500 18604 7528
rect 17460 7488 17466 7500
rect 13556 7460 13584 7488
rect 14185 7463 14243 7469
rect 14185 7460 14197 7463
rect 13556 7432 14197 7460
rect 14185 7429 14197 7432
rect 14231 7429 14243 7463
rect 14185 7423 14243 7429
rect 16758 7420 16764 7472
rect 16816 7460 16822 7472
rect 17129 7463 17187 7469
rect 17129 7460 17141 7463
rect 16816 7432 17141 7460
rect 16816 7420 16822 7432
rect 17129 7429 17141 7432
rect 17175 7460 17187 7463
rect 17865 7463 17923 7469
rect 17865 7460 17877 7463
rect 17175 7432 17877 7460
rect 17175 7429 17187 7432
rect 17129 7423 17187 7429
rect 17865 7429 17877 7432
rect 17911 7429 17923 7463
rect 17865 7423 17923 7429
rect 13725 7395 13783 7401
rect 13725 7392 13737 7395
rect 13464 7364 13737 7392
rect 13725 7361 13737 7364
rect 13771 7361 13783 7395
rect 13906 7392 13912 7404
rect 13867 7364 13912 7392
rect 13725 7355 13783 7361
rect 2884 7296 4476 7324
rect 7837 7327 7895 7333
rect 2593 7287 2651 7293
rect 7837 7293 7849 7327
rect 7883 7324 7895 7327
rect 7926 7324 7932 7336
rect 7883 7296 7932 7324
rect 7883 7293 7895 7296
rect 7837 7287 7895 7293
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7324 9827 7327
rect 10318 7324 10324 7336
rect 9815 7296 10324 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 10318 7284 10324 7296
rect 10376 7324 10382 7336
rect 10502 7324 10508 7336
rect 10376 7296 10508 7324
rect 10376 7284 10382 7296
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 12124 7296 12296 7324
rect 12124 7284 12130 7296
rect 3053 7259 3111 7265
rect 3053 7225 3065 7259
rect 3099 7256 3111 7259
rect 3234 7256 3240 7268
rect 3099 7228 3240 7256
rect 3099 7225 3111 7228
rect 3053 7219 3111 7225
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 3602 7256 3608 7268
rect 3563 7228 3608 7256
rect 3602 7216 3608 7228
rect 3660 7216 3666 7268
rect 566 7148 572 7200
rect 624 7188 630 7200
rect 1857 7191 1915 7197
rect 1857 7188 1869 7191
rect 624 7160 1869 7188
rect 624 7148 630 7160
rect 1857 7157 1869 7160
rect 1903 7188 1915 7191
rect 2314 7188 2320 7200
rect 1903 7160 2320 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 5626 7148 5632 7200
rect 5684 7188 5690 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 5684 7160 5917 7188
rect 5684 7148 5690 7160
rect 5905 7157 5917 7160
rect 5951 7157 5963 7191
rect 5905 7151 5963 7157
rect 6457 7191 6515 7197
rect 6457 7157 6469 7191
rect 6503 7188 6515 7191
rect 6730 7188 6736 7200
rect 6503 7160 6736 7188
rect 6503 7157 6515 7160
rect 6457 7151 6515 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8389 7191 8447 7197
rect 8389 7188 8401 7191
rect 8352 7160 8401 7188
rect 8352 7148 8358 7160
rect 8389 7157 8401 7160
rect 8435 7188 8447 7191
rect 9122 7188 9128 7200
rect 8435 7160 9128 7188
rect 8435 7157 8447 7160
rect 8389 7151 8447 7157
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 12069 7191 12127 7197
rect 12069 7157 12081 7191
rect 12115 7188 12127 7191
rect 12158 7188 12164 7200
rect 12115 7160 12164 7188
rect 12115 7157 12127 7160
rect 12069 7151 12127 7157
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12268 7188 12296 7296
rect 12526 7284 12532 7336
rect 12584 7324 12590 7336
rect 12667 7327 12725 7333
rect 12667 7324 12679 7327
rect 12584 7296 12679 7324
rect 12584 7284 12590 7296
rect 12667 7293 12679 7296
rect 12713 7324 12725 7327
rect 13740 7324 13768 7355
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7392 16727 7395
rect 16850 7392 16856 7404
rect 16715 7364 16856 7392
rect 16715 7361 16727 7364
rect 16669 7355 16727 7361
rect 16850 7352 16856 7364
rect 16908 7392 16914 7404
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16908 7364 16957 7392
rect 16908 7352 16914 7364
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 17954 7392 17960 7404
rect 17915 7364 17960 7392
rect 16945 7355 17003 7361
rect 17954 7352 17960 7364
rect 18012 7352 18018 7404
rect 18156 7401 18184 7500
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 19794 7488 19800 7540
rect 19852 7528 19858 7540
rect 19889 7531 19947 7537
rect 19889 7528 19901 7531
rect 19852 7500 19901 7528
rect 19852 7488 19858 7500
rect 19889 7497 19901 7500
rect 19935 7497 19947 7531
rect 22830 7528 22836 7540
rect 22791 7500 22836 7528
rect 19889 7491 19947 7497
rect 22830 7488 22836 7500
rect 22888 7488 22894 7540
rect 23661 7531 23719 7537
rect 23661 7497 23673 7531
rect 23707 7528 23719 7531
rect 23842 7528 23848 7540
rect 23707 7500 23848 7528
rect 23707 7497 23719 7500
rect 23661 7491 23719 7497
rect 23842 7488 23848 7500
rect 23900 7488 23906 7540
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7361 18199 7395
rect 18322 7392 18328 7404
rect 18283 7364 18328 7392
rect 18141 7355 18199 7361
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7361 18475 7395
rect 18417 7355 18475 7361
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 16482 7324 16488 7336
rect 12713 7296 13124 7324
rect 13740 7296 16488 7324
rect 12713 7293 12725 7296
rect 12667 7287 12725 7293
rect 13096 7265 13124 7296
rect 16482 7284 16488 7296
rect 16540 7324 16546 7336
rect 17034 7324 17040 7336
rect 16540 7296 17040 7324
rect 16540 7284 16546 7296
rect 17034 7284 17040 7296
rect 17092 7324 17098 7336
rect 17221 7327 17279 7333
rect 17221 7324 17233 7327
rect 17092 7296 17233 7324
rect 17092 7284 17098 7296
rect 17221 7293 17233 7296
rect 17267 7293 17279 7327
rect 18432 7324 18460 7355
rect 17221 7287 17279 7293
rect 17696 7296 18460 7324
rect 13081 7259 13139 7265
rect 13081 7225 13093 7259
rect 13127 7256 13139 7259
rect 13446 7256 13452 7268
rect 13127 7228 13452 7256
rect 13127 7225 13139 7228
rect 13081 7219 13139 7225
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 17696 7265 17724 7296
rect 17589 7259 17647 7265
rect 17589 7225 17601 7259
rect 17635 7225 17647 7259
rect 17589 7219 17647 7225
rect 17681 7259 17739 7265
rect 17681 7225 17693 7259
rect 17727 7225 17739 7259
rect 17681 7219 17739 7225
rect 17865 7259 17923 7265
rect 17865 7225 17877 7259
rect 17911 7256 17923 7259
rect 19352 7256 19380 7355
rect 19518 7352 19524 7404
rect 19576 7392 19582 7404
rect 19705 7395 19763 7401
rect 19705 7392 19717 7395
rect 19576 7364 19717 7392
rect 19576 7352 19582 7364
rect 19705 7361 19717 7364
rect 19751 7361 19763 7395
rect 20530 7392 20536 7404
rect 20491 7364 20536 7392
rect 19705 7355 19763 7361
rect 20530 7352 20536 7364
rect 20588 7352 20594 7404
rect 22925 7395 22983 7401
rect 22925 7361 22937 7395
rect 22971 7392 22983 7395
rect 24118 7392 24124 7404
rect 22971 7364 24124 7392
rect 22971 7361 22983 7364
rect 22925 7355 22983 7361
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 24213 7395 24271 7401
rect 24213 7361 24225 7395
rect 24259 7392 24271 7395
rect 24302 7392 24308 7404
rect 24259 7364 24308 7392
rect 24259 7361 24271 7364
rect 24213 7355 24271 7361
rect 24302 7352 24308 7364
rect 24360 7352 24366 7404
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7392 24455 7395
rect 24486 7392 24492 7404
rect 24443 7364 24492 7392
rect 24443 7361 24455 7364
rect 24397 7355 24455 7361
rect 24486 7352 24492 7364
rect 24544 7352 24550 7404
rect 21358 7284 21364 7336
rect 21416 7324 21422 7336
rect 23109 7327 23167 7333
rect 23109 7324 23121 7327
rect 21416 7296 23121 7324
rect 21416 7284 21422 7296
rect 23109 7293 23121 7296
rect 23155 7293 23167 7327
rect 23750 7324 23756 7336
rect 23711 7296 23756 7324
rect 23109 7287 23167 7293
rect 17911 7228 19380 7256
rect 19521 7259 19579 7265
rect 17911 7225 17923 7228
rect 17865 7219 17923 7225
rect 19521 7225 19533 7259
rect 19567 7256 19579 7259
rect 19978 7256 19984 7268
rect 19567 7228 19984 7256
rect 19567 7225 19579 7228
rect 19521 7219 19579 7225
rect 16114 7188 16120 7200
rect 12268 7160 16120 7188
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 17604 7188 17632 7219
rect 19978 7216 19984 7228
rect 20036 7256 20042 7268
rect 20162 7256 20168 7268
rect 20036 7228 20168 7256
rect 20036 7216 20042 7228
rect 20162 7216 20168 7228
rect 20220 7216 20226 7268
rect 23124 7256 23152 7287
rect 23750 7284 23756 7296
rect 23808 7284 23814 7336
rect 23845 7327 23903 7333
rect 23845 7293 23857 7327
rect 23891 7293 23903 7327
rect 23845 7287 23903 7293
rect 23382 7256 23388 7268
rect 23124 7228 23388 7256
rect 23382 7216 23388 7228
rect 23440 7256 23446 7268
rect 23860 7256 23888 7287
rect 23440 7228 23888 7256
rect 23440 7216 23446 7228
rect 18138 7188 18144 7200
rect 17604 7160 18144 7188
rect 18138 7148 18144 7160
rect 18196 7148 18202 7200
rect 20254 7148 20260 7200
rect 20312 7188 20318 7200
rect 20349 7191 20407 7197
rect 20349 7188 20361 7191
rect 20312 7160 20361 7188
rect 20312 7148 20318 7160
rect 20349 7157 20361 7160
rect 20395 7157 20407 7191
rect 20349 7151 20407 7157
rect 22278 7148 22284 7200
rect 22336 7188 22342 7200
rect 22465 7191 22523 7197
rect 22465 7188 22477 7191
rect 22336 7160 22477 7188
rect 22336 7148 22342 7160
rect 22465 7157 22477 7160
rect 22511 7157 22523 7191
rect 22465 7151 22523 7157
rect 22554 7148 22560 7200
rect 22612 7188 22618 7200
rect 23293 7191 23351 7197
rect 23293 7188 23305 7191
rect 22612 7160 23305 7188
rect 22612 7148 22618 7160
rect 23293 7157 23305 7160
rect 23339 7157 23351 7191
rect 23293 7151 23351 7157
rect 24489 7191 24547 7197
rect 24489 7157 24501 7191
rect 24535 7188 24547 7191
rect 24854 7188 24860 7200
rect 24535 7160 24860 7188
rect 24535 7157 24547 7160
rect 24489 7151 24547 7157
rect 24854 7148 24860 7160
rect 24912 7148 24918 7200
rect 1104 7098 26128 7120
rect 1104 7046 5120 7098
rect 5172 7046 5184 7098
rect 5236 7046 5248 7098
rect 5300 7046 5312 7098
rect 5364 7046 5376 7098
rect 5428 7046 13462 7098
rect 13514 7046 13526 7098
rect 13578 7046 13590 7098
rect 13642 7046 13654 7098
rect 13706 7046 13718 7098
rect 13770 7046 21803 7098
rect 21855 7046 21867 7098
rect 21919 7046 21931 7098
rect 21983 7046 21995 7098
rect 22047 7046 22059 7098
rect 22111 7046 26128 7098
rect 1104 7024 26128 7046
rect 12161 6987 12219 6993
rect 12161 6953 12173 6987
rect 12207 6984 12219 6987
rect 12250 6984 12256 6996
rect 12207 6956 12256 6984
rect 12207 6953 12219 6956
rect 12161 6947 12219 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 13170 6984 13176 6996
rect 12406 6956 13176 6984
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 10744 6888 11100 6916
rect 10744 6876 10750 6888
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 4525 6851 4583 6857
rect 4525 6848 4537 6851
rect 4396 6820 4537 6848
rect 4396 6808 4402 6820
rect 4525 6817 4537 6820
rect 4571 6817 4583 6851
rect 4525 6811 4583 6817
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 6454 6848 6460 6860
rect 5684 6820 6224 6848
rect 6415 6820 6460 6848
rect 5684 6808 5690 6820
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6196 6780 6224 6820
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 7006 6848 7012 6860
rect 6871 6820 7012 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 8021 6851 8079 6857
rect 8021 6848 8033 6851
rect 7616 6820 8033 6848
rect 7616 6808 7622 6820
rect 6254 6783 6312 6789
rect 6254 6780 6266 6783
rect 6196 6752 6266 6780
rect 6089 6743 6147 6749
rect 6254 6749 6266 6752
rect 6300 6749 6312 6783
rect 6254 6743 6312 6749
rect 4792 6715 4850 6721
rect 4792 6681 4804 6715
rect 4838 6712 4850 6715
rect 5534 6712 5540 6724
rect 4838 6684 5540 6712
rect 4838 6681 4850 6684
rect 4792 6675 4850 6681
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 6104 6712 6132 6743
rect 6362 6740 6368 6792
rect 6420 6780 6426 6792
rect 6641 6783 6699 6789
rect 6420 6752 6465 6780
rect 6420 6740 6426 6752
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 6730 6780 6736 6792
rect 6687 6752 6736 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 7852 6789 7880 6820
rect 8021 6817 8033 6820
rect 8067 6817 8079 6851
rect 11072 6848 11100 6888
rect 12406 6860 12434 6956
rect 13170 6944 13176 6956
rect 13228 6984 13234 6996
rect 20349 6987 20407 6993
rect 13228 6956 20300 6984
rect 13228 6944 13234 6956
rect 12618 6876 12624 6928
rect 12676 6916 12682 6928
rect 13357 6919 13415 6925
rect 13357 6916 13369 6919
rect 12676 6888 13369 6916
rect 12676 6876 12682 6888
rect 13357 6885 13369 6888
rect 13403 6916 13415 6919
rect 13541 6919 13599 6925
rect 13541 6916 13553 6919
rect 13403 6888 13553 6916
rect 13403 6885 13415 6888
rect 13357 6879 13415 6885
rect 13541 6885 13553 6888
rect 13587 6885 13599 6919
rect 13541 6879 13599 6885
rect 20165 6919 20223 6925
rect 20165 6885 20177 6919
rect 20211 6885 20223 6919
rect 20272 6916 20300 6956
rect 20349 6953 20361 6987
rect 20395 6984 20407 6987
rect 20530 6984 20536 6996
rect 20395 6956 20536 6984
rect 20395 6953 20407 6956
rect 20349 6947 20407 6953
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 23750 6944 23756 6996
rect 23808 6984 23814 6996
rect 24949 6987 25007 6993
rect 24949 6984 24961 6987
rect 23808 6956 24961 6984
rect 23808 6944 23814 6956
rect 24949 6953 24961 6956
rect 24995 6953 25007 6987
rect 24949 6947 25007 6953
rect 21634 6916 21640 6928
rect 20272 6888 21640 6916
rect 20165 6879 20223 6885
rect 12406 6848 12440 6860
rect 11072 6820 12440 6848
rect 8021 6811 8079 6817
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 15470 6848 15476 6860
rect 13136 6820 13308 6848
rect 15431 6820 15476 6848
rect 13136 6808 13142 6820
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 7883 6752 7917 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 10134 6740 10140 6792
rect 10192 6789 10198 6792
rect 10192 6780 10204 6789
rect 10413 6783 10471 6789
rect 10192 6752 10237 6780
rect 10192 6743 10204 6752
rect 10413 6749 10425 6783
rect 10459 6780 10471 6783
rect 10502 6780 10508 6792
rect 10459 6752 10508 6780
rect 10459 6749 10471 6752
rect 10413 6743 10471 6749
rect 10192 6740 10198 6743
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6780 12127 6783
rect 12250 6780 12256 6792
rect 12115 6752 12256 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 13170 6780 13176 6792
rect 13131 6752 13176 6780
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 13280 6789 13308 6820
rect 15470 6808 15476 6820
rect 15528 6848 15534 6860
rect 16298 6848 16304 6860
rect 15528 6820 16304 6848
rect 15528 6808 15534 6820
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 16574 6808 16580 6860
rect 16632 6808 16638 6860
rect 20180 6848 20208 6879
rect 21634 6876 21640 6888
rect 21692 6876 21698 6928
rect 22465 6919 22523 6925
rect 22465 6885 22477 6919
rect 22511 6916 22523 6919
rect 22554 6916 22560 6928
rect 22511 6888 22560 6916
rect 22511 6885 22523 6888
rect 22465 6879 22523 6885
rect 22554 6876 22560 6888
rect 22612 6876 22618 6928
rect 24121 6919 24179 6925
rect 24121 6885 24133 6919
rect 24167 6914 24179 6919
rect 24167 6886 24201 6914
rect 24167 6885 24179 6886
rect 24121 6879 24179 6885
rect 20346 6848 20352 6860
rect 20180 6820 20352 6848
rect 20346 6808 20352 6820
rect 20404 6808 20410 6860
rect 22738 6848 22744 6860
rect 22699 6820 22744 6848
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 24136 6848 24164 6879
rect 24854 6876 24860 6928
rect 24912 6876 24918 6928
rect 24486 6848 24492 6860
rect 24136 6820 24492 6848
rect 24486 6808 24492 6820
rect 24544 6808 24550 6860
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 6914 6712 6920 6724
rect 5644 6684 6040 6712
rect 6104 6684 6920 6712
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 5644 6644 5672 6684
rect 5902 6644 5908 6656
rect 3476 6616 5672 6644
rect 5863 6616 5908 6644
rect 3476 6604 3482 6616
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6012 6644 6040 6684
rect 6914 6672 6920 6684
rect 6972 6672 6978 6724
rect 13280 6712 13308 6743
rect 14182 6740 14188 6792
rect 14240 6780 14246 6792
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 14240 6752 14657 6780
rect 14240 6740 14246 6752
rect 14645 6749 14657 6752
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6780 15347 6783
rect 15654 6780 15660 6792
rect 15335 6752 15660 6780
rect 15335 6749 15347 6752
rect 15289 6743 15347 6749
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6780 16175 6783
rect 16592 6780 16620 6808
rect 16758 6780 16764 6792
rect 16163 6752 16620 6780
rect 16719 6752 16764 6780
rect 16163 6749 16175 6752
rect 16117 6743 16175 6749
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 20959 6783 21017 6789
rect 20959 6749 20971 6783
rect 21005 6780 21017 6783
rect 21266 6780 21272 6792
rect 21005 6752 21128 6780
rect 21227 6752 21272 6780
rect 21005 6749 21017 6752
rect 20959 6743 21017 6749
rect 7024 6684 13308 6712
rect 7024 6644 7052 6684
rect 15838 6672 15844 6724
rect 15896 6712 15902 6724
rect 16390 6712 16396 6724
rect 15896 6684 16396 6712
rect 15896 6672 15902 6684
rect 16390 6672 16396 6684
rect 16448 6712 16454 6724
rect 16577 6715 16635 6721
rect 16577 6712 16589 6715
rect 16448 6684 16589 6712
rect 16448 6672 16454 6684
rect 16577 6681 16589 6684
rect 16623 6681 16635 6715
rect 16577 6675 16635 6681
rect 19058 6672 19064 6724
rect 19116 6712 19122 6724
rect 19889 6715 19947 6721
rect 19889 6712 19901 6715
rect 19116 6684 19901 6712
rect 19116 6672 19122 6684
rect 19889 6681 19901 6684
rect 19935 6712 19947 6715
rect 21100 6712 21128 6752
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6780 21419 6783
rect 21450 6780 21456 6792
rect 21407 6752 21456 6780
rect 21407 6749 21419 6752
rect 21361 6743 21419 6749
rect 21450 6740 21456 6752
rect 21508 6740 21514 6792
rect 23014 6789 23020 6792
rect 23008 6743 23020 6789
rect 23072 6780 23078 6792
rect 24394 6780 24400 6792
rect 23072 6752 23108 6780
rect 24355 6752 24400 6780
rect 23014 6740 23020 6743
rect 23072 6740 23078 6752
rect 24394 6740 24400 6752
rect 24452 6740 24458 6792
rect 24872 6789 24900 6876
rect 24856 6783 24914 6789
rect 24856 6749 24868 6783
rect 24902 6749 24914 6783
rect 24856 6743 24914 6749
rect 21542 6712 21548 6724
rect 19935 6684 20944 6712
rect 21100 6684 21548 6712
rect 19935 6681 19947 6684
rect 19889 6675 19947 6681
rect 7742 6644 7748 6656
rect 6012 6616 7052 6644
rect 7703 6616 7748 6644
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 9030 6644 9036 6656
rect 8991 6616 9036 6644
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 12986 6644 12992 6656
rect 12947 6616 12992 6644
rect 12986 6604 12992 6616
rect 13044 6604 13050 6656
rect 14826 6644 14832 6656
rect 14787 6616 14832 6644
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 14918 6604 14924 6656
rect 14976 6644 14982 6656
rect 14976 6616 15021 6644
rect 14976 6604 14982 6616
rect 15378 6604 15384 6656
rect 15436 6644 15442 6656
rect 15436 6616 15481 6644
rect 15436 6604 15442 6616
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 15749 6647 15807 6653
rect 15749 6644 15761 6647
rect 15620 6616 15761 6644
rect 15620 6604 15626 6616
rect 15749 6613 15761 6616
rect 15795 6613 15807 6647
rect 15749 6607 15807 6613
rect 16209 6647 16267 6653
rect 16209 6613 16221 6647
rect 16255 6644 16267 6647
rect 16758 6644 16764 6656
rect 16255 6616 16764 6644
rect 16255 6613 16267 6616
rect 16209 6607 16267 6613
rect 16758 6604 16764 6616
rect 16816 6604 16822 6656
rect 20806 6644 20812 6656
rect 20767 6616 20812 6644
rect 20806 6604 20812 6616
rect 20864 6604 20870 6656
rect 20916 6644 20944 6684
rect 21542 6672 21548 6684
rect 21600 6672 21606 6724
rect 22097 6715 22155 6721
rect 22097 6681 22109 6715
rect 22143 6712 22155 6715
rect 22370 6712 22376 6724
rect 22143 6684 22376 6712
rect 22143 6681 22155 6684
rect 22097 6675 22155 6681
rect 22112 6644 22140 6675
rect 22370 6672 22376 6684
rect 22428 6672 22434 6724
rect 20916 6616 22140 6644
rect 22557 6647 22615 6653
rect 22557 6613 22569 6647
rect 22603 6644 22615 6647
rect 23290 6644 23296 6656
rect 22603 6616 23296 6644
rect 22603 6613 22615 6616
rect 22557 6607 22615 6613
rect 23290 6604 23296 6616
rect 23348 6604 23354 6656
rect 1104 6554 26128 6576
rect 1104 6502 9291 6554
rect 9343 6502 9355 6554
rect 9407 6502 9419 6554
rect 9471 6502 9483 6554
rect 9535 6502 9547 6554
rect 9599 6502 17632 6554
rect 17684 6502 17696 6554
rect 17748 6502 17760 6554
rect 17812 6502 17824 6554
rect 17876 6502 17888 6554
rect 17940 6502 26128 6554
rect 1104 6480 26128 6502
rect 3329 6443 3387 6449
rect 3329 6440 3341 6443
rect 2746 6412 3341 6440
rect 1857 6375 1915 6381
rect 1857 6341 1869 6375
rect 1903 6372 1915 6375
rect 2746 6372 2774 6412
rect 3329 6409 3341 6412
rect 3375 6409 3387 6443
rect 4157 6443 4215 6449
rect 4157 6440 4169 6443
rect 3329 6403 3387 6409
rect 3896 6412 4169 6440
rect 3234 6372 3240 6384
rect 1903 6344 2452 6372
rect 1903 6341 1915 6344
rect 1857 6335 1915 6341
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6304 2007 6307
rect 2038 6304 2044 6316
rect 1995 6276 2044 6304
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2148 6168 2176 6267
rect 2424 6236 2452 6344
rect 2700 6344 2774 6372
rect 2884 6344 3240 6372
rect 2700 6313 2728 6344
rect 2884 6313 2912 6344
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 3896 6381 3924 6412
rect 4157 6409 4169 6412
rect 4203 6440 4215 6443
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 4203 6412 4629 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 5534 6440 5540 6452
rect 5495 6412 5540 6440
rect 4617 6403 4675 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 9214 6440 9220 6452
rect 8444 6412 9220 6440
rect 8444 6400 8450 6412
rect 9214 6400 9220 6412
rect 9272 6440 9278 6452
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 9272 6412 9413 6440
rect 9272 6400 9278 6412
rect 9401 6409 9413 6412
rect 9447 6409 9459 6443
rect 12434 6440 12440 6452
rect 9401 6403 9459 6409
rect 12406 6400 12440 6440
rect 12492 6400 12498 6452
rect 14182 6440 14188 6452
rect 14143 6412 14188 6440
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 14918 6440 14924 6452
rect 14568 6412 14924 6440
rect 3881 6375 3939 6381
rect 3881 6341 3893 6375
rect 3927 6341 3939 6375
rect 3881 6335 3939 6341
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 4522 6372 4528 6384
rect 4120 6344 4528 6372
rect 4120 6332 4126 6344
rect 4522 6332 4528 6344
rect 4580 6372 4586 6384
rect 4709 6375 4767 6381
rect 4709 6372 4721 6375
rect 4580 6344 4721 6372
rect 4580 6332 4586 6344
rect 4709 6341 4721 6344
rect 4755 6372 4767 6375
rect 6362 6372 6368 6384
rect 4755 6344 5019 6372
rect 4755 6341 4767 6344
rect 4709 6335 4767 6341
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6273 2743 6307
rect 2685 6267 2743 6273
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6273 2927 6307
rect 3050 6304 3056 6316
rect 3011 6276 3056 6304
rect 2869 6267 2927 6273
rect 2884 6236 2912 6267
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 3326 6304 3332 6316
rect 3287 6276 3332 6304
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 3602 6264 3608 6316
rect 3660 6304 3666 6316
rect 3973 6307 4031 6313
rect 3973 6304 3985 6307
rect 3660 6276 3985 6304
rect 3660 6264 3666 6276
rect 3973 6273 3985 6276
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 4893 6307 4951 6313
rect 4893 6304 4905 6307
rect 4212 6276 4905 6304
rect 4212 6264 4218 6276
rect 4893 6273 4905 6276
rect 4939 6273 4951 6307
rect 4991 6304 5019 6344
rect 5184 6344 6368 6372
rect 5184 6313 5212 6344
rect 6362 6332 6368 6344
rect 6420 6332 6426 6384
rect 8288 6375 8346 6381
rect 8288 6341 8300 6375
rect 8334 6372 8346 6375
rect 8478 6372 8484 6384
rect 8334 6344 8484 6372
rect 8334 6341 8346 6344
rect 8288 6335 8346 6341
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 12406 6372 12434 6400
rect 11992 6344 12434 6372
rect 5058 6307 5116 6313
rect 5058 6304 5070 6307
rect 4991 6276 5070 6304
rect 4893 6267 4951 6273
rect 5058 6273 5070 6276
rect 5104 6273 5116 6307
rect 5058 6267 5116 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6304 5503 6307
rect 5810 6304 5816 6316
rect 5491 6276 5816 6304
rect 5491 6273 5503 6276
rect 5445 6267 5503 6273
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 7742 6304 7748 6316
rect 5951 6276 7748 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 11514 6304 11520 6316
rect 7852 6276 11520 6304
rect 2424 6208 2912 6236
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6236 3295 6239
rect 3418 6236 3424 6248
rect 3283 6208 3424 6236
rect 3283 6205 3295 6208
rect 3237 6199 3295 6205
rect 3418 6196 3424 6208
rect 3476 6196 3482 6248
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 6454 6236 6460 6248
rect 5307 6208 6460 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 6454 6196 6460 6208
rect 6512 6196 6518 6248
rect 2685 6171 2743 6177
rect 2685 6168 2697 6171
rect 2148 6140 2697 6168
rect 2685 6137 2697 6140
rect 2731 6137 2743 6171
rect 2685 6131 2743 6137
rect 4338 6128 4344 6180
rect 4396 6168 4402 6180
rect 5721 6171 5779 6177
rect 5721 6168 5733 6171
rect 4396 6140 5733 6168
rect 4396 6128 4402 6140
rect 5721 6137 5733 6140
rect 5767 6168 5779 6171
rect 6362 6168 6368 6180
rect 5767 6140 6368 6168
rect 5767 6137 5779 6140
rect 5721 6131 5779 6137
rect 6362 6128 6368 6140
rect 6420 6128 6426 6180
rect 2314 6100 2320 6112
rect 2275 6072 2320 6100
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 4617 6103 4675 6109
rect 4617 6069 4629 6103
rect 4663 6100 4675 6103
rect 7852 6100 7880 6276
rect 11514 6264 11520 6276
rect 11572 6264 11578 6316
rect 11992 6313 12020 6344
rect 11609 6307 11667 6313
rect 11609 6273 11621 6307
rect 11655 6304 11667 6307
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 11655 6276 11989 6304
rect 11655 6273 11667 6276
rect 11609 6267 11667 6273
rect 11977 6273 11989 6276
rect 12023 6273 12035 6307
rect 12158 6304 12164 6316
rect 12119 6276 12164 6304
rect 11977 6267 12035 6273
rect 12158 6264 12164 6276
rect 12216 6264 12222 6316
rect 7926 6196 7932 6248
rect 7984 6236 7990 6248
rect 8021 6239 8079 6245
rect 8021 6236 8033 6239
rect 7984 6208 8033 6236
rect 7984 6196 7990 6208
rect 8021 6205 8033 6208
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 9950 6196 9956 6248
rect 10008 6236 10014 6248
rect 13906 6236 13912 6248
rect 10008 6208 13912 6236
rect 10008 6196 10014 6208
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 14369 6171 14427 6177
rect 14369 6137 14381 6171
rect 14415 6168 14427 6171
rect 14568 6168 14596 6412
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 15010 6400 15016 6452
rect 15068 6400 15074 6452
rect 16758 6440 16764 6452
rect 16719 6412 16764 6440
rect 16758 6400 16764 6412
rect 16816 6400 16822 6452
rect 18969 6443 19027 6449
rect 18969 6409 18981 6443
rect 19015 6440 19027 6443
rect 19058 6440 19064 6452
rect 19015 6412 19064 6440
rect 19015 6409 19027 6412
rect 18969 6403 19027 6409
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19429 6443 19487 6449
rect 19429 6409 19441 6443
rect 19475 6440 19487 6443
rect 19702 6440 19708 6452
rect 19475 6412 19708 6440
rect 19475 6409 19487 6412
rect 19429 6403 19487 6409
rect 19702 6400 19708 6412
rect 19760 6400 19766 6452
rect 20346 6440 20352 6452
rect 20307 6412 20352 6440
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 20806 6440 20812 6452
rect 20767 6412 20812 6440
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 21174 6400 21180 6452
rect 21232 6400 21238 6452
rect 22097 6443 22155 6449
rect 22097 6409 22109 6443
rect 22143 6409 22155 6443
rect 22097 6403 22155 6409
rect 15028 6372 15056 6400
rect 14752 6344 15056 6372
rect 14752 6313 14780 6344
rect 15102 6332 15108 6384
rect 15160 6372 15166 6384
rect 19518 6372 19524 6384
rect 15160 6344 19524 6372
rect 15160 6332 15166 6344
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6273 14795 6307
rect 14737 6267 14795 6273
rect 14826 6264 14832 6316
rect 14884 6304 14890 6316
rect 14993 6307 15051 6313
rect 14993 6304 15005 6307
rect 14884 6276 15005 6304
rect 14884 6264 14890 6276
rect 14993 6273 15005 6276
rect 15039 6273 15051 6307
rect 14993 6267 15051 6273
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 16485 6307 16543 6313
rect 16485 6304 16497 6307
rect 15804 6276 16497 6304
rect 15804 6264 15810 6276
rect 16485 6273 16497 6276
rect 16531 6273 16543 6307
rect 16485 6267 16543 6273
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 18800 6313 18828 6344
rect 19518 6332 19524 6344
rect 19576 6332 19582 6384
rect 19794 6332 19800 6384
rect 19852 6372 19858 6384
rect 20073 6375 20131 6381
rect 20073 6372 20085 6375
rect 19852 6344 20085 6372
rect 19852 6332 19858 6344
rect 20073 6341 20085 6344
rect 20119 6341 20131 6375
rect 20073 6335 20131 6341
rect 20717 6375 20775 6381
rect 20717 6341 20729 6375
rect 20763 6372 20775 6375
rect 21192 6372 21220 6400
rect 20763 6344 21220 6372
rect 20763 6341 20775 6344
rect 20717 6335 20775 6341
rect 21266 6332 21272 6384
rect 21324 6372 21330 6384
rect 21361 6375 21419 6381
rect 21361 6372 21373 6375
rect 21324 6344 21373 6372
rect 21324 6332 21330 6344
rect 21361 6341 21373 6344
rect 21407 6341 21419 6375
rect 21542 6372 21548 6384
rect 21503 6344 21548 6372
rect 21361 6335 21419 6341
rect 21542 6332 21548 6344
rect 21600 6332 21606 6384
rect 22112 6372 22140 6403
rect 24118 6400 24124 6452
rect 24176 6440 24182 6452
rect 24305 6443 24363 6449
rect 24305 6440 24317 6443
rect 24176 6412 24317 6440
rect 24176 6400 24182 6412
rect 24305 6409 24317 6412
rect 24351 6409 24363 6443
rect 24305 6403 24363 6409
rect 22434 6375 22492 6381
rect 22434 6372 22446 6375
rect 22112 6344 22446 6372
rect 22434 6341 22446 6344
rect 22480 6341 22492 6375
rect 22434 6335 22492 6341
rect 16854 6307 16912 6313
rect 16854 6304 16866 6307
rect 16632 6276 16866 6304
rect 16632 6264 16638 6276
rect 16854 6273 16866 6276
rect 16900 6273 16912 6307
rect 16854 6267 16912 6273
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 19242 6264 19248 6316
rect 19300 6304 19306 6316
rect 19889 6307 19947 6313
rect 19889 6304 19901 6307
rect 19300 6276 19901 6304
rect 19300 6264 19306 6276
rect 19889 6273 19901 6276
rect 19935 6273 19947 6307
rect 19889 6267 19947 6273
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6304 21235 6307
rect 21450 6304 21456 6316
rect 21223 6276 21456 6304
rect 21223 6273 21235 6276
rect 21177 6267 21235 6273
rect 21450 6264 21456 6276
rect 21508 6264 21514 6316
rect 14642 6196 14648 6248
rect 14700 6236 14706 6248
rect 14700 6208 14745 6236
rect 14700 6196 14706 6208
rect 17126 6196 17132 6248
rect 17184 6236 17190 6248
rect 17221 6239 17279 6245
rect 17221 6236 17233 6239
rect 17184 6208 17233 6236
rect 17184 6196 17190 6208
rect 17221 6205 17233 6208
rect 17267 6205 17279 6239
rect 17221 6199 17279 6205
rect 17310 6196 17316 6248
rect 17368 6236 17374 6248
rect 17368 6208 17413 6236
rect 17368 6196 17374 6208
rect 19334 6196 19340 6248
rect 19392 6236 19398 6248
rect 19521 6239 19579 6245
rect 19521 6236 19533 6239
rect 19392 6208 19533 6236
rect 19392 6196 19398 6208
rect 19521 6205 19533 6208
rect 19567 6205 19579 6239
rect 19521 6199 19579 6205
rect 19613 6239 19671 6245
rect 19613 6205 19625 6239
rect 19659 6236 19671 6239
rect 20901 6239 20959 6245
rect 20901 6236 20913 6239
rect 19659 6208 20913 6236
rect 19659 6205 19671 6208
rect 19613 6199 19671 6205
rect 20901 6205 20913 6208
rect 20947 6236 20959 6239
rect 21358 6236 21364 6248
rect 20947 6208 21364 6236
rect 20947 6205 20959 6208
rect 20901 6199 20959 6205
rect 14415 6140 14596 6168
rect 16117 6171 16175 6177
rect 14415 6137 14427 6140
rect 14369 6131 14427 6137
rect 16117 6137 16129 6171
rect 16163 6168 16175 6171
rect 17494 6168 17500 6180
rect 16163 6140 17500 6168
rect 16163 6137 16175 6140
rect 16117 6131 16175 6137
rect 4663 6072 7880 6100
rect 4663 6069 4675 6072
rect 4617 6063 4675 6069
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 8076 6072 11805 6100
rect 8076 6060 8082 6072
rect 11793 6069 11805 6072
rect 11839 6069 11851 6103
rect 11793 6063 11851 6069
rect 12161 6103 12219 6109
rect 12161 6069 12173 6103
rect 12207 6100 12219 6103
rect 12250 6100 12256 6112
rect 12207 6072 12256 6100
rect 12207 6069 12219 6072
rect 12161 6063 12219 6069
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 15654 6060 15660 6112
rect 15712 6100 15718 6112
rect 16132 6100 16160 6131
rect 17494 6128 17500 6140
rect 17552 6128 17558 6180
rect 19628 6168 19656 6199
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 21468 6168 21496 6264
rect 18984 6140 19656 6168
rect 20180 6140 21496 6168
rect 16298 6100 16304 6112
rect 15712 6072 16160 6100
rect 16259 6072 16304 6100
rect 15712 6060 15718 6072
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 18984 6100 19012 6140
rect 16448 6072 19012 6100
rect 16448 6060 16454 6072
rect 19058 6060 19064 6112
rect 19116 6100 19122 6112
rect 19116 6072 19161 6100
rect 19116 6060 19122 6072
rect 19610 6060 19616 6112
rect 19668 6100 19674 6112
rect 20180 6109 20208 6140
rect 20165 6103 20223 6109
rect 20165 6100 20177 6103
rect 19668 6072 20177 6100
rect 19668 6060 19674 6072
rect 20165 6069 20177 6072
rect 20211 6069 20223 6103
rect 21560 6100 21588 6332
rect 21913 6307 21971 6313
rect 21913 6273 21925 6307
rect 21959 6304 21971 6307
rect 22094 6304 22100 6316
rect 21959 6276 22100 6304
rect 21959 6273 21971 6276
rect 21913 6267 21971 6273
rect 22094 6264 22100 6276
rect 22152 6264 22158 6316
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6304 22247 6307
rect 22738 6304 22744 6316
rect 22235 6276 22744 6304
rect 22235 6273 22247 6276
rect 22189 6267 22247 6273
rect 22738 6264 22744 6276
rect 22796 6264 22802 6316
rect 23658 6264 23664 6316
rect 23716 6304 23722 6316
rect 24155 6307 24213 6313
rect 24155 6304 24167 6307
rect 23716 6276 24167 6304
rect 23716 6264 23722 6276
rect 24155 6273 24167 6276
rect 24201 6304 24213 6307
rect 24394 6304 24400 6316
rect 24201 6276 24400 6304
rect 24201 6273 24213 6276
rect 24155 6267 24213 6273
rect 24394 6264 24400 6276
rect 24452 6264 24458 6316
rect 23753 6239 23811 6245
rect 23753 6236 23765 6239
rect 23216 6208 23765 6236
rect 23216 6100 23244 6208
rect 23753 6205 23765 6208
rect 23799 6205 23811 6239
rect 23753 6199 23811 6205
rect 23845 6239 23903 6245
rect 23845 6205 23857 6239
rect 23891 6205 23903 6239
rect 23845 6199 23903 6205
rect 23860 6168 23888 6199
rect 23584 6140 23888 6168
rect 23584 6112 23612 6140
rect 23290 6100 23296 6112
rect 21560 6072 23296 6100
rect 20165 6063 20223 6069
rect 23290 6060 23296 6072
rect 23348 6060 23354 6112
rect 23566 6100 23572 6112
rect 23527 6072 23572 6100
rect 23566 6060 23572 6072
rect 23624 6060 23630 6112
rect 1104 6010 26128 6032
rect 1104 5958 5120 6010
rect 5172 5958 5184 6010
rect 5236 5958 5248 6010
rect 5300 5958 5312 6010
rect 5364 5958 5376 6010
rect 5428 5958 13462 6010
rect 13514 5958 13526 6010
rect 13578 5958 13590 6010
rect 13642 5958 13654 6010
rect 13706 5958 13718 6010
rect 13770 5958 21803 6010
rect 21855 5958 21867 6010
rect 21919 5958 21931 6010
rect 21983 5958 21995 6010
rect 22047 5958 22059 6010
rect 22111 5958 26128 6010
rect 1104 5936 26128 5958
rect 3050 5856 3056 5908
rect 3108 5896 3114 5908
rect 3145 5899 3203 5905
rect 3145 5896 3157 5899
rect 3108 5868 3157 5896
rect 3108 5856 3114 5868
rect 3145 5865 3157 5868
rect 3191 5865 3203 5899
rect 3145 5859 3203 5865
rect 3160 5828 3188 5859
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8444 5868 8677 5896
rect 8444 5856 8450 5868
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 10870 5856 10876 5908
rect 10928 5896 10934 5908
rect 12713 5899 12771 5905
rect 12713 5896 12725 5899
rect 10928 5868 12725 5896
rect 10928 5856 10934 5868
rect 12713 5865 12725 5868
rect 12759 5865 12771 5899
rect 12713 5859 12771 5865
rect 15197 5899 15255 5905
rect 15197 5865 15209 5899
rect 15243 5896 15255 5899
rect 15378 5896 15384 5908
rect 15243 5868 15384 5896
rect 15243 5865 15255 5868
rect 15197 5859 15255 5865
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 16482 5896 16488 5908
rect 15856 5868 16488 5896
rect 3160 5800 7604 5828
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5760 3019 5763
rect 4338 5760 4344 5772
rect 3007 5732 4344 5760
rect 3007 5729 3019 5732
rect 2961 5723 3019 5729
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 2314 5652 2320 5704
rect 2372 5692 2378 5704
rect 2694 5695 2752 5701
rect 2694 5692 2706 5695
rect 2372 5664 2706 5692
rect 2372 5652 2378 5664
rect 2694 5661 2706 5664
rect 2740 5661 2752 5695
rect 2694 5655 2752 5661
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5692 5503 5695
rect 5534 5692 5540 5704
rect 5491 5664 5540 5692
rect 5491 5661 5503 5664
rect 5445 5655 5503 5661
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 6546 5624 6552 5636
rect 5276 5596 6552 5624
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 2038 5556 2044 5568
rect 1627 5528 2044 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5276 5565 5304 5596
rect 6546 5584 6552 5596
rect 6604 5584 6610 5636
rect 5261 5559 5319 5565
rect 5261 5556 5273 5559
rect 4948 5528 5273 5556
rect 4948 5516 4954 5528
rect 5261 5525 5273 5528
rect 5307 5525 5319 5559
rect 5261 5519 5319 5525
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 5905 5559 5963 5565
rect 5905 5556 5917 5559
rect 5776 5528 5917 5556
rect 5776 5516 5782 5528
rect 5905 5525 5917 5528
rect 5951 5556 5963 5559
rect 6270 5556 6276 5568
rect 5951 5528 6276 5556
rect 5951 5525 5963 5528
rect 5905 5519 5963 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 7576 5556 7604 5800
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 7984 5800 9444 5828
rect 7984 5788 7990 5800
rect 8662 5760 8668 5772
rect 8423 5732 8668 5760
rect 8202 5692 8208 5704
rect 8163 5664 8208 5692
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 8423 5701 8451 5732
rect 8662 5720 8668 5732
rect 8720 5720 8726 5772
rect 8389 5695 8451 5701
rect 8389 5661 8401 5695
rect 8435 5661 8451 5695
rect 8389 5660 8451 5661
rect 8389 5655 8447 5660
rect 8479 5652 8485 5704
rect 8537 5692 8543 5704
rect 8754 5692 8760 5704
rect 8537 5664 8581 5692
rect 8715 5664 8760 5692
rect 8537 5652 8543 5664
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 7742 5584 7748 5636
rect 7800 5624 7806 5636
rect 9416 5633 9444 5800
rect 11146 5788 11152 5840
rect 11204 5828 11210 5840
rect 11701 5831 11759 5837
rect 11701 5828 11713 5831
rect 11204 5800 11713 5828
rect 11204 5788 11210 5800
rect 11701 5797 11713 5800
rect 11747 5797 11759 5831
rect 11701 5791 11759 5797
rect 12986 5788 12992 5840
rect 13044 5788 13050 5840
rect 12250 5760 12256 5772
rect 12211 5732 12256 5760
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 13004 5760 13032 5788
rect 15654 5760 15660 5772
rect 12912 5732 14872 5760
rect 15615 5732 15660 5760
rect 11422 5692 11428 5704
rect 11383 5664 11428 5692
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 11514 5652 11520 5704
rect 11572 5692 11578 5704
rect 12912 5701 12940 5732
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11572 5664 12081 5692
rect 11572 5652 11578 5664
rect 12069 5661 12081 5664
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 12986 5652 12992 5704
rect 13044 5692 13050 5704
rect 14844 5701 14872 5732
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 15856 5760 15884 5868
rect 16482 5856 16488 5868
rect 16540 5856 16546 5908
rect 19334 5896 19340 5908
rect 19295 5868 19340 5896
rect 19334 5856 19340 5868
rect 19392 5856 19398 5908
rect 21266 5856 21272 5908
rect 21324 5896 21330 5908
rect 21361 5899 21419 5905
rect 21361 5896 21373 5899
rect 21324 5868 21373 5896
rect 21324 5856 21330 5868
rect 21361 5865 21373 5868
rect 21407 5865 21419 5899
rect 21361 5859 21419 5865
rect 22186 5856 22192 5908
rect 22244 5896 22250 5908
rect 22373 5899 22431 5905
rect 22373 5896 22385 5899
rect 22244 5868 22385 5896
rect 22244 5856 22250 5868
rect 22373 5865 22385 5868
rect 22419 5865 22431 5899
rect 22373 5859 22431 5865
rect 18601 5831 18659 5837
rect 18601 5797 18613 5831
rect 18647 5797 18659 5831
rect 18601 5791 18659 5797
rect 18785 5831 18843 5837
rect 18785 5797 18797 5831
rect 18831 5828 18843 5831
rect 19058 5828 19064 5840
rect 18831 5800 19064 5828
rect 18831 5797 18843 5800
rect 18785 5791 18843 5797
rect 15795 5732 15884 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 14829 5695 14887 5701
rect 13044 5664 13089 5692
rect 13044 5652 13050 5664
rect 14829 5661 14841 5695
rect 14875 5692 14887 5695
rect 15102 5692 15108 5704
rect 14875 5664 15108 5692
rect 14875 5661 14887 5664
rect 14829 5655 14887 5661
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 15347 5695 15405 5701
rect 15347 5661 15359 5695
rect 15393 5692 15405 5695
rect 15393 5664 15608 5692
rect 15393 5661 15405 5664
rect 15347 5655 15405 5661
rect 9217 5627 9275 5633
rect 9217 5624 9229 5627
rect 7800 5596 9229 5624
rect 7800 5584 7806 5596
rect 9217 5593 9229 5596
rect 9263 5593 9275 5627
rect 9217 5587 9275 5593
rect 9401 5627 9459 5633
rect 9401 5593 9413 5627
rect 9447 5624 9459 5627
rect 10502 5624 10508 5636
rect 9447 5596 10508 5624
rect 9447 5593 9459 5596
rect 9401 5587 9459 5593
rect 10502 5584 10508 5596
rect 10560 5584 10566 5636
rect 11882 5624 11888 5636
rect 11440 5596 11888 5624
rect 11440 5556 11468 5596
rect 11882 5584 11888 5596
rect 11940 5584 11946 5636
rect 12161 5627 12219 5633
rect 12161 5593 12173 5627
rect 12207 5624 12219 5627
rect 13081 5627 13139 5633
rect 13081 5624 13093 5627
rect 12207 5596 13093 5624
rect 12207 5593 12219 5596
rect 12161 5587 12219 5593
rect 13081 5593 13093 5596
rect 13127 5593 13139 5627
rect 15580 5624 15608 5664
rect 15838 5652 15844 5704
rect 15896 5692 15902 5704
rect 17310 5692 17316 5704
rect 15896 5664 15941 5692
rect 16040 5664 17316 5692
rect 15896 5652 15902 5664
rect 16040 5624 16068 5664
rect 17310 5652 17316 5664
rect 17368 5692 17374 5704
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 17368 5664 17785 5692
rect 17368 5652 17374 5664
rect 17773 5661 17785 5664
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18616 5692 18644 5791
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 22278 5828 22284 5840
rect 22239 5800 22284 5828
rect 22278 5788 22284 5800
rect 22336 5788 22342 5840
rect 23658 5828 23664 5840
rect 23619 5800 23664 5828
rect 23658 5788 23664 5800
rect 23716 5788 23722 5840
rect 19978 5760 19984 5772
rect 19939 5732 19984 5760
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 21913 5763 21971 5769
rect 21913 5729 21925 5763
rect 21959 5760 21971 5763
rect 22370 5760 22376 5772
rect 21959 5732 22376 5760
rect 21959 5729 21971 5732
rect 21913 5723 21971 5729
rect 22370 5720 22376 5732
rect 22428 5720 22434 5772
rect 18279 5664 18644 5692
rect 19061 5695 19119 5701
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 19061 5661 19073 5695
rect 19107 5692 19119 5695
rect 19150 5692 19156 5704
rect 19107 5664 19156 5692
rect 19107 5661 19119 5664
rect 19061 5655 19119 5661
rect 19150 5652 19156 5664
rect 19208 5652 19214 5704
rect 19487 5695 19545 5701
rect 19487 5661 19499 5695
rect 19533 5692 19545 5695
rect 19610 5692 19616 5704
rect 19533 5664 19616 5692
rect 19533 5661 19545 5664
rect 19487 5655 19545 5661
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 19794 5692 19800 5704
rect 19755 5664 19800 5692
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 20254 5701 20260 5704
rect 19889 5695 19947 5701
rect 19889 5661 19901 5695
rect 19935 5661 19947 5695
rect 20248 5692 20260 5701
rect 20215 5664 20260 5692
rect 19889 5655 19947 5661
rect 20248 5655 20260 5664
rect 15580 5596 16068 5624
rect 16108 5627 16166 5633
rect 13081 5587 13139 5593
rect 16108 5593 16120 5627
rect 16154 5624 16166 5627
rect 16298 5624 16304 5636
rect 16154 5596 16304 5624
rect 16154 5593 16166 5596
rect 16108 5587 16166 5593
rect 16298 5584 16304 5596
rect 16356 5584 16362 5636
rect 16482 5584 16488 5636
rect 16540 5624 16546 5636
rect 17405 5627 17463 5633
rect 17405 5624 17417 5627
rect 16540 5596 17417 5624
rect 16540 5584 16546 5596
rect 17405 5593 17417 5596
rect 17451 5593 17463 5627
rect 17405 5587 17463 5593
rect 17494 5584 17500 5636
rect 17552 5624 17558 5636
rect 17589 5627 17647 5633
rect 17589 5624 17601 5627
rect 17552 5596 17601 5624
rect 17552 5584 17558 5596
rect 17589 5593 17601 5596
rect 17635 5593 17647 5627
rect 17589 5587 17647 5593
rect 19242 5584 19248 5636
rect 19300 5624 19306 5636
rect 19904 5624 19932 5655
rect 20254 5652 20260 5655
rect 20312 5652 20318 5704
rect 23290 5692 23296 5704
rect 23251 5664 23296 5692
rect 23290 5652 23296 5664
rect 23348 5652 23354 5704
rect 23477 5695 23535 5701
rect 23477 5661 23489 5695
rect 23523 5692 23535 5695
rect 23566 5692 23572 5704
rect 23523 5664 23572 5692
rect 23523 5661 23535 5664
rect 23477 5655 23535 5661
rect 23566 5652 23572 5664
rect 23624 5652 23630 5704
rect 19300 5596 19932 5624
rect 19300 5584 19306 5596
rect 11606 5556 11612 5568
rect 7576 5528 11468 5556
rect 11567 5528 11612 5556
rect 11606 5516 11612 5528
rect 11664 5516 11670 5568
rect 14642 5556 14648 5568
rect 14555 5528 14648 5556
rect 14642 5516 14648 5528
rect 14700 5556 14706 5568
rect 15286 5556 15292 5568
rect 14700 5528 15292 5556
rect 14700 5516 14706 5528
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 17126 5516 17132 5568
rect 17184 5556 17190 5568
rect 17221 5559 17279 5565
rect 17221 5556 17233 5559
rect 17184 5528 17233 5556
rect 17184 5516 17190 5528
rect 17221 5525 17233 5528
rect 17267 5525 17279 5559
rect 18414 5556 18420 5568
rect 18375 5528 18420 5556
rect 17221 5519 17279 5525
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 1104 5466 26128 5488
rect 1104 5414 9291 5466
rect 9343 5414 9355 5466
rect 9407 5414 9419 5466
rect 9471 5414 9483 5466
rect 9535 5414 9547 5466
rect 9599 5414 17632 5466
rect 17684 5414 17696 5466
rect 17748 5414 17760 5466
rect 17812 5414 17824 5466
rect 17876 5414 17888 5466
rect 17940 5414 26128 5466
rect 1104 5392 26128 5414
rect 2777 5355 2835 5361
rect 2777 5321 2789 5355
rect 2823 5321 2835 5355
rect 4985 5355 5043 5361
rect 4985 5352 4997 5355
rect 2777 5315 2835 5321
rect 4724 5324 4997 5352
rect 2792 5284 2820 5315
rect 3326 5284 3332 5296
rect 2792 5256 3332 5284
rect 3326 5244 3332 5256
rect 3384 5284 3390 5296
rect 4724 5293 4752 5324
rect 4985 5321 4997 5324
rect 5031 5321 5043 5355
rect 4985 5315 5043 5321
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8478 5352 8484 5364
rect 8168 5324 8484 5352
rect 8168 5312 8174 5324
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 8754 5312 8760 5364
rect 8812 5352 8818 5364
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 8812 5324 9321 5352
rect 8812 5312 8818 5324
rect 9309 5321 9321 5324
rect 9355 5352 9367 5355
rect 9861 5355 9919 5361
rect 9861 5352 9873 5355
rect 9355 5324 9873 5352
rect 9355 5321 9367 5324
rect 9309 5315 9367 5321
rect 9861 5321 9873 5324
rect 9907 5321 9919 5355
rect 9861 5315 9919 5321
rect 11241 5355 11299 5361
rect 11241 5321 11253 5355
rect 11287 5352 11299 5355
rect 11422 5352 11428 5364
rect 11287 5324 11428 5352
rect 11287 5321 11299 5324
rect 11241 5315 11299 5321
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 15657 5355 15715 5361
rect 15657 5321 15669 5355
rect 15703 5352 15715 5355
rect 15746 5352 15752 5364
rect 15703 5324 15752 5352
rect 15703 5321 15715 5324
rect 15657 5315 15715 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16393 5355 16451 5361
rect 16393 5321 16405 5355
rect 16439 5352 16451 5355
rect 16574 5352 16580 5364
rect 16439 5324 16580 5352
rect 16439 5321 16451 5324
rect 16393 5315 16451 5321
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 16942 5312 16948 5364
rect 17000 5352 17006 5364
rect 17129 5355 17187 5361
rect 17129 5352 17141 5355
rect 17000 5324 17141 5352
rect 17000 5312 17006 5324
rect 17129 5321 17141 5324
rect 17175 5321 17187 5355
rect 17129 5315 17187 5321
rect 17218 5312 17224 5364
rect 17276 5352 17282 5364
rect 17276 5324 17321 5352
rect 17276 5312 17282 5324
rect 19794 5312 19800 5364
rect 19852 5352 19858 5364
rect 20257 5355 20315 5361
rect 20257 5352 20269 5355
rect 19852 5324 20269 5352
rect 19852 5312 19858 5324
rect 20257 5321 20269 5324
rect 20303 5321 20315 5355
rect 20257 5315 20315 5321
rect 4617 5287 4675 5293
rect 4617 5284 4629 5287
rect 3384 5256 4629 5284
rect 3384 5244 3390 5256
rect 4617 5253 4629 5256
rect 4663 5253 4675 5287
rect 4617 5247 4675 5253
rect 4709 5287 4767 5293
rect 4709 5253 4721 5287
rect 4755 5253 4767 5287
rect 4709 5247 4767 5253
rect 5353 5287 5411 5293
rect 5353 5253 5365 5287
rect 5399 5284 5411 5287
rect 5442 5284 5448 5296
rect 5399 5256 5448 5284
rect 5399 5253 5411 5256
rect 5353 5247 5411 5253
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 8018 5284 8024 5296
rect 6012 5256 8024 5284
rect 3878 5216 3884 5228
rect 3936 5225 3942 5228
rect 3848 5188 3884 5216
rect 3878 5176 3884 5188
rect 3936 5179 3948 5225
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 4338 5216 4344 5228
rect 4203 5188 4344 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 3936 5176 3942 5179
rect 4338 5176 4344 5188
rect 4396 5176 4402 5228
rect 4520 5219 4578 5225
rect 4520 5185 4532 5219
rect 4566 5216 4578 5219
rect 4890 5216 4896 5228
rect 4566 5188 4752 5216
rect 4851 5188 4896 5216
rect 4566 5185 4578 5188
rect 4520 5179 4578 5185
rect 4724 5080 4752 5188
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 6012 5225 6040 5256
rect 8018 5244 8024 5256
rect 8076 5244 8082 5296
rect 8202 5293 8208 5296
rect 8196 5284 8208 5293
rect 8163 5256 8208 5284
rect 8196 5247 8208 5256
rect 8202 5244 8208 5247
rect 8260 5244 8266 5296
rect 9214 5244 9220 5296
rect 9272 5284 9278 5296
rect 9953 5287 10011 5293
rect 9953 5284 9965 5287
rect 9272 5256 9965 5284
rect 9272 5244 9278 5256
rect 9953 5253 9965 5256
rect 9999 5253 10011 5287
rect 9953 5247 10011 5253
rect 10781 5287 10839 5293
rect 10781 5253 10793 5287
rect 10827 5284 10839 5287
rect 10870 5284 10876 5296
rect 10827 5256 10876 5284
rect 10827 5253 10839 5256
rect 10781 5247 10839 5253
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 11606 5244 11612 5296
rect 11664 5284 11670 5296
rect 11762 5287 11820 5293
rect 11762 5284 11774 5287
rect 11664 5256 11774 5284
rect 11664 5244 11670 5256
rect 11762 5253 11774 5256
rect 11808 5253 11820 5287
rect 11762 5247 11820 5253
rect 12618 5244 12624 5296
rect 12676 5284 12682 5296
rect 13265 5287 13323 5293
rect 13265 5284 13277 5287
rect 12676 5256 13277 5284
rect 12676 5244 12682 5256
rect 13265 5253 13277 5256
rect 13311 5253 13323 5287
rect 16482 5284 16488 5296
rect 13265 5247 13323 5253
rect 16040 5256 16488 5284
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5185 6055 5219
rect 6362 5216 6368 5228
rect 6323 5188 6368 5216
rect 5997 5179 6055 5185
rect 4798 5108 4804 5160
rect 4856 5148 4862 5160
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 4856 5120 5457 5148
rect 4856 5108 4862 5120
rect 5445 5117 5457 5120
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5718 5148 5724 5160
rect 5675 5120 5724 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 6012 5080 6040 5179
rect 6362 5176 6368 5188
rect 6420 5176 6426 5228
rect 6638 5225 6644 5228
rect 6632 5179 6644 5225
rect 6696 5216 6702 5228
rect 7926 5216 7932 5228
rect 6696 5188 6732 5216
rect 7887 5188 7932 5216
rect 6638 5176 6644 5179
rect 6696 5176 6702 5188
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 8478 5216 8484 5228
rect 8036 5188 8484 5216
rect 8036 5148 8064 5188
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 10560 5188 11529 5216
rect 10560 5176 10566 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 12986 5216 12992 5228
rect 12899 5188 12992 5216
rect 11517 5179 11575 5185
rect 4724 5052 6040 5080
rect 7760 5120 8064 5148
rect 10137 5151 10195 5157
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 4341 5015 4399 5021
rect 4341 5012 4353 5015
rect 3936 4984 4353 5012
rect 3936 4972 3942 4984
rect 4341 4981 4353 4984
rect 4387 4981 4399 5015
rect 5810 5012 5816 5024
rect 5771 4984 5816 5012
rect 4341 4975 4399 4981
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 6270 5012 6276 5024
rect 6227 4984 6276 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 7760 5021 7788 5120
rect 10137 5117 10149 5151
rect 10183 5148 10195 5151
rect 10183 5120 10456 5148
rect 10183 5117 10195 5120
rect 10137 5111 10195 5117
rect 7745 5015 7803 5021
rect 7745 5012 7757 5015
rect 7524 4984 7757 5012
rect 7524 4972 7530 4984
rect 7745 4981 7757 4984
rect 7791 4981 7803 5015
rect 7745 4975 7803 4981
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 10428 5021 10456 5120
rect 11146 5080 11152 5092
rect 11107 5052 11152 5080
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 9493 5015 9551 5021
rect 9493 5012 9505 5015
rect 7892 4984 9505 5012
rect 7892 4972 7898 4984
rect 9493 4981 9505 4984
rect 9539 4981 9551 5015
rect 9493 4975 9551 4981
rect 10413 5015 10471 5021
rect 10413 4981 10425 5015
rect 10459 5012 10471 5015
rect 10594 5012 10600 5024
rect 10459 4984 10600 5012
rect 10459 4981 10471 4984
rect 10413 4975 10471 4981
rect 10594 4972 10600 4984
rect 10652 5012 10658 5024
rect 12526 5012 12532 5024
rect 10652 4984 12532 5012
rect 10652 4972 10658 4984
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 12802 4972 12808 5024
rect 12860 5012 12866 5024
rect 12912 5021 12940 5188
rect 12986 5176 12992 5188
rect 13044 5216 13050 5228
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 13044 5188 13093 5216
rect 13044 5176 13050 5188
rect 13081 5185 13093 5188
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 16040 5225 16068 5256
rect 16482 5244 16488 5256
rect 16540 5244 16546 5296
rect 17144 5256 17908 5284
rect 17144 5228 17172 5256
rect 16025 5219 16083 5225
rect 15528 5188 15976 5216
rect 15528 5176 15534 5188
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5148 15255 5151
rect 15286 5148 15292 5160
rect 15243 5120 15292 5148
rect 15243 5117 15255 5120
rect 15197 5111 15255 5117
rect 15286 5108 15292 5120
rect 15344 5148 15350 5160
rect 15746 5148 15752 5160
rect 15344 5120 15752 5148
rect 15344 5108 15350 5120
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 15948 5148 15976 5188
rect 16025 5185 16037 5219
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 16209 5219 16267 5225
rect 16209 5185 16221 5219
rect 16255 5216 16267 5219
rect 17126 5216 17132 5228
rect 16255 5188 17132 5216
rect 16255 5185 16267 5188
rect 16209 5179 16267 5185
rect 17126 5176 17132 5188
rect 17184 5176 17190 5228
rect 17236 5188 17356 5216
rect 17236 5148 17264 5188
rect 17328 5157 17356 5188
rect 17402 5176 17408 5228
rect 17460 5216 17466 5228
rect 17880 5225 17908 5256
rect 18414 5244 18420 5296
rect 18472 5284 18478 5296
rect 19122 5287 19180 5293
rect 19122 5284 19134 5287
rect 18472 5256 19134 5284
rect 18472 5244 18478 5256
rect 19122 5253 19134 5256
rect 19168 5253 19180 5287
rect 19122 5247 19180 5253
rect 17589 5219 17647 5225
rect 17589 5216 17601 5219
rect 17460 5188 17601 5216
rect 17460 5176 17466 5188
rect 17589 5185 17601 5188
rect 17635 5185 17647 5219
rect 17589 5179 17647 5185
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 15948 5120 17264 5148
rect 17313 5151 17371 5157
rect 17313 5117 17325 5151
rect 17359 5117 17371 5151
rect 17678 5148 17684 5160
rect 17639 5120 17684 5148
rect 17313 5111 17371 5117
rect 17678 5108 17684 5120
rect 17736 5108 17742 5160
rect 18874 5148 18880 5160
rect 18835 5120 18880 5148
rect 18874 5108 18880 5120
rect 18932 5108 18938 5160
rect 13449 5083 13507 5089
rect 13449 5049 13461 5083
rect 13495 5080 13507 5083
rect 13814 5080 13820 5092
rect 13495 5052 13820 5080
rect 13495 5049 13507 5052
rect 13449 5043 13507 5049
rect 13814 5040 13820 5052
rect 13872 5040 13878 5092
rect 15562 5080 15568 5092
rect 15523 5052 15568 5080
rect 15562 5040 15568 5052
rect 15620 5040 15626 5092
rect 16224 5052 17540 5080
rect 16224 5021 16252 5052
rect 17512 5024 17540 5052
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 12860 4984 12909 5012
rect 12860 4972 12866 4984
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 12897 4975 12955 4981
rect 16209 5015 16267 5021
rect 16209 4981 16221 5015
rect 16255 4981 16267 5015
rect 16758 5012 16764 5024
rect 16719 4984 16764 5012
rect 16209 4975 16267 4981
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 17494 4972 17500 5024
rect 17552 5012 17558 5024
rect 17589 5015 17647 5021
rect 17589 5012 17601 5015
rect 17552 4984 17601 5012
rect 17552 4972 17558 4984
rect 17589 4981 17601 4984
rect 17635 4981 17647 5015
rect 18046 5012 18052 5024
rect 18007 4984 18052 5012
rect 17589 4975 17647 4981
rect 18046 4972 18052 4984
rect 18104 5012 18110 5024
rect 19242 5012 19248 5024
rect 18104 4984 19248 5012
rect 18104 4972 18110 4984
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 1104 4922 26128 4944
rect 1104 4870 5120 4922
rect 5172 4870 5184 4922
rect 5236 4870 5248 4922
rect 5300 4870 5312 4922
rect 5364 4870 5376 4922
rect 5428 4870 13462 4922
rect 13514 4870 13526 4922
rect 13578 4870 13590 4922
rect 13642 4870 13654 4922
rect 13706 4870 13718 4922
rect 13770 4870 21803 4922
rect 21855 4870 21867 4922
rect 21919 4870 21931 4922
rect 21983 4870 21995 4922
rect 22047 4870 22059 4922
rect 22111 4870 26128 4922
rect 1104 4848 26128 4870
rect 4246 4808 4252 4820
rect 3896 4780 4252 4808
rect 3896 4681 3924 4780
rect 4246 4768 4252 4780
rect 4304 4768 4310 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5442 4808 5448 4820
rect 5307 4780 5448 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 5810 4768 5816 4820
rect 5868 4808 5874 4820
rect 6365 4811 6423 4817
rect 6365 4808 6377 4811
rect 5868 4780 6377 4808
rect 5868 4768 5874 4780
rect 6365 4777 6377 4780
rect 6411 4777 6423 4811
rect 6365 4771 6423 4777
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 6825 4811 6883 4817
rect 6825 4808 6837 4811
rect 6696 4780 6837 4808
rect 6696 4768 6702 4780
rect 6825 4777 6837 4780
rect 6871 4777 6883 4811
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 6825 4771 6883 4777
rect 6932 4780 7849 4808
rect 6546 4740 6552 4752
rect 6459 4712 6552 4740
rect 6546 4700 6552 4712
rect 6604 4740 6610 4752
rect 6932 4740 6960 4780
rect 7837 4777 7849 4780
rect 7883 4808 7895 4811
rect 8386 4808 8392 4820
rect 7883 4780 8392 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 8662 4768 8668 4820
rect 8720 4808 8726 4820
rect 8757 4811 8815 4817
rect 8757 4808 8769 4811
rect 8720 4780 8769 4808
rect 8720 4768 8726 4780
rect 8757 4777 8769 4780
rect 8803 4777 8815 4811
rect 10594 4808 10600 4820
rect 10555 4780 10600 4808
rect 8757 4771 8815 4777
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 13998 4768 14004 4820
rect 14056 4808 14062 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 14056 4780 14105 4808
rect 14056 4768 14062 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14093 4771 14151 4777
rect 17218 4768 17224 4820
rect 17276 4808 17282 4820
rect 17589 4811 17647 4817
rect 17589 4808 17601 4811
rect 17276 4780 17601 4808
rect 17276 4768 17282 4780
rect 17589 4777 17601 4780
rect 17635 4777 17647 4811
rect 17589 4771 17647 4777
rect 6604 4712 6960 4740
rect 6604 4700 6610 4712
rect 7650 4700 7656 4752
rect 7708 4700 7714 4752
rect 9033 4743 9091 4749
rect 9033 4740 9045 4743
rect 8036 4712 9045 4740
rect 3881 4675 3939 4681
rect 3881 4641 3893 4675
rect 3927 4641 3939 4675
rect 5902 4672 5908 4684
rect 5863 4644 5908 4672
rect 3881 4635 3939 4641
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 6089 4675 6147 4681
rect 6089 4641 6101 4675
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 2038 4604 2044 4616
rect 1999 4576 2044 4604
rect 2038 4564 2044 4576
rect 2096 4564 2102 4616
rect 6104 4604 6132 4635
rect 6270 4604 6276 4616
rect 6104 4576 6276 4604
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6564 4613 6592 4700
rect 7466 4672 7472 4684
rect 6656 4644 7472 4672
rect 6656 4613 6684 4644
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 7668 4672 7696 4700
rect 7576 4644 7696 4672
rect 7929 4675 7987 4681
rect 7576 4613 7604 4644
rect 7929 4641 7941 4675
rect 7975 4672 7987 4675
rect 8036 4672 8064 4712
rect 9033 4709 9045 4712
rect 9079 4740 9091 4743
rect 9214 4740 9220 4752
rect 9079 4712 9220 4740
rect 9079 4709 9091 4712
rect 9033 4703 9091 4709
rect 9214 4700 9220 4712
rect 9272 4700 9278 4752
rect 11057 4743 11115 4749
rect 11057 4709 11069 4743
rect 11103 4740 11115 4743
rect 11333 4743 11391 4749
rect 11333 4740 11345 4743
rect 11103 4712 11345 4740
rect 11103 4709 11115 4712
rect 11057 4703 11115 4709
rect 11333 4709 11345 4712
rect 11379 4709 11391 4743
rect 15470 4740 15476 4752
rect 11333 4703 11391 4709
rect 13556 4712 15476 4740
rect 8202 4672 8208 4684
rect 7975 4644 8064 4672
rect 8163 4644 8208 4672
rect 7975 4641 7987 4644
rect 7929 4635 7987 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4672 8355 4675
rect 8570 4672 8576 4684
rect 8343 4644 8576 4672
rect 8343 4641 8355 4644
rect 8297 4635 8355 4641
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4672 10747 4675
rect 10870 4672 10876 4684
rect 10735 4644 10876 4672
rect 10735 4641 10747 4644
rect 10689 4635 10747 4641
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 11977 4675 12035 4681
rect 11977 4641 11989 4675
rect 12023 4672 12035 4675
rect 12250 4672 12256 4684
rect 12023 4644 12256 4672
rect 12023 4641 12035 4644
rect 11977 4635 12035 4641
rect 12250 4632 12256 4644
rect 12308 4672 12314 4684
rect 13556 4681 13584 4712
rect 12713 4675 12771 4681
rect 12713 4672 12725 4675
rect 12308 4644 12725 4672
rect 12308 4632 12314 4644
rect 12713 4641 12725 4644
rect 12759 4672 12771 4675
rect 13541 4675 13599 4681
rect 13541 4672 13553 4675
rect 12759 4644 13553 4672
rect 12759 4641 12771 4644
rect 12713 4635 12771 4641
rect 13541 4641 13553 4644
rect 13587 4641 13599 4675
rect 15102 4672 15108 4684
rect 13541 4635 13599 4641
rect 14108 4644 15108 4672
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 7561 4607 7619 4613
rect 7055 4576 7236 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 4148 4539 4206 4545
rect 4148 4505 4160 4539
rect 4194 4536 4206 4539
rect 4798 4536 4804 4548
rect 4194 4508 4804 4536
rect 4194 4505 4206 4508
rect 4148 4499 4206 4505
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 4982 4428 4988 4480
rect 5040 4468 5046 4480
rect 5445 4471 5503 4477
rect 5445 4468 5457 4471
rect 5040 4440 5457 4468
rect 5040 4428 5046 4440
rect 5445 4437 5457 4440
rect 5491 4437 5503 4471
rect 5445 4431 5503 4437
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 5813 4471 5871 4477
rect 5813 4468 5825 4471
rect 5776 4440 5825 4468
rect 5776 4428 5782 4440
rect 5813 4437 5825 4440
rect 5859 4437 5871 4471
rect 7098 4468 7104 4480
rect 7059 4440 7104 4468
rect 5813 4431 5871 4437
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 7208 4468 7236 4576
rect 7561 4573 7573 4607
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 7742 4604 7748 4616
rect 7699 4576 7748 4604
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 7742 4564 7748 4576
rect 7800 4604 7806 4616
rect 8110 4604 8116 4616
rect 7800 4576 8116 4604
rect 7800 4564 7806 4576
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 8478 4604 8484 4616
rect 8435 4576 8484 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4604 10471 4607
rect 10502 4604 10508 4616
rect 10459 4576 10508 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 11514 4564 11520 4616
rect 11572 4604 11578 4616
rect 11701 4607 11759 4613
rect 11701 4604 11713 4607
rect 11572 4576 11713 4604
rect 11572 4564 11578 4576
rect 11701 4573 11713 4576
rect 11747 4604 11759 4607
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 11747 4576 12541 4604
rect 11747 4573 11759 4576
rect 11701 4567 11759 4573
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 12529 4567 12587 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13814 4564 13820 4616
rect 13872 4604 13878 4616
rect 14108 4613 14136 4644
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 15396 4681 15424 4712
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 16117 4743 16175 4749
rect 16117 4709 16129 4743
rect 16163 4740 16175 4743
rect 16758 4740 16764 4752
rect 16163 4712 16764 4740
rect 16163 4709 16175 4712
rect 16117 4703 16175 4709
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 16945 4743 17003 4749
rect 16945 4709 16957 4743
rect 16991 4740 17003 4743
rect 17678 4740 17684 4752
rect 16991 4712 17684 4740
rect 16991 4709 17003 4712
rect 16945 4703 17003 4709
rect 17678 4700 17684 4712
rect 17736 4700 17742 4752
rect 15381 4675 15439 4681
rect 15381 4641 15393 4675
rect 15427 4641 15439 4675
rect 15381 4635 15439 4641
rect 16574 4632 16580 4684
rect 16632 4672 16638 4684
rect 17037 4675 17095 4681
rect 17037 4672 17049 4675
rect 16632 4644 17049 4672
rect 16632 4632 16638 4644
rect 17037 4641 17049 4644
rect 17083 4641 17095 4675
rect 17037 4635 17095 4641
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13872 4576 14105 4604
rect 13872 4564 13878 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14093 4567 14151 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 15194 4604 15200 4616
rect 15155 4576 15200 4604
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4573 17187 4607
rect 17129 4567 17187 4573
rect 17496 4607 17554 4613
rect 17496 4573 17508 4607
rect 17542 4604 17554 4607
rect 18046 4604 18052 4616
rect 17542 4576 18052 4604
rect 17542 4573 17554 4576
rect 17496 4567 17554 4573
rect 7377 4539 7435 4545
rect 7377 4505 7389 4539
rect 7423 4536 7435 4539
rect 10146 4539 10204 4545
rect 10146 4536 10158 4539
rect 7423 4508 10158 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 10146 4505 10158 4508
rect 10192 4505 10204 4539
rect 10146 4499 10204 4505
rect 12621 4539 12679 4545
rect 12621 4505 12633 4539
rect 12667 4536 12679 4539
rect 14366 4536 14372 4548
rect 12667 4508 14372 4536
rect 12667 4505 12679 4508
rect 12621 4499 12679 4505
rect 14366 4496 14372 4508
rect 14424 4496 14430 4548
rect 15746 4536 15752 4548
rect 15707 4508 15752 4536
rect 15746 4496 15752 4508
rect 15804 4496 15810 4548
rect 16574 4536 16580 4548
rect 16535 4508 16580 4536
rect 16574 4496 16580 4508
rect 16632 4496 16638 4548
rect 16758 4536 16764 4548
rect 16719 4508 16764 4536
rect 16758 4496 16764 4508
rect 16816 4536 16822 4548
rect 17144 4536 17172 4567
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 16816 4508 17172 4536
rect 16816 4496 16822 4508
rect 8018 4468 8024 4480
rect 7208 4440 8024 4468
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 11149 4471 11207 4477
rect 11149 4437 11161 4471
rect 11195 4468 11207 4471
rect 11514 4468 11520 4480
rect 11195 4440 11520 4468
rect 11195 4437 11207 4440
rect 11149 4431 11207 4437
rect 11514 4428 11520 4440
rect 11572 4428 11578 4480
rect 11793 4471 11851 4477
rect 11793 4437 11805 4471
rect 11839 4468 11851 4471
rect 12066 4468 12072 4480
rect 11839 4440 12072 4468
rect 11839 4437 11851 4440
rect 11793 4431 11851 4437
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 12158 4428 12164 4480
rect 12216 4468 12222 4480
rect 12216 4440 12261 4468
rect 12216 4428 12222 4440
rect 12710 4428 12716 4480
rect 12768 4468 12774 4480
rect 12989 4471 13047 4477
rect 12989 4468 13001 4471
rect 12768 4440 13001 4468
rect 12768 4428 12774 4440
rect 12989 4437 13001 4440
rect 13035 4437 13047 4471
rect 12989 4431 13047 4437
rect 13449 4471 13507 4477
rect 13449 4437 13461 4471
rect 13495 4468 13507 4471
rect 14090 4468 14096 4480
rect 13495 4440 14096 4468
rect 13495 4437 13507 4440
rect 13449 4431 13507 4437
rect 14090 4428 14096 4440
rect 14148 4428 14154 4480
rect 14458 4468 14464 4480
rect 14419 4440 14464 4468
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 14829 4471 14887 4477
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 14918 4468 14924 4480
rect 14875 4440 14924 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15286 4428 15292 4480
rect 15344 4468 15350 4480
rect 16209 4471 16267 4477
rect 15344 4440 15389 4468
rect 15344 4428 15350 4440
rect 16209 4437 16221 4471
rect 16255 4468 16267 4471
rect 17126 4468 17132 4480
rect 16255 4440 17132 4468
rect 16255 4437 16267 4440
rect 16209 4431 16267 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 1104 4378 26128 4400
rect 1104 4326 9291 4378
rect 9343 4326 9355 4378
rect 9407 4326 9419 4378
rect 9471 4326 9483 4378
rect 9535 4326 9547 4378
rect 9599 4326 17632 4378
rect 17684 4326 17696 4378
rect 17748 4326 17760 4378
rect 17812 4326 17824 4378
rect 17876 4326 17888 4378
rect 17940 4326 26128 4378
rect 1104 4304 26128 4326
rect 4798 4264 4804 4276
rect 4759 4236 4804 4264
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 5810 4224 5816 4276
rect 5868 4224 5874 4276
rect 5905 4267 5963 4273
rect 5905 4233 5917 4267
rect 5951 4264 5963 4267
rect 5994 4264 6000 4276
rect 5951 4236 6000 4264
rect 5951 4233 5963 4236
rect 5905 4227 5963 4233
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 7742 4264 7748 4276
rect 7703 4236 7748 4264
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 9214 4264 9220 4276
rect 9175 4236 9220 4264
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 9769 4267 9827 4273
rect 9769 4264 9781 4267
rect 9646 4236 9781 4264
rect 5828 4196 5856 4224
rect 5276 4168 5856 4196
rect 6733 4199 6791 4205
rect 4982 4128 4988 4140
rect 4943 4100 4988 4128
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5276 4128 5304 4168
rect 6733 4165 6745 4199
rect 6779 4196 6791 4199
rect 7466 4196 7472 4208
rect 6779 4168 7472 4196
rect 6779 4165 6791 4168
rect 6733 4159 6791 4165
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 8202 4196 8208 4208
rect 8115 4168 8208 4196
rect 8202 4156 8208 4168
rect 8260 4196 8266 4208
rect 8260 4168 8708 4196
rect 8260 4156 8266 4168
rect 5123 4100 5304 4128
rect 5353 4131 5411 4137
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5353 4097 5365 4131
rect 5399 4128 5411 4131
rect 5442 4128 5448 4140
rect 5399 4100 5448 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6086 4128 6092 4140
rect 5859 4100 6092 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 6328 4100 7052 4128
rect 6328 4088 6334 4100
rect 5261 4063 5319 4069
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 5534 4060 5540 4072
rect 5307 4032 5540 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4060 6055 4063
rect 6288 4060 6316 4088
rect 6043 4032 6316 4060
rect 6043 4029 6055 4032
rect 5997 4023 6055 4029
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 7024 4069 7052 4100
rect 7098 4088 7104 4140
rect 7156 4128 7162 4140
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 7156 4100 7205 4128
rect 7156 4088 7162 4100
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 7929 4131 7987 4137
rect 7929 4097 7941 4131
rect 7975 4128 7987 4131
rect 8018 4128 8024 4140
rect 7975 4100 8024 4128
rect 7975 4097 7987 4100
rect 7929 4091 7987 4097
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6788 4032 6837 4060
rect 6788 4020 6794 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 7055 4032 7573 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 7561 4029 7573 4032
rect 7607 4060 7619 4063
rect 7650 4060 7656 4072
rect 7607 4032 7656 4060
rect 7607 4029 7619 4032
rect 7561 4023 7619 4029
rect 7650 4020 7656 4032
rect 7708 4060 7714 4072
rect 8220 4060 8248 4156
rect 8386 4128 8392 4140
rect 8347 4100 8392 4128
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 7708 4032 8248 4060
rect 7708 4020 7714 4032
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 8680 4069 8708 4168
rect 9030 4088 9036 4140
rect 9088 4128 9094 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9088 4100 9321 4128
rect 9088 4088 9094 4100
rect 9309 4097 9321 4100
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8352 4032 8493 4060
rect 8352 4020 8358 4032
rect 8481 4029 8493 4032
rect 8527 4029 8539 4063
rect 8481 4023 8539 4029
rect 8665 4063 8723 4069
rect 8665 4029 8677 4063
rect 8711 4060 8723 4063
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 8711 4032 9505 4060
rect 8711 4029 8723 4032
rect 8665 4023 8723 4029
rect 9493 4029 9505 4032
rect 9539 4060 9551 4063
rect 9646 4060 9674 4236
rect 9769 4233 9781 4236
rect 9815 4264 9827 4267
rect 9953 4267 10011 4273
rect 9953 4264 9965 4267
rect 9815 4236 9965 4264
rect 9815 4233 9827 4236
rect 9769 4227 9827 4233
rect 9953 4233 9965 4236
rect 9999 4264 10011 4267
rect 10594 4264 10600 4276
rect 9999 4236 10600 4264
rect 9999 4233 10011 4236
rect 9953 4227 10011 4233
rect 10594 4224 10600 4236
rect 10652 4224 10658 4276
rect 14274 4264 14280 4276
rect 14235 4236 14280 4264
rect 14274 4224 14280 4236
rect 14332 4224 14338 4276
rect 10689 4199 10747 4205
rect 10689 4165 10701 4199
rect 10735 4196 10747 4199
rect 10781 4199 10839 4205
rect 10781 4196 10793 4199
rect 10735 4168 10793 4196
rect 10735 4165 10747 4168
rect 10689 4159 10747 4165
rect 10781 4165 10793 4168
rect 10827 4196 10839 4199
rect 10870 4196 10876 4208
rect 10827 4168 10876 4196
rect 10827 4165 10839 4168
rect 10781 4159 10839 4165
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 12066 4196 12072 4208
rect 12027 4168 12072 4196
rect 12066 4156 12072 4168
rect 12124 4156 12130 4208
rect 13814 4196 13820 4208
rect 12406 4168 13820 4196
rect 11514 4128 11520 4140
rect 11475 4100 11520 4128
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 12311 4131 12369 4137
rect 12311 4097 12323 4131
rect 12357 4128 12369 4131
rect 12406 4128 12434 4168
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 13998 4156 14004 4208
rect 14056 4196 14062 4208
rect 14056 4168 15056 4196
rect 14056 4156 14062 4168
rect 12618 4128 12624 4140
rect 12357 4100 12434 4128
rect 12579 4100 12624 4128
rect 12357 4097 12369 4100
rect 12311 4091 12369 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4128 12771 4131
rect 12802 4128 12808 4140
rect 12759 4100 12808 4128
rect 12759 4097 12771 4100
rect 12713 4091 12771 4097
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 13170 4137 13176 4140
rect 13164 4091 13176 4137
rect 13228 4128 13234 4140
rect 13228 4100 13264 4128
rect 13170 4088 13176 4091
rect 13228 4088 13234 4100
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 15028 4137 15056 4168
rect 15102 4156 15108 4208
rect 15160 4196 15166 4208
rect 15197 4199 15255 4205
rect 15197 4196 15209 4199
rect 15160 4168 15209 4196
rect 15160 4156 15166 4168
rect 15197 4165 15209 4168
rect 15243 4165 15255 4199
rect 15197 4159 15255 4165
rect 15286 4156 15292 4208
rect 15344 4196 15350 4208
rect 15749 4199 15807 4205
rect 15749 4196 15761 4199
rect 15344 4168 15761 4196
rect 15344 4156 15350 4168
rect 15749 4165 15761 4168
rect 15795 4165 15807 4199
rect 16482 4196 16488 4208
rect 15749 4159 15807 4165
rect 16224 4168 16488 4196
rect 14461 4131 14519 4137
rect 14461 4128 14473 4131
rect 14424 4100 14473 4128
rect 14424 4088 14430 4100
rect 14461 4097 14473 4100
rect 14507 4097 14519 4131
rect 14461 4091 14519 4097
rect 14703 4131 14761 4137
rect 14703 4097 14715 4131
rect 14749 4097 14761 4131
rect 14703 4091 14761 4097
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4128 15071 4131
rect 15381 4131 15439 4137
rect 15381 4128 15393 4131
rect 15059 4100 15393 4128
rect 15059 4097 15071 4100
rect 15013 4091 15071 4097
rect 15381 4097 15393 4100
rect 15427 4097 15439 4131
rect 15381 4091 15439 4097
rect 15991 4131 16049 4137
rect 15991 4097 16003 4131
rect 16037 4128 16049 4131
rect 16224 4128 16252 4168
rect 16482 4156 16488 4168
rect 16540 4156 16546 4208
rect 16853 4199 16911 4205
rect 16853 4196 16865 4199
rect 16592 4168 16865 4196
rect 16592 4140 16620 4168
rect 16853 4165 16865 4168
rect 16899 4165 16911 4199
rect 17402 4196 17408 4208
rect 16853 4159 16911 4165
rect 16960 4168 17408 4196
rect 16037 4100 16252 4128
rect 16301 4131 16359 4137
rect 16037 4097 16049 4100
rect 15991 4091 16049 4097
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 16574 4128 16580 4140
rect 16347 4100 16580 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 12158 4060 12164 4072
rect 9539 4032 9674 4060
rect 11072 4032 12164 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 5552 3992 5580 4020
rect 7098 3992 7104 4004
rect 5552 3964 7104 3992
rect 7098 3952 7104 3964
rect 7156 3952 7162 4004
rect 7377 3995 7435 4001
rect 7377 3961 7389 3995
rect 7423 3992 7435 3995
rect 8202 3992 8208 4004
rect 7423 3964 8208 3992
rect 7423 3961 7435 3964
rect 7377 3955 7435 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 10413 3995 10471 4001
rect 10413 3961 10425 3995
rect 10459 3992 10471 3995
rect 11072 3992 11100 4032
rect 12158 4020 12164 4032
rect 12216 4020 12222 4072
rect 12897 4063 12955 4069
rect 12897 4029 12909 4063
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 10459 3964 11100 3992
rect 11149 3995 11207 4001
rect 10459 3961 10471 3964
rect 10413 3955 10471 3961
rect 11149 3961 11161 3995
rect 11195 3992 11207 3995
rect 11195 3964 11928 3992
rect 11195 3961 11207 3964
rect 11149 3955 11207 3961
rect 5442 3924 5448 3936
rect 5403 3896 5448 3924
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 5868 3896 6377 3924
rect 5868 3884 5874 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8294 3924 8300 3936
rect 8067 3896 8300 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8478 3884 8484 3936
rect 8536 3924 8542 3936
rect 8849 3927 8907 3933
rect 8849 3924 8861 3927
rect 8536 3896 8861 3924
rect 8536 3884 8542 3896
rect 8849 3893 8861 3896
rect 8895 3893 8907 3927
rect 8849 3887 8907 3893
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3924 10287 3927
rect 11054 3924 11060 3936
rect 10275 3896 11060 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11238 3924 11244 3936
rect 11199 3896 11244 3924
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 11701 3927 11759 3933
rect 11701 3893 11713 3927
rect 11747 3924 11759 3927
rect 11790 3924 11796 3936
rect 11747 3896 11796 3924
rect 11747 3893 11759 3896
rect 11701 3887 11759 3893
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 11900 3924 11928 3964
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 12912 3992 12940 4023
rect 14718 4004 14746 4091
rect 16574 4088 16580 4100
rect 16632 4088 16638 4140
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4128 16727 4131
rect 16960 4128 16988 4168
rect 17402 4156 17408 4168
rect 17460 4156 17466 4208
rect 22738 4196 22744 4208
rect 22020 4168 22744 4196
rect 17126 4128 17132 4140
rect 16715 4100 16988 4128
rect 17087 4100 17132 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 15102 4060 15108 4072
rect 15063 4032 15108 4060
rect 15102 4020 15108 4032
rect 15160 4020 15166 4072
rect 16393 4063 16451 4069
rect 16393 4029 16405 4063
rect 16439 4029 16451 4063
rect 16393 4023 16451 4029
rect 14718 3992 14740 4004
rect 12400 3964 12940 3992
rect 14647 3964 14740 3992
rect 12400 3952 12406 3964
rect 14734 3952 14740 3964
rect 14792 3992 14798 4004
rect 15565 3995 15623 4001
rect 15565 3992 15577 3995
rect 14792 3964 15577 3992
rect 14792 3952 14798 3964
rect 15565 3961 15577 3964
rect 15611 3961 15623 3995
rect 15565 3955 15623 3961
rect 16408 3992 16436 4023
rect 16684 3992 16712 4091
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 22020 4137 22048 4168
rect 22738 4156 22744 4168
rect 22796 4156 22802 4208
rect 22278 4137 22284 4140
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 22272 4091 22284 4137
rect 22336 4128 22342 4140
rect 22336 4100 22372 4128
rect 22278 4088 22284 4091
rect 22336 4088 22342 4100
rect 16408 3964 16712 3992
rect 12710 3924 12716 3936
rect 11900 3896 12716 3924
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 14458 3884 14464 3936
rect 14516 3924 14522 3936
rect 16408 3924 16436 3964
rect 17126 3952 17132 4004
rect 17184 3992 17190 4004
rect 18230 3992 18236 4004
rect 17184 3964 18236 3992
rect 17184 3952 17190 3964
rect 18230 3952 18236 3964
rect 18288 3952 18294 4004
rect 23106 3952 23112 4004
rect 23164 3992 23170 4004
rect 23385 3995 23443 4001
rect 23385 3992 23397 3995
rect 23164 3964 23397 3992
rect 23164 3952 23170 3964
rect 23385 3961 23397 3964
rect 23431 3961 23443 3995
rect 23385 3955 23443 3961
rect 14516 3896 16436 3924
rect 14516 3884 14522 3896
rect 16482 3884 16488 3936
rect 16540 3924 16546 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 16540 3896 16957 3924
rect 16540 3884 16546 3896
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 17310 3924 17316 3936
rect 17271 3896 17316 3924
rect 16945 3887 17003 3893
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 1104 3834 26128 3856
rect 1104 3782 5120 3834
rect 5172 3782 5184 3834
rect 5236 3782 5248 3834
rect 5300 3782 5312 3834
rect 5364 3782 5376 3834
rect 5428 3782 13462 3834
rect 13514 3782 13526 3834
rect 13578 3782 13590 3834
rect 13642 3782 13654 3834
rect 13706 3782 13718 3834
rect 13770 3782 21803 3834
rect 21855 3782 21867 3834
rect 21919 3782 21931 3834
rect 21983 3782 21995 3834
rect 22047 3782 22059 3834
rect 22111 3782 26128 3834
rect 1104 3760 26128 3782
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 5626 3720 5632 3732
rect 4120 3692 5632 3720
rect 4120 3680 4126 3692
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 5813 3723 5871 3729
rect 5813 3720 5825 3723
rect 5776 3692 5825 3720
rect 5776 3680 5782 3692
rect 5813 3689 5825 3692
rect 5859 3689 5871 3723
rect 7650 3720 7656 3732
rect 7611 3692 7656 3720
rect 5813 3683 5871 3689
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 10042 3720 10048 3732
rect 8904 3692 10048 3720
rect 8904 3680 8910 3692
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 11885 3723 11943 3729
rect 11885 3720 11897 3723
rect 10428 3692 11897 3720
rect 2133 3655 2191 3661
rect 2133 3621 2145 3655
rect 2179 3652 2191 3655
rect 2774 3652 2780 3664
rect 2179 3624 2780 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 2774 3612 2780 3624
rect 2832 3612 2838 3664
rect 8386 3652 8392 3664
rect 8128 3624 8392 3652
rect 4338 3544 4344 3596
rect 4396 3584 4402 3596
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 4396 3556 4445 3584
rect 4396 3544 4402 3556
rect 4433 3553 4445 3556
rect 4479 3553 4491 3587
rect 4433 3547 4491 3553
rect 7469 3587 7527 3593
rect 7469 3553 7481 3587
rect 7515 3584 7527 3587
rect 7926 3584 7932 3596
rect 7515 3556 7932 3584
rect 7515 3553 7527 3556
rect 7469 3547 7527 3553
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 8128 3593 8156 3624
rect 8386 3612 8392 3624
rect 8444 3652 8450 3664
rect 9033 3655 9091 3661
rect 9033 3652 9045 3655
rect 8444 3624 9045 3652
rect 8444 3612 8450 3624
rect 9033 3621 9045 3624
rect 9079 3621 9091 3655
rect 9033 3615 9091 3621
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 8202 3544 8208 3596
rect 8260 3584 8266 3596
rect 10428 3584 10456 3692
rect 11885 3689 11897 3692
rect 11931 3720 11943 3723
rect 13262 3720 13268 3732
rect 11931 3692 13268 3720
rect 11931 3689 11943 3692
rect 11885 3683 11943 3689
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 13725 3723 13783 3729
rect 13725 3689 13737 3723
rect 13771 3720 13783 3723
rect 13998 3720 14004 3732
rect 13771 3692 14004 3720
rect 13771 3689 13783 3692
rect 13725 3683 13783 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 15010 3720 15016 3732
rect 14608 3692 15016 3720
rect 14608 3680 14614 3692
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 15838 3720 15844 3732
rect 15120 3692 15844 3720
rect 14090 3652 14096 3664
rect 14051 3624 14096 3652
rect 14090 3612 14096 3624
rect 14148 3612 14154 3664
rect 15120 3593 15148 3692
rect 15838 3680 15844 3692
rect 15896 3720 15902 3732
rect 18874 3720 18880 3732
rect 15896 3692 18880 3720
rect 15896 3680 15902 3692
rect 16485 3655 16543 3661
rect 16485 3621 16497 3655
rect 16531 3652 16543 3655
rect 16574 3652 16580 3664
rect 16531 3624 16580 3652
rect 16531 3621 16543 3624
rect 16485 3615 16543 3621
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 16758 3652 16764 3664
rect 16719 3624 16764 3652
rect 16758 3612 16764 3624
rect 16816 3612 16822 3664
rect 18156 3593 18184 3692
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 22278 3720 22284 3732
rect 22239 3692 22284 3720
rect 22278 3680 22284 3692
rect 22336 3680 22342 3732
rect 15105 3587 15163 3593
rect 15105 3584 15117 3587
rect 8260 3556 8305 3584
rect 10336 3556 10456 3584
rect 14200 3556 15117 3584
rect 8260 3544 8266 3556
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3516 2375 3519
rect 2501 3519 2559 3525
rect 2501 3516 2513 3519
rect 2363 3488 2513 3516
rect 2363 3485 2375 3488
rect 2317 3479 2375 3485
rect 2501 3485 2513 3488
rect 2547 3516 2559 3519
rect 2547 3488 7604 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 3786 3448 3792 3460
rect 1728 3420 3792 3448
rect 1728 3408 1734 3420
rect 3786 3408 3792 3420
rect 3844 3408 3850 3460
rect 4700 3451 4758 3457
rect 4700 3417 4712 3451
rect 4746 3448 4758 3451
rect 4798 3448 4804 3460
rect 4746 3420 4804 3448
rect 4746 3417 4758 3420
rect 4700 3411 4758 3417
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 5994 3408 6000 3460
rect 6052 3448 6058 3460
rect 7202 3451 7260 3457
rect 7202 3448 7214 3451
rect 6052 3420 7214 3448
rect 6052 3408 6058 3420
rect 7202 3417 7214 3420
rect 7248 3417 7260 3451
rect 7576 3448 7604 3488
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 7800 3488 8401 3516
rect 7800 3476 7806 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8536 3488 8581 3516
rect 8536 3476 8542 3488
rect 8665 3451 8723 3457
rect 7576 3420 8064 3448
rect 7202 3411 7260 3417
rect 6086 3380 6092 3392
rect 6047 3352 6092 3380
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 8036 3380 8064 3420
rect 8665 3417 8677 3451
rect 8711 3448 8723 3451
rect 10146 3451 10204 3457
rect 10146 3448 10158 3451
rect 8711 3420 10158 3448
rect 8711 3417 8723 3420
rect 8665 3411 8723 3417
rect 10146 3417 10158 3420
rect 10192 3417 10204 3451
rect 10146 3411 10204 3417
rect 10336 3380 10364 3556
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3516 10471 3519
rect 10502 3516 10508 3528
rect 10459 3488 10508 3516
rect 10459 3485 10471 3488
rect 10413 3479 10471 3485
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 10778 3525 10784 3528
rect 10772 3479 10784 3525
rect 10836 3516 10842 3528
rect 10836 3488 10872 3516
rect 10778 3476 10784 3479
rect 10836 3476 10842 3488
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 11112 3488 12081 3516
rect 11112 3476 11118 3488
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 12342 3516 12348 3528
rect 12255 3488 12348 3516
rect 12069 3479 12127 3485
rect 12342 3476 12348 3488
rect 12400 3516 12406 3528
rect 14200 3516 14228 3556
rect 15105 3553 15117 3556
rect 15151 3553 15163 3587
rect 15105 3547 15163 3553
rect 18141 3587 18199 3593
rect 18141 3553 18153 3587
rect 18187 3553 18199 3587
rect 18141 3547 18199 3553
rect 12400 3488 14228 3516
rect 14335 3519 14393 3525
rect 12400 3476 12406 3488
rect 14335 3485 14347 3519
rect 14381 3516 14393 3519
rect 14458 3516 14464 3528
rect 14381 3488 14464 3516
rect 14381 3485 14393 3488
rect 14335 3479 14393 3485
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14625 3519 14683 3525
rect 14625 3516 14637 3519
rect 14567 3488 14637 3516
rect 12590 3451 12648 3457
rect 12590 3448 12602 3451
rect 12268 3420 12602 3448
rect 12268 3389 12296 3420
rect 12590 3417 12602 3420
rect 12636 3417 12648 3451
rect 14567 3448 14595 3488
rect 14625 3485 14637 3488
rect 14671 3485 14683 3519
rect 14625 3479 14683 3485
rect 14730 3519 14788 3525
rect 14730 3485 14742 3519
rect 14776 3485 14788 3519
rect 14730 3479 14788 3485
rect 12590 3411 12648 3417
rect 14292 3420 14595 3448
rect 14292 3392 14320 3420
rect 14757 3392 14785 3479
rect 14826 3476 14832 3528
rect 14884 3516 14890 3528
rect 14884 3488 14929 3516
rect 14884 3476 14890 3488
rect 17310 3476 17316 3528
rect 17368 3516 17374 3528
rect 17874 3519 17932 3525
rect 17874 3516 17886 3519
rect 17368 3488 17886 3516
rect 17368 3476 17374 3488
rect 17874 3485 17886 3488
rect 17920 3485 17932 3519
rect 17874 3479 17932 3485
rect 21821 3519 21879 3525
rect 21821 3485 21833 3519
rect 21867 3516 21879 3519
rect 22465 3519 22523 3525
rect 22465 3516 22477 3519
rect 21867 3488 22477 3516
rect 21867 3485 21879 3488
rect 21821 3479 21879 3485
rect 22465 3485 22477 3488
rect 22511 3485 22523 3519
rect 23106 3516 23112 3528
rect 23067 3488 23112 3516
rect 22465 3479 22523 3485
rect 23106 3476 23112 3488
rect 23164 3476 23170 3528
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 24360 3488 24409 3516
rect 24360 3476 24366 3488
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 25041 3519 25099 3525
rect 25041 3485 25053 3519
rect 25087 3516 25099 3519
rect 25498 3516 25504 3528
rect 25087 3488 25504 3516
rect 25087 3485 25099 3488
rect 25041 3479 25099 3485
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 15350 3451 15408 3457
rect 15350 3448 15362 3451
rect 15212 3420 15362 3448
rect 8036 3352 10364 3380
rect 12253 3383 12311 3389
rect 12253 3349 12265 3383
rect 12299 3349 12311 3383
rect 12253 3343 12311 3349
rect 14274 3340 14280 3392
rect 14332 3340 14338 3392
rect 14734 3340 14740 3392
rect 14792 3340 14798 3392
rect 15013 3383 15071 3389
rect 15013 3349 15025 3383
rect 15059 3380 15071 3383
rect 15212 3380 15240 3420
rect 15350 3417 15362 3420
rect 15396 3417 15408 3451
rect 15350 3411 15408 3417
rect 16114 3408 16120 3460
rect 16172 3448 16178 3460
rect 21726 3448 21732 3460
rect 16172 3420 21732 3448
rect 16172 3408 16178 3420
rect 21726 3408 21732 3420
rect 21784 3408 21790 3460
rect 22005 3451 22063 3457
rect 22005 3417 22017 3451
rect 22051 3417 22063 3451
rect 22005 3411 22063 3417
rect 22189 3451 22247 3457
rect 22189 3417 22201 3451
rect 22235 3417 22247 3451
rect 22189 3411 22247 3417
rect 21634 3380 21640 3392
rect 15059 3352 15240 3380
rect 21547 3352 21640 3380
rect 15059 3349 15071 3352
rect 15013 3343 15071 3349
rect 21634 3340 21640 3352
rect 21692 3380 21698 3392
rect 22020 3380 22048 3411
rect 21692 3352 22048 3380
rect 22204 3380 22232 3411
rect 22646 3380 22652 3392
rect 22204 3352 22652 3380
rect 21692 3340 21698 3352
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 1104 3290 26128 3312
rect 1104 3238 9291 3290
rect 9343 3238 9355 3290
rect 9407 3238 9419 3290
rect 9471 3238 9483 3290
rect 9535 3238 9547 3290
rect 9599 3238 17632 3290
rect 17684 3238 17696 3290
rect 17748 3238 17760 3290
rect 17812 3238 17824 3290
rect 17876 3238 17888 3290
rect 17940 3238 26128 3290
rect 1104 3216 26128 3238
rect 4798 3176 4804 3188
rect 4759 3148 4804 3176
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 5994 3176 6000 3188
rect 5955 3148 6000 3176
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6270 3136 6276 3188
rect 6328 3176 6334 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 6328 3148 6377 3176
rect 6328 3136 6334 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 7466 3176 7472 3188
rect 7427 3148 7472 3176
rect 6365 3139 6423 3145
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12434 3176 12440 3188
rect 12032 3148 12440 3176
rect 12032 3136 12038 3148
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 12897 3179 12955 3185
rect 12897 3176 12909 3179
rect 12676 3148 12909 3176
rect 12676 3136 12682 3148
rect 12897 3145 12909 3148
rect 12943 3145 12955 3179
rect 12897 3139 12955 3145
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 13265 3179 13323 3185
rect 13265 3176 13277 3179
rect 13228 3148 13277 3176
rect 13228 3136 13234 3148
rect 13265 3145 13277 3148
rect 13311 3145 13323 3179
rect 14826 3176 14832 3188
rect 14787 3148 14832 3176
rect 13265 3139 13323 3145
rect 14826 3136 14832 3148
rect 14884 3136 14890 3188
rect 22370 3176 22376 3188
rect 14936 3148 22376 3176
rect 5442 3108 5448 3120
rect 5000 3080 5448 3108
rect 5000 3049 5028 3080
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 5902 3108 5908 3120
rect 5736 3080 5908 3108
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3009 5043 3043
rect 4985 3003 5043 3009
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 5626 3040 5632 3052
rect 5399 3012 5632 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 5092 2904 5120 3003
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 5736 3049 5764 3080
rect 5902 3068 5908 3080
rect 5960 3068 5966 3120
rect 11238 3068 11244 3120
rect 11296 3108 11302 3120
rect 11296 3080 13124 3108
rect 11296 3068 11302 3080
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 8570 3040 8576 3052
rect 8628 3049 8634 3052
rect 5868 3012 5913 3040
rect 8540 3012 8576 3040
rect 5868 3000 5874 3012
rect 8570 3000 8576 3012
rect 8628 3003 8640 3049
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 10502 3040 10508 3052
rect 8895 3012 10508 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 8628 3000 8634 3003
rect 10502 3000 10508 3012
rect 10560 3040 10566 3052
rect 11790 3049 11796 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 10560 3012 11529 3040
rect 10560 3000 10566 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11784 3040 11796 3049
rect 11751 3012 11796 3040
rect 11517 3003 11575 3009
rect 11784 3003 11796 3012
rect 11790 3000 11796 3003
rect 11848 3000 11854 3052
rect 13096 3049 13124 3080
rect 13906 3068 13912 3120
rect 13964 3108 13970 3120
rect 14936 3108 14964 3148
rect 22370 3136 22376 3148
rect 22428 3136 22434 3188
rect 13964 3080 14964 3108
rect 15289 3111 15347 3117
rect 13964 3068 13970 3080
rect 15289 3077 15301 3111
rect 15335 3108 15347 3111
rect 15746 3108 15752 3120
rect 15335 3080 15752 3108
rect 15335 3077 15347 3080
rect 15289 3071 15347 3077
rect 15746 3068 15752 3080
rect 15804 3068 15810 3120
rect 22186 3108 22192 3120
rect 22066 3080 22192 3108
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3009 13139 3043
rect 13081 3003 13139 3009
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 22066 3040 22094 3080
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 13320 3012 22094 3040
rect 13320 3000 13326 3012
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2972 5503 2975
rect 6086 2972 6092 2984
rect 5491 2944 6092 2972
rect 5491 2941 5503 2944
rect 5445 2935 5503 2941
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 19518 2972 19524 2984
rect 15068 2944 19524 2972
rect 15068 2932 15074 2944
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 5902 2904 5908 2916
rect 5092 2876 5908 2904
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 14918 2904 14924 2916
rect 6288 2876 6960 2904
rect 14879 2876 14924 2904
rect 5261 2839 5319 2845
rect 5261 2805 5273 2839
rect 5307 2836 5319 2839
rect 5537 2839 5595 2845
rect 5537 2836 5549 2839
rect 5307 2808 5549 2836
rect 5307 2805 5319 2808
rect 5261 2799 5319 2805
rect 5537 2805 5549 2808
rect 5583 2836 5595 2839
rect 6288 2836 6316 2876
rect 5583 2808 6316 2836
rect 6932 2836 6960 2876
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 8202 2836 8208 2848
rect 6932 2808 8208 2836
rect 5583 2805 5595 2808
rect 5537 2799 5595 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 16022 2836 16028 2848
rect 14792 2808 16028 2836
rect 14792 2796 14798 2808
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 1104 2746 26128 2768
rect 1104 2694 5120 2746
rect 5172 2694 5184 2746
rect 5236 2694 5248 2746
rect 5300 2694 5312 2746
rect 5364 2694 5376 2746
rect 5428 2694 13462 2746
rect 13514 2694 13526 2746
rect 13578 2694 13590 2746
rect 13642 2694 13654 2746
rect 13706 2694 13718 2746
rect 13770 2694 21803 2746
rect 21855 2694 21867 2746
rect 21919 2694 21931 2746
rect 21983 2694 21995 2746
rect 22047 2694 22059 2746
rect 22111 2694 26128 2746
rect 1104 2672 26128 2694
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8202 2632 8208 2644
rect 8067 2604 8208 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 8570 2632 8576 2644
rect 8527 2604 8576 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 7929 2499 7987 2505
rect 7929 2496 7941 2499
rect 7524 2468 7941 2496
rect 7524 2456 7530 2468
rect 7929 2465 7941 2468
rect 7975 2465 7987 2499
rect 7929 2459 7987 2465
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 7800 2400 8217 2428
rect 7800 2388 7806 2400
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 8352 2400 8397 2428
rect 8352 2388 8358 2400
rect 1104 2202 26128 2224
rect 1104 2150 9291 2202
rect 9343 2150 9355 2202
rect 9407 2150 9419 2202
rect 9471 2150 9483 2202
rect 9535 2150 9547 2202
rect 9599 2150 17632 2202
rect 17684 2150 17696 2202
rect 17748 2150 17760 2202
rect 17812 2150 17824 2202
rect 17876 2150 17888 2202
rect 17940 2150 26128 2202
rect 1104 2128 26128 2150
rect 3142 1300 3148 1352
rect 3200 1340 3206 1352
rect 12894 1340 12900 1352
rect 3200 1312 12900 1340
rect 3200 1300 3206 1312
rect 12894 1300 12900 1312
rect 12952 1300 12958 1352
<< via1 >>
rect 26240 28475 26292 28484
rect 26240 28441 26249 28475
rect 26249 28441 26283 28475
rect 26283 28441 26292 28475
rect 26240 28432 26292 28441
rect 9291 27174 9343 27226
rect 9355 27174 9407 27226
rect 9419 27174 9471 27226
rect 9483 27174 9535 27226
rect 9547 27174 9599 27226
rect 17632 27174 17684 27226
rect 17696 27174 17748 27226
rect 17760 27174 17812 27226
rect 17824 27174 17876 27226
rect 17888 27174 17940 27226
rect 5120 26630 5172 26682
rect 5184 26630 5236 26682
rect 5248 26630 5300 26682
rect 5312 26630 5364 26682
rect 5376 26630 5428 26682
rect 13462 26630 13514 26682
rect 13526 26630 13578 26682
rect 13590 26630 13642 26682
rect 13654 26630 13706 26682
rect 13718 26630 13770 26682
rect 21803 26630 21855 26682
rect 21867 26630 21919 26682
rect 21931 26630 21983 26682
rect 21995 26630 22047 26682
rect 22059 26630 22111 26682
rect 12348 26528 12400 26580
rect 11796 26367 11848 26376
rect 11796 26333 11805 26367
rect 11805 26333 11839 26367
rect 11839 26333 11848 26367
rect 11796 26324 11848 26333
rect 12348 26324 12400 26376
rect 13820 26324 13872 26376
rect 14372 26324 14424 26376
rect 12716 26299 12768 26308
rect 12716 26265 12725 26299
rect 12725 26265 12759 26299
rect 12759 26265 12768 26299
rect 12716 26256 12768 26265
rect 14188 26256 14240 26308
rect 14556 26299 14608 26308
rect 14556 26265 14565 26299
rect 14565 26265 14599 26299
rect 14599 26265 14608 26299
rect 14556 26256 14608 26265
rect 12348 26231 12400 26240
rect 12348 26197 12357 26231
rect 12357 26197 12391 26231
rect 12391 26197 12400 26231
rect 12348 26188 12400 26197
rect 15476 26299 15528 26308
rect 15476 26265 15485 26299
rect 15485 26265 15519 26299
rect 15519 26265 15528 26299
rect 15476 26256 15528 26265
rect 16396 26256 16448 26308
rect 16580 26256 16632 26308
rect 16672 26299 16724 26308
rect 16672 26265 16681 26299
rect 16681 26265 16715 26299
rect 16715 26265 16724 26299
rect 16672 26256 16724 26265
rect 9291 26086 9343 26138
rect 9355 26086 9407 26138
rect 9419 26086 9471 26138
rect 9483 26086 9535 26138
rect 9547 26086 9599 26138
rect 17632 26086 17684 26138
rect 17696 26086 17748 26138
rect 17760 26086 17812 26138
rect 17824 26086 17876 26138
rect 17888 26086 17940 26138
rect 572 25984 624 26036
rect 11612 25984 11664 26036
rect 12716 25984 12768 26036
rect 15476 25984 15528 26036
rect 7932 25891 7984 25900
rect 7932 25857 7966 25891
rect 7966 25857 7984 25891
rect 11060 25891 11112 25900
rect 7932 25848 7984 25857
rect 11060 25857 11069 25891
rect 11069 25857 11103 25891
rect 11103 25857 11112 25891
rect 11060 25848 11112 25857
rect 11152 25891 11204 25900
rect 11152 25857 11161 25891
rect 11161 25857 11195 25891
rect 11195 25857 11204 25891
rect 11152 25848 11204 25857
rect 6920 25780 6972 25832
rect 13176 25848 13228 25900
rect 14924 25891 14976 25900
rect 14924 25857 14958 25891
rect 14958 25857 14976 25891
rect 14924 25848 14976 25857
rect 16488 25848 16540 25900
rect 21732 25848 21784 25900
rect 23112 25891 23164 25900
rect 23112 25857 23121 25891
rect 23121 25857 23155 25891
rect 23155 25857 23164 25891
rect 23112 25848 23164 25857
rect 25504 25848 25556 25900
rect 14648 25823 14700 25832
rect 14648 25789 14657 25823
rect 14657 25789 14691 25823
rect 14691 25789 14700 25823
rect 14648 25780 14700 25789
rect 16396 25780 16448 25832
rect 16120 25712 16172 25764
rect 7196 25644 7248 25696
rect 7564 25644 7616 25696
rect 8852 25644 8904 25696
rect 10692 25644 10744 25696
rect 14464 25687 14516 25696
rect 14464 25653 14473 25687
rect 14473 25653 14507 25687
rect 14507 25653 14516 25687
rect 14464 25644 14516 25653
rect 16580 25644 16632 25696
rect 19248 25644 19300 25696
rect 5120 25542 5172 25594
rect 5184 25542 5236 25594
rect 5248 25542 5300 25594
rect 5312 25542 5364 25594
rect 5376 25542 5428 25594
rect 13462 25542 13514 25594
rect 13526 25542 13578 25594
rect 13590 25542 13642 25594
rect 13654 25542 13706 25594
rect 13718 25542 13770 25594
rect 21803 25542 21855 25594
rect 21867 25542 21919 25594
rect 21931 25542 21983 25594
rect 21995 25542 22047 25594
rect 22059 25542 22111 25594
rect 6920 25440 6972 25492
rect 7196 25372 7248 25424
rect 7288 25304 7340 25356
rect 7104 25236 7156 25288
rect 7564 25236 7616 25288
rect 7840 25236 7892 25288
rect 8208 25304 8260 25356
rect 13176 25440 13228 25492
rect 14372 25483 14424 25492
rect 14372 25449 14381 25483
rect 14381 25449 14415 25483
rect 14415 25449 14424 25483
rect 14372 25440 14424 25449
rect 16580 25440 16632 25492
rect 16764 25440 16816 25492
rect 11796 25415 11848 25424
rect 10416 25347 10468 25356
rect 10416 25313 10425 25347
rect 10425 25313 10459 25347
rect 10459 25313 10468 25347
rect 10416 25304 10468 25313
rect 10692 25279 10744 25288
rect 10692 25245 10726 25279
rect 10726 25245 10744 25279
rect 6644 25168 6696 25220
rect 7196 25211 7248 25220
rect 7196 25177 7205 25211
rect 7205 25177 7239 25211
rect 7239 25177 7248 25211
rect 7196 25168 7248 25177
rect 7380 25211 7432 25220
rect 7380 25177 7389 25211
rect 7389 25177 7423 25211
rect 7423 25177 7432 25211
rect 7380 25168 7432 25177
rect 8116 25211 8168 25220
rect 8116 25177 8125 25211
rect 8125 25177 8159 25211
rect 8159 25177 8168 25211
rect 8116 25168 8168 25177
rect 9220 25168 9272 25220
rect 10692 25236 10744 25245
rect 11796 25381 11805 25415
rect 11805 25381 11839 25415
rect 11839 25381 11848 25415
rect 11796 25372 11848 25381
rect 12348 25304 12400 25356
rect 12624 25347 12676 25356
rect 12624 25313 12633 25347
rect 12633 25313 12667 25347
rect 12667 25313 12676 25347
rect 12624 25304 12676 25313
rect 12808 25279 12860 25288
rect 12808 25245 12817 25279
rect 12817 25245 12851 25279
rect 12851 25245 12860 25279
rect 12808 25236 12860 25245
rect 14188 25372 14240 25424
rect 14464 25304 14516 25356
rect 14648 25304 14700 25356
rect 25044 25347 25096 25356
rect 25044 25313 25053 25347
rect 25053 25313 25087 25347
rect 25087 25313 25096 25347
rect 25044 25304 25096 25313
rect 13820 25279 13872 25288
rect 13820 25245 13829 25279
rect 13829 25245 13863 25279
rect 13863 25245 13872 25279
rect 13820 25236 13872 25245
rect 14096 25279 14148 25288
rect 14096 25245 14105 25279
rect 14105 25245 14139 25279
rect 14139 25245 14148 25279
rect 14096 25236 14148 25245
rect 15016 25279 15068 25288
rect 15016 25245 15025 25279
rect 15025 25245 15059 25279
rect 15059 25245 15068 25279
rect 15016 25236 15068 25245
rect 18328 25279 18380 25288
rect 18328 25245 18337 25279
rect 18337 25245 18371 25279
rect 18371 25245 18380 25279
rect 18328 25236 18380 25245
rect 13176 25211 13228 25220
rect 13176 25177 13185 25211
rect 13185 25177 13219 25211
rect 13219 25177 13228 25211
rect 13176 25168 13228 25177
rect 15108 25168 15160 25220
rect 8392 25100 8444 25152
rect 11704 25100 11756 25152
rect 11980 25143 12032 25152
rect 11980 25109 11989 25143
rect 11989 25109 12023 25143
rect 12023 25109 12032 25143
rect 11980 25100 12032 25109
rect 12348 25143 12400 25152
rect 12348 25109 12357 25143
rect 12357 25109 12391 25143
rect 12391 25109 12400 25143
rect 12348 25100 12400 25109
rect 14464 25100 14516 25152
rect 14832 25143 14884 25152
rect 14832 25109 14841 25143
rect 14841 25109 14875 25143
rect 14875 25109 14884 25143
rect 14832 25100 14884 25109
rect 16856 25168 16908 25220
rect 16396 25100 16448 25152
rect 9291 24998 9343 25050
rect 9355 24998 9407 25050
rect 9419 24998 9471 25050
rect 9483 24998 9535 25050
rect 9547 24998 9599 25050
rect 17632 24998 17684 25050
rect 17696 24998 17748 25050
rect 17760 24998 17812 25050
rect 17824 24998 17876 25050
rect 17888 24998 17940 25050
rect 7840 24896 7892 24948
rect 7932 24896 7984 24948
rect 8116 24896 8168 24948
rect 1676 24828 1728 24880
rect 2688 24828 2740 24880
rect 6736 24803 6788 24812
rect 6736 24769 6745 24803
rect 6745 24769 6779 24803
rect 6779 24769 6788 24803
rect 7104 24803 7156 24812
rect 6736 24760 6788 24769
rect 7104 24769 7113 24803
rect 7113 24769 7147 24803
rect 7147 24769 7156 24803
rect 7104 24760 7156 24769
rect 7288 24803 7340 24812
rect 7288 24769 7297 24803
rect 7297 24769 7331 24803
rect 7331 24769 7340 24803
rect 7288 24760 7340 24769
rect 7748 24828 7800 24880
rect 8484 24828 8536 24880
rect 7196 24692 7248 24744
rect 8208 24760 8260 24812
rect 12164 24896 12216 24948
rect 13176 24896 13228 24948
rect 10968 24871 11020 24880
rect 10968 24837 11002 24871
rect 11002 24837 11020 24871
rect 10968 24828 11020 24837
rect 14372 24896 14424 24948
rect 16856 24896 16908 24948
rect 14280 24871 14332 24880
rect 14280 24837 14289 24871
rect 14289 24837 14323 24871
rect 14323 24837 14332 24871
rect 14280 24828 14332 24837
rect 15384 24828 15436 24880
rect 16488 24828 16540 24880
rect 9220 24803 9272 24812
rect 9220 24769 9229 24803
rect 9229 24769 9263 24803
rect 9263 24769 9272 24803
rect 9220 24760 9272 24769
rect 7840 24692 7892 24744
rect 8760 24692 8812 24744
rect 11060 24760 11112 24812
rect 11336 24803 11388 24812
rect 11336 24769 11345 24803
rect 11345 24769 11379 24803
rect 11379 24769 11388 24803
rect 11336 24760 11388 24769
rect 11704 24760 11756 24812
rect 13268 24760 13320 24812
rect 13360 24760 13412 24812
rect 14096 24760 14148 24812
rect 14556 24760 14608 24812
rect 14832 24760 14884 24812
rect 15568 24803 15620 24812
rect 7840 24556 7892 24608
rect 8116 24556 8168 24608
rect 11888 24692 11940 24744
rect 12164 24735 12216 24744
rect 12164 24701 12173 24735
rect 12173 24701 12207 24735
rect 12207 24701 12216 24735
rect 12164 24692 12216 24701
rect 12624 24692 12676 24744
rect 14004 24735 14056 24744
rect 14004 24701 14013 24735
rect 14013 24701 14047 24735
rect 14047 24701 14056 24735
rect 15568 24769 15577 24803
rect 15577 24769 15611 24803
rect 15611 24769 15620 24803
rect 15568 24760 15620 24769
rect 16120 24803 16172 24812
rect 16120 24769 16129 24803
rect 16129 24769 16172 24803
rect 16120 24760 16172 24769
rect 16396 24803 16448 24812
rect 16396 24769 16405 24803
rect 16405 24769 16439 24803
rect 16439 24769 16448 24803
rect 16396 24760 16448 24769
rect 14004 24692 14056 24701
rect 12348 24624 12400 24676
rect 14924 24624 14976 24676
rect 15660 24692 15712 24744
rect 16580 24692 16632 24744
rect 17040 24803 17092 24812
rect 17040 24769 17083 24803
rect 17083 24769 17092 24803
rect 17040 24760 17092 24769
rect 16764 24735 16816 24744
rect 16764 24701 16773 24735
rect 16773 24701 16807 24735
rect 16807 24701 16816 24735
rect 16764 24692 16816 24701
rect 10508 24556 10560 24608
rect 12532 24599 12584 24608
rect 12532 24565 12541 24599
rect 12541 24565 12575 24599
rect 12575 24565 12584 24599
rect 12532 24556 12584 24565
rect 14556 24556 14608 24608
rect 16304 24556 16356 24608
rect 5120 24454 5172 24506
rect 5184 24454 5236 24506
rect 5248 24454 5300 24506
rect 5312 24454 5364 24506
rect 5376 24454 5428 24506
rect 13462 24454 13514 24506
rect 13526 24454 13578 24506
rect 13590 24454 13642 24506
rect 13654 24454 13706 24506
rect 13718 24454 13770 24506
rect 21803 24454 21855 24506
rect 21867 24454 21919 24506
rect 21931 24454 21983 24506
rect 21995 24454 22047 24506
rect 22059 24454 22111 24506
rect 2136 24395 2188 24404
rect 2136 24361 2145 24395
rect 2145 24361 2179 24395
rect 2179 24361 2188 24395
rect 2136 24352 2188 24361
rect 6368 24352 6420 24404
rect 7104 24352 7156 24404
rect 7288 24352 7340 24404
rect 7564 24352 7616 24404
rect 7840 24284 7892 24336
rect 8116 24284 8168 24336
rect 8392 24259 8444 24268
rect 8392 24225 8401 24259
rect 8401 24225 8435 24259
rect 8435 24225 8444 24259
rect 8392 24216 8444 24225
rect 8760 24216 8812 24268
rect 3792 24148 3844 24200
rect 7380 24148 7432 24200
rect 8024 24148 8076 24200
rect 10416 24259 10468 24268
rect 10416 24225 10425 24259
rect 10425 24225 10459 24259
rect 10459 24225 10468 24259
rect 10416 24216 10468 24225
rect 11152 24352 11204 24404
rect 11980 24352 12032 24404
rect 12532 24395 12584 24404
rect 12532 24361 12541 24395
rect 12541 24361 12575 24395
rect 12575 24361 12584 24395
rect 12532 24352 12584 24361
rect 12808 24352 12860 24404
rect 14004 24352 14056 24404
rect 14556 24395 14608 24404
rect 14556 24361 14565 24395
rect 14565 24361 14599 24395
rect 14599 24361 14608 24395
rect 14556 24352 14608 24361
rect 15016 24352 15068 24404
rect 15568 24352 15620 24404
rect 10876 24216 10928 24268
rect 13360 24216 13412 24268
rect 16304 24259 16356 24268
rect 16304 24225 16313 24259
rect 16313 24225 16347 24259
rect 16347 24225 16356 24259
rect 16304 24216 16356 24225
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 5264 24080 5316 24132
rect 5908 24080 5960 24132
rect 6828 24080 6880 24132
rect 6736 24012 6788 24064
rect 7564 24012 7616 24064
rect 8392 24080 8444 24132
rect 10140 24123 10192 24132
rect 10140 24089 10158 24123
rect 10158 24089 10192 24123
rect 10140 24080 10192 24089
rect 11244 24148 11296 24200
rect 11336 24148 11388 24200
rect 12348 24148 12400 24200
rect 15108 24191 15160 24200
rect 11152 24080 11204 24132
rect 7932 24055 7984 24064
rect 7932 24021 7941 24055
rect 7941 24021 7975 24055
rect 7975 24021 7984 24055
rect 7932 24012 7984 24021
rect 8944 24012 8996 24064
rect 10600 24055 10652 24064
rect 10600 24021 10609 24055
rect 10609 24021 10643 24055
rect 10643 24021 10652 24055
rect 10600 24012 10652 24021
rect 12256 24012 12308 24064
rect 14188 24123 14240 24132
rect 14188 24089 14197 24123
rect 14197 24089 14231 24123
rect 14231 24089 14240 24123
rect 14188 24080 14240 24089
rect 14464 24080 14516 24132
rect 15108 24157 15117 24191
rect 15117 24157 15151 24191
rect 15151 24157 15160 24191
rect 15108 24148 15160 24157
rect 18328 24148 18380 24200
rect 18880 24148 18932 24200
rect 19248 24191 19300 24200
rect 19248 24157 19257 24191
rect 19257 24157 19291 24191
rect 19291 24157 19300 24191
rect 19248 24148 19300 24157
rect 19524 24148 19576 24200
rect 17040 24080 17092 24132
rect 18604 24080 18656 24132
rect 20444 24080 20496 24132
rect 16028 24012 16080 24064
rect 16580 24012 16632 24064
rect 18512 24012 18564 24064
rect 19616 24055 19668 24064
rect 19616 24021 19625 24055
rect 19625 24021 19659 24055
rect 19659 24021 19668 24055
rect 19616 24012 19668 24021
rect 9291 23910 9343 23962
rect 9355 23910 9407 23962
rect 9419 23910 9471 23962
rect 9483 23910 9535 23962
rect 9547 23910 9599 23962
rect 17632 23910 17684 23962
rect 17696 23910 17748 23962
rect 17760 23910 17812 23962
rect 17824 23910 17876 23962
rect 17888 23910 17940 23962
rect 5264 23851 5316 23860
rect 5264 23817 5273 23851
rect 5273 23817 5307 23851
rect 5307 23817 5316 23851
rect 5264 23808 5316 23817
rect 5908 23851 5960 23860
rect 5908 23817 5917 23851
rect 5917 23817 5951 23851
rect 5951 23817 5960 23851
rect 5908 23808 5960 23817
rect 8024 23851 8076 23860
rect 8024 23817 8033 23851
rect 8033 23817 8067 23851
rect 8067 23817 8076 23851
rect 8024 23808 8076 23817
rect 8208 23808 8260 23860
rect 7288 23740 7340 23792
rect 5816 23604 5868 23656
rect 6368 23672 6420 23724
rect 6644 23715 6696 23724
rect 6644 23681 6653 23715
rect 6653 23681 6687 23715
rect 6687 23681 6696 23715
rect 6644 23672 6696 23681
rect 7932 23740 7984 23792
rect 7748 23672 7800 23724
rect 8024 23672 8076 23724
rect 7656 23647 7708 23656
rect 7656 23613 7665 23647
rect 7665 23613 7699 23647
rect 7699 23613 7708 23647
rect 8392 23808 8444 23860
rect 10140 23851 10192 23860
rect 10140 23817 10149 23851
rect 10149 23817 10183 23851
rect 10183 23817 10192 23851
rect 10140 23808 10192 23817
rect 11244 23808 11296 23860
rect 9772 23740 9824 23792
rect 8668 23715 8720 23724
rect 7656 23604 7708 23613
rect 8024 23536 8076 23588
rect 6736 23511 6788 23520
rect 6736 23477 6745 23511
rect 6745 23477 6779 23511
rect 6779 23477 6788 23511
rect 6736 23468 6788 23477
rect 8668 23681 8677 23715
rect 8677 23681 8711 23715
rect 8711 23681 8720 23715
rect 8668 23672 8720 23681
rect 8760 23715 8812 23724
rect 8760 23681 8769 23715
rect 8769 23681 8803 23715
rect 8803 23681 8812 23715
rect 8944 23715 8996 23724
rect 8760 23672 8812 23681
rect 8944 23681 8953 23715
rect 8953 23681 8987 23715
rect 8987 23681 8996 23715
rect 8944 23672 8996 23681
rect 8484 23647 8536 23656
rect 8484 23613 8493 23647
rect 8493 23613 8527 23647
rect 8527 23613 8536 23647
rect 9128 23672 9180 23724
rect 10140 23715 10192 23724
rect 10140 23681 10149 23715
rect 10149 23681 10183 23715
rect 10183 23681 10192 23715
rect 10140 23672 10192 23681
rect 10968 23740 11020 23792
rect 11060 23715 11112 23724
rect 8484 23604 8536 23613
rect 9864 23647 9916 23656
rect 9864 23613 9873 23647
rect 9873 23613 9907 23647
rect 9907 23613 9916 23647
rect 11060 23681 11069 23715
rect 11069 23681 11103 23715
rect 11103 23681 11112 23715
rect 11060 23672 11112 23681
rect 11520 23715 11572 23724
rect 11520 23681 11529 23715
rect 11529 23681 11563 23715
rect 11563 23681 11572 23715
rect 11520 23672 11572 23681
rect 11888 23808 11940 23860
rect 12256 23851 12308 23860
rect 12256 23817 12265 23851
rect 12265 23817 12299 23851
rect 12299 23817 12308 23851
rect 12256 23808 12308 23817
rect 13268 23851 13320 23860
rect 13268 23817 13277 23851
rect 13277 23817 13311 23851
rect 13311 23817 13320 23851
rect 13268 23808 13320 23817
rect 17040 23851 17092 23860
rect 17040 23817 17049 23851
rect 17049 23817 17083 23851
rect 17083 23817 17092 23851
rect 17040 23808 17092 23817
rect 15108 23740 15160 23792
rect 16028 23740 16080 23792
rect 18052 23740 18104 23792
rect 13268 23672 13320 23724
rect 17500 23715 17552 23724
rect 17500 23681 17509 23715
rect 17509 23681 17543 23715
rect 17543 23681 17552 23715
rect 17500 23672 17552 23681
rect 18972 23808 19024 23860
rect 18512 23740 18564 23792
rect 18604 23672 18656 23724
rect 19156 23715 19208 23724
rect 19156 23681 19190 23715
rect 19190 23681 19208 23715
rect 20444 23715 20496 23724
rect 19156 23672 19208 23681
rect 20444 23681 20453 23715
rect 20453 23681 20487 23715
rect 20487 23681 20496 23715
rect 20444 23672 20496 23681
rect 12624 23647 12676 23656
rect 9864 23604 9916 23613
rect 12624 23613 12633 23647
rect 12633 23613 12667 23647
rect 12667 23613 12676 23647
rect 12624 23604 12676 23613
rect 14464 23604 14516 23656
rect 16396 23604 16448 23656
rect 8852 23511 8904 23520
rect 8852 23477 8861 23511
rect 8861 23477 8895 23511
rect 8895 23477 8904 23511
rect 8852 23468 8904 23477
rect 8944 23468 8996 23520
rect 10600 23511 10652 23520
rect 10600 23477 10609 23511
rect 10609 23477 10643 23511
rect 10643 23477 10652 23511
rect 10600 23468 10652 23477
rect 10968 23468 11020 23520
rect 11152 23468 11204 23520
rect 15660 23511 15712 23520
rect 15660 23477 15669 23511
rect 15669 23477 15703 23511
rect 15703 23477 15712 23511
rect 15660 23468 15712 23477
rect 18512 23604 18564 23656
rect 18880 23647 18932 23656
rect 18880 23613 18889 23647
rect 18889 23613 18923 23647
rect 18923 23613 18932 23647
rect 18880 23604 18932 23613
rect 19248 23468 19300 23520
rect 19524 23468 19576 23520
rect 5120 23366 5172 23418
rect 5184 23366 5236 23418
rect 5248 23366 5300 23418
rect 5312 23366 5364 23418
rect 5376 23366 5428 23418
rect 13462 23366 13514 23418
rect 13526 23366 13578 23418
rect 13590 23366 13642 23418
rect 13654 23366 13706 23418
rect 13718 23366 13770 23418
rect 21803 23366 21855 23418
rect 21867 23366 21919 23418
rect 21931 23366 21983 23418
rect 21995 23366 22047 23418
rect 22059 23366 22111 23418
rect 5816 23264 5868 23316
rect 7748 23264 7800 23316
rect 8116 23264 8168 23316
rect 8484 23307 8536 23316
rect 8484 23273 8493 23307
rect 8493 23273 8527 23307
rect 8527 23273 8536 23307
rect 8484 23264 8536 23273
rect 14188 23307 14240 23316
rect 14188 23273 14197 23307
rect 14197 23273 14231 23307
rect 14231 23273 14240 23307
rect 14188 23264 14240 23273
rect 16580 23307 16632 23316
rect 16580 23273 16589 23307
rect 16589 23273 16623 23307
rect 16623 23273 16632 23307
rect 16580 23264 16632 23273
rect 7748 23128 7800 23180
rect 8760 23196 8812 23248
rect 11520 23196 11572 23248
rect 16028 23196 16080 23248
rect 18512 23196 18564 23248
rect 18880 23196 18932 23248
rect 2136 23103 2188 23112
rect 2136 23069 2145 23103
rect 2145 23069 2179 23103
rect 2179 23069 2188 23103
rect 2136 23060 2188 23069
rect 6736 23060 6788 23112
rect 7380 23103 7432 23112
rect 7380 23069 7389 23103
rect 7389 23069 7423 23103
rect 7423 23069 7432 23103
rect 7380 23060 7432 23069
rect 7656 23103 7708 23112
rect 7656 23069 7665 23103
rect 7665 23069 7699 23103
rect 7699 23069 7708 23103
rect 7656 23060 7708 23069
rect 8300 23128 8352 23180
rect 7104 22992 7156 23044
rect 8208 23060 8260 23112
rect 8576 23060 8628 23112
rect 16672 23128 16724 23180
rect 9772 23103 9824 23112
rect 8300 23035 8352 23044
rect 8300 23001 8309 23035
rect 8309 23001 8343 23035
rect 8343 23001 8352 23035
rect 8300 22992 8352 23001
rect 9220 22992 9272 23044
rect 9772 23069 9781 23103
rect 9781 23069 9815 23103
rect 9815 23069 9824 23103
rect 9772 23060 9824 23069
rect 9864 23103 9916 23112
rect 9864 23069 9873 23103
rect 9873 23069 9907 23103
rect 9907 23069 9916 23103
rect 13268 23103 13320 23112
rect 9864 23060 9916 23069
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 13268 23060 13320 23069
rect 18696 23128 18748 23180
rect 19340 23128 19392 23180
rect 10048 23035 10100 23044
rect 10048 23001 10057 23035
rect 10057 23001 10091 23035
rect 10091 23001 10100 23035
rect 10048 22992 10100 23001
rect 11888 22992 11940 23044
rect 14648 23035 14700 23044
rect 14648 23001 14657 23035
rect 14657 23001 14691 23035
rect 14691 23001 14700 23035
rect 14648 22992 14700 23001
rect 16856 22992 16908 23044
rect 18052 22992 18104 23044
rect 19892 23060 19944 23112
rect 19340 22992 19392 23044
rect 19984 22992 20036 23044
rect 6276 22924 6328 22976
rect 6644 22924 6696 22976
rect 7012 22967 7064 22976
rect 7012 22933 7021 22967
rect 7021 22933 7055 22967
rect 7055 22933 7064 22967
rect 7012 22924 7064 22933
rect 8576 22924 8628 22976
rect 8760 22924 8812 22976
rect 9772 22924 9824 22976
rect 10784 22924 10836 22976
rect 11336 22924 11388 22976
rect 12624 22924 12676 22976
rect 13360 22924 13412 22976
rect 14556 22967 14608 22976
rect 14556 22933 14565 22967
rect 14565 22933 14599 22967
rect 14599 22933 14608 22967
rect 14556 22924 14608 22933
rect 16120 22967 16172 22976
rect 16120 22933 16129 22967
rect 16129 22933 16163 22967
rect 16163 22933 16172 22967
rect 16120 22924 16172 22933
rect 16212 22967 16264 22976
rect 16212 22933 16221 22967
rect 16221 22933 16255 22967
rect 16255 22933 16264 22967
rect 16212 22924 16264 22933
rect 19156 22924 19208 22976
rect 19708 22967 19760 22976
rect 19708 22933 19717 22967
rect 19717 22933 19751 22967
rect 19751 22933 19760 22967
rect 20352 23060 20404 23112
rect 23388 23060 23440 23112
rect 19708 22924 19760 22933
rect 20260 22924 20312 22976
rect 22192 22992 22244 23044
rect 22100 22924 22152 22976
rect 23204 22924 23256 22976
rect 23480 22967 23532 22976
rect 23480 22933 23489 22967
rect 23489 22933 23523 22967
rect 23523 22933 23532 22967
rect 23480 22924 23532 22933
rect 9291 22822 9343 22874
rect 9355 22822 9407 22874
rect 9419 22822 9471 22874
rect 9483 22822 9535 22874
rect 9547 22822 9599 22874
rect 17632 22822 17684 22874
rect 17696 22822 17748 22874
rect 17760 22822 17812 22874
rect 17824 22822 17876 22874
rect 17888 22822 17940 22874
rect 7012 22720 7064 22772
rect 7380 22720 7432 22772
rect 8300 22763 8352 22772
rect 8300 22729 8309 22763
rect 8309 22729 8343 22763
rect 8343 22729 8352 22763
rect 8300 22720 8352 22729
rect 10140 22720 10192 22772
rect 14280 22720 14332 22772
rect 16120 22720 16172 22772
rect 17500 22763 17552 22772
rect 17500 22729 17509 22763
rect 17509 22729 17543 22763
rect 17543 22729 17552 22763
rect 17500 22720 17552 22729
rect 7104 22652 7156 22704
rect 3976 22584 4028 22636
rect 7840 22627 7892 22636
rect 7840 22593 7849 22627
rect 7849 22593 7883 22627
rect 7883 22593 7892 22627
rect 7840 22584 7892 22593
rect 8392 22627 8444 22636
rect 8392 22593 8401 22627
rect 8401 22593 8435 22627
rect 8435 22593 8444 22627
rect 8392 22584 8444 22593
rect 8576 22627 8628 22636
rect 8576 22593 8585 22627
rect 8585 22593 8619 22627
rect 8619 22593 8628 22627
rect 8576 22584 8628 22593
rect 8760 22627 8812 22636
rect 8760 22593 8769 22627
rect 8769 22593 8803 22627
rect 8803 22593 8812 22627
rect 8760 22584 8812 22593
rect 9220 22627 9272 22636
rect 9220 22593 9229 22627
rect 9229 22593 9263 22627
rect 9263 22593 9272 22627
rect 9220 22584 9272 22593
rect 9772 22584 9824 22636
rect 10692 22627 10744 22636
rect 10692 22593 10701 22627
rect 10701 22593 10735 22627
rect 10735 22593 10744 22627
rect 10692 22584 10744 22593
rect 11888 22627 11940 22636
rect 11888 22593 11897 22627
rect 11897 22593 11931 22627
rect 11931 22593 11940 22627
rect 11888 22584 11940 22593
rect 13360 22584 13412 22636
rect 14096 22627 14148 22636
rect 4344 22516 4396 22568
rect 9128 22516 9180 22568
rect 10140 22559 10192 22568
rect 10140 22525 10149 22559
rect 10149 22525 10183 22559
rect 10183 22525 10192 22559
rect 10140 22516 10192 22525
rect 10324 22559 10376 22568
rect 10324 22525 10333 22559
rect 10333 22525 10367 22559
rect 10367 22525 10376 22559
rect 10324 22516 10376 22525
rect 10600 22516 10652 22568
rect 14096 22593 14105 22627
rect 14105 22593 14139 22627
rect 14139 22593 14148 22627
rect 14096 22584 14148 22593
rect 15200 22584 15252 22636
rect 17408 22652 17460 22704
rect 19708 22720 19760 22772
rect 19892 22720 19944 22772
rect 22192 22763 22244 22772
rect 22192 22729 22201 22763
rect 22201 22729 22235 22763
rect 22235 22729 22244 22763
rect 22192 22720 22244 22729
rect 24860 22720 24912 22772
rect 17776 22652 17828 22704
rect 8208 22448 8260 22500
rect 3700 22380 3752 22432
rect 6828 22380 6880 22432
rect 9496 22423 9548 22432
rect 9496 22389 9505 22423
rect 9505 22389 9539 22423
rect 9539 22389 9548 22423
rect 9496 22380 9548 22389
rect 9772 22380 9824 22432
rect 10692 22448 10744 22500
rect 13912 22516 13964 22568
rect 14556 22516 14608 22568
rect 14832 22559 14884 22568
rect 14832 22525 14841 22559
rect 14841 22525 14875 22559
rect 14875 22525 14884 22559
rect 14832 22516 14884 22525
rect 15844 22559 15896 22568
rect 15844 22525 15853 22559
rect 15853 22525 15887 22559
rect 15887 22525 15896 22559
rect 15844 22516 15896 22525
rect 16672 22584 16724 22636
rect 18696 22627 18748 22636
rect 15384 22491 15436 22500
rect 10324 22380 10376 22432
rect 10416 22380 10468 22432
rect 12348 22380 12400 22432
rect 13084 22380 13136 22432
rect 15384 22457 15393 22491
rect 15393 22457 15427 22491
rect 15427 22457 15436 22491
rect 15384 22448 15436 22457
rect 16948 22559 17000 22568
rect 16948 22525 16957 22559
rect 16957 22525 16991 22559
rect 16991 22525 17000 22559
rect 16948 22516 17000 22525
rect 18696 22593 18705 22627
rect 18705 22593 18739 22627
rect 18739 22593 18748 22627
rect 18696 22584 18748 22593
rect 18972 22627 19024 22636
rect 18972 22593 18981 22627
rect 18981 22593 19015 22627
rect 19015 22593 19024 22627
rect 18972 22584 19024 22593
rect 19616 22652 19668 22704
rect 19708 22627 19760 22636
rect 19708 22593 19717 22627
rect 19717 22593 19751 22627
rect 19751 22593 19760 22627
rect 19708 22584 19760 22593
rect 17408 22491 17460 22500
rect 17408 22457 17417 22491
rect 17417 22457 17451 22491
rect 17451 22457 17460 22491
rect 17408 22448 17460 22457
rect 19524 22516 19576 22568
rect 20352 22627 20404 22636
rect 20352 22593 20361 22627
rect 20361 22593 20395 22627
rect 20395 22593 20404 22627
rect 20352 22584 20404 22593
rect 20720 22584 20772 22636
rect 22284 22584 22336 22636
rect 22652 22627 22704 22636
rect 22652 22593 22661 22627
rect 22661 22593 22695 22627
rect 22695 22593 22704 22627
rect 22652 22584 22704 22593
rect 23204 22627 23256 22636
rect 23204 22593 23213 22627
rect 23213 22593 23247 22627
rect 23247 22593 23256 22627
rect 23204 22584 23256 22593
rect 23664 22584 23716 22636
rect 23940 22584 23992 22636
rect 24676 22584 24728 22636
rect 20904 22516 20956 22568
rect 21088 22559 21140 22568
rect 21088 22525 21097 22559
rect 21097 22525 21131 22559
rect 21131 22525 21140 22559
rect 21088 22516 21140 22525
rect 23020 22516 23072 22568
rect 24400 22559 24452 22568
rect 18788 22448 18840 22500
rect 19340 22448 19392 22500
rect 19708 22448 19760 22500
rect 13820 22380 13872 22432
rect 16396 22423 16448 22432
rect 16396 22389 16405 22423
rect 16405 22389 16439 22423
rect 16439 22389 16448 22423
rect 16396 22380 16448 22389
rect 16856 22380 16908 22432
rect 17776 22380 17828 22432
rect 18512 22423 18564 22432
rect 18512 22389 18521 22423
rect 18521 22389 18555 22423
rect 18555 22389 18564 22423
rect 18512 22380 18564 22389
rect 22376 22380 22428 22432
rect 24400 22525 24409 22559
rect 24409 22525 24443 22559
rect 24443 22525 24452 22559
rect 24400 22516 24452 22525
rect 23848 22380 23900 22432
rect 5120 22278 5172 22330
rect 5184 22278 5236 22330
rect 5248 22278 5300 22330
rect 5312 22278 5364 22330
rect 5376 22278 5428 22330
rect 13462 22278 13514 22330
rect 13526 22278 13578 22330
rect 13590 22278 13642 22330
rect 13654 22278 13706 22330
rect 13718 22278 13770 22330
rect 21803 22278 21855 22330
rect 21867 22278 21919 22330
rect 21931 22278 21983 22330
rect 21995 22278 22047 22330
rect 22059 22278 22111 22330
rect 7656 22176 7708 22228
rect 8116 22176 8168 22228
rect 9496 22219 9548 22228
rect 5816 22108 5868 22160
rect 6276 22108 6328 22160
rect 9496 22185 9505 22219
rect 9505 22185 9539 22219
rect 9539 22185 9548 22219
rect 9496 22176 9548 22185
rect 10140 22176 10192 22228
rect 13360 22176 13412 22228
rect 14096 22219 14148 22228
rect 14096 22185 14105 22219
rect 14105 22185 14139 22219
rect 14139 22185 14148 22219
rect 14096 22176 14148 22185
rect 6920 22040 6972 22092
rect 9956 22108 10008 22160
rect 13912 22108 13964 22160
rect 15200 22176 15252 22228
rect 16212 22219 16264 22228
rect 16212 22185 16221 22219
rect 16221 22185 16255 22219
rect 16255 22185 16264 22219
rect 16212 22176 16264 22185
rect 16948 22176 17000 22228
rect 20260 22176 20312 22228
rect 21088 22176 21140 22228
rect 22376 22176 22428 22228
rect 24860 22219 24912 22228
rect 24860 22185 24869 22219
rect 24869 22185 24903 22219
rect 24903 22185 24912 22219
rect 24860 22176 24912 22185
rect 16120 22108 16172 22160
rect 2780 21972 2832 22024
rect 3792 22015 3844 22024
rect 3792 21981 3801 22015
rect 3801 21981 3835 22015
rect 3835 21981 3844 22015
rect 3792 21972 3844 21981
rect 4804 21972 4856 22024
rect 3240 21904 3292 21956
rect 4160 21904 4212 21956
rect 3332 21879 3384 21888
rect 3332 21845 3341 21879
rect 3341 21845 3375 21879
rect 3375 21845 3384 21879
rect 3332 21836 3384 21845
rect 4344 21836 4396 21888
rect 5356 21836 5408 21888
rect 6644 21972 6696 22024
rect 8300 21972 8352 22024
rect 8576 21972 8628 22024
rect 10692 22040 10744 22092
rect 10784 22040 10836 22092
rect 6000 21904 6052 21956
rect 8484 21904 8536 21956
rect 9680 22015 9732 22024
rect 9680 21981 9689 22015
rect 9689 21981 9723 22015
rect 9723 21981 9732 22015
rect 9864 22015 9916 22024
rect 9680 21972 9732 21981
rect 9864 21981 9873 22015
rect 9873 21981 9907 22015
rect 9907 21981 9916 22015
rect 9864 21972 9916 21981
rect 10416 22015 10468 22024
rect 10416 21981 10425 22015
rect 10425 21981 10459 22015
rect 10459 21981 10468 22015
rect 10416 21972 10468 21981
rect 11244 22015 11296 22024
rect 11244 21981 11253 22015
rect 11253 21981 11287 22015
rect 11287 21981 11296 22015
rect 11244 21972 11296 21981
rect 13360 22015 13412 22024
rect 11612 21904 11664 21956
rect 12256 21904 12308 21956
rect 6368 21836 6420 21888
rect 8208 21836 8260 21888
rect 8668 21879 8720 21888
rect 8668 21845 8677 21879
rect 8677 21845 8711 21879
rect 8711 21845 8720 21879
rect 8668 21836 8720 21845
rect 9864 21836 9916 21888
rect 9956 21836 10008 21888
rect 11336 21836 11388 21888
rect 12072 21836 12124 21888
rect 13360 21981 13369 22015
rect 13369 21981 13403 22015
rect 13403 21981 13412 22015
rect 13360 21972 13412 21981
rect 14556 22040 14608 22092
rect 16396 22040 16448 22092
rect 15200 22015 15252 22024
rect 15200 21981 15209 22015
rect 15209 21981 15243 22015
rect 15243 21981 15252 22015
rect 15200 21972 15252 21981
rect 15384 22015 15436 22024
rect 15384 21981 15393 22015
rect 15393 21981 15427 22015
rect 15427 21981 15436 22015
rect 16764 22108 16816 22160
rect 22284 22151 22336 22160
rect 22284 22117 22293 22151
rect 22293 22117 22327 22151
rect 22327 22117 22336 22151
rect 22284 22108 22336 22117
rect 23020 22108 23072 22160
rect 16856 22083 16908 22092
rect 16856 22049 16865 22083
rect 16865 22049 16899 22083
rect 16899 22049 16908 22083
rect 16856 22040 16908 22049
rect 23848 22083 23900 22092
rect 23848 22049 23857 22083
rect 23857 22049 23891 22083
rect 23891 22049 23900 22083
rect 23848 22040 23900 22049
rect 15384 21972 15436 21981
rect 19708 21972 19760 22024
rect 24676 22015 24728 22024
rect 24676 21981 24685 22015
rect 24685 21981 24719 22015
rect 24719 21981 24728 22015
rect 24676 21972 24728 21981
rect 15476 21904 15528 21956
rect 15844 21947 15896 21956
rect 15844 21913 15853 21947
rect 15853 21913 15887 21947
rect 15887 21913 15896 21947
rect 15844 21904 15896 21913
rect 17040 21947 17092 21956
rect 17040 21913 17049 21947
rect 17049 21913 17083 21947
rect 17083 21913 17092 21947
rect 17040 21904 17092 21913
rect 14464 21879 14516 21888
rect 14464 21845 14473 21879
rect 14473 21845 14507 21879
rect 14507 21845 14516 21879
rect 14464 21836 14516 21845
rect 14556 21879 14608 21888
rect 14556 21845 14565 21879
rect 14565 21845 14599 21879
rect 14599 21845 14608 21879
rect 15016 21879 15068 21888
rect 14556 21836 14608 21845
rect 15016 21845 15025 21879
rect 15025 21845 15059 21879
rect 15059 21845 15068 21879
rect 15016 21836 15068 21845
rect 15200 21836 15252 21888
rect 15752 21879 15804 21888
rect 15752 21845 15761 21879
rect 15761 21845 15795 21879
rect 15795 21845 15804 21879
rect 15752 21836 15804 21845
rect 23480 21904 23532 21956
rect 24032 21904 24084 21956
rect 23572 21836 23624 21888
rect 23756 21879 23808 21888
rect 23756 21845 23765 21879
rect 23765 21845 23799 21879
rect 23799 21845 23808 21879
rect 23756 21836 23808 21845
rect 23848 21836 23900 21888
rect 25044 21879 25096 21888
rect 25044 21845 25053 21879
rect 25053 21845 25087 21879
rect 25087 21845 25096 21879
rect 25044 21836 25096 21845
rect 9291 21734 9343 21786
rect 9355 21734 9407 21786
rect 9419 21734 9471 21786
rect 9483 21734 9535 21786
rect 9547 21734 9599 21786
rect 17632 21734 17684 21786
rect 17696 21734 17748 21786
rect 17760 21734 17812 21786
rect 17824 21734 17876 21786
rect 17888 21734 17940 21786
rect 3240 21675 3292 21684
rect 3240 21641 3249 21675
rect 3249 21641 3283 21675
rect 3283 21641 3292 21675
rect 3240 21632 3292 21641
rect 4804 21632 4856 21684
rect 5816 21675 5868 21684
rect 5816 21641 5825 21675
rect 5825 21641 5859 21675
rect 5859 21641 5868 21675
rect 5816 21632 5868 21641
rect 5908 21632 5960 21684
rect 3976 21564 4028 21616
rect 3240 21496 3292 21548
rect 4436 21496 4488 21548
rect 5356 21539 5408 21548
rect 5356 21505 5374 21539
rect 5374 21505 5408 21539
rect 5356 21496 5408 21505
rect 3700 21471 3752 21480
rect 3700 21437 3709 21471
rect 3709 21437 3743 21471
rect 3743 21437 3752 21471
rect 3700 21428 3752 21437
rect 3884 21428 3936 21480
rect 5724 21428 5776 21480
rect 6460 21496 6512 21548
rect 6368 21471 6420 21480
rect 6368 21437 6377 21471
rect 6377 21437 6411 21471
rect 6411 21437 6420 21471
rect 6368 21428 6420 21437
rect 7564 21632 7616 21684
rect 10784 21632 10836 21684
rect 11152 21675 11204 21684
rect 11152 21641 11161 21675
rect 11161 21641 11195 21675
rect 11195 21641 11204 21675
rect 11152 21632 11204 21641
rect 11612 21675 11664 21684
rect 11612 21641 11621 21675
rect 11621 21641 11655 21675
rect 11655 21641 11664 21675
rect 11612 21632 11664 21641
rect 7012 21539 7064 21548
rect 7012 21505 7021 21539
rect 7021 21505 7055 21539
rect 7055 21505 7064 21539
rect 7012 21496 7064 21505
rect 7656 21539 7708 21548
rect 7656 21505 7665 21539
rect 7665 21505 7699 21539
rect 7699 21505 7708 21539
rect 7656 21496 7708 21505
rect 7748 21496 7800 21548
rect 8024 21428 8076 21480
rect 8668 21428 8720 21480
rect 8944 21428 8996 21480
rect 9680 21539 9732 21548
rect 9680 21505 9689 21539
rect 9689 21505 9723 21539
rect 9723 21505 9732 21539
rect 9680 21496 9732 21505
rect 9956 21496 10008 21548
rect 9772 21428 9824 21480
rect 10140 21539 10192 21548
rect 10140 21505 10149 21539
rect 10149 21505 10183 21539
rect 10183 21505 10192 21539
rect 10140 21496 10192 21505
rect 12164 21632 12216 21684
rect 14556 21632 14608 21684
rect 14832 21632 14884 21684
rect 15752 21632 15804 21684
rect 24676 21632 24728 21684
rect 12256 21539 12308 21548
rect 6828 21360 6880 21412
rect 7012 21360 7064 21412
rect 7564 21360 7616 21412
rect 8300 21360 8352 21412
rect 9128 21360 9180 21412
rect 10876 21428 10928 21480
rect 4620 21292 4672 21344
rect 7104 21335 7156 21344
rect 7104 21301 7113 21335
rect 7113 21301 7147 21335
rect 7147 21301 7156 21335
rect 7104 21292 7156 21301
rect 7840 21292 7892 21344
rect 8668 21292 8720 21344
rect 10140 21292 10192 21344
rect 11152 21360 11204 21412
rect 12256 21505 12265 21539
rect 12265 21505 12299 21539
rect 12299 21505 12308 21539
rect 12256 21496 12308 21505
rect 12900 21496 12952 21548
rect 13084 21539 13136 21548
rect 13084 21505 13093 21539
rect 13093 21505 13127 21539
rect 13127 21505 13136 21539
rect 13084 21496 13136 21505
rect 13820 21539 13872 21548
rect 13268 21428 13320 21480
rect 13820 21505 13829 21539
rect 13829 21505 13863 21539
rect 13863 21505 13872 21539
rect 13820 21496 13872 21505
rect 10416 21292 10468 21344
rect 13820 21292 13872 21344
rect 15016 21496 15068 21548
rect 15384 21564 15436 21616
rect 20904 21564 20956 21616
rect 21732 21564 21784 21616
rect 22192 21564 22244 21616
rect 22468 21564 22520 21616
rect 17684 21496 17736 21548
rect 19156 21496 19208 21548
rect 23480 21564 23532 21616
rect 25044 21564 25096 21616
rect 23388 21539 23440 21548
rect 18880 21428 18932 21480
rect 23388 21505 23397 21539
rect 23397 21505 23431 21539
rect 23431 21505 23440 21539
rect 23388 21496 23440 21505
rect 15476 21360 15528 21412
rect 16396 21360 16448 21412
rect 17132 21360 17184 21412
rect 18420 21360 18472 21412
rect 18328 21292 18380 21344
rect 23664 21292 23716 21344
rect 24032 21292 24084 21344
rect 24584 21292 24636 21344
rect 5120 21190 5172 21242
rect 5184 21190 5236 21242
rect 5248 21190 5300 21242
rect 5312 21190 5364 21242
rect 5376 21190 5428 21242
rect 13462 21190 13514 21242
rect 13526 21190 13578 21242
rect 13590 21190 13642 21242
rect 13654 21190 13706 21242
rect 13718 21190 13770 21242
rect 21803 21190 21855 21242
rect 21867 21190 21919 21242
rect 21931 21190 21983 21242
rect 21995 21190 22047 21242
rect 22059 21190 22111 21242
rect 3976 21131 4028 21140
rect 3976 21097 3985 21131
rect 3985 21097 4019 21131
rect 4019 21097 4028 21131
rect 3976 21088 4028 21097
rect 4160 21131 4212 21140
rect 4160 21097 4169 21131
rect 4169 21097 4203 21131
rect 4203 21097 4212 21131
rect 4160 21088 4212 21097
rect 4620 21131 4672 21140
rect 4620 21097 4629 21131
rect 4629 21097 4663 21131
rect 4663 21097 4672 21131
rect 4620 21088 4672 21097
rect 4436 21020 4488 21072
rect 6644 21088 6696 21140
rect 7748 21088 7800 21140
rect 3240 20927 3292 20936
rect 3240 20893 3249 20927
rect 3249 20893 3283 20927
rect 3283 20893 3292 20927
rect 3240 20884 3292 20893
rect 4068 20884 4120 20936
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 4436 20927 4488 20936
rect 4436 20893 4445 20927
rect 4445 20893 4479 20927
rect 4479 20893 4488 20927
rect 4712 20995 4764 21004
rect 4712 20961 4721 20995
rect 4721 20961 4755 20995
rect 4755 20961 4764 20995
rect 4712 20952 4764 20961
rect 6828 21020 6880 21072
rect 7656 21020 7708 21072
rect 8944 21088 8996 21140
rect 11888 21088 11940 21140
rect 17684 21131 17736 21140
rect 17684 21097 17693 21131
rect 17693 21097 17727 21131
rect 17727 21097 17736 21131
rect 17684 21088 17736 21097
rect 23296 21088 23348 21140
rect 23848 21088 23900 21140
rect 23940 21131 23992 21140
rect 23940 21097 23949 21131
rect 23949 21097 23983 21131
rect 23983 21097 23992 21131
rect 23940 21088 23992 21097
rect 24400 21088 24452 21140
rect 6644 20952 6696 21004
rect 4436 20884 4488 20893
rect 5816 20884 5868 20936
rect 6368 20927 6420 20936
rect 6368 20893 6377 20927
rect 6377 20893 6411 20927
rect 6411 20893 6420 20927
rect 6368 20884 6420 20893
rect 6460 20884 6512 20936
rect 8208 20952 8260 21004
rect 8576 20995 8628 21004
rect 8576 20961 8585 20995
rect 8585 20961 8619 20995
rect 8619 20961 8628 20995
rect 8576 20952 8628 20961
rect 6920 20884 6972 20936
rect 7472 20927 7524 20936
rect 7472 20893 7481 20927
rect 7481 20893 7515 20927
rect 7515 20893 7524 20927
rect 7472 20884 7524 20893
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 7656 20884 7708 20893
rect 8024 20927 8076 20936
rect 8024 20893 8033 20927
rect 8033 20893 8067 20927
rect 8067 20893 8076 20927
rect 8024 20884 8076 20893
rect 8392 20927 8444 20936
rect 8392 20893 8401 20927
rect 8401 20893 8435 20927
rect 8435 20893 8444 20927
rect 8392 20884 8444 20893
rect 9772 21020 9824 21072
rect 10416 21020 10468 21072
rect 11152 21020 11204 21072
rect 14464 21020 14516 21072
rect 14924 21020 14976 21072
rect 25044 21020 25096 21072
rect 9864 20952 9916 21004
rect 18052 20952 18104 21004
rect 9956 20927 10008 20936
rect 4620 20816 4672 20868
rect 3792 20748 3844 20800
rect 5632 20816 5684 20868
rect 8668 20859 8720 20868
rect 5540 20748 5592 20800
rect 8668 20825 8677 20859
rect 8677 20825 8711 20859
rect 8711 20825 8720 20859
rect 8668 20816 8720 20825
rect 8300 20748 8352 20800
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 10140 20927 10192 20936
rect 10140 20893 10149 20927
rect 10149 20893 10183 20927
rect 10183 20893 10192 20927
rect 10140 20884 10192 20893
rect 10876 20884 10928 20936
rect 14832 20927 14884 20936
rect 14832 20893 14841 20927
rect 14841 20893 14875 20927
rect 14875 20893 14884 20927
rect 14832 20884 14884 20893
rect 16488 20884 16540 20936
rect 18328 20884 18380 20936
rect 18512 20884 18564 20936
rect 21732 20952 21784 21004
rect 22376 20927 22428 20936
rect 11060 20859 11112 20868
rect 11060 20825 11069 20859
rect 11069 20825 11103 20859
rect 11103 20825 11112 20859
rect 11060 20816 11112 20825
rect 15292 20859 15344 20868
rect 15292 20825 15301 20859
rect 15301 20825 15335 20859
rect 15335 20825 15344 20859
rect 15292 20816 15344 20825
rect 18972 20816 19024 20868
rect 10784 20748 10836 20800
rect 11336 20748 11388 20800
rect 14464 20748 14516 20800
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 18696 20748 18748 20800
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 22836 20927 22888 20936
rect 22836 20893 22845 20927
rect 22845 20893 22879 20927
rect 22879 20893 22888 20927
rect 22836 20884 22888 20893
rect 23664 20884 23716 20936
rect 24584 20927 24636 20936
rect 24584 20893 24593 20927
rect 24593 20893 24627 20927
rect 24627 20893 24636 20927
rect 24584 20884 24636 20893
rect 20168 20816 20220 20868
rect 23848 20816 23900 20868
rect 19524 20791 19576 20800
rect 19524 20757 19533 20791
rect 19533 20757 19567 20791
rect 19567 20757 19576 20791
rect 19524 20748 19576 20757
rect 20260 20748 20312 20800
rect 20536 20748 20588 20800
rect 21456 20748 21508 20800
rect 21548 20748 21600 20800
rect 9291 20646 9343 20698
rect 9355 20646 9407 20698
rect 9419 20646 9471 20698
rect 9483 20646 9535 20698
rect 9547 20646 9599 20698
rect 17632 20646 17684 20698
rect 17696 20646 17748 20698
rect 17760 20646 17812 20698
rect 17824 20646 17876 20698
rect 17888 20646 17940 20698
rect 4436 20587 4488 20596
rect 4436 20553 4445 20587
rect 4445 20553 4479 20587
rect 4479 20553 4488 20587
rect 4436 20544 4488 20553
rect 4712 20544 4764 20596
rect 1492 20408 1544 20460
rect 2780 20476 2832 20528
rect 3884 20451 3936 20460
rect 3884 20417 3893 20451
rect 3893 20417 3927 20451
rect 3927 20417 3936 20451
rect 3884 20408 3936 20417
rect 5448 20451 5500 20460
rect 5448 20417 5457 20451
rect 5457 20417 5491 20451
rect 5491 20417 5500 20451
rect 5448 20408 5500 20417
rect 3792 20383 3844 20392
rect 3792 20349 3801 20383
rect 3801 20349 3835 20383
rect 3835 20349 3844 20383
rect 3792 20340 3844 20349
rect 4160 20272 4212 20324
rect 7012 20544 7064 20596
rect 7656 20544 7708 20596
rect 8576 20544 8628 20596
rect 9956 20587 10008 20596
rect 9956 20553 9965 20587
rect 9965 20553 9999 20587
rect 9999 20553 10008 20587
rect 9956 20544 10008 20553
rect 11336 20587 11388 20596
rect 11336 20553 11345 20587
rect 11345 20553 11379 20587
rect 11379 20553 11388 20587
rect 11336 20544 11388 20553
rect 11980 20544 12032 20596
rect 12348 20544 12400 20596
rect 15292 20544 15344 20596
rect 18052 20587 18104 20596
rect 18052 20553 18061 20587
rect 18061 20553 18095 20587
rect 18095 20553 18104 20587
rect 18052 20544 18104 20553
rect 5724 20451 5776 20460
rect 5724 20417 5733 20451
rect 5733 20417 5767 20451
rect 5767 20417 5776 20451
rect 5724 20408 5776 20417
rect 6920 20476 6972 20528
rect 9864 20451 9916 20460
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 10876 20451 10928 20460
rect 10876 20417 10885 20451
rect 10885 20417 10919 20451
rect 10919 20417 10928 20451
rect 10876 20408 10928 20417
rect 11152 20451 11204 20460
rect 11152 20417 11161 20451
rect 11161 20417 11195 20451
rect 11195 20417 11204 20451
rect 11152 20408 11204 20417
rect 11244 20408 11296 20460
rect 14648 20476 14700 20528
rect 16488 20476 16540 20528
rect 6368 20383 6420 20392
rect 6368 20349 6377 20383
rect 6377 20349 6411 20383
rect 6411 20349 6420 20383
rect 6368 20340 6420 20349
rect 14464 20451 14516 20460
rect 14464 20417 14498 20451
rect 14498 20417 14516 20451
rect 14464 20408 14516 20417
rect 15200 20408 15252 20460
rect 18512 20476 18564 20528
rect 16396 20340 16448 20392
rect 18604 20451 18656 20460
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 19064 20451 19116 20460
rect 19064 20417 19073 20451
rect 19073 20417 19107 20451
rect 19107 20417 19116 20451
rect 19064 20408 19116 20417
rect 22376 20544 22428 20596
rect 19248 20476 19300 20528
rect 19892 20408 19944 20460
rect 21548 20476 21600 20528
rect 22468 20476 22520 20528
rect 23664 20476 23716 20528
rect 21456 20451 21508 20460
rect 21456 20417 21465 20451
rect 21465 20417 21499 20451
rect 21499 20417 21508 20451
rect 21456 20408 21508 20417
rect 24308 20451 24360 20460
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24308 20408 24360 20417
rect 24492 20451 24544 20460
rect 24492 20417 24501 20451
rect 24501 20417 24535 20451
rect 24535 20417 24544 20451
rect 24492 20408 24544 20417
rect 3148 20204 3200 20256
rect 7104 20204 7156 20256
rect 8300 20204 8352 20256
rect 11336 20204 11388 20256
rect 12900 20247 12952 20256
rect 12900 20213 12909 20247
rect 12909 20213 12943 20247
rect 12943 20213 12952 20247
rect 12900 20204 12952 20213
rect 15844 20247 15896 20256
rect 15844 20213 15853 20247
rect 15853 20213 15887 20247
rect 15887 20213 15896 20247
rect 15844 20204 15896 20213
rect 18236 20340 18288 20392
rect 18696 20383 18748 20392
rect 18696 20349 18705 20383
rect 18705 20349 18739 20383
rect 18739 20349 18748 20383
rect 18696 20340 18748 20349
rect 18420 20204 18472 20256
rect 18880 20204 18932 20256
rect 19432 20315 19484 20324
rect 19432 20281 19441 20315
rect 19441 20281 19475 20315
rect 19475 20281 19484 20315
rect 19432 20272 19484 20281
rect 20536 20340 20588 20392
rect 21548 20383 21600 20392
rect 21548 20349 21557 20383
rect 21557 20349 21591 20383
rect 21591 20349 21600 20383
rect 21548 20340 21600 20349
rect 24952 20340 25004 20392
rect 19616 20204 19668 20256
rect 24308 20272 24360 20324
rect 23848 20204 23900 20256
rect 24584 20247 24636 20256
rect 24584 20213 24593 20247
rect 24593 20213 24627 20247
rect 24627 20213 24636 20247
rect 24584 20204 24636 20213
rect 5120 20102 5172 20154
rect 5184 20102 5236 20154
rect 5248 20102 5300 20154
rect 5312 20102 5364 20154
rect 5376 20102 5428 20154
rect 13462 20102 13514 20154
rect 13526 20102 13578 20154
rect 13590 20102 13642 20154
rect 13654 20102 13706 20154
rect 13718 20102 13770 20154
rect 21803 20102 21855 20154
rect 21867 20102 21919 20154
rect 21931 20102 21983 20154
rect 21995 20102 22047 20154
rect 22059 20102 22111 20154
rect 1492 19907 1544 19916
rect 1492 19873 1501 19907
rect 1501 19873 1535 19907
rect 1535 19873 1544 19907
rect 1492 19864 1544 19873
rect 3148 19839 3200 19848
rect 3148 19805 3157 19839
rect 3157 19805 3191 19839
rect 3191 19805 3200 19839
rect 3148 19796 3200 19805
rect 4068 20000 4120 20052
rect 3884 19932 3936 19984
rect 4160 19839 4212 19848
rect 4160 19805 4169 19839
rect 4169 19805 4203 19839
rect 4203 19805 4212 19839
rect 4160 19796 4212 19805
rect 5724 20000 5776 20052
rect 6276 20043 6328 20052
rect 6276 20009 6285 20043
rect 6285 20009 6319 20043
rect 6319 20009 6328 20043
rect 6276 20000 6328 20009
rect 11060 20000 11112 20052
rect 11520 19932 11572 19984
rect 8116 19864 8168 19916
rect 14832 20000 14884 20052
rect 16396 20000 16448 20052
rect 16488 20000 16540 20052
rect 18420 20043 18472 20052
rect 12900 19864 12952 19916
rect 4436 19728 4488 19780
rect 10968 19796 11020 19848
rect 4252 19660 4304 19712
rect 7104 19660 7156 19712
rect 7288 19703 7340 19712
rect 7288 19669 7297 19703
rect 7297 19669 7331 19703
rect 7331 19669 7340 19703
rect 7288 19660 7340 19669
rect 8300 19660 8352 19712
rect 11336 19796 11388 19848
rect 11612 19728 11664 19780
rect 11704 19660 11756 19712
rect 12256 19839 12308 19848
rect 12256 19805 12265 19839
rect 12265 19805 12299 19839
rect 12299 19805 12308 19839
rect 12256 19796 12308 19805
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 12348 19728 12400 19780
rect 15844 19932 15896 19984
rect 18420 20009 18429 20043
rect 18429 20009 18463 20043
rect 18463 20009 18472 20043
rect 18420 20000 18472 20009
rect 18972 20043 19024 20052
rect 18972 20009 18981 20043
rect 18981 20009 19015 20043
rect 19015 20009 19024 20043
rect 18972 20000 19024 20009
rect 19616 20043 19668 20052
rect 19616 20009 19625 20043
rect 19625 20009 19659 20043
rect 19659 20009 19668 20043
rect 19616 20000 19668 20009
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 19432 19932 19484 19984
rect 15660 19864 15712 19916
rect 13820 19796 13872 19848
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 16028 19796 16080 19848
rect 16948 19864 17000 19916
rect 22836 19864 22888 19916
rect 24308 19932 24360 19984
rect 25320 19932 25372 19984
rect 20812 19839 20864 19848
rect 20812 19805 20821 19839
rect 20821 19805 20855 19839
rect 20855 19805 20864 19839
rect 20812 19796 20864 19805
rect 21548 19796 21600 19848
rect 22744 19796 22796 19848
rect 23296 19839 23348 19848
rect 15292 19728 15344 19780
rect 16856 19728 16908 19780
rect 18052 19771 18104 19780
rect 18052 19737 18061 19771
rect 18061 19737 18095 19771
rect 18095 19737 18104 19771
rect 18052 19728 18104 19737
rect 21456 19728 21508 19780
rect 12164 19660 12216 19712
rect 12624 19703 12676 19712
rect 12624 19669 12633 19703
rect 12633 19669 12667 19703
rect 12667 19669 12676 19703
rect 12624 19660 12676 19669
rect 16580 19703 16632 19712
rect 16580 19669 16589 19703
rect 16589 19669 16623 19703
rect 16623 19669 16632 19703
rect 16580 19660 16632 19669
rect 17408 19660 17460 19712
rect 19524 19660 19576 19712
rect 20536 19703 20588 19712
rect 20536 19669 20545 19703
rect 20545 19669 20579 19703
rect 20579 19669 20588 19703
rect 20536 19660 20588 19669
rect 21180 19660 21232 19712
rect 22468 19728 22520 19780
rect 23296 19805 23305 19839
rect 23305 19805 23339 19839
rect 23339 19805 23348 19839
rect 23296 19796 23348 19805
rect 23848 19839 23900 19848
rect 23848 19805 23857 19839
rect 23857 19805 23900 19839
rect 23848 19796 23900 19805
rect 24492 19796 24544 19848
rect 24952 19839 25004 19848
rect 24952 19805 24961 19839
rect 24961 19805 24995 19839
rect 24995 19805 25004 19839
rect 24952 19796 25004 19805
rect 25044 19839 25096 19848
rect 25044 19805 25053 19839
rect 25053 19805 25087 19839
rect 25087 19805 25096 19839
rect 25044 19796 25096 19805
rect 23940 19728 23992 19780
rect 24216 19660 24268 19712
rect 9291 19558 9343 19610
rect 9355 19558 9407 19610
rect 9419 19558 9471 19610
rect 9483 19558 9535 19610
rect 9547 19558 9599 19610
rect 17632 19558 17684 19610
rect 17696 19558 17748 19610
rect 17760 19558 17812 19610
rect 17824 19558 17876 19610
rect 17888 19558 17940 19610
rect 3884 19456 3936 19508
rect 4344 19456 4396 19508
rect 5632 19456 5684 19508
rect 6276 19456 6328 19508
rect 8208 19456 8260 19508
rect 1492 19320 1544 19372
rect 6000 19388 6052 19440
rect 6368 19388 6420 19440
rect 4160 19320 4212 19372
rect 4344 19363 4396 19372
rect 4344 19329 4353 19363
rect 4353 19329 4387 19363
rect 4387 19329 4396 19363
rect 4344 19320 4396 19329
rect 5540 19320 5592 19372
rect 6644 19320 6696 19372
rect 7012 19320 7064 19372
rect 4252 19295 4304 19304
rect 4252 19261 4261 19295
rect 4261 19261 4295 19295
rect 4295 19261 4304 19295
rect 4252 19252 4304 19261
rect 5816 19252 5868 19304
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 7288 19252 7340 19304
rect 8208 19320 8260 19372
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 11152 19456 11204 19508
rect 11060 19363 11112 19372
rect 11060 19329 11069 19363
rect 11069 19329 11103 19363
rect 11103 19329 11112 19363
rect 11060 19320 11112 19329
rect 11336 19363 11388 19372
rect 11336 19329 11345 19363
rect 11345 19329 11379 19363
rect 11379 19329 11388 19363
rect 11336 19320 11388 19329
rect 11704 19363 11756 19372
rect 5448 19184 5500 19236
rect 7104 19184 7156 19236
rect 7472 19227 7524 19236
rect 7472 19193 7481 19227
rect 7481 19193 7515 19227
rect 7515 19193 7524 19227
rect 7472 19184 7524 19193
rect 6460 19159 6512 19168
rect 6460 19125 6469 19159
rect 6469 19125 6503 19159
rect 6503 19125 6512 19159
rect 6460 19116 6512 19125
rect 6828 19116 6880 19168
rect 11244 19184 11296 19236
rect 11704 19329 11712 19363
rect 11712 19329 11746 19363
rect 11746 19329 11756 19363
rect 11704 19320 11756 19329
rect 12256 19456 12308 19508
rect 14096 19499 14148 19508
rect 14096 19465 14105 19499
rect 14105 19465 14139 19499
rect 14139 19465 14148 19499
rect 14096 19456 14148 19465
rect 15292 19456 15344 19508
rect 18696 19499 18748 19508
rect 18696 19465 18705 19499
rect 18705 19465 18739 19499
rect 18739 19465 18748 19499
rect 18696 19456 18748 19465
rect 19524 19499 19576 19508
rect 19524 19465 19533 19499
rect 19533 19465 19567 19499
rect 19567 19465 19576 19499
rect 19524 19456 19576 19465
rect 20444 19456 20496 19508
rect 21180 19456 21232 19508
rect 21456 19499 21508 19508
rect 21456 19465 21465 19499
rect 21465 19465 21499 19499
rect 21499 19465 21508 19499
rect 21456 19456 21508 19465
rect 22744 19499 22796 19508
rect 22744 19465 22753 19499
rect 22753 19465 22787 19499
rect 22787 19465 22796 19499
rect 22744 19456 22796 19465
rect 12164 19320 12216 19372
rect 11612 19184 11664 19236
rect 11888 19184 11940 19236
rect 12624 19388 12676 19440
rect 14372 19388 14424 19440
rect 18052 19388 18104 19440
rect 16028 19363 16080 19372
rect 16028 19329 16037 19363
rect 16037 19329 16071 19363
rect 16071 19329 16080 19363
rect 16028 19320 16080 19329
rect 18880 19388 18932 19440
rect 19616 19388 19668 19440
rect 18328 19320 18380 19372
rect 12532 19252 12584 19304
rect 12624 19252 12676 19304
rect 15660 19252 15712 19304
rect 19064 19320 19116 19372
rect 19708 19363 19760 19372
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 20996 19363 21048 19372
rect 20996 19329 21005 19363
rect 21005 19329 21039 19363
rect 21039 19329 21048 19363
rect 20996 19320 21048 19329
rect 22468 19388 22520 19440
rect 20904 19252 20956 19304
rect 21272 19295 21324 19304
rect 21272 19261 21281 19295
rect 21281 19261 21315 19295
rect 21315 19261 21324 19295
rect 21272 19252 21324 19261
rect 23848 19456 23900 19508
rect 24952 19456 25004 19508
rect 23572 19431 23624 19440
rect 23572 19397 23590 19431
rect 23590 19397 23624 19431
rect 23572 19388 23624 19397
rect 23204 19363 23256 19372
rect 23204 19329 23213 19363
rect 23213 19329 23247 19363
rect 23247 19329 23256 19363
rect 25412 19388 25464 19440
rect 23204 19320 23256 19329
rect 25228 19320 25280 19372
rect 14740 19184 14792 19236
rect 17960 19184 18012 19236
rect 8300 19116 8352 19168
rect 12164 19159 12216 19168
rect 12164 19125 12173 19159
rect 12173 19125 12207 19159
rect 12207 19125 12216 19159
rect 12164 19116 12216 19125
rect 16580 19116 16632 19168
rect 22192 19184 22244 19236
rect 22836 19252 22888 19304
rect 24032 19252 24084 19304
rect 20536 19116 20588 19168
rect 21272 19116 21324 19168
rect 22284 19116 22336 19168
rect 23296 19116 23348 19168
rect 23480 19116 23532 19168
rect 5120 19014 5172 19066
rect 5184 19014 5236 19066
rect 5248 19014 5300 19066
rect 5312 19014 5364 19066
rect 5376 19014 5428 19066
rect 13462 19014 13514 19066
rect 13526 19014 13578 19066
rect 13590 19014 13642 19066
rect 13654 19014 13706 19066
rect 13718 19014 13770 19066
rect 21803 19014 21855 19066
rect 21867 19014 21919 19066
rect 21931 19014 21983 19066
rect 21995 19014 22047 19066
rect 22059 19014 22111 19066
rect 4896 18912 4948 18964
rect 5908 18912 5960 18964
rect 6828 18912 6880 18964
rect 8484 18912 8536 18964
rect 10692 18912 10744 18964
rect 16580 18912 16632 18964
rect 17224 18912 17276 18964
rect 21732 18912 21784 18964
rect 22192 18955 22244 18964
rect 22192 18921 22201 18955
rect 22201 18921 22235 18955
rect 22235 18921 22244 18955
rect 22192 18912 22244 18921
rect 5632 18844 5684 18896
rect 11612 18844 11664 18896
rect 17132 18887 17184 18896
rect 17132 18853 17141 18887
rect 17141 18853 17175 18887
rect 17175 18853 17184 18887
rect 20628 18887 20680 18896
rect 17132 18844 17184 18853
rect 20628 18853 20637 18887
rect 20637 18853 20671 18887
rect 20671 18853 20680 18887
rect 20628 18844 20680 18853
rect 23664 18912 23716 18964
rect 25228 18955 25280 18964
rect 25228 18921 25237 18955
rect 25237 18921 25271 18955
rect 25271 18921 25280 18955
rect 25228 18912 25280 18921
rect 4252 18708 4304 18760
rect 5632 18751 5684 18760
rect 5632 18717 5641 18751
rect 5641 18717 5675 18751
rect 5675 18717 5684 18751
rect 5632 18708 5684 18717
rect 6460 18708 6512 18760
rect 7196 18751 7248 18760
rect 7196 18717 7205 18751
rect 7205 18717 7239 18751
rect 7239 18717 7248 18751
rect 7196 18708 7248 18717
rect 11152 18708 11204 18760
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 12624 18708 12676 18760
rect 13360 18708 13412 18760
rect 15108 18708 15160 18760
rect 19616 18708 19668 18760
rect 20812 18751 20864 18760
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 23204 18776 23256 18828
rect 23940 18819 23992 18828
rect 23940 18785 23949 18819
rect 23949 18785 23983 18819
rect 23983 18785 23992 18819
rect 23940 18776 23992 18785
rect 5172 18640 5224 18692
rect 7104 18640 7156 18692
rect 7472 18683 7524 18692
rect 7472 18649 7506 18683
rect 7506 18649 7524 18683
rect 7472 18640 7524 18649
rect 10508 18640 10560 18692
rect 12164 18640 12216 18692
rect 15568 18640 15620 18692
rect 17040 18640 17092 18692
rect 20444 18683 20496 18692
rect 20444 18649 20462 18683
rect 20462 18649 20496 18683
rect 20444 18640 20496 18649
rect 21088 18683 21140 18692
rect 21088 18649 21122 18683
rect 21122 18649 21140 18683
rect 21088 18640 21140 18649
rect 3792 18572 3844 18624
rect 6828 18572 6880 18624
rect 6920 18572 6972 18624
rect 7656 18572 7708 18624
rect 8392 18572 8444 18624
rect 11336 18615 11388 18624
rect 11336 18581 11345 18615
rect 11345 18581 11379 18615
rect 11379 18581 11388 18615
rect 11336 18572 11388 18581
rect 11980 18572 12032 18624
rect 12532 18572 12584 18624
rect 14832 18572 14884 18624
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 16396 18615 16448 18624
rect 16396 18581 16405 18615
rect 16405 18581 16439 18615
rect 16439 18581 16448 18615
rect 16396 18572 16448 18581
rect 16672 18572 16724 18624
rect 16948 18572 17000 18624
rect 17224 18572 17276 18624
rect 17500 18572 17552 18624
rect 18236 18572 18288 18624
rect 21364 18572 21416 18624
rect 23572 18640 23624 18692
rect 24216 18776 24268 18828
rect 25136 18640 25188 18692
rect 23480 18615 23532 18624
rect 23480 18581 23489 18615
rect 23489 18581 23523 18615
rect 23523 18581 23532 18615
rect 23480 18572 23532 18581
rect 23848 18615 23900 18624
rect 23848 18581 23857 18615
rect 23857 18581 23891 18615
rect 23891 18581 23900 18615
rect 23848 18572 23900 18581
rect 24216 18572 24268 18624
rect 25412 18751 25464 18760
rect 25412 18717 25421 18751
rect 25421 18717 25455 18751
rect 25455 18717 25464 18751
rect 25412 18708 25464 18717
rect 9291 18470 9343 18522
rect 9355 18470 9407 18522
rect 9419 18470 9471 18522
rect 9483 18470 9535 18522
rect 9547 18470 9599 18522
rect 17632 18470 17684 18522
rect 17696 18470 17748 18522
rect 17760 18470 17812 18522
rect 17824 18470 17876 18522
rect 17888 18470 17940 18522
rect 3700 18368 3752 18420
rect 3240 18300 3292 18352
rect 3148 18232 3200 18284
rect 3792 18275 3844 18284
rect 3240 18207 3292 18216
rect 3240 18173 3249 18207
rect 3249 18173 3283 18207
rect 3283 18173 3292 18207
rect 3240 18164 3292 18173
rect 3792 18241 3801 18275
rect 3801 18241 3835 18275
rect 3835 18241 3844 18275
rect 3792 18232 3844 18241
rect 4252 18275 4304 18284
rect 4252 18241 4261 18275
rect 4261 18241 4295 18275
rect 4295 18241 4304 18275
rect 4252 18232 4304 18241
rect 5540 18368 5592 18420
rect 4804 18275 4856 18284
rect 2872 18139 2924 18148
rect 2872 18105 2881 18139
rect 2881 18105 2915 18139
rect 2915 18105 2924 18139
rect 2872 18096 2924 18105
rect 4344 18164 4396 18216
rect 4804 18241 4812 18275
rect 4812 18241 4846 18275
rect 4846 18241 4856 18275
rect 4804 18232 4856 18241
rect 4896 18275 4948 18284
rect 4896 18241 4905 18275
rect 4905 18241 4939 18275
rect 4939 18241 4948 18275
rect 5172 18275 5224 18284
rect 4896 18232 4948 18241
rect 5172 18241 5181 18275
rect 5181 18241 5215 18275
rect 5215 18241 5224 18275
rect 5172 18232 5224 18241
rect 5724 18368 5776 18420
rect 5448 18275 5500 18284
rect 5448 18241 5463 18275
rect 5463 18241 5497 18275
rect 5497 18241 5500 18275
rect 5448 18232 5500 18241
rect 5908 18232 5960 18284
rect 7748 18368 7800 18420
rect 8576 18368 8628 18420
rect 13820 18368 13872 18420
rect 14740 18411 14792 18420
rect 14740 18377 14749 18411
rect 14749 18377 14783 18411
rect 14783 18377 14792 18411
rect 14740 18368 14792 18377
rect 14832 18368 14884 18420
rect 15568 18411 15620 18420
rect 7196 18300 7248 18352
rect 7840 18300 7892 18352
rect 8116 18343 8168 18352
rect 8116 18309 8125 18343
rect 8125 18309 8159 18343
rect 8159 18309 8168 18343
rect 8116 18300 8168 18309
rect 8392 18300 8444 18352
rect 9680 18343 9732 18352
rect 9680 18309 9689 18343
rect 9689 18309 9723 18343
rect 9723 18309 9732 18343
rect 9680 18300 9732 18309
rect 11244 18300 11296 18352
rect 15568 18377 15577 18411
rect 15577 18377 15611 18411
rect 15611 18377 15620 18411
rect 15568 18368 15620 18377
rect 16672 18368 16724 18420
rect 20812 18368 20864 18420
rect 21088 18368 21140 18420
rect 21364 18411 21416 18420
rect 21364 18377 21373 18411
rect 21373 18377 21407 18411
rect 21407 18377 21416 18411
rect 21364 18368 21416 18377
rect 21732 18368 21784 18420
rect 22284 18411 22336 18420
rect 22284 18377 22293 18411
rect 22293 18377 22327 18411
rect 22327 18377 22336 18411
rect 22284 18368 22336 18377
rect 16396 18300 16448 18352
rect 21272 18300 21324 18352
rect 5816 18207 5868 18216
rect 5816 18173 5825 18207
rect 5825 18173 5859 18207
rect 5859 18173 5868 18207
rect 5816 18164 5868 18173
rect 11612 18232 11664 18284
rect 11888 18275 11940 18284
rect 10784 18164 10836 18216
rect 11888 18241 11897 18275
rect 11897 18241 11931 18275
rect 11931 18241 11940 18275
rect 11888 18232 11940 18241
rect 12072 18275 12124 18284
rect 12072 18241 12081 18275
rect 12081 18241 12115 18275
rect 12115 18241 12124 18275
rect 12072 18232 12124 18241
rect 13360 18275 13412 18284
rect 13360 18241 13369 18275
rect 13369 18241 13403 18275
rect 13403 18241 13412 18275
rect 13360 18232 13412 18241
rect 13452 18232 13504 18284
rect 4528 18096 4580 18148
rect 5448 18096 5500 18148
rect 5540 18096 5592 18148
rect 3792 18028 3844 18080
rect 5816 18028 5868 18080
rect 12900 18096 12952 18148
rect 7748 18071 7800 18080
rect 7748 18037 7757 18071
rect 7757 18037 7791 18071
rect 7791 18037 7800 18071
rect 7748 18028 7800 18037
rect 8300 18071 8352 18080
rect 8300 18037 8309 18071
rect 8309 18037 8343 18071
rect 8343 18037 8352 18071
rect 8300 18028 8352 18037
rect 12164 18071 12216 18080
rect 12164 18037 12173 18071
rect 12173 18037 12207 18071
rect 12207 18037 12216 18071
rect 12164 18028 12216 18037
rect 13084 18028 13136 18080
rect 15292 18207 15344 18216
rect 15292 18173 15301 18207
rect 15301 18173 15335 18207
rect 15335 18173 15344 18207
rect 15292 18164 15344 18173
rect 16580 18232 16632 18284
rect 16948 18275 17000 18284
rect 16948 18241 16957 18275
rect 16957 18241 16991 18275
rect 16991 18241 17000 18275
rect 16948 18232 17000 18241
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 18052 18232 18104 18284
rect 18144 18232 18196 18284
rect 18420 18275 18472 18284
rect 18420 18241 18429 18275
rect 18429 18241 18463 18275
rect 18463 18241 18472 18275
rect 18420 18232 18472 18241
rect 20628 18232 20680 18284
rect 20904 18232 20956 18284
rect 16396 18164 16448 18216
rect 17500 18164 17552 18216
rect 22560 18232 22612 18284
rect 24216 18368 24268 18420
rect 25320 18368 25372 18420
rect 24584 18300 24636 18352
rect 24032 18207 24084 18216
rect 15108 18096 15160 18148
rect 17408 18139 17460 18148
rect 17408 18105 17417 18139
rect 17417 18105 17451 18139
rect 17451 18105 17460 18139
rect 17408 18096 17460 18105
rect 24032 18173 24041 18207
rect 24041 18173 24075 18207
rect 24075 18173 24084 18207
rect 24032 18164 24084 18173
rect 16948 18028 17000 18080
rect 19248 18096 19300 18148
rect 20812 18096 20864 18148
rect 19064 18028 19116 18080
rect 5120 17926 5172 17978
rect 5184 17926 5236 17978
rect 5248 17926 5300 17978
rect 5312 17926 5364 17978
rect 5376 17926 5428 17978
rect 13462 17926 13514 17978
rect 13526 17926 13578 17978
rect 13590 17926 13642 17978
rect 13654 17926 13706 17978
rect 13718 17926 13770 17978
rect 21803 17926 21855 17978
rect 21867 17926 21919 17978
rect 21931 17926 21983 17978
rect 21995 17926 22047 17978
rect 22059 17926 22111 17978
rect 5448 17824 5500 17876
rect 4068 17756 4120 17808
rect 12532 17824 12584 17876
rect 12900 17867 12952 17876
rect 12900 17833 12909 17867
rect 12909 17833 12943 17867
rect 12943 17833 12952 17867
rect 12900 17824 12952 17833
rect 13360 17824 13412 17876
rect 10508 17799 10560 17808
rect 10508 17765 10517 17799
rect 10517 17765 10551 17799
rect 10551 17765 10560 17799
rect 10508 17756 10560 17765
rect 3792 17688 3844 17740
rect 5448 17688 5500 17740
rect 2044 17663 2096 17672
rect 2044 17629 2053 17663
rect 2053 17629 2087 17663
rect 2087 17629 2096 17663
rect 2044 17620 2096 17629
rect 2780 17552 2832 17604
rect 2964 17552 3016 17604
rect 4160 17595 4212 17604
rect 4160 17561 4169 17595
rect 4169 17561 4203 17595
rect 4203 17561 4212 17595
rect 4160 17552 4212 17561
rect 5540 17663 5592 17672
rect 4620 17552 4672 17604
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 5632 17620 5684 17672
rect 5816 17620 5868 17672
rect 7840 17620 7892 17672
rect 11336 17756 11388 17808
rect 13176 17756 13228 17808
rect 10968 17731 11020 17740
rect 10968 17697 10977 17731
rect 10977 17697 11011 17731
rect 11011 17697 11020 17731
rect 10968 17688 11020 17697
rect 12716 17688 12768 17740
rect 15936 17824 15988 17876
rect 16856 17824 16908 17876
rect 18052 17867 18104 17876
rect 18052 17833 18061 17867
rect 18061 17833 18095 17867
rect 18095 17833 18104 17867
rect 18052 17824 18104 17833
rect 18604 17824 18656 17876
rect 14464 17756 14516 17808
rect 17132 17756 17184 17808
rect 6092 17552 6144 17604
rect 6828 17552 6880 17604
rect 10692 17663 10744 17672
rect 10692 17629 10701 17663
rect 10701 17629 10735 17663
rect 10735 17629 10744 17663
rect 10692 17620 10744 17629
rect 11520 17663 11572 17672
rect 9864 17552 9916 17604
rect 10508 17552 10560 17604
rect 3884 17484 3936 17536
rect 4528 17484 4580 17536
rect 4896 17484 4948 17536
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7104 17484 7156 17493
rect 10232 17484 10284 17536
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 12164 17620 12216 17672
rect 12624 17620 12676 17672
rect 13084 17663 13136 17672
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 13268 17663 13320 17672
rect 13268 17629 13276 17663
rect 13276 17629 13310 17663
rect 13310 17629 13320 17663
rect 13268 17620 13320 17629
rect 13820 17620 13872 17672
rect 14740 17663 14792 17672
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 11612 17484 11664 17536
rect 14556 17484 14608 17536
rect 16948 17688 17000 17740
rect 19248 17688 19300 17740
rect 17224 17620 17276 17672
rect 15108 17552 15160 17604
rect 17960 17620 18012 17672
rect 19064 17663 19116 17672
rect 19064 17629 19073 17663
rect 19073 17629 19107 17663
rect 19107 17629 19116 17663
rect 19064 17620 19116 17629
rect 19156 17620 19208 17672
rect 23388 17620 23440 17672
rect 17132 17484 17184 17536
rect 17316 17484 17368 17536
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 19616 17527 19668 17536
rect 19616 17493 19625 17527
rect 19625 17493 19659 17527
rect 19659 17493 19668 17527
rect 19616 17484 19668 17493
rect 9291 17382 9343 17434
rect 9355 17382 9407 17434
rect 9419 17382 9471 17434
rect 9483 17382 9535 17434
rect 9547 17382 9599 17434
rect 17632 17382 17684 17434
rect 17696 17382 17748 17434
rect 17760 17382 17812 17434
rect 17824 17382 17876 17434
rect 17888 17382 17940 17434
rect 3976 17280 4028 17332
rect 4160 17280 4212 17332
rect 2044 17212 2096 17264
rect 4068 17212 4120 17264
rect 9036 17280 9088 17332
rect 9680 17323 9732 17332
rect 9680 17289 9689 17323
rect 9689 17289 9723 17323
rect 9723 17289 9732 17323
rect 9680 17280 9732 17289
rect 9864 17323 9916 17332
rect 9864 17289 9873 17323
rect 9873 17289 9907 17323
rect 9907 17289 9916 17323
rect 9864 17280 9916 17289
rect 2964 17076 3016 17128
rect 5724 17144 5776 17196
rect 3424 17008 3476 17060
rect 4712 16940 4764 16992
rect 8852 17187 8904 17196
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 6276 16940 6328 16992
rect 8852 17153 8861 17187
rect 8861 17153 8895 17187
rect 8895 17153 8904 17187
rect 8852 17144 8904 17153
rect 9036 17187 9088 17196
rect 9036 17153 9045 17187
rect 9045 17153 9079 17187
rect 9079 17153 9088 17187
rect 9036 17144 9088 17153
rect 9312 17144 9364 17196
rect 9680 17144 9732 17196
rect 9956 17187 10008 17196
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 10048 17144 10100 17196
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 10784 17187 10836 17196
rect 10784 17153 10792 17187
rect 10792 17153 10826 17187
rect 10826 17153 10836 17187
rect 10784 17144 10836 17153
rect 13268 17280 13320 17332
rect 15936 17280 15988 17332
rect 18052 17323 18104 17332
rect 18052 17289 18061 17323
rect 18061 17289 18095 17323
rect 18095 17289 18104 17323
rect 18052 17280 18104 17289
rect 19156 17280 19208 17332
rect 19616 17280 19668 17332
rect 20904 17280 20956 17332
rect 12532 17212 12584 17264
rect 14004 17212 14056 17264
rect 18236 17255 18288 17264
rect 18236 17221 18245 17255
rect 18245 17221 18279 17255
rect 18279 17221 18288 17255
rect 18236 17212 18288 17221
rect 19432 17212 19484 17264
rect 21548 17212 21600 17264
rect 11244 17144 11296 17196
rect 16764 17144 16816 17196
rect 17408 17144 17460 17196
rect 18512 17187 18564 17196
rect 18512 17153 18521 17187
rect 18521 17153 18555 17187
rect 18555 17153 18564 17187
rect 18512 17144 18564 17153
rect 19708 17144 19760 17196
rect 19800 17144 19852 17196
rect 22192 17144 22244 17196
rect 24216 17187 24268 17196
rect 24216 17153 24225 17187
rect 24225 17153 24259 17187
rect 24259 17153 24268 17187
rect 24216 17144 24268 17153
rect 10968 17119 11020 17128
rect 10968 17085 10977 17119
rect 10977 17085 11011 17119
rect 11011 17085 11020 17119
rect 10968 17076 11020 17085
rect 11520 17119 11572 17128
rect 11520 17085 11529 17119
rect 11529 17085 11563 17119
rect 11563 17085 11572 17119
rect 11520 17076 11572 17085
rect 16672 17119 16724 17128
rect 16672 17085 16681 17119
rect 16681 17085 16715 17119
rect 16715 17085 16724 17119
rect 16672 17076 16724 17085
rect 18144 17076 18196 17128
rect 19432 17119 19484 17128
rect 7840 17008 7892 17060
rect 19432 17085 19441 17119
rect 19441 17085 19475 17119
rect 19475 17085 19484 17119
rect 19432 17076 19484 17085
rect 19524 17119 19576 17128
rect 19524 17085 19533 17119
rect 19533 17085 19567 17119
rect 19567 17085 19576 17119
rect 19524 17076 19576 17085
rect 25412 17008 25464 17060
rect 7564 16940 7616 16992
rect 9036 16940 9088 16992
rect 10048 16940 10100 16992
rect 14280 16940 14332 16992
rect 19800 16940 19852 16992
rect 20720 16940 20772 16992
rect 21732 16940 21784 16992
rect 23204 16940 23256 16992
rect 24492 16983 24544 16992
rect 24492 16949 24501 16983
rect 24501 16949 24535 16983
rect 24535 16949 24544 16983
rect 24492 16940 24544 16949
rect 5120 16838 5172 16890
rect 5184 16838 5236 16890
rect 5248 16838 5300 16890
rect 5312 16838 5364 16890
rect 5376 16838 5428 16890
rect 13462 16838 13514 16890
rect 13526 16838 13578 16890
rect 13590 16838 13642 16890
rect 13654 16838 13706 16890
rect 13718 16838 13770 16890
rect 21803 16838 21855 16890
rect 21867 16838 21919 16890
rect 21931 16838 21983 16890
rect 21995 16838 22047 16890
rect 22059 16838 22111 16890
rect 3424 16736 3476 16788
rect 2044 16600 2096 16652
rect 5632 16736 5684 16788
rect 8852 16736 8904 16788
rect 9312 16736 9364 16788
rect 10140 16736 10192 16788
rect 10784 16736 10836 16788
rect 2872 16532 2924 16584
rect 2964 16532 3016 16584
rect 14556 16736 14608 16788
rect 16764 16779 16816 16788
rect 16764 16745 16773 16779
rect 16773 16745 16807 16779
rect 16807 16745 16816 16779
rect 16764 16736 16816 16745
rect 17040 16736 17092 16788
rect 17224 16668 17276 16720
rect 18512 16736 18564 16788
rect 19248 16736 19300 16788
rect 14556 16643 14608 16652
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 4068 16532 4120 16584
rect 3792 16464 3844 16516
rect 4436 16532 4488 16584
rect 4896 16575 4948 16584
rect 4896 16541 4930 16575
rect 4930 16541 4948 16575
rect 4896 16532 4948 16541
rect 7840 16532 7892 16584
rect 14556 16609 14565 16643
rect 14565 16609 14599 16643
rect 14599 16609 14608 16643
rect 14556 16600 14608 16609
rect 9036 16532 9088 16584
rect 10416 16532 10468 16584
rect 11704 16532 11756 16584
rect 15844 16532 15896 16584
rect 4804 16464 4856 16516
rect 8024 16464 8076 16516
rect 8392 16507 8444 16516
rect 8392 16473 8401 16507
rect 8401 16473 8435 16507
rect 8435 16473 8444 16507
rect 8392 16464 8444 16473
rect 8484 16464 8536 16516
rect 11796 16464 11848 16516
rect 13084 16464 13136 16516
rect 14832 16507 14884 16516
rect 14832 16473 14866 16507
rect 14866 16473 14884 16507
rect 14832 16464 14884 16473
rect 15292 16464 15344 16516
rect 16028 16464 16080 16516
rect 17316 16643 17368 16652
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 16396 16575 16448 16584
rect 16396 16541 16405 16575
rect 16405 16541 16439 16575
rect 16439 16541 16448 16575
rect 16396 16532 16448 16541
rect 17408 16575 17460 16584
rect 3700 16396 3752 16448
rect 4620 16396 4672 16448
rect 6092 16396 6144 16448
rect 6828 16396 6880 16448
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 10140 16396 10192 16448
rect 14372 16396 14424 16448
rect 14740 16396 14792 16448
rect 17408 16541 17417 16575
rect 17417 16541 17451 16575
rect 17451 16541 17460 16575
rect 17408 16532 17460 16541
rect 18144 16668 18196 16720
rect 19340 16668 19392 16720
rect 19616 16779 19668 16788
rect 19616 16745 19625 16779
rect 19625 16745 19659 16779
rect 19659 16745 19668 16779
rect 25596 16779 25648 16788
rect 19616 16736 19668 16745
rect 25596 16745 25605 16779
rect 25605 16745 25639 16779
rect 25639 16745 25648 16779
rect 25596 16736 25648 16745
rect 17960 16600 18012 16652
rect 18236 16600 18288 16652
rect 18512 16600 18564 16652
rect 19708 16600 19760 16652
rect 19524 16532 19576 16584
rect 19800 16575 19852 16584
rect 19800 16541 19809 16575
rect 19809 16541 19843 16575
rect 19843 16541 19852 16575
rect 19800 16532 19852 16541
rect 20720 16575 20772 16584
rect 20720 16541 20729 16575
rect 20729 16541 20763 16575
rect 20763 16541 20772 16575
rect 20720 16532 20772 16541
rect 21548 16643 21600 16652
rect 21548 16609 21557 16643
rect 21557 16609 21591 16643
rect 21591 16609 21600 16643
rect 21548 16600 21600 16609
rect 23204 16643 23256 16652
rect 21732 16532 21784 16584
rect 23204 16609 23213 16643
rect 23213 16609 23247 16643
rect 23247 16609 23256 16643
rect 23204 16600 23256 16609
rect 24492 16643 24544 16652
rect 24492 16609 24501 16643
rect 24501 16609 24535 16643
rect 24535 16609 24544 16643
rect 24492 16600 24544 16609
rect 24676 16643 24728 16652
rect 24676 16609 24685 16643
rect 24685 16609 24719 16643
rect 24719 16609 24728 16643
rect 24676 16600 24728 16609
rect 18052 16464 18104 16516
rect 22100 16507 22152 16516
rect 22100 16473 22109 16507
rect 22109 16473 22143 16507
rect 22143 16473 22152 16507
rect 22836 16532 22888 16584
rect 22100 16464 22152 16473
rect 22928 16464 22980 16516
rect 23664 16464 23716 16516
rect 24952 16464 25004 16516
rect 18328 16396 18380 16448
rect 19432 16396 19484 16448
rect 19892 16439 19944 16448
rect 19892 16405 19901 16439
rect 19901 16405 19935 16439
rect 19935 16405 19944 16439
rect 19892 16396 19944 16405
rect 20260 16439 20312 16448
rect 20260 16405 20269 16439
rect 20269 16405 20303 16439
rect 20303 16405 20312 16439
rect 20260 16396 20312 16405
rect 21180 16396 21232 16448
rect 22560 16439 22612 16448
rect 22560 16405 22569 16439
rect 22569 16405 22603 16439
rect 22603 16405 22612 16439
rect 22560 16396 22612 16405
rect 22652 16439 22704 16448
rect 22652 16405 22661 16439
rect 22661 16405 22695 16439
rect 22695 16405 22704 16439
rect 23020 16439 23072 16448
rect 22652 16396 22704 16405
rect 23020 16405 23029 16439
rect 23029 16405 23063 16439
rect 23063 16405 23072 16439
rect 23020 16396 23072 16405
rect 23756 16396 23808 16448
rect 24584 16396 24636 16448
rect 24860 16396 24912 16448
rect 25136 16439 25188 16448
rect 25136 16405 25145 16439
rect 25145 16405 25179 16439
rect 25179 16405 25188 16439
rect 25136 16396 25188 16405
rect 9291 16294 9343 16346
rect 9355 16294 9407 16346
rect 9419 16294 9471 16346
rect 9483 16294 9535 16346
rect 9547 16294 9599 16346
rect 17632 16294 17684 16346
rect 17696 16294 17748 16346
rect 17760 16294 17812 16346
rect 17824 16294 17876 16346
rect 17888 16294 17940 16346
rect 3240 16192 3292 16244
rect 4068 16192 4120 16244
rect 8300 16192 8352 16244
rect 2780 16124 2832 16176
rect 9956 16235 10008 16244
rect 9956 16201 9965 16235
rect 9965 16201 9999 16235
rect 9999 16201 10008 16235
rect 9956 16192 10008 16201
rect 3332 16124 3384 16176
rect 8024 16124 8076 16176
rect 9312 16124 9364 16176
rect 9404 16124 9456 16176
rect 13084 16235 13136 16244
rect 13084 16201 13093 16235
rect 13093 16201 13127 16235
rect 13127 16201 13136 16235
rect 13084 16192 13136 16201
rect 14004 16235 14056 16244
rect 14004 16201 14013 16235
rect 14013 16201 14047 16235
rect 14047 16201 14056 16235
rect 14004 16192 14056 16201
rect 14832 16235 14884 16244
rect 14832 16201 14841 16235
rect 14841 16201 14875 16235
rect 14875 16201 14884 16235
rect 14832 16192 14884 16201
rect 19248 16192 19300 16244
rect 4620 16056 4672 16108
rect 8116 16099 8168 16108
rect 8116 16065 8150 16099
rect 8150 16065 8168 16099
rect 8116 16056 8168 16065
rect 9588 16099 9640 16108
rect 9588 16065 9597 16099
rect 9597 16065 9631 16099
rect 9631 16065 9640 16099
rect 9588 16056 9640 16065
rect 10232 16099 10284 16108
rect 3792 15988 3844 16040
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 12348 16124 12400 16176
rect 13820 16124 13872 16176
rect 14096 16124 14148 16176
rect 12532 16056 12584 16108
rect 12900 16056 12952 16108
rect 14188 16099 14240 16108
rect 12716 16031 12768 16040
rect 3884 15920 3936 15972
rect 9312 15920 9364 15972
rect 12716 15997 12725 16031
rect 12725 15997 12759 16031
rect 12759 15997 12768 16031
rect 12716 15988 12768 15997
rect 3516 15852 3568 15904
rect 7380 15852 7432 15904
rect 8760 15852 8812 15904
rect 12440 15920 12492 15972
rect 13176 15988 13228 16040
rect 10876 15852 10928 15904
rect 12348 15852 12400 15904
rect 12624 15852 12676 15904
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 14004 15988 14056 16040
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 14740 16099 14792 16108
rect 14740 16065 14749 16099
rect 14749 16065 14783 16099
rect 14783 16065 14792 16099
rect 14740 16056 14792 16065
rect 14648 15988 14700 16040
rect 15936 16099 15988 16108
rect 15936 16065 15945 16099
rect 15945 16065 15979 16099
rect 15979 16065 15988 16099
rect 15936 16056 15988 16065
rect 16028 16031 16080 16040
rect 16028 15997 16037 16031
rect 16037 15997 16071 16031
rect 16071 15997 16080 16031
rect 16028 15988 16080 15997
rect 16396 15988 16448 16040
rect 16672 16031 16724 16040
rect 16672 15997 16681 16031
rect 16681 15997 16715 16031
rect 16715 15997 16724 16031
rect 16672 15988 16724 15997
rect 15844 15920 15896 15972
rect 14372 15852 14424 15904
rect 20812 16192 20864 16244
rect 21180 16235 21232 16244
rect 21180 16201 21189 16235
rect 21189 16201 21223 16235
rect 21223 16201 21232 16235
rect 21180 16192 21232 16201
rect 21272 16235 21324 16244
rect 21272 16201 21281 16235
rect 21281 16201 21315 16235
rect 21315 16201 21324 16235
rect 21272 16192 21324 16201
rect 21456 16192 21508 16244
rect 22836 16192 22888 16244
rect 23020 16192 23072 16244
rect 23848 16192 23900 16244
rect 24860 16235 24912 16244
rect 24860 16201 24869 16235
rect 24869 16201 24903 16235
rect 24903 16201 24912 16235
rect 24860 16192 24912 16201
rect 24952 16235 25004 16244
rect 24952 16201 24961 16235
rect 24961 16201 24995 16235
rect 24995 16201 25004 16235
rect 25412 16235 25464 16244
rect 24952 16192 25004 16201
rect 25412 16201 25421 16235
rect 25421 16201 25455 16235
rect 25455 16201 25464 16235
rect 25412 16192 25464 16201
rect 20904 16124 20956 16176
rect 24124 16124 24176 16176
rect 21088 16056 21140 16108
rect 21640 16056 21692 16108
rect 24308 16056 24360 16108
rect 22560 16031 22612 16040
rect 18972 15852 19024 15904
rect 20996 15920 21048 15972
rect 22560 15997 22569 16031
rect 22569 15997 22603 16031
rect 22603 15997 22612 16031
rect 22560 15988 22612 15997
rect 22744 16031 22796 16040
rect 22744 15997 22753 16031
rect 22753 15997 22787 16031
rect 22787 15997 22796 16031
rect 22744 15988 22796 15997
rect 23204 15988 23256 16040
rect 23480 15988 23532 16040
rect 25228 15988 25280 16040
rect 23756 15920 23808 15972
rect 25504 16031 25556 16040
rect 25504 15997 25513 16031
rect 25513 15997 25547 16031
rect 25547 15997 25556 16031
rect 25504 15988 25556 15997
rect 22652 15852 22704 15904
rect 23664 15852 23716 15904
rect 5120 15750 5172 15802
rect 5184 15750 5236 15802
rect 5248 15750 5300 15802
rect 5312 15750 5364 15802
rect 5376 15750 5428 15802
rect 13462 15750 13514 15802
rect 13526 15750 13578 15802
rect 13590 15750 13642 15802
rect 13654 15750 13706 15802
rect 13718 15750 13770 15802
rect 21803 15750 21855 15802
rect 21867 15750 21919 15802
rect 21931 15750 21983 15802
rect 21995 15750 22047 15802
rect 22059 15750 22111 15802
rect 3792 15512 3844 15564
rect 3056 15444 3108 15496
rect 3240 15487 3292 15496
rect 3240 15453 3249 15487
rect 3249 15453 3283 15487
rect 3283 15453 3292 15487
rect 3240 15444 3292 15453
rect 2780 15419 2832 15428
rect 2780 15385 2789 15419
rect 2789 15385 2823 15419
rect 2823 15385 2832 15419
rect 3516 15487 3568 15496
rect 3516 15453 3525 15487
rect 3525 15453 3559 15487
rect 3559 15453 3568 15487
rect 4804 15648 4856 15700
rect 6552 15648 6604 15700
rect 8484 15648 8536 15700
rect 9036 15648 9088 15700
rect 10324 15648 10376 15700
rect 10508 15648 10560 15700
rect 12348 15691 12400 15700
rect 7840 15580 7892 15632
rect 5632 15555 5684 15564
rect 5632 15521 5641 15555
rect 5641 15521 5675 15555
rect 5675 15521 5684 15555
rect 5632 15512 5684 15521
rect 8116 15512 8168 15564
rect 11612 15580 11664 15632
rect 3516 15444 3568 15453
rect 4068 15444 4120 15496
rect 2780 15376 2832 15385
rect 4252 15376 4304 15428
rect 6276 15376 6328 15428
rect 8024 15444 8076 15496
rect 8484 15487 8536 15496
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 7288 15308 7340 15360
rect 7932 15308 7984 15360
rect 8484 15308 8536 15360
rect 9404 15444 9456 15496
rect 12348 15657 12357 15691
rect 12357 15657 12391 15691
rect 12391 15657 12400 15691
rect 12348 15648 12400 15657
rect 14464 15648 14516 15700
rect 16028 15648 16080 15700
rect 19248 15648 19300 15700
rect 19984 15691 20036 15700
rect 19984 15657 19993 15691
rect 19993 15657 20027 15691
rect 20027 15657 20036 15691
rect 19984 15648 20036 15657
rect 20260 15648 20312 15700
rect 21088 15648 21140 15700
rect 22744 15648 22796 15700
rect 22928 15691 22980 15700
rect 22928 15657 22937 15691
rect 22937 15657 22971 15691
rect 22971 15657 22980 15691
rect 22928 15648 22980 15657
rect 24216 15648 24268 15700
rect 24308 15648 24360 15700
rect 25228 15691 25280 15700
rect 25228 15657 25237 15691
rect 25237 15657 25271 15691
rect 25271 15657 25280 15691
rect 25228 15648 25280 15657
rect 15936 15580 15988 15632
rect 12440 15512 12492 15564
rect 11152 15444 11204 15496
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 13268 15512 13320 15564
rect 9772 15376 9824 15428
rect 10600 15376 10652 15428
rect 11060 15376 11112 15428
rect 11520 15351 11572 15360
rect 11520 15317 11529 15351
rect 11529 15317 11563 15351
rect 11563 15317 11572 15351
rect 12440 15376 12492 15428
rect 13636 15487 13688 15496
rect 13636 15453 13645 15487
rect 13645 15453 13679 15487
rect 13679 15453 13688 15487
rect 13636 15444 13688 15453
rect 21456 15580 21508 15632
rect 24768 15580 24820 15632
rect 25504 15623 25556 15632
rect 19248 15512 19300 15564
rect 20536 15512 20588 15564
rect 20720 15512 20772 15564
rect 21548 15512 21600 15564
rect 22560 15512 22612 15564
rect 23480 15555 23532 15564
rect 23480 15521 23489 15555
rect 23489 15521 23523 15555
rect 23523 15521 23532 15555
rect 23480 15512 23532 15521
rect 23756 15555 23808 15564
rect 23756 15521 23765 15555
rect 23765 15521 23799 15555
rect 23799 15521 23808 15555
rect 23756 15512 23808 15521
rect 25504 15589 25513 15623
rect 25513 15589 25547 15623
rect 25547 15589 25556 15623
rect 25504 15580 25556 15589
rect 18696 15487 18748 15496
rect 18696 15453 18705 15487
rect 18705 15453 18739 15487
rect 18739 15453 18748 15487
rect 18696 15444 18748 15453
rect 20168 15487 20220 15496
rect 20168 15453 20177 15487
rect 20177 15453 20211 15487
rect 20211 15453 20220 15487
rect 20168 15444 20220 15453
rect 20996 15444 21048 15496
rect 22652 15487 22704 15496
rect 22652 15453 22661 15487
rect 22661 15453 22695 15487
rect 22695 15453 22704 15487
rect 22652 15444 22704 15453
rect 23664 15444 23716 15496
rect 24032 15444 24084 15496
rect 24584 15444 24636 15496
rect 25412 15487 25464 15496
rect 25412 15453 25421 15487
rect 25421 15453 25455 15487
rect 25455 15453 25464 15487
rect 25412 15444 25464 15453
rect 18236 15419 18288 15428
rect 18236 15385 18245 15419
rect 18245 15385 18279 15419
rect 18279 15385 18288 15419
rect 18236 15376 18288 15385
rect 18328 15376 18380 15428
rect 18604 15419 18656 15428
rect 18604 15385 18613 15419
rect 18613 15385 18647 15419
rect 18647 15385 18656 15419
rect 18604 15376 18656 15385
rect 11520 15308 11572 15317
rect 15200 15308 15252 15360
rect 18512 15308 18564 15360
rect 19616 15351 19668 15360
rect 19616 15317 19625 15351
rect 19625 15317 19659 15351
rect 19659 15317 19668 15351
rect 19616 15308 19668 15317
rect 20536 15308 20588 15360
rect 23388 15351 23440 15360
rect 23388 15317 23397 15351
rect 23397 15317 23431 15351
rect 23431 15317 23440 15351
rect 24216 15376 24268 15428
rect 23388 15308 23440 15317
rect 24676 15308 24728 15360
rect 9291 15206 9343 15258
rect 9355 15206 9407 15258
rect 9419 15206 9471 15258
rect 9483 15206 9535 15258
rect 9547 15206 9599 15258
rect 17632 15206 17684 15258
rect 17696 15206 17748 15258
rect 17760 15206 17812 15258
rect 17824 15206 17876 15258
rect 17888 15206 17940 15258
rect 3056 15104 3108 15156
rect 4252 15147 4304 15156
rect 4252 15113 4261 15147
rect 4261 15113 4295 15147
rect 4295 15113 4304 15147
rect 4252 15104 4304 15113
rect 4712 15147 4764 15156
rect 4712 15113 4721 15147
rect 4721 15113 4755 15147
rect 4755 15113 4764 15147
rect 4712 15104 4764 15113
rect 2780 15036 2832 15088
rect 8668 15104 8720 15156
rect 10600 15147 10652 15156
rect 10600 15113 10609 15147
rect 10609 15113 10643 15147
rect 10643 15113 10652 15147
rect 10600 15104 10652 15113
rect 14188 15104 14240 15156
rect 16120 15104 16172 15156
rect 18144 15104 18196 15156
rect 18788 15147 18840 15156
rect 18788 15113 18797 15147
rect 18797 15113 18831 15147
rect 18831 15113 18840 15147
rect 18788 15104 18840 15113
rect 19616 15104 19668 15156
rect 20168 15104 20220 15156
rect 20628 15104 20680 15156
rect 21272 15147 21324 15156
rect 21272 15113 21281 15147
rect 21281 15113 21315 15147
rect 21315 15113 21324 15147
rect 21272 15104 21324 15113
rect 23388 15104 23440 15156
rect 25412 15104 25464 15156
rect 2964 15011 3016 15020
rect 2964 14977 2973 15011
rect 2973 14977 3007 15011
rect 3007 14977 3016 15011
rect 2964 14968 3016 14977
rect 2688 14764 2740 14816
rect 3516 14968 3568 15020
rect 3608 15011 3660 15020
rect 3608 14977 3616 15011
rect 3616 14977 3650 15011
rect 3650 14977 3660 15011
rect 3608 14968 3660 14977
rect 4620 15011 4672 15020
rect 3240 14900 3292 14952
rect 3792 14943 3844 14952
rect 3792 14909 3801 14943
rect 3801 14909 3835 14943
rect 3835 14909 3844 14943
rect 3792 14900 3844 14909
rect 4620 14977 4629 15011
rect 4629 14977 4663 15011
rect 4663 14977 4672 15011
rect 4620 14968 4672 14977
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 7840 15036 7892 15088
rect 6920 15011 6972 15020
rect 6920 14977 6954 15011
rect 6954 14977 6972 15011
rect 6920 14968 6972 14977
rect 8576 14968 8628 15020
rect 10232 15036 10284 15088
rect 12992 15036 13044 15088
rect 19984 15036 20036 15088
rect 24768 15079 24820 15088
rect 24768 15045 24777 15079
rect 24777 15045 24811 15079
rect 24811 15045 24820 15079
rect 24768 15036 24820 15045
rect 9128 14968 9180 15020
rect 10140 15011 10192 15020
rect 10140 14977 10148 15011
rect 10148 14977 10182 15011
rect 10182 14977 10192 15011
rect 10140 14968 10192 14977
rect 10324 15011 10376 15020
rect 10324 14977 10333 15011
rect 10333 14977 10367 15011
rect 10367 14977 10376 15011
rect 10324 14968 10376 14977
rect 11520 14968 11572 15020
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 12900 14968 12952 14977
rect 13820 14968 13872 15020
rect 15108 14968 15160 15020
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 16764 14968 16816 15020
rect 4528 14900 4580 14952
rect 10876 14900 10928 14952
rect 14556 14900 14608 14952
rect 18144 14900 18196 14952
rect 19064 14900 19116 14952
rect 19524 15011 19576 15020
rect 19524 14977 19533 15011
rect 19533 14977 19567 15011
rect 19567 14977 19576 15011
rect 19524 14968 19576 14977
rect 20536 14968 20588 15020
rect 20812 15011 20864 15020
rect 20812 14977 20821 15011
rect 20821 14977 20855 15011
rect 20855 14977 20864 15011
rect 20812 14968 20864 14977
rect 21088 15011 21140 15020
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 23296 15011 23348 15020
rect 20720 14900 20772 14952
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 23664 14968 23716 15020
rect 23756 14968 23808 15020
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 5540 14832 5592 14884
rect 14740 14875 14792 14884
rect 4068 14807 4120 14816
rect 4068 14773 4077 14807
rect 4077 14773 4111 14807
rect 4111 14773 4120 14807
rect 4068 14764 4120 14773
rect 6552 14764 6604 14816
rect 14740 14841 14749 14875
rect 14749 14841 14783 14875
rect 14783 14841 14792 14875
rect 14740 14832 14792 14841
rect 8024 14807 8076 14816
rect 8024 14773 8033 14807
rect 8033 14773 8067 14807
rect 8067 14773 8076 14807
rect 8024 14764 8076 14773
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 11520 14764 11572 14816
rect 12900 14764 12952 14816
rect 14188 14807 14240 14816
rect 14188 14773 14197 14807
rect 14197 14773 14231 14807
rect 14231 14773 14240 14807
rect 14188 14764 14240 14773
rect 14924 14764 14976 14816
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 19524 14832 19576 14884
rect 16396 14764 16448 14773
rect 18144 14764 18196 14816
rect 19616 14807 19668 14816
rect 19616 14773 19625 14807
rect 19625 14773 19659 14807
rect 19659 14773 19668 14807
rect 19616 14764 19668 14773
rect 21088 14764 21140 14816
rect 23664 14807 23716 14816
rect 23664 14773 23673 14807
rect 23673 14773 23707 14807
rect 23707 14773 23716 14807
rect 23664 14764 23716 14773
rect 5120 14662 5172 14714
rect 5184 14662 5236 14714
rect 5248 14662 5300 14714
rect 5312 14662 5364 14714
rect 5376 14662 5428 14714
rect 13462 14662 13514 14714
rect 13526 14662 13578 14714
rect 13590 14662 13642 14714
rect 13654 14662 13706 14714
rect 13718 14662 13770 14714
rect 21803 14662 21855 14714
rect 21867 14662 21919 14714
rect 21931 14662 21983 14714
rect 21995 14662 22047 14714
rect 22059 14662 22111 14714
rect 2412 14560 2464 14612
rect 3056 14467 3108 14476
rect 5540 14560 5592 14612
rect 6092 14560 6144 14612
rect 6276 14603 6328 14612
rect 6276 14569 6285 14603
rect 6285 14569 6319 14603
rect 6319 14569 6328 14603
rect 6276 14560 6328 14569
rect 3056 14433 3070 14467
rect 3070 14433 3104 14467
rect 3104 14433 3108 14467
rect 3056 14424 3108 14433
rect 5908 14467 5960 14476
rect 5908 14433 5917 14467
rect 5917 14433 5951 14467
rect 5951 14433 5960 14467
rect 5908 14424 5960 14433
rect 2872 14356 2924 14408
rect 2964 14399 3016 14408
rect 2964 14365 2973 14399
rect 2973 14365 3007 14399
rect 3007 14365 3016 14399
rect 2964 14356 3016 14365
rect 3148 14399 3200 14408
rect 3148 14365 3158 14399
rect 3158 14365 3192 14399
rect 3192 14365 3200 14399
rect 3148 14356 3200 14365
rect 4068 14399 4120 14408
rect 4068 14365 4102 14399
rect 4102 14365 4120 14399
rect 4068 14356 4120 14365
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 3516 14288 3568 14340
rect 5908 14288 5960 14340
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 6644 14492 6696 14544
rect 7012 14560 7064 14612
rect 7288 14603 7340 14612
rect 7288 14569 7297 14603
rect 7297 14569 7331 14603
rect 7331 14569 7340 14603
rect 7288 14560 7340 14569
rect 7380 14560 7432 14612
rect 8116 14603 8168 14612
rect 8116 14569 8125 14603
rect 8125 14569 8159 14603
rect 8159 14569 8168 14603
rect 8116 14560 8168 14569
rect 8392 14560 8444 14612
rect 8668 14603 8720 14612
rect 8668 14569 8677 14603
rect 8677 14569 8711 14603
rect 8711 14569 8720 14603
rect 8668 14560 8720 14569
rect 6736 14467 6788 14476
rect 6736 14433 6745 14467
rect 6745 14433 6779 14467
rect 6779 14433 6788 14467
rect 6736 14424 6788 14433
rect 7196 14492 7248 14544
rect 7104 14424 7156 14476
rect 7840 14467 7892 14476
rect 7840 14433 7849 14467
rect 7849 14433 7883 14467
rect 7883 14433 7892 14467
rect 7840 14424 7892 14433
rect 8024 14356 8076 14408
rect 8116 14356 8168 14408
rect 8760 14399 8812 14408
rect 8760 14365 8763 14399
rect 8763 14365 8797 14399
rect 8797 14365 8812 14399
rect 11060 14560 11112 14612
rect 8760 14356 8812 14365
rect 7288 14288 7340 14340
rect 8208 14288 8260 14340
rect 11152 14424 11204 14476
rect 11980 14467 12032 14476
rect 11612 14399 11664 14408
rect 2688 14263 2740 14272
rect 2688 14229 2697 14263
rect 2697 14229 2731 14263
rect 2731 14229 2740 14263
rect 2688 14220 2740 14229
rect 3424 14220 3476 14272
rect 8668 14220 8720 14272
rect 8852 14220 8904 14272
rect 11612 14365 11621 14399
rect 11621 14365 11655 14399
rect 11655 14365 11664 14399
rect 11612 14356 11664 14365
rect 11980 14433 11989 14467
rect 11989 14433 12023 14467
rect 12023 14433 12032 14467
rect 11980 14424 12032 14433
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 13820 14560 13872 14612
rect 14280 14560 14332 14612
rect 15108 14560 15160 14612
rect 16028 14560 16080 14612
rect 14464 14467 14516 14476
rect 14464 14433 14473 14467
rect 14473 14433 14507 14467
rect 14507 14433 14516 14467
rect 14464 14424 14516 14433
rect 14648 14424 14700 14476
rect 15936 14492 15988 14544
rect 15384 14467 15436 14476
rect 15384 14433 15393 14467
rect 15393 14433 15427 14467
rect 15427 14433 15436 14467
rect 15384 14424 15436 14433
rect 15660 14424 15712 14476
rect 16764 14560 16816 14612
rect 19432 14560 19484 14612
rect 21088 14560 21140 14612
rect 18696 14535 18748 14544
rect 18696 14501 18705 14535
rect 18705 14501 18739 14535
rect 18739 14501 18748 14535
rect 18696 14492 18748 14501
rect 20812 14492 20864 14544
rect 23296 14492 23348 14544
rect 18328 14424 18380 14476
rect 19616 14467 19668 14476
rect 19616 14433 19625 14467
rect 19625 14433 19659 14467
rect 19659 14433 19668 14467
rect 19616 14424 19668 14433
rect 20260 14424 20312 14476
rect 23020 14424 23072 14476
rect 23664 14424 23716 14476
rect 24216 14467 24268 14476
rect 11888 14356 11940 14365
rect 13084 14356 13136 14408
rect 10784 14220 10836 14272
rect 14096 14356 14148 14408
rect 14280 14356 14332 14408
rect 14924 14356 14976 14408
rect 15200 14399 15252 14408
rect 15200 14365 15208 14399
rect 15208 14365 15242 14399
rect 15242 14365 15252 14399
rect 15568 14399 15620 14408
rect 15200 14356 15252 14365
rect 15568 14365 15577 14399
rect 15577 14365 15611 14399
rect 15611 14365 15620 14399
rect 15568 14356 15620 14365
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 15936 14288 15988 14340
rect 17960 14356 18012 14408
rect 16488 14288 16540 14340
rect 18236 14356 18288 14408
rect 20076 14399 20128 14408
rect 20076 14365 20085 14399
rect 20085 14365 20119 14399
rect 20119 14365 20128 14399
rect 20076 14356 20128 14365
rect 20444 14399 20496 14408
rect 20444 14365 20453 14399
rect 20453 14365 20487 14399
rect 20487 14365 20496 14399
rect 20444 14356 20496 14365
rect 18604 14288 18656 14340
rect 19248 14288 19300 14340
rect 19708 14288 19760 14340
rect 23572 14399 23624 14408
rect 23572 14365 23581 14399
rect 23581 14365 23615 14399
rect 23615 14365 23624 14399
rect 24216 14433 24225 14467
rect 24225 14433 24259 14467
rect 24259 14433 24268 14467
rect 24216 14424 24268 14433
rect 23572 14356 23624 14365
rect 24308 14356 24360 14408
rect 23756 14288 23808 14340
rect 14004 14220 14056 14272
rect 14280 14220 14332 14272
rect 15016 14220 15068 14272
rect 17408 14220 17460 14272
rect 20812 14220 20864 14272
rect 21180 14220 21232 14272
rect 23204 14220 23256 14272
rect 24676 14220 24728 14272
rect 9291 14118 9343 14170
rect 9355 14118 9407 14170
rect 9419 14118 9471 14170
rect 9483 14118 9535 14170
rect 9547 14118 9599 14170
rect 17632 14118 17684 14170
rect 17696 14118 17748 14170
rect 17760 14118 17812 14170
rect 17824 14118 17876 14170
rect 17888 14118 17940 14170
rect 2964 14016 3016 14068
rect 3608 14016 3660 14068
rect 3792 14016 3844 14068
rect 5632 14016 5684 14068
rect 5908 14059 5960 14068
rect 5908 14025 5917 14059
rect 5917 14025 5951 14059
rect 5951 14025 5960 14059
rect 5908 14016 5960 14025
rect 6000 14016 6052 14068
rect 6828 14059 6880 14068
rect 6828 14025 6837 14059
rect 6837 14025 6871 14059
rect 6871 14025 6880 14059
rect 6828 14016 6880 14025
rect 7656 14059 7708 14068
rect 7656 14025 7665 14059
rect 7665 14025 7699 14059
rect 7699 14025 7708 14059
rect 7656 14016 7708 14025
rect 8116 14059 8168 14068
rect 8116 14025 8125 14059
rect 8125 14025 8159 14059
rect 8159 14025 8168 14059
rect 8116 14016 8168 14025
rect 11152 14059 11204 14068
rect 11152 14025 11161 14059
rect 11161 14025 11195 14059
rect 11195 14025 11204 14059
rect 11152 14016 11204 14025
rect 11612 14016 11664 14068
rect 11888 14016 11940 14068
rect 12256 14016 12308 14068
rect 12992 14016 13044 14068
rect 15200 14016 15252 14068
rect 15844 14016 15896 14068
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 4896 13948 4948 14000
rect 3332 13923 3384 13932
rect 3332 13889 3342 13923
rect 3342 13889 3376 13923
rect 3376 13889 3384 13923
rect 3332 13880 3384 13889
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 3700 13880 3752 13932
rect 4712 13923 4764 13932
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 5724 13923 5776 13958
rect 5724 13906 5725 13923
rect 5725 13906 5759 13923
rect 5759 13906 5776 13923
rect 8392 13948 8444 14000
rect 9220 13948 9272 14000
rect 3056 13812 3108 13864
rect 4344 13855 4396 13864
rect 4344 13821 4353 13855
rect 4353 13821 4387 13855
rect 4387 13821 4396 13855
rect 4344 13812 4396 13821
rect 4528 13812 4580 13864
rect 2780 13787 2832 13796
rect 2780 13753 2789 13787
rect 2789 13753 2823 13787
rect 2823 13753 2832 13787
rect 2780 13744 2832 13753
rect 4160 13744 4212 13796
rect 5448 13744 5500 13796
rect 6552 13880 6604 13932
rect 7288 13880 7340 13932
rect 8300 13880 8352 13932
rect 8668 13923 8720 13932
rect 8668 13889 8677 13923
rect 8677 13889 8711 13923
rect 8711 13889 8720 13923
rect 8668 13880 8720 13889
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 7656 13812 7708 13864
rect 7840 13812 7892 13864
rect 8852 13880 8904 13932
rect 9680 13948 9732 14000
rect 14096 13948 14148 14000
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 8944 13812 8996 13821
rect 9956 13880 10008 13932
rect 11796 13923 11848 13932
rect 11796 13889 11830 13923
rect 11830 13889 11848 13923
rect 13084 13923 13136 13932
rect 11796 13880 11848 13889
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 13176 13880 13228 13932
rect 14740 13880 14792 13932
rect 15660 13948 15712 14000
rect 16488 14016 16540 14068
rect 17224 14016 17276 14068
rect 18328 14016 18380 14068
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 19248 14016 19300 14068
rect 20076 14016 20128 14068
rect 23296 14059 23348 14068
rect 23296 14025 23305 14059
rect 23305 14025 23339 14059
rect 23339 14025 23348 14059
rect 23296 14016 23348 14025
rect 24584 14016 24636 14068
rect 15568 13880 15620 13932
rect 17592 13880 17644 13932
rect 18420 13880 18472 13932
rect 19064 13923 19116 13932
rect 19064 13889 19073 13923
rect 19073 13889 19107 13923
rect 19107 13889 19116 13923
rect 19064 13880 19116 13889
rect 19432 13923 19484 13932
rect 19432 13889 19441 13923
rect 19441 13889 19475 13923
rect 19475 13889 19484 13923
rect 19432 13880 19484 13889
rect 11520 13855 11572 13864
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 9312 13744 9364 13796
rect 9588 13744 9640 13796
rect 6184 13719 6236 13728
rect 6184 13685 6193 13719
rect 6193 13685 6227 13719
rect 6227 13685 6236 13719
rect 6184 13676 6236 13685
rect 6920 13676 6972 13728
rect 9956 13719 10008 13728
rect 9956 13685 9965 13719
rect 9965 13685 9999 13719
rect 9999 13685 10008 13719
rect 9956 13676 10008 13685
rect 14004 13676 14056 13728
rect 14556 13676 14608 13728
rect 17408 13812 17460 13864
rect 19984 13948 20036 14000
rect 19616 13880 19668 13932
rect 20352 13923 20404 13932
rect 20352 13889 20361 13923
rect 20361 13889 20395 13923
rect 20395 13889 20404 13923
rect 20352 13880 20404 13889
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20812 13923 20864 13932
rect 20444 13880 20496 13889
rect 20812 13889 20821 13923
rect 20821 13889 20855 13923
rect 20855 13889 20864 13923
rect 20812 13880 20864 13889
rect 21180 13880 21232 13932
rect 21364 13880 21416 13932
rect 23204 13923 23256 13932
rect 23204 13889 23213 13923
rect 23213 13889 23247 13923
rect 23247 13889 23256 13923
rect 23204 13880 23256 13889
rect 23664 13948 23716 14000
rect 23572 13923 23624 13932
rect 23572 13889 23581 13923
rect 23581 13889 23615 13923
rect 23615 13889 23624 13923
rect 23572 13880 23624 13889
rect 23848 13880 23900 13932
rect 24308 13923 24360 13932
rect 24308 13889 24317 13923
rect 24317 13889 24351 13923
rect 24351 13889 24360 13923
rect 24308 13880 24360 13889
rect 17224 13787 17276 13796
rect 17224 13753 17233 13787
rect 17233 13753 17267 13787
rect 17267 13753 17276 13787
rect 17224 13744 17276 13753
rect 17316 13719 17368 13728
rect 17316 13685 17325 13719
rect 17325 13685 17359 13719
rect 17359 13685 17368 13719
rect 17316 13676 17368 13685
rect 18144 13719 18196 13728
rect 18144 13685 18153 13719
rect 18153 13685 18187 13719
rect 18187 13685 18196 13719
rect 18144 13676 18196 13685
rect 23756 13855 23808 13864
rect 23756 13821 23765 13855
rect 23765 13821 23799 13855
rect 23799 13821 23808 13855
rect 23756 13812 23808 13821
rect 21456 13787 21508 13796
rect 21456 13753 21465 13787
rect 21465 13753 21499 13787
rect 21499 13753 21508 13787
rect 21456 13744 21508 13753
rect 22192 13787 22244 13796
rect 22192 13753 22201 13787
rect 22201 13753 22235 13787
rect 22235 13753 22244 13787
rect 22192 13744 22244 13753
rect 23940 13787 23992 13796
rect 23940 13753 23949 13787
rect 23949 13753 23983 13787
rect 23983 13753 23992 13787
rect 23940 13744 23992 13753
rect 23572 13676 23624 13728
rect 24032 13676 24084 13728
rect 5120 13574 5172 13626
rect 5184 13574 5236 13626
rect 5248 13574 5300 13626
rect 5312 13574 5364 13626
rect 5376 13574 5428 13626
rect 13462 13574 13514 13626
rect 13526 13574 13578 13626
rect 13590 13574 13642 13626
rect 13654 13574 13706 13626
rect 13718 13574 13770 13626
rect 21803 13574 21855 13626
rect 21867 13574 21919 13626
rect 21931 13574 21983 13626
rect 21995 13574 22047 13626
rect 22059 13574 22111 13626
rect 3148 13472 3200 13524
rect 4160 13472 4212 13524
rect 6184 13472 6236 13524
rect 7104 13472 7156 13524
rect 8668 13472 8720 13524
rect 8852 13472 8904 13524
rect 3976 13336 4028 13388
rect 4344 13379 4396 13388
rect 4344 13345 4353 13379
rect 4353 13345 4387 13379
rect 4387 13345 4396 13379
rect 4344 13336 4396 13345
rect 1676 13268 1728 13320
rect 2412 13268 2464 13320
rect 4712 13268 4764 13320
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 2688 13243 2740 13252
rect 2688 13209 2706 13243
rect 2706 13209 2740 13243
rect 2688 13200 2740 13209
rect 7012 13404 7064 13456
rect 9036 13404 9088 13456
rect 9220 13404 9272 13456
rect 5908 13379 5960 13388
rect 5908 13345 5917 13379
rect 5917 13345 5951 13379
rect 5951 13345 5960 13379
rect 5908 13336 5960 13345
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 5816 13311 5868 13320
rect 5816 13277 5825 13311
rect 5825 13277 5859 13311
rect 5859 13277 5868 13311
rect 5816 13268 5868 13277
rect 6184 13311 6236 13320
rect 6184 13277 6193 13311
rect 6193 13277 6227 13311
rect 6227 13277 6236 13311
rect 7380 13336 7432 13388
rect 7656 13379 7708 13388
rect 7656 13345 7665 13379
rect 7665 13345 7699 13379
rect 7699 13345 7708 13379
rect 7656 13336 7708 13345
rect 11152 13472 11204 13524
rect 11060 13404 11112 13456
rect 10876 13379 10928 13388
rect 6184 13268 6236 13277
rect 6644 13311 6696 13320
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 6920 13268 6972 13320
rect 7104 13268 7156 13320
rect 7748 13268 7800 13320
rect 9036 13268 9088 13320
rect 10876 13345 10885 13379
rect 10885 13345 10919 13379
rect 10919 13345 10928 13379
rect 10876 13336 10928 13345
rect 2872 13132 2924 13184
rect 3976 13132 4028 13184
rect 5540 13175 5592 13184
rect 5540 13141 5549 13175
rect 5549 13141 5583 13175
rect 5583 13141 5592 13175
rect 5540 13132 5592 13141
rect 6460 13132 6512 13184
rect 8852 13200 8904 13252
rect 9404 13277 9450 13298
rect 9450 13277 9456 13298
rect 9404 13246 9456 13277
rect 9128 13132 9180 13184
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 9956 13268 10008 13320
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 11152 13268 11204 13320
rect 10140 13200 10192 13252
rect 10048 13175 10100 13184
rect 10048 13141 10057 13175
rect 10057 13141 10091 13175
rect 10091 13141 10100 13175
rect 10048 13132 10100 13141
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 10876 13200 10928 13252
rect 11796 13472 11848 13524
rect 14648 13515 14700 13524
rect 11796 13336 11848 13388
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 12256 13404 12308 13456
rect 12532 13404 12584 13456
rect 13176 13404 13228 13456
rect 11612 13268 11664 13277
rect 12624 13336 12676 13388
rect 14648 13481 14657 13515
rect 14657 13481 14691 13515
rect 14691 13481 14700 13515
rect 14648 13472 14700 13481
rect 17500 13472 17552 13524
rect 20352 13472 20404 13524
rect 21364 13472 21416 13524
rect 21548 13472 21600 13524
rect 23664 13472 23716 13524
rect 24124 13472 24176 13524
rect 14096 13447 14148 13456
rect 14096 13413 14105 13447
rect 14105 13413 14139 13447
rect 14139 13413 14148 13447
rect 14096 13404 14148 13413
rect 23388 13404 23440 13456
rect 17592 13379 17644 13388
rect 17592 13345 17601 13379
rect 17601 13345 17635 13379
rect 17635 13345 17644 13379
rect 17592 13336 17644 13345
rect 17684 13379 17736 13388
rect 17684 13345 17693 13379
rect 17693 13345 17727 13379
rect 17727 13345 17736 13379
rect 18420 13379 18472 13388
rect 17684 13336 17736 13345
rect 18420 13345 18429 13379
rect 18429 13345 18463 13379
rect 18463 13345 18472 13379
rect 18420 13336 18472 13345
rect 19340 13336 19392 13388
rect 20352 13336 20404 13388
rect 21456 13336 21508 13388
rect 13084 13268 13136 13320
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 14464 13311 14516 13320
rect 13544 13268 13596 13277
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 17316 13268 17368 13320
rect 18144 13268 18196 13320
rect 20444 13268 20496 13320
rect 21272 13268 21324 13320
rect 21916 13311 21968 13320
rect 14280 13243 14332 13252
rect 11336 13132 11388 13184
rect 11612 13132 11664 13184
rect 11796 13132 11848 13184
rect 12256 13132 12308 13184
rect 13636 13175 13688 13184
rect 13636 13141 13645 13175
rect 13645 13141 13679 13175
rect 13679 13141 13688 13175
rect 13636 13132 13688 13141
rect 14280 13209 14289 13243
rect 14289 13209 14323 13243
rect 14323 13209 14332 13243
rect 14280 13200 14332 13209
rect 14556 13200 14608 13252
rect 21916 13277 21925 13311
rect 21925 13277 21959 13311
rect 21959 13277 21968 13311
rect 23848 13336 23900 13388
rect 23940 13336 23992 13388
rect 21916 13268 21968 13277
rect 23664 13311 23716 13320
rect 22008 13243 22060 13252
rect 14924 13175 14976 13184
rect 14924 13141 14933 13175
rect 14933 13141 14967 13175
rect 14967 13141 14976 13175
rect 14924 13132 14976 13141
rect 17132 13175 17184 13184
rect 17132 13141 17141 13175
rect 17141 13141 17175 13175
rect 17175 13141 17184 13175
rect 17132 13132 17184 13141
rect 17960 13175 18012 13184
rect 17960 13141 17969 13175
rect 17969 13141 18003 13175
rect 18003 13141 18012 13175
rect 17960 13132 18012 13141
rect 20352 13175 20404 13184
rect 20352 13141 20361 13175
rect 20361 13141 20395 13175
rect 20395 13141 20404 13175
rect 20352 13132 20404 13141
rect 20904 13132 20956 13184
rect 22008 13209 22017 13243
rect 22017 13209 22051 13243
rect 22051 13209 22060 13243
rect 22008 13200 22060 13209
rect 22468 13200 22520 13252
rect 23664 13277 23673 13311
rect 23673 13277 23707 13311
rect 23707 13277 23716 13311
rect 23664 13268 23716 13277
rect 24308 13200 24360 13252
rect 22928 13132 22980 13184
rect 23756 13132 23808 13184
rect 9291 13030 9343 13082
rect 9355 13030 9407 13082
rect 9419 13030 9471 13082
rect 9483 13030 9535 13082
rect 9547 13030 9599 13082
rect 17632 13030 17684 13082
rect 17696 13030 17748 13082
rect 17760 13030 17812 13082
rect 17824 13030 17876 13082
rect 17888 13030 17940 13082
rect 2964 12928 3016 12980
rect 3332 12928 3384 12980
rect 5448 12928 5500 12980
rect 5632 12928 5684 12980
rect 6184 12928 6236 12980
rect 7380 12928 7432 12980
rect 9036 12928 9088 12980
rect 9680 12971 9732 12980
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 10140 12928 10192 12980
rect 10692 12928 10744 12980
rect 10876 12928 10928 12980
rect 14096 12928 14148 12980
rect 2780 12860 2832 12912
rect 3884 12903 3936 12912
rect 3884 12869 3893 12903
rect 3893 12869 3927 12903
rect 3927 12869 3936 12903
rect 3884 12860 3936 12869
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 5540 12792 5592 12844
rect 8668 12860 8720 12912
rect 6460 12792 6512 12844
rect 9864 12860 9916 12912
rect 10600 12860 10652 12912
rect 1676 12724 1728 12776
rect 4344 12724 4396 12776
rect 8668 12724 8720 12776
rect 8944 12724 8996 12776
rect 10048 12792 10100 12844
rect 11520 12792 11572 12844
rect 11612 12724 11664 12776
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 12440 12792 12492 12844
rect 12992 12792 13044 12844
rect 13636 12792 13688 12844
rect 15936 12860 15988 12912
rect 18144 12928 18196 12980
rect 18788 12928 18840 12980
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 21272 12928 21324 12980
rect 21640 12928 21692 12980
rect 22376 12860 22428 12912
rect 15016 12835 15068 12844
rect 15016 12801 15025 12835
rect 15025 12801 15059 12835
rect 15059 12801 15068 12835
rect 15016 12792 15068 12801
rect 15568 12792 15620 12844
rect 18420 12835 18472 12844
rect 18420 12801 18429 12835
rect 18429 12801 18463 12835
rect 18463 12801 18472 12835
rect 18420 12792 18472 12801
rect 19064 12792 19116 12844
rect 20812 12792 20864 12844
rect 21916 12792 21968 12844
rect 24124 12928 24176 12980
rect 22928 12860 22980 12912
rect 23848 12792 23900 12844
rect 24124 12792 24176 12844
rect 13268 12724 13320 12776
rect 17500 12724 17552 12776
rect 19340 12724 19392 12776
rect 19800 12724 19852 12776
rect 21456 12724 21508 12776
rect 21640 12724 21692 12776
rect 22008 12724 22060 12776
rect 9128 12699 9180 12708
rect 9128 12665 9137 12699
rect 9137 12665 9171 12699
rect 9171 12665 9180 12699
rect 9128 12656 9180 12665
rect 11336 12656 11388 12708
rect 12440 12656 12492 12708
rect 12716 12656 12768 12708
rect 22468 12656 22520 12708
rect 24124 12656 24176 12708
rect 8484 12588 8536 12640
rect 10324 12588 10376 12640
rect 11428 12588 11480 12640
rect 11888 12588 11940 12640
rect 12256 12588 12308 12640
rect 12532 12631 12584 12640
rect 12532 12597 12541 12631
rect 12541 12597 12575 12631
rect 12575 12597 12584 12631
rect 12532 12588 12584 12597
rect 13084 12588 13136 12640
rect 14924 12588 14976 12640
rect 21088 12588 21140 12640
rect 22652 12631 22704 12640
rect 22652 12597 22661 12631
rect 22661 12597 22695 12631
rect 22695 12597 22704 12631
rect 22652 12588 22704 12597
rect 22836 12631 22888 12640
rect 22836 12597 22845 12631
rect 22845 12597 22879 12631
rect 22879 12597 22888 12631
rect 23756 12631 23808 12640
rect 22836 12588 22888 12597
rect 23756 12597 23765 12631
rect 23765 12597 23799 12631
rect 23799 12597 23808 12631
rect 23756 12588 23808 12597
rect 5120 12486 5172 12538
rect 5184 12486 5236 12538
rect 5248 12486 5300 12538
rect 5312 12486 5364 12538
rect 5376 12486 5428 12538
rect 13462 12486 13514 12538
rect 13526 12486 13578 12538
rect 13590 12486 13642 12538
rect 13654 12486 13706 12538
rect 13718 12486 13770 12538
rect 21803 12486 21855 12538
rect 21867 12486 21919 12538
rect 21931 12486 21983 12538
rect 21995 12486 22047 12538
rect 22059 12486 22111 12538
rect 7932 12384 7984 12436
rect 9220 12384 9272 12436
rect 9588 12384 9640 12436
rect 8300 12316 8352 12368
rect 9036 12316 9088 12368
rect 8392 12248 8444 12300
rect 11152 12384 11204 12436
rect 11612 12384 11664 12436
rect 12624 12384 12676 12436
rect 6552 12180 6604 12232
rect 8668 12180 8720 12232
rect 9036 12180 9088 12232
rect 9220 12180 9272 12232
rect 9588 12180 9640 12232
rect 9772 12180 9824 12232
rect 10876 12248 10928 12300
rect 11336 12291 11388 12300
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11336 12257 11345 12291
rect 11345 12257 11379 12291
rect 11379 12257 11388 12291
rect 11336 12248 11388 12257
rect 11612 12223 11664 12232
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 12072 12180 12124 12232
rect 6828 12044 6880 12096
rect 7748 12044 7800 12096
rect 9036 12087 9088 12096
rect 9036 12053 9045 12087
rect 9045 12053 9079 12087
rect 9079 12053 9088 12087
rect 9036 12044 9088 12053
rect 10416 12044 10468 12096
rect 10876 12087 10928 12096
rect 10876 12053 10885 12087
rect 10885 12053 10919 12087
rect 10919 12053 10928 12087
rect 10876 12044 10928 12053
rect 12256 12112 12308 12164
rect 12624 12248 12676 12300
rect 23572 12384 23624 12436
rect 15752 12316 15804 12368
rect 16764 12316 16816 12368
rect 17224 12316 17276 12368
rect 17500 12316 17552 12368
rect 18420 12359 18472 12368
rect 18420 12325 18429 12359
rect 18429 12325 18463 12359
rect 18463 12325 18472 12359
rect 18420 12316 18472 12325
rect 15568 12248 15620 12300
rect 16580 12248 16632 12300
rect 20352 12316 20404 12368
rect 20812 12359 20864 12368
rect 20812 12325 20821 12359
rect 20821 12325 20855 12359
rect 20855 12325 20864 12359
rect 20812 12316 20864 12325
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 15108 12223 15160 12232
rect 15108 12189 15116 12223
rect 15116 12189 15150 12223
rect 15150 12189 15160 12223
rect 15108 12180 15160 12189
rect 12808 12112 12860 12164
rect 15936 12180 15988 12232
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 19800 12291 19852 12300
rect 19800 12257 19809 12291
rect 19809 12257 19843 12291
rect 19843 12257 19852 12291
rect 19800 12248 19852 12257
rect 21456 12291 21508 12300
rect 21456 12257 21465 12291
rect 21465 12257 21499 12291
rect 21499 12257 21508 12291
rect 21456 12248 21508 12257
rect 24124 12316 24176 12368
rect 21916 12248 21968 12300
rect 23664 12248 23716 12300
rect 11612 12044 11664 12096
rect 11796 12044 11848 12096
rect 13268 12044 13320 12096
rect 15384 12112 15436 12164
rect 15476 12044 15528 12096
rect 16672 12044 16724 12096
rect 18328 12180 18380 12232
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 18604 12223 18656 12232
rect 18604 12189 18613 12223
rect 18613 12189 18647 12223
rect 18647 12189 18656 12223
rect 18604 12180 18656 12189
rect 18788 12112 18840 12164
rect 19340 12112 19392 12164
rect 21640 12180 21692 12232
rect 22560 12223 22612 12232
rect 22560 12189 22569 12223
rect 22569 12189 22603 12223
rect 22603 12189 22612 12223
rect 22560 12180 22612 12189
rect 24584 12180 24636 12232
rect 20444 12112 20496 12164
rect 21916 12155 21968 12164
rect 21916 12121 21925 12155
rect 21925 12121 21959 12155
rect 21959 12121 21968 12155
rect 21916 12112 21968 12121
rect 19064 12044 19116 12096
rect 19616 12087 19668 12096
rect 19616 12053 19625 12087
rect 19625 12053 19659 12087
rect 19659 12053 19668 12087
rect 19616 12044 19668 12053
rect 20904 12087 20956 12096
rect 20904 12053 20913 12087
rect 20913 12053 20947 12087
rect 20947 12053 20956 12087
rect 20904 12044 20956 12053
rect 20996 12044 21048 12096
rect 21364 12087 21416 12096
rect 21364 12053 21373 12087
rect 21373 12053 21407 12087
rect 21407 12053 21416 12087
rect 21364 12044 21416 12053
rect 22100 12044 22152 12096
rect 22192 12087 22244 12096
rect 22192 12053 22201 12087
rect 22201 12053 22235 12087
rect 22235 12053 22244 12087
rect 22192 12044 22244 12053
rect 22836 12044 22888 12096
rect 23664 12087 23716 12096
rect 23664 12053 23673 12087
rect 23673 12053 23707 12087
rect 23707 12053 23716 12087
rect 24124 12087 24176 12096
rect 23664 12044 23716 12053
rect 24124 12053 24133 12087
rect 24133 12053 24167 12087
rect 24167 12053 24176 12087
rect 24124 12044 24176 12053
rect 24400 12087 24452 12096
rect 24400 12053 24409 12087
rect 24409 12053 24443 12087
rect 24443 12053 24452 12087
rect 24400 12044 24452 12053
rect 9291 11942 9343 11994
rect 9355 11942 9407 11994
rect 9419 11942 9471 11994
rect 9483 11942 9535 11994
rect 9547 11942 9599 11994
rect 17632 11942 17684 11994
rect 17696 11942 17748 11994
rect 17760 11942 17812 11994
rect 17824 11942 17876 11994
rect 17888 11942 17940 11994
rect 3240 11883 3292 11892
rect 3240 11849 3249 11883
rect 3249 11849 3283 11883
rect 3283 11849 3292 11883
rect 3240 11840 3292 11849
rect 8944 11840 8996 11892
rect 16856 11883 16908 11892
rect 1768 11704 1820 11756
rect 2596 11704 2648 11756
rect 4712 11772 4764 11824
rect 7196 11772 7248 11824
rect 3148 11747 3200 11756
rect 3148 11713 3157 11747
rect 3157 11713 3191 11747
rect 3191 11713 3200 11747
rect 3148 11704 3200 11713
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 7748 11704 7800 11756
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 3792 11636 3844 11688
rect 8392 11704 8444 11756
rect 8668 11704 8720 11756
rect 8852 11704 8904 11756
rect 8944 11704 8996 11756
rect 3424 11568 3476 11620
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 6000 11500 6052 11552
rect 6920 11500 6972 11552
rect 9036 11636 9088 11688
rect 15200 11772 15252 11824
rect 16396 11772 16448 11824
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 18144 11883 18196 11892
rect 18144 11849 18153 11883
rect 18153 11849 18187 11883
rect 18187 11849 18196 11883
rect 18144 11840 18196 11849
rect 18512 11840 18564 11892
rect 11796 11747 11848 11756
rect 11796 11713 11830 11747
rect 11830 11713 11848 11747
rect 11796 11704 11848 11713
rect 12072 11704 12124 11756
rect 11520 11679 11572 11688
rect 11520 11645 11529 11679
rect 11529 11645 11563 11679
rect 11563 11645 11572 11679
rect 11520 11636 11572 11645
rect 9220 11568 9272 11620
rect 9036 11500 9088 11552
rect 10600 11500 10652 11552
rect 12624 11500 12676 11552
rect 15660 11704 15712 11756
rect 16672 11747 16724 11756
rect 16672 11713 16681 11747
rect 16681 11713 16715 11747
rect 16715 11713 16724 11747
rect 16672 11704 16724 11713
rect 13176 11636 13228 11688
rect 14004 11636 14056 11688
rect 14464 11636 14516 11688
rect 15016 11679 15068 11688
rect 15016 11645 15025 11679
rect 15025 11645 15059 11679
rect 15059 11645 15068 11679
rect 15016 11636 15068 11645
rect 18328 11772 18380 11824
rect 17316 11704 17368 11756
rect 17500 11679 17552 11688
rect 17500 11645 17509 11679
rect 17509 11645 17543 11679
rect 17543 11645 17552 11679
rect 17500 11636 17552 11645
rect 18788 11747 18840 11756
rect 18788 11713 18797 11747
rect 18797 11713 18831 11747
rect 18831 11713 18840 11747
rect 18788 11704 18840 11713
rect 18880 11636 18932 11688
rect 19524 11840 19576 11892
rect 19616 11840 19668 11892
rect 19892 11840 19944 11892
rect 21916 11840 21968 11892
rect 23572 11840 23624 11892
rect 24400 11840 24452 11892
rect 19708 11772 19760 11824
rect 20536 11772 20588 11824
rect 21732 11772 21784 11824
rect 24584 11772 24636 11824
rect 19340 11704 19392 11756
rect 20444 11747 20496 11756
rect 20444 11713 20453 11747
rect 20453 11713 20487 11747
rect 20487 11713 20496 11747
rect 20444 11704 20496 11713
rect 20720 11704 20772 11756
rect 21548 11704 21600 11756
rect 21456 11679 21508 11688
rect 21456 11645 21465 11679
rect 21465 11645 21499 11679
rect 21499 11645 21508 11679
rect 21456 11636 21508 11645
rect 22192 11636 22244 11688
rect 22376 11679 22428 11688
rect 22376 11645 22385 11679
rect 22385 11645 22419 11679
rect 22419 11645 22428 11679
rect 22376 11636 22428 11645
rect 22468 11568 22520 11620
rect 23664 11636 23716 11688
rect 24308 11679 24360 11688
rect 24308 11645 24317 11679
rect 24317 11645 24351 11679
rect 24351 11645 24360 11679
rect 24308 11636 24360 11645
rect 14004 11500 14056 11552
rect 14188 11500 14240 11552
rect 14648 11500 14700 11552
rect 16120 11500 16172 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 17224 11500 17276 11552
rect 20720 11500 20772 11552
rect 21272 11500 21324 11552
rect 23204 11500 23256 11552
rect 23848 11500 23900 11552
rect 5120 11398 5172 11450
rect 5184 11398 5236 11450
rect 5248 11398 5300 11450
rect 5312 11398 5364 11450
rect 5376 11398 5428 11450
rect 13462 11398 13514 11450
rect 13526 11398 13578 11450
rect 13590 11398 13642 11450
rect 13654 11398 13706 11450
rect 13718 11398 13770 11450
rect 21803 11398 21855 11450
rect 21867 11398 21919 11450
rect 21931 11398 21983 11450
rect 21995 11398 22047 11450
rect 22059 11398 22111 11450
rect 1768 11339 1820 11348
rect 1768 11305 1777 11339
rect 1777 11305 1811 11339
rect 1811 11305 1820 11339
rect 1768 11296 1820 11305
rect 6828 11296 6880 11348
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 8760 11339 8812 11348
rect 8760 11305 8769 11339
rect 8769 11305 8803 11339
rect 8803 11305 8812 11339
rect 8760 11296 8812 11305
rect 9220 11296 9272 11348
rect 6736 11271 6788 11280
rect 6736 11237 6745 11271
rect 6745 11237 6779 11271
rect 6779 11237 6788 11271
rect 6736 11228 6788 11237
rect 8300 11271 8352 11280
rect 8300 11237 8309 11271
rect 8309 11237 8343 11271
rect 8343 11237 8352 11271
rect 8300 11228 8352 11237
rect 4712 11160 4764 11212
rect 8944 11203 8996 11212
rect 1676 10956 1728 11008
rect 3332 11135 3384 11144
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 3332 11092 3384 11101
rect 3056 10956 3108 11008
rect 4896 11092 4948 11144
rect 6736 11092 6788 11144
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9036 11092 9088 11144
rect 5632 11067 5684 11076
rect 5632 11033 5666 11067
rect 5666 11033 5684 11067
rect 5632 11024 5684 11033
rect 5816 11024 5868 11076
rect 5724 10956 5776 11008
rect 8668 11024 8720 11076
rect 10600 11296 10652 11348
rect 15660 11339 15712 11348
rect 13268 11228 13320 11280
rect 13452 11228 13504 11280
rect 14096 11228 14148 11280
rect 15108 11228 15160 11280
rect 15292 11228 15344 11280
rect 14280 11160 14332 11212
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 18328 11339 18380 11348
rect 18328 11305 18337 11339
rect 18337 11305 18371 11339
rect 18371 11305 18380 11339
rect 18328 11296 18380 11305
rect 20444 11296 20496 11348
rect 20996 11339 21048 11348
rect 20996 11305 21005 11339
rect 21005 11305 21039 11339
rect 21039 11305 21048 11339
rect 20996 11296 21048 11305
rect 22192 11296 22244 11348
rect 16580 11228 16632 11280
rect 11980 11092 12032 11144
rect 12440 11092 12492 11144
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 13176 11135 13228 11144
rect 13176 11101 13184 11135
rect 13184 11101 13218 11135
rect 13218 11101 13228 11135
rect 13176 11092 13228 11101
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 13452 11092 13504 11144
rect 12808 11024 12860 11076
rect 8300 10956 8352 11008
rect 10232 10956 10284 11008
rect 10600 10956 10652 11008
rect 14188 11092 14240 11144
rect 14004 11024 14056 11076
rect 14096 11067 14148 11076
rect 14096 11033 14105 11067
rect 14105 11033 14139 11067
rect 14139 11033 14148 11067
rect 15752 11160 15804 11212
rect 15200 11135 15252 11144
rect 15200 11101 15208 11135
rect 15208 11101 15242 11135
rect 15242 11101 15252 11135
rect 15200 11092 15252 11101
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 15936 11092 15988 11144
rect 16120 11092 16172 11144
rect 16488 11092 16540 11144
rect 16856 11160 16908 11212
rect 17500 11228 17552 11280
rect 18880 11228 18932 11280
rect 18788 11160 18840 11212
rect 19340 11228 19392 11280
rect 21180 11160 21232 11212
rect 22376 11228 22428 11280
rect 23296 11228 23348 11280
rect 24308 11160 24360 11212
rect 24676 11160 24728 11212
rect 14096 11024 14148 11033
rect 14648 11067 14700 11076
rect 14648 11033 14657 11067
rect 14657 11033 14691 11067
rect 14691 11033 14700 11067
rect 14648 11024 14700 11033
rect 14832 11067 14884 11076
rect 14832 11033 14841 11067
rect 14841 11033 14875 11067
rect 14875 11033 14884 11067
rect 14832 11024 14884 11033
rect 16856 11024 16908 11076
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 19616 11135 19668 11144
rect 18420 11092 18472 11101
rect 19616 11101 19625 11135
rect 19625 11101 19659 11135
rect 19659 11101 19668 11135
rect 19616 11092 19668 11101
rect 20536 11092 20588 11144
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 23204 11135 23256 11144
rect 23204 11101 23213 11135
rect 23213 11101 23247 11135
rect 23247 11101 23256 11135
rect 23204 11092 23256 11101
rect 23572 11092 23624 11144
rect 16580 10956 16632 11008
rect 22836 10999 22888 11008
rect 22836 10965 22845 10999
rect 22845 10965 22879 10999
rect 22879 10965 22888 10999
rect 22836 10956 22888 10965
rect 24768 10999 24820 11008
rect 24768 10965 24777 10999
rect 24777 10965 24811 10999
rect 24811 10965 24820 10999
rect 24768 10956 24820 10965
rect 9291 10854 9343 10906
rect 9355 10854 9407 10906
rect 9419 10854 9471 10906
rect 9483 10854 9535 10906
rect 9547 10854 9599 10906
rect 17632 10854 17684 10906
rect 17696 10854 17748 10906
rect 17760 10854 17812 10906
rect 17824 10854 17876 10906
rect 17888 10854 17940 10906
rect 5816 10752 5868 10804
rect 7196 10795 7248 10804
rect 7196 10761 7205 10795
rect 7205 10761 7239 10795
rect 7239 10761 7248 10795
rect 7196 10752 7248 10761
rect 8668 10752 8720 10804
rect 2504 10684 2556 10736
rect 3148 10684 3200 10736
rect 4252 10684 4304 10736
rect 3424 10659 3476 10668
rect 3424 10625 3433 10659
rect 3433 10625 3467 10659
rect 3467 10625 3476 10659
rect 3424 10616 3476 10625
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 4160 10616 4212 10668
rect 4528 10659 4580 10668
rect 4528 10625 4536 10659
rect 4536 10625 4570 10659
rect 4570 10625 4580 10659
rect 4528 10616 4580 10625
rect 4988 10684 5040 10736
rect 5632 10684 5684 10736
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 5448 10616 5500 10668
rect 5724 10659 5776 10668
rect 5724 10625 5734 10659
rect 5734 10625 5768 10659
rect 5768 10625 5776 10659
rect 7748 10684 7800 10736
rect 5724 10616 5776 10625
rect 6828 10616 6880 10668
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 8300 10684 8352 10736
rect 9496 10684 9548 10736
rect 12808 10684 12860 10736
rect 14004 10684 14056 10736
rect 15568 10752 15620 10804
rect 17040 10795 17092 10804
rect 17040 10761 17049 10795
rect 17049 10761 17083 10795
rect 17083 10761 17092 10795
rect 17040 10752 17092 10761
rect 17500 10752 17552 10804
rect 19340 10795 19392 10804
rect 18328 10684 18380 10736
rect 8116 10659 8168 10668
rect 8116 10625 8150 10659
rect 8150 10625 8168 10659
rect 8116 10616 8168 10625
rect 8944 10616 8996 10668
rect 9680 10659 9732 10668
rect 9680 10625 9714 10659
rect 9714 10625 9732 10659
rect 9680 10616 9732 10625
rect 1676 10548 1728 10600
rect 3608 10591 3660 10600
rect 3608 10557 3617 10591
rect 3617 10557 3651 10591
rect 3651 10557 3660 10591
rect 3608 10548 3660 10557
rect 2872 10480 2924 10532
rect 4344 10480 4396 10532
rect 6000 10548 6052 10600
rect 7472 10548 7524 10600
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 4528 10412 4580 10464
rect 6092 10412 6144 10464
rect 8208 10412 8260 10464
rect 14464 10616 14516 10668
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 15476 10659 15528 10668
rect 15476 10625 15519 10659
rect 15519 10625 15528 10659
rect 15476 10616 15528 10625
rect 15016 10591 15068 10600
rect 13452 10480 13504 10532
rect 11980 10412 12032 10464
rect 13084 10412 13136 10464
rect 15016 10557 15025 10591
rect 15025 10557 15059 10591
rect 15059 10557 15068 10591
rect 15016 10548 15068 10557
rect 15200 10591 15252 10600
rect 15200 10557 15209 10591
rect 15209 10557 15243 10591
rect 15243 10557 15252 10591
rect 15200 10548 15252 10557
rect 19340 10761 19349 10795
rect 19349 10761 19383 10795
rect 19383 10761 19392 10795
rect 19340 10752 19392 10761
rect 23480 10752 23532 10804
rect 24768 10752 24820 10804
rect 19616 10684 19668 10736
rect 23664 10684 23716 10736
rect 24676 10684 24728 10736
rect 18420 10480 18472 10532
rect 19708 10455 19760 10464
rect 19708 10421 19717 10455
rect 19717 10421 19751 10455
rect 19751 10421 19760 10455
rect 19708 10412 19760 10421
rect 5120 10310 5172 10362
rect 5184 10310 5236 10362
rect 5248 10310 5300 10362
rect 5312 10310 5364 10362
rect 5376 10310 5428 10362
rect 13462 10310 13514 10362
rect 13526 10310 13578 10362
rect 13590 10310 13642 10362
rect 13654 10310 13706 10362
rect 13718 10310 13770 10362
rect 21803 10310 21855 10362
rect 21867 10310 21919 10362
rect 21931 10310 21983 10362
rect 21995 10310 22047 10362
rect 22059 10310 22111 10362
rect 3332 10208 3384 10260
rect 7288 10208 7340 10260
rect 8116 10208 8168 10260
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 3424 10140 3476 10192
rect 9680 10208 9732 10260
rect 13360 10208 13412 10260
rect 13912 10251 13964 10260
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 15476 10208 15528 10260
rect 2872 10115 2924 10124
rect 2872 10081 2881 10115
rect 2881 10081 2915 10115
rect 2915 10081 2924 10115
rect 2872 10072 2924 10081
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 3792 10072 3844 10124
rect 4344 10115 4396 10124
rect 3240 10004 3292 10056
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 4712 10072 4764 10124
rect 4252 10047 4304 10056
rect 4252 10013 4261 10047
rect 4261 10013 4295 10047
rect 4295 10013 4304 10047
rect 4528 10047 4580 10056
rect 4252 10004 4304 10013
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 8760 10072 8812 10124
rect 8208 10004 8260 10056
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 8484 10047 8536 10056
rect 8484 10013 8494 10047
rect 8494 10013 8528 10047
rect 8528 10013 8536 10047
rect 8668 10047 8720 10056
rect 8484 10004 8536 10013
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 9128 10047 9180 10056
rect 9128 10013 9136 10047
rect 9136 10013 9170 10047
rect 9170 10013 9180 10047
rect 9128 10004 9180 10013
rect 10600 10140 10652 10192
rect 23112 10183 23164 10192
rect 9864 10115 9916 10124
rect 9864 10081 9873 10115
rect 9873 10081 9907 10115
rect 9907 10081 9916 10115
rect 14188 10115 14240 10124
rect 9864 10072 9916 10081
rect 14188 10081 14197 10115
rect 14197 10081 14231 10115
rect 14231 10081 14240 10115
rect 14188 10072 14240 10081
rect 15108 10072 15160 10124
rect 21456 10115 21508 10124
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 9496 10047 9548 10056
rect 4620 9936 4672 9988
rect 5540 9936 5592 9988
rect 3792 9911 3844 9920
rect 3792 9877 3801 9911
rect 3801 9877 3835 9911
rect 3835 9877 3844 9911
rect 3792 9868 3844 9877
rect 4160 9868 4212 9920
rect 4528 9868 4580 9920
rect 5632 9868 5684 9920
rect 8024 9936 8076 9988
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 14096 10047 14148 10056
rect 9680 9936 9732 9988
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 20720 10047 20772 10056
rect 20720 10013 20729 10047
rect 20729 10013 20763 10047
rect 20763 10013 20772 10047
rect 20720 10004 20772 10013
rect 20904 10004 20956 10056
rect 23112 10149 23121 10183
rect 23121 10149 23155 10183
rect 23155 10149 23164 10183
rect 23112 10140 23164 10149
rect 24584 10047 24636 10056
rect 24584 10013 24594 10047
rect 24594 10013 24628 10047
rect 24628 10013 24636 10047
rect 24952 10047 25004 10056
rect 24584 10004 24636 10013
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 25596 10004 25648 10056
rect 7012 9868 7064 9920
rect 9128 9868 9180 9920
rect 9864 9868 9916 9920
rect 22100 9936 22152 9988
rect 22652 9936 22704 9988
rect 24400 9979 24452 9988
rect 24400 9945 24409 9979
rect 24409 9945 24443 9979
rect 24443 9945 24452 9979
rect 24400 9936 24452 9945
rect 15200 9868 15252 9920
rect 15476 9868 15528 9920
rect 20536 9911 20588 9920
rect 20536 9877 20545 9911
rect 20545 9877 20579 9911
rect 20579 9877 20588 9911
rect 20536 9868 20588 9877
rect 20812 9911 20864 9920
rect 20812 9877 20821 9911
rect 20821 9877 20855 9911
rect 20855 9877 20864 9911
rect 20812 9868 20864 9877
rect 22284 9868 22336 9920
rect 23204 9868 23256 9920
rect 9291 9766 9343 9818
rect 9355 9766 9407 9818
rect 9419 9766 9471 9818
rect 9483 9766 9535 9818
rect 9547 9766 9599 9818
rect 17632 9766 17684 9818
rect 17696 9766 17748 9818
rect 17760 9766 17812 9818
rect 17824 9766 17876 9818
rect 17888 9766 17940 9818
rect 2780 9664 2832 9716
rect 5632 9707 5684 9716
rect 2320 9596 2372 9648
rect 3056 9596 3108 9648
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 3240 9528 3292 9580
rect 4068 9596 4120 9648
rect 4344 9596 4396 9648
rect 5632 9673 5641 9707
rect 5641 9673 5675 9707
rect 5675 9673 5684 9707
rect 5632 9664 5684 9673
rect 6736 9664 6788 9716
rect 9680 9664 9732 9716
rect 9772 9664 9824 9716
rect 13360 9664 13412 9716
rect 13912 9664 13964 9716
rect 14372 9664 14424 9716
rect 15568 9664 15620 9716
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 4804 9528 4856 9580
rect 5540 9596 5592 9648
rect 2596 9392 2648 9444
rect 1952 9324 2004 9376
rect 2780 9324 2832 9376
rect 3148 9392 3200 9444
rect 3884 9460 3936 9512
rect 4252 9460 4304 9512
rect 8576 9528 8628 9580
rect 8852 9528 8904 9580
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10784 9596 10836 9648
rect 17960 9639 18012 9648
rect 7012 9460 7064 9512
rect 7104 9460 7156 9512
rect 8484 9460 8536 9512
rect 4436 9392 4488 9444
rect 4712 9392 4764 9444
rect 8668 9392 8720 9444
rect 10232 9435 10284 9444
rect 10232 9401 10241 9435
rect 10241 9401 10275 9435
rect 10275 9401 10284 9435
rect 10232 9392 10284 9401
rect 3700 9367 3752 9376
rect 3700 9333 3709 9367
rect 3709 9333 3743 9367
rect 3743 9333 3752 9367
rect 3700 9324 3752 9333
rect 4528 9367 4580 9376
rect 4528 9333 4537 9367
rect 4537 9333 4571 9367
rect 4571 9333 4580 9367
rect 4528 9324 4580 9333
rect 4804 9324 4856 9376
rect 5448 9324 5500 9376
rect 7932 9324 7984 9376
rect 8116 9367 8168 9376
rect 8116 9333 8125 9367
rect 8125 9333 8159 9367
rect 8159 9333 8168 9367
rect 8116 9324 8168 9333
rect 8208 9324 8260 9376
rect 12164 9528 12216 9580
rect 13360 9528 13412 9580
rect 14188 9528 14240 9580
rect 15476 9571 15528 9580
rect 15476 9537 15485 9571
rect 15485 9537 15519 9571
rect 15519 9537 15528 9571
rect 15476 9528 15528 9537
rect 17316 9571 17368 9580
rect 17316 9537 17325 9571
rect 17325 9537 17359 9571
rect 17359 9537 17368 9571
rect 17316 9528 17368 9537
rect 17960 9605 17969 9639
rect 17969 9605 18003 9639
rect 18003 9605 18012 9639
rect 17960 9596 18012 9605
rect 21088 9596 21140 9648
rect 20628 9528 20680 9580
rect 21732 9596 21784 9648
rect 23112 9664 23164 9716
rect 24952 9664 25004 9716
rect 22192 9596 22244 9648
rect 24400 9596 24452 9648
rect 21548 9528 21600 9580
rect 14004 9460 14056 9512
rect 16672 9460 16724 9512
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 19800 9503 19852 9512
rect 13912 9392 13964 9444
rect 14924 9392 14976 9444
rect 17224 9392 17276 9444
rect 17960 9392 18012 9444
rect 19800 9469 19809 9503
rect 19809 9469 19843 9503
rect 19843 9469 19852 9503
rect 19800 9460 19852 9469
rect 20904 9503 20956 9512
rect 20904 9469 20913 9503
rect 20913 9469 20947 9503
rect 20947 9469 20956 9503
rect 20904 9460 20956 9469
rect 23480 9528 23532 9580
rect 25596 9571 25648 9580
rect 25596 9537 25605 9571
rect 25605 9537 25639 9571
rect 25639 9537 25648 9571
rect 25596 9528 25648 9537
rect 23296 9460 23348 9512
rect 23388 9503 23440 9512
rect 23388 9469 23397 9503
rect 23397 9469 23431 9503
rect 23431 9469 23440 9503
rect 23664 9503 23716 9512
rect 23388 9460 23440 9469
rect 23664 9469 23673 9503
rect 23673 9469 23707 9503
rect 23707 9469 23716 9503
rect 23664 9460 23716 9469
rect 21456 9392 21508 9444
rect 10692 9324 10744 9376
rect 11888 9324 11940 9376
rect 12256 9324 12308 9376
rect 14464 9324 14516 9376
rect 15292 9324 15344 9376
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 20720 9324 20772 9376
rect 21364 9367 21416 9376
rect 21364 9333 21373 9367
rect 21373 9333 21407 9367
rect 21407 9333 21416 9367
rect 21364 9324 21416 9333
rect 22928 9324 22980 9376
rect 24584 9324 24636 9376
rect 5120 9222 5172 9274
rect 5184 9222 5236 9274
rect 5248 9222 5300 9274
rect 5312 9222 5364 9274
rect 5376 9222 5428 9274
rect 13462 9222 13514 9274
rect 13526 9222 13578 9274
rect 13590 9222 13642 9274
rect 13654 9222 13706 9274
rect 13718 9222 13770 9274
rect 21803 9222 21855 9274
rect 21867 9222 21919 9274
rect 21931 9222 21983 9274
rect 21995 9222 22047 9274
rect 22059 9222 22111 9274
rect 3608 9120 3660 9172
rect 11060 9120 11112 9172
rect 13360 9120 13412 9172
rect 14004 9120 14056 9172
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 10968 9052 11020 9104
rect 3884 9027 3936 9036
rect 3884 8993 3893 9027
rect 3893 8993 3927 9027
rect 3927 8993 3936 9027
rect 3884 8984 3936 8993
rect 3976 8984 4028 9036
rect 7104 8984 7156 9036
rect 8484 8984 8536 9036
rect 9036 8984 9088 9036
rect 13912 9052 13964 9104
rect 1952 8959 2004 8968
rect 1952 8925 1986 8959
rect 1986 8925 2004 8959
rect 1952 8916 2004 8925
rect 3056 8916 3108 8968
rect 3700 8916 3752 8968
rect 3240 8848 3292 8900
rect 8300 8916 8352 8968
rect 8852 8916 8904 8968
rect 10876 8916 10928 8968
rect 12256 8959 12308 8968
rect 8024 8848 8076 8900
rect 8944 8891 8996 8900
rect 6920 8780 6972 8832
rect 8944 8857 8953 8891
rect 8953 8857 8987 8891
rect 8987 8857 8996 8891
rect 8944 8848 8996 8857
rect 9220 8848 9272 8900
rect 11152 8848 11204 8900
rect 11612 8848 11664 8900
rect 12256 8925 12265 8959
rect 12265 8925 12299 8959
rect 12299 8925 12308 8959
rect 12256 8916 12308 8925
rect 12624 8916 12676 8968
rect 14004 8984 14056 9036
rect 14372 9027 14424 9036
rect 14372 8993 14381 9027
rect 14381 8993 14415 9027
rect 14415 8993 14424 9027
rect 14372 8984 14424 8993
rect 15200 9052 15252 9104
rect 17040 9120 17092 9172
rect 20076 9163 20128 9172
rect 20076 9129 20085 9163
rect 20085 9129 20119 9163
rect 20119 9129 20128 9163
rect 20076 9120 20128 9129
rect 17960 8984 18012 9036
rect 19340 8984 19392 9036
rect 21456 9120 21508 9172
rect 23480 9120 23532 9172
rect 22284 9095 22336 9104
rect 22008 8984 22060 9036
rect 22284 9061 22293 9095
rect 22293 9061 22327 9095
rect 22327 9061 22336 9095
rect 22284 9052 22336 9061
rect 23388 8984 23440 9036
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 13360 8916 13412 8968
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 19064 8916 19116 8968
rect 15016 8848 15068 8900
rect 15292 8891 15344 8900
rect 15292 8857 15301 8891
rect 15301 8857 15335 8891
rect 15335 8857 15344 8891
rect 15292 8848 15344 8857
rect 8576 8780 8628 8832
rect 11796 8780 11848 8832
rect 13176 8780 13228 8832
rect 13360 8823 13412 8832
rect 13360 8789 13369 8823
rect 13369 8789 13403 8823
rect 13403 8789 13412 8823
rect 13360 8780 13412 8789
rect 15568 8848 15620 8900
rect 15844 8848 15896 8900
rect 20260 8959 20312 8968
rect 20260 8925 20269 8959
rect 20269 8925 20312 8959
rect 20260 8916 20312 8925
rect 20628 8959 20680 8968
rect 20628 8925 20637 8959
rect 20637 8925 20671 8959
rect 20671 8925 20680 8959
rect 20628 8916 20680 8925
rect 19984 8848 20036 8900
rect 15660 8823 15712 8832
rect 15660 8789 15669 8823
rect 15669 8789 15703 8823
rect 15703 8789 15712 8823
rect 15660 8780 15712 8789
rect 17408 8780 17460 8832
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 20168 8780 20220 8832
rect 20996 8891 21048 8900
rect 20996 8857 21030 8891
rect 21030 8857 21048 8891
rect 20996 8848 21048 8857
rect 21732 8916 21784 8968
rect 22928 8959 22980 8968
rect 22928 8925 22937 8959
rect 22937 8925 22971 8959
rect 22971 8925 22980 8959
rect 22928 8916 22980 8925
rect 23204 8959 23256 8968
rect 23204 8925 23213 8959
rect 23213 8925 23247 8959
rect 23247 8925 23256 8959
rect 23204 8916 23256 8925
rect 23756 8916 23808 8968
rect 22744 8848 22796 8900
rect 24860 8916 24912 8968
rect 25228 8916 25280 8968
rect 25596 8848 25648 8900
rect 23480 8823 23532 8832
rect 23480 8789 23489 8823
rect 23489 8789 23523 8823
rect 23523 8789 23532 8823
rect 23480 8780 23532 8789
rect 9291 8678 9343 8730
rect 9355 8678 9407 8730
rect 9419 8678 9471 8730
rect 9483 8678 9535 8730
rect 9547 8678 9599 8730
rect 17632 8678 17684 8730
rect 17696 8678 17748 8730
rect 17760 8678 17812 8730
rect 17824 8678 17876 8730
rect 17888 8678 17940 8730
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 3884 8576 3936 8628
rect 6092 8619 6144 8628
rect 3056 8483 3108 8492
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 8576 8576 8628 8628
rect 9036 8619 9088 8628
rect 9036 8585 9045 8619
rect 9045 8585 9079 8619
rect 9079 8585 9088 8619
rect 9036 8576 9088 8585
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 11612 8619 11664 8628
rect 11612 8585 11621 8619
rect 11621 8585 11655 8619
rect 11655 8585 11664 8619
rect 11612 8576 11664 8585
rect 12348 8576 12400 8628
rect 13360 8619 13412 8628
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 4068 8440 4120 8492
rect 4160 8440 4212 8492
rect 5356 8440 5408 8492
rect 5908 8440 5960 8492
rect 6920 8508 6972 8560
rect 7012 8508 7064 8560
rect 7932 8508 7984 8560
rect 10968 8508 11020 8560
rect 3240 8304 3292 8356
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 5632 8372 5684 8381
rect 6368 8372 6420 8424
rect 6736 8372 6788 8424
rect 6000 8347 6052 8356
rect 3148 8279 3200 8288
rect 3148 8245 3157 8279
rect 3157 8245 3191 8279
rect 3191 8245 3200 8279
rect 3148 8236 3200 8245
rect 3332 8236 3384 8288
rect 4344 8236 4396 8288
rect 6000 8313 6009 8347
rect 6009 8313 6043 8347
rect 6043 8313 6052 8347
rect 6000 8304 6052 8313
rect 6644 8304 6696 8356
rect 8484 8483 8536 8492
rect 8484 8449 8494 8483
rect 8494 8449 8528 8483
rect 8528 8449 8536 8483
rect 8668 8483 8720 8492
rect 8484 8440 8536 8449
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 11888 8551 11940 8560
rect 11888 8517 11897 8551
rect 11897 8517 11931 8551
rect 11931 8517 11940 8551
rect 11888 8508 11940 8517
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 14004 8619 14056 8628
rect 14004 8585 14013 8619
rect 14013 8585 14047 8619
rect 14047 8585 14056 8619
rect 14004 8576 14056 8585
rect 15016 8619 15068 8628
rect 15016 8585 15025 8619
rect 15025 8585 15059 8619
rect 15059 8585 15068 8619
rect 15016 8576 15068 8585
rect 15844 8619 15896 8628
rect 15844 8585 15853 8619
rect 15853 8585 15887 8619
rect 15887 8585 15896 8619
rect 15844 8576 15896 8585
rect 8208 8372 8260 8424
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 10232 8415 10284 8424
rect 8392 8372 8444 8381
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 10876 8415 10928 8424
rect 10232 8372 10284 8381
rect 9220 8304 9272 8356
rect 10600 8304 10652 8356
rect 10876 8381 10885 8415
rect 10885 8381 10919 8415
rect 10919 8381 10928 8415
rect 10876 8372 10928 8381
rect 11612 8372 11664 8424
rect 11796 8415 11848 8424
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 13912 8508 13964 8560
rect 14832 8508 14884 8560
rect 12716 8440 12768 8492
rect 17132 8576 17184 8628
rect 18052 8576 18104 8628
rect 21548 8619 21600 8628
rect 21548 8585 21557 8619
rect 21557 8585 21591 8619
rect 21591 8585 21600 8619
rect 21548 8576 21600 8585
rect 25228 8619 25280 8628
rect 25228 8585 25237 8619
rect 25237 8585 25271 8619
rect 25271 8585 25280 8619
rect 25228 8576 25280 8585
rect 19340 8508 19392 8560
rect 19800 8508 19852 8560
rect 16304 8440 16356 8492
rect 10784 8304 10836 8356
rect 10968 8236 11020 8288
rect 13268 8372 13320 8424
rect 14004 8372 14056 8424
rect 16488 8415 16540 8424
rect 16488 8381 16497 8415
rect 16497 8381 16531 8415
rect 16531 8381 16540 8415
rect 16488 8372 16540 8381
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 17960 8440 18012 8492
rect 18604 8440 18656 8492
rect 19524 8483 19576 8492
rect 19524 8449 19534 8483
rect 19534 8449 19568 8483
rect 19568 8449 19576 8483
rect 20168 8483 20220 8492
rect 19524 8440 19576 8449
rect 20168 8449 20177 8483
rect 20177 8449 20211 8483
rect 20211 8449 20220 8483
rect 20168 8440 20220 8449
rect 20536 8508 20588 8560
rect 21732 8508 21784 8560
rect 22008 8551 22060 8560
rect 22008 8517 22017 8551
rect 22017 8517 22051 8551
rect 22051 8517 22060 8551
rect 22008 8508 22060 8517
rect 22928 8508 22980 8560
rect 13360 8304 13412 8356
rect 17868 8372 17920 8424
rect 19892 8415 19944 8424
rect 19892 8381 19901 8415
rect 19901 8381 19935 8415
rect 19935 8381 19944 8415
rect 19892 8372 19944 8381
rect 19984 8415 20036 8424
rect 19984 8381 19993 8415
rect 19993 8381 20027 8415
rect 20027 8381 20036 8415
rect 19984 8372 20036 8381
rect 20168 8304 20220 8356
rect 22744 8440 22796 8492
rect 23664 8440 23716 8492
rect 23940 8440 23992 8492
rect 22652 8372 22704 8424
rect 23480 8372 23532 8424
rect 12532 8279 12584 8288
rect 12532 8245 12541 8279
rect 12541 8245 12575 8279
rect 12575 8245 12584 8279
rect 12532 8236 12584 8245
rect 23664 8236 23716 8288
rect 5120 8134 5172 8186
rect 5184 8134 5236 8186
rect 5248 8134 5300 8186
rect 5312 8134 5364 8186
rect 5376 8134 5428 8186
rect 13462 8134 13514 8186
rect 13526 8134 13578 8186
rect 13590 8134 13642 8186
rect 13654 8134 13706 8186
rect 13718 8134 13770 8186
rect 21803 8134 21855 8186
rect 21867 8134 21919 8186
rect 21931 8134 21983 8186
rect 21995 8134 22047 8186
rect 22059 8134 22111 8186
rect 3056 8032 3108 8084
rect 3792 7896 3844 7948
rect 4344 7939 4396 7948
rect 2136 7760 2188 7812
rect 3056 7828 3108 7880
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 5632 8032 5684 8084
rect 6460 8075 6512 8084
rect 6460 8041 6469 8075
rect 6469 8041 6503 8075
rect 6503 8041 6512 8075
rect 6460 8032 6512 8041
rect 6736 8075 6788 8084
rect 6736 8041 6745 8075
rect 6745 8041 6779 8075
rect 6779 8041 6788 8075
rect 6736 8032 6788 8041
rect 7012 8032 7064 8084
rect 7840 8032 7892 8084
rect 8116 8032 8168 8084
rect 9036 8032 9088 8084
rect 9864 8075 9916 8084
rect 9864 8041 9873 8075
rect 9873 8041 9907 8075
rect 9907 8041 9916 8075
rect 9864 8032 9916 8041
rect 10968 8032 11020 8084
rect 7104 7896 7156 7948
rect 8300 7964 8352 8016
rect 9128 7964 9180 8016
rect 11704 8007 11756 8016
rect 4804 7828 4856 7880
rect 4344 7760 4396 7812
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 7012 7828 7064 7837
rect 7840 7871 7892 7880
rect 6000 7760 6052 7812
rect 3424 7692 3476 7744
rect 3792 7692 3844 7744
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 5908 7692 5960 7744
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 7932 7828 7984 7880
rect 8300 7828 8352 7880
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 9036 7828 9088 7880
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 11704 7973 11713 8007
rect 11713 7973 11747 8007
rect 11747 7973 11756 8007
rect 11704 7964 11756 7973
rect 12164 7896 12216 7948
rect 13268 7896 13320 7948
rect 13452 7896 13504 7948
rect 9220 7828 9272 7837
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 10600 7871 10652 7880
rect 10600 7837 10634 7871
rect 10634 7837 10652 7871
rect 10600 7828 10652 7837
rect 11060 7828 11112 7880
rect 10140 7760 10192 7812
rect 12256 7828 12308 7880
rect 13820 7896 13872 7948
rect 15016 7828 15068 7880
rect 17132 8032 17184 8084
rect 17316 8075 17368 8084
rect 17316 8041 17325 8075
rect 17325 8041 17359 8075
rect 17359 8041 17368 8075
rect 17316 8032 17368 8041
rect 19340 8032 19392 8084
rect 17224 8007 17276 8016
rect 17224 7973 17233 8007
rect 17233 7973 17267 8007
rect 17267 7973 17276 8007
rect 17224 7964 17276 7973
rect 19984 8032 20036 8084
rect 20996 8032 21048 8084
rect 23940 8032 23992 8084
rect 20812 8007 20864 8016
rect 16396 7896 16448 7948
rect 19892 7896 19944 7948
rect 17408 7828 17460 7880
rect 20812 7973 20821 8007
rect 20821 7973 20855 8007
rect 20855 7973 20864 8007
rect 20812 7964 20864 7973
rect 12348 7760 12400 7812
rect 8300 7692 8352 7744
rect 8484 7735 8536 7744
rect 8484 7701 8493 7735
rect 8493 7701 8527 7735
rect 8527 7701 8536 7735
rect 8484 7692 8536 7701
rect 9220 7692 9272 7744
rect 12624 7692 12676 7744
rect 12808 7735 12860 7744
rect 12808 7701 12817 7735
rect 12817 7701 12851 7735
rect 12851 7701 12860 7735
rect 13268 7760 13320 7812
rect 14004 7760 14056 7812
rect 13176 7735 13228 7744
rect 12808 7692 12860 7701
rect 13176 7701 13185 7735
rect 13185 7701 13219 7735
rect 13219 7701 13228 7735
rect 13176 7692 13228 7701
rect 13912 7692 13964 7744
rect 17040 7760 17092 7812
rect 17500 7760 17552 7812
rect 20260 7828 20312 7880
rect 18328 7692 18380 7744
rect 19524 7692 19576 7744
rect 19800 7692 19852 7744
rect 23296 7871 23348 7880
rect 23296 7837 23305 7871
rect 23305 7837 23339 7871
rect 23339 7837 23348 7871
rect 23296 7828 23348 7837
rect 23664 7871 23716 7880
rect 23664 7837 23673 7871
rect 23673 7837 23707 7871
rect 23707 7837 23716 7871
rect 23664 7828 23716 7837
rect 23020 7692 23072 7744
rect 9291 7590 9343 7642
rect 9355 7590 9407 7642
rect 9419 7590 9471 7642
rect 9483 7590 9535 7642
rect 9547 7590 9599 7642
rect 17632 7590 17684 7642
rect 17696 7590 17748 7642
rect 17760 7590 17812 7642
rect 17824 7590 17876 7642
rect 17888 7590 17940 7642
rect 2136 7531 2188 7540
rect 2136 7497 2145 7531
rect 2145 7497 2179 7531
rect 2179 7497 2188 7531
rect 2136 7488 2188 7497
rect 4804 7488 4856 7540
rect 8300 7488 8352 7540
rect 9036 7488 9088 7540
rect 11612 7531 11664 7540
rect 11612 7497 11621 7531
rect 11621 7497 11655 7531
rect 11655 7497 11664 7531
rect 12532 7531 12584 7540
rect 11612 7488 11664 7497
rect 12532 7497 12541 7531
rect 12541 7497 12575 7531
rect 12575 7497 12584 7531
rect 12532 7488 12584 7497
rect 3424 7463 3476 7472
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 3424 7429 3433 7463
rect 3433 7429 3467 7463
rect 3467 7429 3476 7463
rect 3424 7420 3476 7429
rect 4712 7420 4764 7472
rect 2320 7352 2372 7361
rect 3056 7352 3108 7404
rect 3332 7352 3384 7404
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 10968 7420 11020 7472
rect 12808 7420 12860 7472
rect 7012 7352 7064 7404
rect 9220 7352 9272 7404
rect 11060 7352 11112 7404
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 13268 7395 13320 7404
rect 13268 7361 13277 7395
rect 13277 7361 13311 7395
rect 13311 7361 13320 7395
rect 13268 7352 13320 7361
rect 13544 7531 13596 7540
rect 13544 7497 13553 7531
rect 13553 7497 13587 7531
rect 13587 7497 13596 7531
rect 14004 7531 14056 7540
rect 13544 7488 13596 7497
rect 14004 7497 14013 7531
rect 14013 7497 14047 7531
rect 14047 7497 14056 7531
rect 14004 7488 14056 7497
rect 17408 7488 17460 7540
rect 18604 7531 18656 7540
rect 16764 7420 16816 7472
rect 13912 7395 13964 7404
rect 7932 7284 7984 7336
rect 10324 7284 10376 7336
rect 10508 7284 10560 7336
rect 12072 7284 12124 7336
rect 3240 7216 3292 7268
rect 3608 7259 3660 7268
rect 3608 7225 3617 7259
rect 3617 7225 3651 7259
rect 3651 7225 3660 7259
rect 3608 7216 3660 7225
rect 572 7148 624 7200
rect 2320 7148 2372 7200
rect 5632 7148 5684 7200
rect 6736 7148 6788 7200
rect 8300 7148 8352 7200
rect 9128 7148 9180 7200
rect 12164 7148 12216 7200
rect 12532 7284 12584 7336
rect 13912 7361 13921 7395
rect 13921 7361 13955 7395
rect 13955 7361 13964 7395
rect 13912 7352 13964 7361
rect 16856 7352 16908 7404
rect 17960 7395 18012 7404
rect 17960 7361 17969 7395
rect 17969 7361 18003 7395
rect 18003 7361 18012 7395
rect 17960 7352 18012 7361
rect 18604 7497 18613 7531
rect 18613 7497 18647 7531
rect 18647 7497 18656 7531
rect 18604 7488 18656 7497
rect 19800 7488 19852 7540
rect 22836 7531 22888 7540
rect 22836 7497 22845 7531
rect 22845 7497 22879 7531
rect 22879 7497 22888 7531
rect 22836 7488 22888 7497
rect 23848 7488 23900 7540
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 16488 7284 16540 7336
rect 17040 7284 17092 7336
rect 13452 7216 13504 7268
rect 19524 7352 19576 7404
rect 20536 7395 20588 7404
rect 20536 7361 20545 7395
rect 20545 7361 20579 7395
rect 20579 7361 20588 7395
rect 20536 7352 20588 7361
rect 24124 7352 24176 7404
rect 24308 7352 24360 7404
rect 24492 7352 24544 7404
rect 21364 7284 21416 7336
rect 23756 7327 23808 7336
rect 16120 7148 16172 7200
rect 19984 7216 20036 7268
rect 20168 7216 20220 7268
rect 23756 7293 23765 7327
rect 23765 7293 23799 7327
rect 23799 7293 23808 7327
rect 23756 7284 23808 7293
rect 23388 7216 23440 7268
rect 18144 7148 18196 7200
rect 20260 7148 20312 7200
rect 22284 7148 22336 7200
rect 22560 7148 22612 7200
rect 24860 7148 24912 7200
rect 5120 7046 5172 7098
rect 5184 7046 5236 7098
rect 5248 7046 5300 7098
rect 5312 7046 5364 7098
rect 5376 7046 5428 7098
rect 13462 7046 13514 7098
rect 13526 7046 13578 7098
rect 13590 7046 13642 7098
rect 13654 7046 13706 7098
rect 13718 7046 13770 7098
rect 21803 7046 21855 7098
rect 21867 7046 21919 7098
rect 21931 7046 21983 7098
rect 21995 7046 22047 7098
rect 22059 7046 22111 7098
rect 12256 6944 12308 6996
rect 10692 6876 10744 6928
rect 4344 6808 4396 6860
rect 5632 6808 5684 6860
rect 6460 6851 6512 6860
rect 6460 6817 6469 6851
rect 6469 6817 6503 6851
rect 6503 6817 6512 6851
rect 6460 6808 6512 6817
rect 7012 6808 7064 6860
rect 7564 6808 7616 6860
rect 5540 6672 5592 6724
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 6736 6740 6788 6792
rect 13176 6944 13228 6996
rect 12624 6876 12676 6928
rect 20536 6944 20588 6996
rect 23756 6944 23808 6996
rect 12440 6808 12492 6860
rect 13084 6808 13136 6860
rect 15476 6851 15528 6860
rect 10140 6783 10192 6792
rect 10140 6749 10158 6783
rect 10158 6749 10192 6783
rect 10140 6740 10192 6749
rect 10508 6740 10560 6792
rect 12256 6740 12308 6792
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 15476 6817 15485 6851
rect 15485 6817 15519 6851
rect 15519 6817 15528 6851
rect 16304 6851 16356 6860
rect 15476 6808 15528 6817
rect 16304 6817 16313 6851
rect 16313 6817 16347 6851
rect 16347 6817 16356 6851
rect 16304 6808 16356 6817
rect 16580 6808 16632 6860
rect 21640 6876 21692 6928
rect 22560 6876 22612 6928
rect 20352 6808 20404 6860
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 22744 6808 22796 6817
rect 24860 6876 24912 6928
rect 24492 6851 24544 6860
rect 24492 6817 24501 6851
rect 24501 6817 24535 6851
rect 24535 6817 24544 6851
rect 24492 6808 24544 6817
rect 3424 6604 3476 6656
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 6920 6672 6972 6724
rect 14188 6740 14240 6792
rect 15660 6740 15712 6792
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 21272 6783 21324 6792
rect 15844 6672 15896 6724
rect 16396 6672 16448 6724
rect 19064 6672 19116 6724
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 21456 6740 21508 6792
rect 23020 6783 23072 6792
rect 23020 6749 23054 6783
rect 23054 6749 23072 6783
rect 24400 6783 24452 6792
rect 23020 6740 23072 6749
rect 24400 6749 24409 6783
rect 24409 6749 24443 6783
rect 24443 6749 24452 6783
rect 24400 6740 24452 6749
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 7748 6604 7800 6613
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 12992 6647 13044 6656
rect 12992 6613 13001 6647
rect 13001 6613 13035 6647
rect 13035 6613 13044 6647
rect 12992 6604 13044 6613
rect 14832 6647 14884 6656
rect 14832 6613 14841 6647
rect 14841 6613 14875 6647
rect 14875 6613 14884 6647
rect 14832 6604 14884 6613
rect 14924 6647 14976 6656
rect 14924 6613 14933 6647
rect 14933 6613 14967 6647
rect 14967 6613 14976 6647
rect 14924 6604 14976 6613
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 15568 6604 15620 6656
rect 16764 6604 16816 6656
rect 20812 6647 20864 6656
rect 20812 6613 20821 6647
rect 20821 6613 20855 6647
rect 20855 6613 20864 6647
rect 20812 6604 20864 6613
rect 21548 6672 21600 6724
rect 22376 6672 22428 6724
rect 23296 6604 23348 6656
rect 9291 6502 9343 6554
rect 9355 6502 9407 6554
rect 9419 6502 9471 6554
rect 9483 6502 9535 6554
rect 9547 6502 9599 6554
rect 17632 6502 17684 6554
rect 17696 6502 17748 6554
rect 17760 6502 17812 6554
rect 17824 6502 17876 6554
rect 17888 6502 17940 6554
rect 2044 6264 2096 6316
rect 3240 6332 3292 6384
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 8392 6400 8444 6452
rect 9220 6400 9272 6452
rect 12440 6400 12492 6452
rect 14188 6443 14240 6452
rect 14188 6409 14197 6443
rect 14197 6409 14231 6443
rect 14231 6409 14240 6443
rect 14188 6400 14240 6409
rect 4068 6332 4120 6384
rect 4528 6332 4580 6384
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 3608 6264 3660 6316
rect 4160 6264 4212 6316
rect 6368 6332 6420 6384
rect 8484 6332 8536 6384
rect 5816 6264 5868 6316
rect 7748 6264 7800 6316
rect 3424 6196 3476 6248
rect 6460 6196 6512 6248
rect 4344 6128 4396 6180
rect 6368 6128 6420 6180
rect 2320 6103 2372 6112
rect 2320 6069 2329 6103
rect 2329 6069 2363 6103
rect 2363 6069 2372 6103
rect 2320 6060 2372 6069
rect 11520 6264 11572 6316
rect 12164 6307 12216 6316
rect 12164 6273 12173 6307
rect 12173 6273 12207 6307
rect 12207 6273 12216 6307
rect 12164 6264 12216 6273
rect 7932 6196 7984 6248
rect 9956 6196 10008 6248
rect 13912 6196 13964 6248
rect 14924 6400 14976 6452
rect 15016 6400 15068 6452
rect 16764 6443 16816 6452
rect 16764 6409 16773 6443
rect 16773 6409 16807 6443
rect 16807 6409 16816 6443
rect 16764 6400 16816 6409
rect 19064 6400 19116 6452
rect 19708 6400 19760 6452
rect 20352 6443 20404 6452
rect 20352 6409 20361 6443
rect 20361 6409 20395 6443
rect 20395 6409 20404 6443
rect 20352 6400 20404 6409
rect 20812 6443 20864 6452
rect 20812 6409 20821 6443
rect 20821 6409 20855 6443
rect 20855 6409 20864 6443
rect 20812 6400 20864 6409
rect 21180 6400 21232 6452
rect 15108 6332 15160 6384
rect 14832 6264 14884 6316
rect 15752 6264 15804 6316
rect 16580 6264 16632 6316
rect 19524 6332 19576 6384
rect 19800 6332 19852 6384
rect 21272 6332 21324 6384
rect 21548 6375 21600 6384
rect 21548 6341 21557 6375
rect 21557 6341 21591 6375
rect 21591 6341 21600 6375
rect 21548 6332 21600 6341
rect 24124 6400 24176 6452
rect 19248 6264 19300 6316
rect 21456 6264 21508 6316
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 17132 6196 17184 6248
rect 17316 6239 17368 6248
rect 17316 6205 17325 6239
rect 17325 6205 17359 6239
rect 17359 6205 17368 6239
rect 17316 6196 17368 6205
rect 19340 6196 19392 6248
rect 8024 6060 8076 6112
rect 12256 6060 12308 6112
rect 15660 6060 15712 6112
rect 17500 6128 17552 6180
rect 21364 6196 21416 6248
rect 16304 6103 16356 6112
rect 16304 6069 16313 6103
rect 16313 6069 16347 6103
rect 16347 6069 16356 6103
rect 16304 6060 16356 6069
rect 16396 6060 16448 6112
rect 19064 6103 19116 6112
rect 19064 6069 19073 6103
rect 19073 6069 19107 6103
rect 19107 6069 19116 6103
rect 19064 6060 19116 6069
rect 19616 6060 19668 6112
rect 22100 6264 22152 6316
rect 22744 6264 22796 6316
rect 23664 6264 23716 6316
rect 24400 6264 24452 6316
rect 23296 6060 23348 6112
rect 23572 6103 23624 6112
rect 23572 6069 23581 6103
rect 23581 6069 23615 6103
rect 23615 6069 23624 6103
rect 23572 6060 23624 6069
rect 5120 5958 5172 6010
rect 5184 5958 5236 6010
rect 5248 5958 5300 6010
rect 5312 5958 5364 6010
rect 5376 5958 5428 6010
rect 13462 5958 13514 6010
rect 13526 5958 13578 6010
rect 13590 5958 13642 6010
rect 13654 5958 13706 6010
rect 13718 5958 13770 6010
rect 21803 5958 21855 6010
rect 21867 5958 21919 6010
rect 21931 5958 21983 6010
rect 21995 5958 22047 6010
rect 22059 5958 22111 6010
rect 3056 5856 3108 5908
rect 8392 5856 8444 5908
rect 10876 5856 10928 5908
rect 15384 5856 15436 5908
rect 4344 5720 4396 5772
rect 2320 5652 2372 5704
rect 5540 5652 5592 5704
rect 2044 5516 2096 5568
rect 4896 5516 4948 5568
rect 6552 5584 6604 5636
rect 5724 5516 5776 5568
rect 6276 5516 6328 5568
rect 7932 5788 7984 5840
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 8668 5720 8720 5772
rect 8485 5695 8537 5704
rect 8485 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8537 5695
rect 8760 5695 8812 5704
rect 8485 5652 8537 5661
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 7748 5584 7800 5636
rect 11152 5788 11204 5840
rect 12992 5788 13044 5840
rect 12256 5763 12308 5772
rect 12256 5729 12265 5763
rect 12265 5729 12299 5763
rect 12299 5729 12308 5763
rect 12256 5720 12308 5729
rect 15660 5763 15712 5772
rect 11428 5695 11480 5704
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 11520 5652 11572 5704
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 16488 5856 16540 5908
rect 19340 5899 19392 5908
rect 19340 5865 19349 5899
rect 19349 5865 19383 5899
rect 19383 5865 19392 5899
rect 19340 5856 19392 5865
rect 21272 5856 21324 5908
rect 22192 5856 22244 5908
rect 12992 5652 13044 5661
rect 15108 5652 15160 5704
rect 10508 5584 10560 5636
rect 11888 5584 11940 5636
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 17316 5652 17368 5704
rect 19064 5788 19116 5840
rect 22284 5831 22336 5840
rect 22284 5797 22293 5831
rect 22293 5797 22327 5831
rect 22327 5797 22336 5831
rect 22284 5788 22336 5797
rect 23664 5831 23716 5840
rect 23664 5797 23673 5831
rect 23673 5797 23707 5831
rect 23707 5797 23716 5831
rect 23664 5788 23716 5797
rect 19984 5763 20036 5772
rect 19984 5729 19993 5763
rect 19993 5729 20027 5763
rect 20027 5729 20036 5763
rect 19984 5720 20036 5729
rect 22376 5720 22428 5772
rect 19156 5652 19208 5704
rect 19616 5652 19668 5704
rect 19800 5695 19852 5704
rect 19800 5661 19809 5695
rect 19809 5661 19843 5695
rect 19843 5661 19852 5695
rect 19800 5652 19852 5661
rect 20260 5695 20312 5704
rect 20260 5661 20294 5695
rect 20294 5661 20312 5695
rect 16304 5584 16356 5636
rect 16488 5584 16540 5636
rect 17500 5584 17552 5636
rect 19248 5584 19300 5636
rect 20260 5652 20312 5661
rect 23296 5695 23348 5704
rect 23296 5661 23305 5695
rect 23305 5661 23339 5695
rect 23339 5661 23348 5695
rect 23296 5652 23348 5661
rect 23572 5652 23624 5704
rect 11612 5559 11664 5568
rect 11612 5525 11621 5559
rect 11621 5525 11655 5559
rect 11655 5525 11664 5559
rect 11612 5516 11664 5525
rect 14648 5559 14700 5568
rect 14648 5525 14657 5559
rect 14657 5525 14691 5559
rect 14691 5525 14700 5559
rect 14648 5516 14700 5525
rect 15292 5516 15344 5568
rect 17132 5516 17184 5568
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 9291 5414 9343 5466
rect 9355 5414 9407 5466
rect 9419 5414 9471 5466
rect 9483 5414 9535 5466
rect 9547 5414 9599 5466
rect 17632 5414 17684 5466
rect 17696 5414 17748 5466
rect 17760 5414 17812 5466
rect 17824 5414 17876 5466
rect 17888 5414 17940 5466
rect 3332 5244 3384 5296
rect 8116 5312 8168 5364
rect 8484 5312 8536 5364
rect 8760 5312 8812 5364
rect 11428 5312 11480 5364
rect 15752 5312 15804 5364
rect 16580 5312 16632 5364
rect 16948 5312 17000 5364
rect 17224 5355 17276 5364
rect 17224 5321 17233 5355
rect 17233 5321 17267 5355
rect 17267 5321 17276 5355
rect 17224 5312 17276 5321
rect 19800 5312 19852 5364
rect 5448 5244 5500 5296
rect 3884 5219 3936 5228
rect 3884 5185 3902 5219
rect 3902 5185 3936 5219
rect 3884 5176 3936 5185
rect 4344 5176 4396 5228
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 8024 5244 8076 5296
rect 8208 5287 8260 5296
rect 8208 5253 8242 5287
rect 8242 5253 8260 5287
rect 8208 5244 8260 5253
rect 9220 5244 9272 5296
rect 10876 5244 10928 5296
rect 11612 5244 11664 5296
rect 12624 5244 12676 5296
rect 6368 5219 6420 5228
rect 4804 5108 4856 5160
rect 5724 5108 5776 5160
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 6644 5219 6696 5228
rect 6644 5185 6678 5219
rect 6678 5185 6696 5219
rect 7932 5219 7984 5228
rect 6644 5176 6696 5185
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 8484 5176 8536 5228
rect 10508 5176 10560 5228
rect 3884 4972 3936 5024
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 5816 4972 5868 4981
rect 6276 4972 6328 5024
rect 7472 4972 7524 5024
rect 7840 4972 7892 5024
rect 11152 5083 11204 5092
rect 11152 5049 11161 5083
rect 11161 5049 11195 5083
rect 11195 5049 11204 5083
rect 11152 5040 11204 5049
rect 10600 4972 10652 5024
rect 12532 4972 12584 5024
rect 12808 4972 12860 5024
rect 12992 5176 13044 5228
rect 15476 5176 15528 5228
rect 16488 5244 16540 5296
rect 15292 5108 15344 5160
rect 15752 5108 15804 5160
rect 17132 5176 17184 5228
rect 17408 5176 17460 5228
rect 18420 5244 18472 5296
rect 17684 5151 17736 5160
rect 17684 5117 17693 5151
rect 17693 5117 17727 5151
rect 17727 5117 17736 5151
rect 17684 5108 17736 5117
rect 18880 5151 18932 5160
rect 18880 5117 18889 5151
rect 18889 5117 18923 5151
rect 18923 5117 18932 5151
rect 18880 5108 18932 5117
rect 13820 5040 13872 5092
rect 15568 5083 15620 5092
rect 15568 5049 15577 5083
rect 15577 5049 15611 5083
rect 15611 5049 15620 5083
rect 15568 5040 15620 5049
rect 16764 5015 16816 5024
rect 16764 4981 16773 5015
rect 16773 4981 16807 5015
rect 16807 4981 16816 5015
rect 16764 4972 16816 4981
rect 17500 4972 17552 5024
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 19248 4972 19300 5024
rect 5120 4870 5172 4922
rect 5184 4870 5236 4922
rect 5248 4870 5300 4922
rect 5312 4870 5364 4922
rect 5376 4870 5428 4922
rect 13462 4870 13514 4922
rect 13526 4870 13578 4922
rect 13590 4870 13642 4922
rect 13654 4870 13706 4922
rect 13718 4870 13770 4922
rect 21803 4870 21855 4922
rect 21867 4870 21919 4922
rect 21931 4870 21983 4922
rect 21995 4870 22047 4922
rect 22059 4870 22111 4922
rect 4252 4768 4304 4820
rect 5448 4768 5500 4820
rect 5816 4768 5868 4820
rect 6644 4768 6696 4820
rect 6552 4700 6604 4752
rect 8392 4768 8444 4820
rect 8668 4768 8720 4820
rect 10600 4811 10652 4820
rect 10600 4777 10609 4811
rect 10609 4777 10643 4811
rect 10643 4777 10652 4811
rect 10600 4768 10652 4777
rect 14004 4768 14056 4820
rect 17224 4768 17276 4820
rect 7656 4700 7708 4752
rect 5908 4675 5960 4684
rect 5908 4641 5917 4675
rect 5917 4641 5951 4675
rect 5951 4641 5960 4675
rect 5908 4632 5960 4641
rect 2044 4607 2096 4616
rect 2044 4573 2053 4607
rect 2053 4573 2087 4607
rect 2087 4573 2096 4607
rect 2044 4564 2096 4573
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 7472 4632 7524 4684
rect 9220 4700 9272 4752
rect 8208 4675 8260 4684
rect 8208 4641 8217 4675
rect 8217 4641 8251 4675
rect 8251 4641 8260 4675
rect 8208 4632 8260 4641
rect 8576 4632 8628 4684
rect 10876 4632 10928 4684
rect 12256 4632 12308 4684
rect 4804 4496 4856 4548
rect 4988 4428 5040 4480
rect 5724 4428 5776 4480
rect 7104 4471 7156 4480
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 7748 4564 7800 4616
rect 8116 4564 8168 4616
rect 8484 4564 8536 4616
rect 10508 4564 10560 4616
rect 11520 4564 11572 4616
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13820 4564 13872 4616
rect 15108 4632 15160 4684
rect 15476 4700 15528 4752
rect 16764 4700 16816 4752
rect 17684 4700 17736 4752
rect 16580 4632 16632 4684
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 15200 4607 15252 4616
rect 15200 4573 15209 4607
rect 15209 4573 15243 4607
rect 15243 4573 15252 4607
rect 15200 4564 15252 4573
rect 14372 4496 14424 4548
rect 15752 4539 15804 4548
rect 15752 4505 15761 4539
rect 15761 4505 15795 4539
rect 15795 4505 15804 4539
rect 15752 4496 15804 4505
rect 16580 4539 16632 4548
rect 16580 4505 16589 4539
rect 16589 4505 16623 4539
rect 16623 4505 16632 4539
rect 16580 4496 16632 4505
rect 16764 4539 16816 4548
rect 16764 4505 16773 4539
rect 16773 4505 16807 4539
rect 16807 4505 16816 4539
rect 18052 4564 18104 4616
rect 16764 4496 16816 4505
rect 8024 4428 8076 4480
rect 11520 4428 11572 4480
rect 12072 4428 12124 4480
rect 12164 4471 12216 4480
rect 12164 4437 12173 4471
rect 12173 4437 12207 4471
rect 12207 4437 12216 4471
rect 12164 4428 12216 4437
rect 12716 4428 12768 4480
rect 14096 4428 14148 4480
rect 14464 4471 14516 4480
rect 14464 4437 14473 4471
rect 14473 4437 14507 4471
rect 14507 4437 14516 4471
rect 14464 4428 14516 4437
rect 14924 4428 14976 4480
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 17132 4428 17184 4480
rect 9291 4326 9343 4378
rect 9355 4326 9407 4378
rect 9419 4326 9471 4378
rect 9483 4326 9535 4378
rect 9547 4326 9599 4378
rect 17632 4326 17684 4378
rect 17696 4326 17748 4378
rect 17760 4326 17812 4378
rect 17824 4326 17876 4378
rect 17888 4326 17940 4378
rect 4804 4267 4856 4276
rect 4804 4233 4813 4267
rect 4813 4233 4847 4267
rect 4847 4233 4856 4267
rect 4804 4224 4856 4233
rect 5816 4224 5868 4276
rect 6000 4224 6052 4276
rect 7748 4267 7800 4276
rect 7748 4233 7757 4267
rect 7757 4233 7791 4267
rect 7791 4233 7800 4267
rect 7748 4224 7800 4233
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 7472 4156 7524 4208
rect 8208 4156 8260 4208
rect 5448 4088 5500 4140
rect 6092 4088 6144 4140
rect 6276 4088 6328 4140
rect 5540 4020 5592 4072
rect 6736 4020 6788 4072
rect 7104 4088 7156 4140
rect 8024 4088 8076 4140
rect 7656 4020 7708 4072
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 8300 4020 8352 4072
rect 9036 4088 9088 4140
rect 10600 4224 10652 4276
rect 14280 4267 14332 4276
rect 14280 4233 14289 4267
rect 14289 4233 14323 4267
rect 14323 4233 14332 4267
rect 14280 4224 14332 4233
rect 10876 4156 10928 4208
rect 12072 4199 12124 4208
rect 12072 4165 12081 4199
rect 12081 4165 12115 4199
rect 12115 4165 12124 4199
rect 12072 4156 12124 4165
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 13820 4156 13872 4208
rect 14004 4156 14056 4208
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 12808 4088 12860 4140
rect 13176 4131 13228 4140
rect 13176 4097 13210 4131
rect 13210 4097 13228 4131
rect 13176 4088 13228 4097
rect 14372 4088 14424 4140
rect 15108 4156 15160 4208
rect 15292 4156 15344 4208
rect 16488 4156 16540 4208
rect 7104 3952 7156 4004
rect 8208 3952 8260 4004
rect 12164 4020 12216 4072
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 5816 3884 5868 3936
rect 8300 3884 8352 3936
rect 8484 3884 8536 3936
rect 11060 3884 11112 3936
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 11796 3884 11848 3936
rect 12348 3952 12400 4004
rect 16580 4088 16632 4140
rect 17408 4156 17460 4208
rect 17132 4131 17184 4140
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 14740 3952 14792 4004
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 22744 4156 22796 4208
rect 22284 4131 22336 4140
rect 22284 4097 22318 4131
rect 22318 4097 22336 4131
rect 22284 4088 22336 4097
rect 12716 3884 12768 3936
rect 14464 3884 14516 3936
rect 17132 3952 17184 4004
rect 18236 3952 18288 4004
rect 23112 3952 23164 4004
rect 16488 3884 16540 3936
rect 17316 3927 17368 3936
rect 17316 3893 17325 3927
rect 17325 3893 17359 3927
rect 17359 3893 17368 3927
rect 17316 3884 17368 3893
rect 5120 3782 5172 3834
rect 5184 3782 5236 3834
rect 5248 3782 5300 3834
rect 5312 3782 5364 3834
rect 5376 3782 5428 3834
rect 13462 3782 13514 3834
rect 13526 3782 13578 3834
rect 13590 3782 13642 3834
rect 13654 3782 13706 3834
rect 13718 3782 13770 3834
rect 21803 3782 21855 3834
rect 21867 3782 21919 3834
rect 21931 3782 21983 3834
rect 21995 3782 22047 3834
rect 22059 3782 22111 3834
rect 4068 3680 4120 3732
rect 5632 3680 5684 3732
rect 5724 3680 5776 3732
rect 7656 3723 7708 3732
rect 7656 3689 7665 3723
rect 7665 3689 7699 3723
rect 7699 3689 7708 3723
rect 7656 3680 7708 3689
rect 8852 3680 8904 3732
rect 10048 3680 10100 3732
rect 2780 3612 2832 3664
rect 4344 3544 4396 3596
rect 7932 3544 7984 3596
rect 8392 3612 8444 3664
rect 8208 3587 8260 3596
rect 8208 3553 8217 3587
rect 8217 3553 8251 3587
rect 8251 3553 8260 3587
rect 13268 3680 13320 3732
rect 14004 3680 14056 3732
rect 14556 3680 14608 3732
rect 15016 3680 15068 3732
rect 14096 3655 14148 3664
rect 14096 3621 14105 3655
rect 14105 3621 14139 3655
rect 14139 3621 14148 3655
rect 14096 3612 14148 3621
rect 15844 3680 15896 3732
rect 16580 3612 16632 3664
rect 16764 3655 16816 3664
rect 16764 3621 16773 3655
rect 16773 3621 16807 3655
rect 16807 3621 16816 3655
rect 16764 3612 16816 3621
rect 18880 3680 18932 3732
rect 22284 3723 22336 3732
rect 22284 3689 22293 3723
rect 22293 3689 22327 3723
rect 22327 3689 22336 3723
rect 22284 3680 22336 3689
rect 8208 3544 8260 3553
rect 1676 3408 1728 3460
rect 3792 3408 3844 3460
rect 4804 3408 4856 3460
rect 6000 3408 6052 3460
rect 7748 3476 7800 3528
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 6092 3383 6144 3392
rect 6092 3349 6101 3383
rect 6101 3349 6135 3383
rect 6135 3349 6144 3383
rect 6092 3340 6144 3349
rect 10508 3519 10560 3528
rect 10508 3485 10517 3519
rect 10517 3485 10551 3519
rect 10551 3485 10560 3519
rect 10508 3476 10560 3485
rect 10784 3519 10836 3528
rect 10784 3485 10818 3519
rect 10818 3485 10836 3519
rect 10784 3476 10836 3485
rect 11060 3476 11112 3528
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 14464 3476 14516 3528
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 17316 3476 17368 3528
rect 23112 3519 23164 3528
rect 23112 3485 23121 3519
rect 23121 3485 23155 3519
rect 23155 3485 23164 3519
rect 23112 3476 23164 3485
rect 24308 3476 24360 3528
rect 25504 3476 25556 3528
rect 14280 3340 14332 3392
rect 14740 3340 14792 3392
rect 16120 3408 16172 3460
rect 21732 3408 21784 3460
rect 21640 3383 21692 3392
rect 21640 3349 21649 3383
rect 21649 3349 21683 3383
rect 21683 3349 21692 3383
rect 22652 3383 22704 3392
rect 21640 3340 21692 3349
rect 22652 3349 22661 3383
rect 22661 3349 22695 3383
rect 22695 3349 22704 3383
rect 22652 3340 22704 3349
rect 9291 3238 9343 3290
rect 9355 3238 9407 3290
rect 9419 3238 9471 3290
rect 9483 3238 9535 3290
rect 9547 3238 9599 3290
rect 17632 3238 17684 3290
rect 17696 3238 17748 3290
rect 17760 3238 17812 3290
rect 17824 3238 17876 3290
rect 17888 3238 17940 3290
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 6000 3179 6052 3188
rect 6000 3145 6009 3179
rect 6009 3145 6043 3179
rect 6043 3145 6052 3179
rect 6000 3136 6052 3145
rect 6276 3136 6328 3188
rect 7472 3179 7524 3188
rect 7472 3145 7481 3179
rect 7481 3145 7515 3179
rect 7515 3145 7524 3179
rect 7472 3136 7524 3145
rect 11980 3136 12032 3188
rect 12440 3136 12492 3188
rect 12624 3136 12676 3188
rect 13176 3136 13228 3188
rect 14832 3179 14884 3188
rect 14832 3145 14841 3179
rect 14841 3145 14875 3179
rect 14875 3145 14884 3179
rect 14832 3136 14884 3145
rect 5448 3068 5500 3120
rect 5632 3000 5684 3052
rect 5908 3068 5960 3120
rect 11244 3068 11296 3120
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 8576 3043 8628 3052
rect 5816 3000 5868 3009
rect 8576 3009 8594 3043
rect 8594 3009 8628 3043
rect 8576 3000 8628 3009
rect 10508 3000 10560 3052
rect 11796 3043 11848 3052
rect 11796 3009 11830 3043
rect 11830 3009 11848 3043
rect 11796 3000 11848 3009
rect 13912 3068 13964 3120
rect 22376 3136 22428 3188
rect 15752 3068 15804 3120
rect 13268 3000 13320 3052
rect 22192 3068 22244 3120
rect 6092 2932 6144 2984
rect 15016 2932 15068 2984
rect 19524 2932 19576 2984
rect 5908 2864 5960 2916
rect 14924 2907 14976 2916
rect 14924 2873 14933 2907
rect 14933 2873 14967 2907
rect 14967 2873 14976 2907
rect 14924 2864 14976 2873
rect 8208 2796 8260 2848
rect 14740 2796 14792 2848
rect 16028 2796 16080 2848
rect 5120 2694 5172 2746
rect 5184 2694 5236 2746
rect 5248 2694 5300 2746
rect 5312 2694 5364 2746
rect 5376 2694 5428 2746
rect 13462 2694 13514 2746
rect 13526 2694 13578 2746
rect 13590 2694 13642 2746
rect 13654 2694 13706 2746
rect 13718 2694 13770 2746
rect 21803 2694 21855 2746
rect 21867 2694 21919 2746
rect 21931 2694 21983 2746
rect 21995 2694 22047 2746
rect 22059 2694 22111 2746
rect 8208 2592 8260 2644
rect 8576 2592 8628 2644
rect 7472 2456 7524 2508
rect 7748 2388 7800 2440
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 9291 2150 9343 2202
rect 9355 2150 9407 2202
rect 9419 2150 9471 2202
rect 9483 2150 9535 2202
rect 9547 2150 9599 2202
rect 17632 2150 17684 2202
rect 17696 2150 17748 2202
rect 17760 2150 17812 2202
rect 17824 2150 17876 2202
rect 17888 2150 17940 2202
rect 3148 1300 3200 1352
rect 12900 1300 12952 1352
<< metal2 >>
rect 570 28642 626 29442
rect 1674 28642 1730 29442
rect 2870 28642 2926 29442
rect 3528 28750 4016 28778
rect 584 26042 612 28642
rect 572 26036 624 26042
rect 572 25978 624 25984
rect 1688 24886 1716 28642
rect 1676 24880 1728 24886
rect 1676 24822 1728 24828
rect 2688 24880 2740 24886
rect 2688 24822 2740 24828
rect 2134 24440 2190 24449
rect 2134 24375 2136 24384
rect 2188 24375 2190 24384
rect 2136 24346 2188 24352
rect 2136 23112 2188 23118
rect 2134 23080 2136 23089
rect 2188 23080 2190 23089
rect 2134 23015 2190 23024
rect 1492 20460 1544 20466
rect 1492 20402 1544 20408
rect 1504 19922 1532 20402
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 1504 19378 1532 19858
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 2056 17270 2084 17614
rect 2044 17264 2096 17270
rect 2044 17206 2096 17212
rect 2056 16658 2084 17206
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2700 14822 2728 24822
rect 2884 22094 2912 28642
rect 2884 22066 3096 22094
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2792 20534 2820 21966
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2872 18148 2924 18154
rect 2872 18090 2924 18096
rect 2780 17604 2832 17610
rect 2780 17546 2832 17552
rect 2792 16182 2820 17546
rect 2884 16590 2912 18090
rect 2964 17604 3016 17610
rect 2964 17546 3016 17552
rect 2976 17134 3004 17546
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2976 16590 3004 17070
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2780 16176 2832 16182
rect 2780 16118 2832 16124
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 2792 15094 2820 15370
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2976 15026 3004 16526
rect 3068 15502 3096 22066
rect 3240 21956 3292 21962
rect 3240 21898 3292 21904
rect 3252 21690 3280 21898
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3344 21570 3372 21830
rect 3252 21554 3372 21570
rect 3240 21548 3372 21554
rect 3292 21542 3372 21548
rect 3240 21490 3292 21496
rect 3252 20942 3280 21490
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 3160 19854 3188 20198
rect 3252 20074 3280 20878
rect 3252 20046 3372 20074
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3160 18290 3188 19790
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 3252 18222 3280 18294
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3252 16250 3280 18158
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3344 16182 3372 20046
rect 3424 17060 3476 17066
rect 3424 17002 3476 17008
rect 3436 16794 3464 17002
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 3528 15910 3556 28750
rect 3988 28642 4016 28750
rect 4066 28642 4122 29442
rect 5262 28642 5318 29442
rect 5736 28750 6408 28778
rect 3988 28614 4108 28642
rect 5120 26684 5428 26704
rect 5120 26682 5126 26684
rect 5182 26682 5206 26684
rect 5262 26682 5286 26684
rect 5342 26682 5366 26684
rect 5422 26682 5428 26684
rect 5182 26630 5184 26682
rect 5364 26630 5366 26682
rect 5120 26628 5126 26630
rect 5182 26628 5206 26630
rect 5262 26628 5286 26630
rect 5342 26628 5366 26630
rect 5422 26628 5428 26630
rect 5120 26608 5428 26628
rect 5120 25596 5428 25616
rect 5120 25594 5126 25596
rect 5182 25594 5206 25596
rect 5262 25594 5286 25596
rect 5342 25594 5366 25596
rect 5422 25594 5428 25596
rect 5182 25542 5184 25594
rect 5364 25542 5366 25594
rect 5120 25540 5126 25542
rect 5182 25540 5206 25542
rect 5262 25540 5286 25542
rect 5342 25540 5366 25542
rect 5422 25540 5428 25542
rect 5120 25520 5428 25540
rect 5120 24508 5428 24528
rect 5120 24506 5126 24508
rect 5182 24506 5206 24508
rect 5262 24506 5286 24508
rect 5342 24506 5366 24508
rect 5422 24506 5428 24508
rect 5182 24454 5184 24506
rect 5364 24454 5366 24506
rect 5120 24452 5126 24454
rect 5182 24452 5206 24454
rect 5262 24452 5286 24454
rect 5342 24452 5366 24454
rect 5422 24452 5428 24454
rect 5120 24432 5428 24452
rect 3792 24200 3844 24206
rect 3792 24142 3844 24148
rect 3700 22432 3752 22438
rect 3700 22374 3752 22380
rect 3712 21486 3740 22374
rect 3804 22030 3832 24142
rect 5264 24132 5316 24138
rect 5264 24074 5316 24080
rect 5276 23866 5304 24074
rect 5264 23860 5316 23866
rect 5264 23802 5316 23808
rect 5120 23420 5428 23440
rect 5120 23418 5126 23420
rect 5182 23418 5206 23420
rect 5262 23418 5286 23420
rect 5342 23418 5366 23420
rect 5422 23418 5428 23420
rect 5182 23366 5184 23418
rect 5364 23366 5366 23418
rect 5120 23364 5126 23366
rect 5182 23364 5206 23366
rect 5262 23364 5286 23366
rect 5342 23364 5366 23366
rect 5422 23364 5428 23366
rect 5120 23344 5428 23364
rect 3976 22636 4028 22642
rect 3976 22578 4028 22584
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 3988 21622 4016 22578
rect 4344 22568 4396 22574
rect 4344 22510 4396 22516
rect 4160 21956 4212 21962
rect 4160 21898 4212 21904
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 3700 21480 3752 21486
rect 3700 21422 3752 21428
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 3792 20800 3844 20806
rect 3792 20742 3844 20748
rect 3804 20398 3832 20742
rect 3896 20466 3924 21422
rect 3988 21146 4016 21558
rect 4172 21146 4200 21898
rect 4356 21894 4384 22510
rect 5120 22332 5428 22352
rect 5120 22330 5126 22332
rect 5182 22330 5206 22332
rect 5262 22330 5286 22332
rect 5342 22330 5366 22332
rect 5422 22330 5428 22332
rect 5182 22278 5184 22330
rect 5364 22278 5366 22330
rect 5120 22276 5126 22278
rect 5182 22276 5206 22278
rect 5262 22276 5286 22278
rect 5342 22276 5366 22278
rect 5422 22276 5428 22278
rect 5120 22256 5428 22276
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 4160 21140 4212 21146
rect 4160 21082 4212 21088
rect 4356 20942 4384 21830
rect 4816 21690 4844 21966
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4436 21548 4488 21554
rect 4436 21490 4488 21496
rect 4448 21078 4476 21490
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4632 21146 4660 21286
rect 4620 21140 4672 21146
rect 4620 21082 4672 21088
rect 4436 21072 4488 21078
rect 4436 21014 4488 21020
rect 4448 20942 4476 21014
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3896 19990 3924 20402
rect 4080 20058 4108 20878
rect 4448 20602 4476 20878
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 3884 19984 3936 19990
rect 3884 19926 3936 19932
rect 3896 19514 3924 19926
rect 4172 19854 4200 20266
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 4172 19378 4200 19790
rect 4436 19780 4488 19786
rect 4436 19722 4488 19728
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4264 19310 4292 19654
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4356 19378 4384 19450
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3712 16454 3740 18362
rect 3804 18290 3832 18566
rect 4264 18290 4292 18702
rect 3792 18284 3844 18290
rect 3792 18226 3844 18232
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 3792 18080 3844 18086
rect 3792 18022 3844 18028
rect 3804 17746 3832 18022
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3792 17740 3844 17746
rect 3792 17682 3844 17688
rect 3804 16522 3832 17682
rect 3884 17536 3936 17542
rect 4080 17513 4108 17750
rect 4160 17604 4212 17610
rect 4160 17546 4212 17552
rect 3884 17478 3936 17484
rect 4066 17504 4122 17513
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 3240 15496 3292 15502
rect 3516 15496 3568 15502
rect 3240 15438 3292 15444
rect 3344 15456 3516 15484
rect 3068 15162 3096 15438
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 3252 14958 3280 15438
rect 3240 14952 3292 14958
rect 3068 14900 3240 14906
rect 3068 14894 3292 14900
rect 3068 14878 3280 14894
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2424 13326 2452 14554
rect 3068 14482 3096 14878
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 1688 12782 1716 13262
rect 2700 13258 2728 14214
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 2792 12918 2820 13738
rect 2884 13190 2912 14350
rect 2976 14074 3004 14350
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2976 12986 3004 13874
rect 3068 13870 3096 14418
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3160 13530 3188 14350
rect 3344 14328 3372 15456
rect 3516 15438 3568 15444
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3422 14648 3478 14657
rect 3422 14583 3478 14592
rect 3252 14300 3372 14328
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 11014 1716 12718
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 1780 11354 1808 11698
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1688 10606 1716 10950
rect 2516 10742 2544 11494
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1688 9042 1716 10542
rect 2608 10062 2636 11698
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2792 10146 2820 11630
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2700 10130 2820 10146
rect 2884 10130 2912 10474
rect 2688 10124 2820 10130
rect 2740 10118 2820 10124
rect 2688 10066 2740 10072
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2608 9738 2636 9998
rect 2608 9710 2728 9738
rect 2792 9722 2820 10118
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2700 9602 2728 9710
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1964 8974 1992 9318
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 2148 7546 2176 7754
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2332 7410 2360 9590
rect 2700 9574 2820 9602
rect 2884 9586 2912 10066
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 2608 8634 2636 9386
rect 2792 9382 2820 9574
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2976 9432 3004 12922
rect 3252 11898 3280 14300
rect 3436 14278 3464 14583
rect 3528 14346 3556 14962
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3528 13938 3556 14282
rect 3620 14074 3648 14962
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3712 13938 3740 16390
rect 3804 16046 3832 16458
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3896 15978 3924 17478
rect 4066 17439 4122 17448
rect 4172 17338 4200 17546
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 3988 16590 4016 17274
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4080 16590 4108 17206
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3804 14958 3832 15506
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3804 14074 3832 14894
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3344 12986 3372 13874
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3896 12918 3924 15914
rect 3988 13394 4016 16526
rect 4080 16250 4108 16526
rect 4356 16436 4384 18158
rect 4448 16590 4476 19722
rect 4528 18148 4580 18154
rect 4528 18090 4580 18096
rect 4540 17542 4568 18090
rect 4632 17610 4660 20810
rect 4724 20602 4752 20946
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 4816 18290 4844 21626
rect 5368 21554 5396 21830
rect 5736 21570 5764 28750
rect 6380 28642 6408 28750
rect 6458 28642 6514 29442
rect 7654 28642 7710 29442
rect 8850 28642 8906 29442
rect 10046 28642 10102 29442
rect 11242 28642 11298 29442
rect 11348 28750 12112 28778
rect 11348 28642 11376 28750
rect 6380 28614 6500 28642
rect 6920 25832 6972 25838
rect 6920 25774 6972 25780
rect 6932 25498 6960 25774
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7564 25696 7616 25702
rect 7564 25638 7616 25644
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 6644 25220 6696 25226
rect 6644 25162 6696 25168
rect 6368 24404 6420 24410
rect 6368 24346 6420 24352
rect 5908 24132 5960 24138
rect 5908 24074 5960 24080
rect 5920 23866 5948 24074
rect 5908 23860 5960 23866
rect 5908 23802 5960 23808
rect 6380 23730 6408 24346
rect 6656 23730 6684 25162
rect 6932 24834 6960 25434
rect 7208 25430 7236 25638
rect 7196 25424 7248 25430
rect 7196 25366 7248 25372
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6840 24806 6960 24834
rect 7116 24818 7144 25230
rect 7208 25226 7236 25366
rect 7288 25356 7340 25362
rect 7288 25298 7340 25304
rect 7196 25220 7248 25226
rect 7196 25162 7248 25168
rect 7300 24818 7328 25298
rect 7576 25294 7604 25638
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7380 25220 7432 25226
rect 7380 25162 7432 25168
rect 7104 24812 7156 24818
rect 6748 24070 6776 24754
rect 6840 24138 6868 24806
rect 7104 24754 7156 24760
rect 7288 24812 7340 24818
rect 7288 24754 7340 24760
rect 7116 24410 7144 24754
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 7104 24404 7156 24410
rect 7208 24392 7236 24686
rect 7288 24404 7340 24410
rect 7208 24364 7288 24392
rect 7104 24346 7156 24352
rect 7288 24346 7340 24352
rect 6828 24132 6880 24138
rect 6828 24074 6880 24080
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6368 23724 6420 23730
rect 6368 23666 6420 23672
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 5816 23656 5868 23662
rect 5816 23598 5868 23604
rect 5828 23322 5856 23598
rect 5816 23316 5868 23322
rect 5816 23258 5868 23264
rect 6656 22982 6684 23666
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6748 23118 6776 23462
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 6288 22166 6316 22918
rect 6840 22438 6868 24074
rect 7116 23050 7144 24346
rect 7392 24206 7420 25162
rect 7668 24834 7696 28642
rect 11256 28614 11376 28642
rect 9291 27228 9599 27248
rect 9291 27226 9297 27228
rect 9353 27226 9377 27228
rect 9433 27226 9457 27228
rect 9513 27226 9537 27228
rect 9593 27226 9599 27228
rect 9353 27174 9355 27226
rect 9535 27174 9537 27226
rect 9291 27172 9297 27174
rect 9353 27172 9377 27174
rect 9433 27172 9457 27174
rect 9513 27172 9537 27174
rect 9593 27172 9599 27174
rect 9291 27152 9599 27172
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 9291 26140 9599 26160
rect 9291 26138 9297 26140
rect 9353 26138 9377 26140
rect 9433 26138 9457 26140
rect 9513 26138 9537 26140
rect 9593 26138 9599 26140
rect 9353 26086 9355 26138
rect 9535 26086 9537 26138
rect 9291 26084 9297 26086
rect 9353 26084 9377 26086
rect 9433 26084 9457 26086
rect 9513 26084 9537 26086
rect 9593 26084 9599 26086
rect 9291 26064 9599 26084
rect 11612 26036 11664 26042
rect 11612 25978 11664 25984
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 11060 25900 11112 25906
rect 11060 25842 11112 25848
rect 11152 25900 11204 25906
rect 11152 25842 11204 25848
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 7852 24954 7880 25230
rect 7944 24954 7972 25842
rect 8852 25696 8904 25702
rect 8852 25638 8904 25644
rect 10692 25696 10744 25702
rect 10692 25638 10744 25644
rect 8208 25356 8260 25362
rect 8208 25298 8260 25304
rect 8116 25220 8168 25226
rect 8116 25162 8168 25168
rect 8128 24954 8156 25162
rect 7840 24948 7892 24954
rect 7840 24890 7892 24896
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 8116 24948 8168 24954
rect 8116 24890 8168 24896
rect 7484 24806 7696 24834
rect 7748 24880 7800 24886
rect 7748 24822 7800 24828
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 7104 23044 7156 23050
rect 7104 22986 7156 22992
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 7024 22778 7052 22918
rect 7012 22772 7064 22778
rect 7012 22714 7064 22720
rect 7116 22710 7144 22986
rect 7104 22704 7156 22710
rect 7104 22646 7156 22652
rect 6828 22432 6880 22438
rect 6828 22374 6880 22380
rect 5816 22160 5868 22166
rect 5816 22102 5868 22108
rect 6276 22160 6328 22166
rect 6276 22102 6328 22108
rect 5828 21690 5856 22102
rect 6000 21956 6052 21962
rect 6000 21898 6052 21904
rect 6012 21729 6040 21898
rect 5998 21720 6054 21729
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5908 21684 5960 21690
rect 5998 21655 6054 21664
rect 5908 21626 5960 21632
rect 5356 21548 5408 21554
rect 5736 21542 5856 21570
rect 5356 21490 5408 21496
rect 5724 21480 5776 21486
rect 5644 21428 5724 21434
rect 5644 21422 5776 21428
rect 5644 21406 5764 21422
rect 5120 21244 5428 21264
rect 5120 21242 5126 21244
rect 5182 21242 5206 21244
rect 5262 21242 5286 21244
rect 5342 21242 5366 21244
rect 5422 21242 5428 21244
rect 5182 21190 5184 21242
rect 5364 21190 5366 21242
rect 5120 21188 5126 21190
rect 5182 21188 5206 21190
rect 5262 21188 5286 21190
rect 5342 21188 5366 21190
rect 5422 21188 5428 21190
rect 5120 21168 5428 21188
rect 5644 20874 5672 21406
rect 5828 21162 5856 21542
rect 5736 21134 5856 21162
rect 5632 20868 5684 20874
rect 5632 20810 5684 20816
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5552 20482 5580 20742
rect 5460 20466 5580 20482
rect 5448 20460 5580 20466
rect 5500 20454 5580 20460
rect 5448 20402 5500 20408
rect 5120 20156 5428 20176
rect 5120 20154 5126 20156
rect 5182 20154 5206 20156
rect 5262 20154 5286 20156
rect 5342 20154 5366 20156
rect 5422 20154 5428 20156
rect 5182 20102 5184 20154
rect 5364 20102 5366 20154
rect 5120 20100 5126 20102
rect 5182 20100 5206 20102
rect 5262 20100 5286 20102
rect 5342 20100 5366 20102
rect 5422 20100 5428 20102
rect 5120 20080 5428 20100
rect 5552 19378 5580 20454
rect 5644 19938 5672 20810
rect 5736 20618 5764 21134
rect 5920 21026 5948 21626
rect 5828 20998 5948 21026
rect 5828 20942 5856 20998
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5736 20590 6224 20618
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5736 20058 5764 20402
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5644 19910 5764 19938
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 5120 19068 5428 19088
rect 5120 19066 5126 19068
rect 5182 19066 5206 19068
rect 5262 19066 5286 19068
rect 5342 19066 5366 19068
rect 5422 19066 5428 19068
rect 5182 19014 5184 19066
rect 5364 19014 5366 19066
rect 5120 19012 5126 19014
rect 5182 19012 5206 19014
rect 5262 19012 5286 19014
rect 5342 19012 5366 19014
rect 5422 19012 5428 19014
rect 5120 18992 5428 19012
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 4908 18290 4936 18906
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 5184 18290 5212 18634
rect 5460 18290 5488 19178
rect 5644 18902 5672 19450
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 5172 18284 5224 18290
rect 5172 18226 5224 18232
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5552 18154 5580 18362
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5120 17980 5428 18000
rect 5120 17978 5126 17980
rect 5182 17978 5206 17980
rect 5262 17978 5286 17980
rect 5342 17978 5366 17980
rect 5422 17978 5428 17980
rect 5182 17926 5184 17978
rect 5364 17926 5366 17978
rect 5120 17924 5126 17926
rect 5182 17924 5206 17926
rect 5262 17924 5286 17926
rect 5342 17924 5366 17926
rect 5422 17924 5428 17926
rect 5120 17904 5428 17924
rect 5460 17882 5488 18090
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5460 17746 5488 17818
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5552 17678 5580 18090
rect 5644 17678 5672 18702
rect 5736 18426 5764 19910
rect 6000 19440 6052 19446
rect 6000 19382 6052 19388
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5828 18222 5856 19246
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 5920 18290 5948 18906
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5828 17678 5856 18022
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 4620 17604 4672 17610
rect 4620 17546 4672 17552
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4540 16436 4568 17478
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4620 16448 4672 16454
rect 4356 16408 4476 16436
rect 4540 16408 4620 16436
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4066 16144 4122 16153
rect 4066 16079 4122 16088
rect 4080 15502 4108 16079
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4264 15162 4292 15370
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4080 14414 4108 14758
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 4172 13530 4200 13738
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4356 13394 4384 13806
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 3988 12434 4016 13126
rect 4356 12782 4384 13330
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 3528 12406 4016 12434
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 3068 9761 3096 10950
rect 3160 10742 3188 11698
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3148 10736 3200 10742
rect 3148 10678 3200 10684
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3252 10062 3280 10406
rect 3344 10266 3372 11086
rect 3436 10674 3464 11562
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3436 10198 3464 10610
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3054 9752 3110 9761
rect 3054 9687 3110 9696
rect 3068 9654 3096 9687
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3252 9586 3280 9998
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 2884 9404 3004 9432
rect 3148 9444 3200 9450
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2332 7206 2360 7346
rect 572 7200 624 7206
rect 572 7142 624 7148
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 584 800 612 7142
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2056 5574 2084 6258
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2332 5710 2360 6054
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2056 4622 2084 5510
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 2056 3505 2084 4558
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2042 3496 2098 3505
rect 1676 3460 1728 3466
rect 2042 3431 2098 3440
rect 1676 3402 1728 3408
rect 1688 800 1716 3402
rect 2792 2145 2820 3606
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 2884 800 2912 9404
rect 3148 9386 3200 9392
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3068 8498 3096 8910
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3068 8090 3096 8434
rect 3160 8294 3188 9386
rect 3252 8906 3280 9522
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3252 8498 3280 8842
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3068 7886 3096 8026
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3068 7410 3096 7822
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3252 7274 3280 8298
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 7410 3372 8230
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3436 7478 3464 7686
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3344 7290 3372 7346
rect 3240 7268 3292 7274
rect 3344 7262 3464 7290
rect 3240 7210 3292 7216
rect 3252 6390 3280 7210
rect 3436 6662 3464 7262
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3068 5914 3096 6258
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3344 5302 3372 6258
rect 3436 6254 3464 6598
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 3528 4865 3556 12406
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3804 10674 3832 11630
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3620 10062 3648 10542
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3620 9178 3648 9998
rect 3804 9926 3832 10066
rect 4172 9926 4200 10610
rect 4264 10062 4292 10678
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 4356 10130 4384 10474
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3712 8974 3740 9318
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3804 7954 3832 9862
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3896 9042 3924 9454
rect 3974 9072 4030 9081
rect 3884 9036 3936 9042
rect 3974 9007 3976 9016
rect 3884 8978 3936 8984
rect 4028 9007 4030 9016
rect 3976 8978 4028 8984
rect 3896 8634 3924 8978
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 4080 8498 4108 9590
rect 4264 9518 4292 9998
rect 4356 9654 4384 10066
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4448 9450 4476 16408
rect 4620 16390 4672 16396
rect 4632 16114 4660 16390
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4724 15162 4752 16934
rect 4908 16590 4936 17478
rect 5120 16892 5428 16912
rect 5120 16890 5126 16892
rect 5182 16890 5206 16892
rect 5262 16890 5286 16892
rect 5342 16890 5366 16892
rect 5422 16890 5428 16892
rect 5182 16838 5184 16890
rect 5364 16838 5366 16890
rect 5120 16836 5126 16838
rect 5182 16836 5206 16838
rect 5262 16836 5286 16838
rect 5342 16836 5366 16838
rect 5422 16836 5428 16838
rect 5120 16816 5428 16836
rect 5644 16794 5672 17614
rect 5724 17196 5776 17202
rect 6012 17184 6040 19382
rect 6092 17604 6144 17610
rect 6092 17546 6144 17552
rect 5776 17156 6040 17184
rect 5724 17138 5776 17144
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4804 16516 4856 16522
rect 4804 16458 4856 16464
rect 4816 15706 4844 16458
rect 5120 15804 5428 15824
rect 5120 15802 5126 15804
rect 5182 15802 5206 15804
rect 5262 15802 5286 15804
rect 5342 15802 5366 15804
rect 5422 15802 5428 15804
rect 5182 15750 5184 15802
rect 5364 15750 5366 15802
rect 5120 15748 5126 15750
rect 5182 15748 5206 15750
rect 5262 15748 5286 15750
rect 5342 15748 5366 15750
rect 5422 15748 5428 15750
rect 5120 15728 5428 15748
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 5644 15570 5672 16730
rect 6104 16454 6132 17546
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4540 13870 4568 14894
rect 4528 13864 4580 13870
rect 4526 13832 4528 13841
rect 4580 13832 4582 13841
rect 4526 13767 4582 13776
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4540 10470 4568 10610
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4632 10282 4660 14962
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5120 14716 5428 14736
rect 5120 14714 5126 14716
rect 5182 14714 5206 14716
rect 5262 14714 5286 14716
rect 5342 14714 5366 14716
rect 5422 14714 5428 14716
rect 5182 14662 5184 14714
rect 5364 14662 5366 14714
rect 5120 14660 5126 14662
rect 5182 14660 5206 14662
rect 5262 14660 5286 14662
rect 5342 14660 5366 14662
rect 5422 14660 5428 14662
rect 5120 14640 5428 14660
rect 5552 14618 5580 14826
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 6092 14612 6144 14618
rect 6196 14600 6224 20590
rect 6288 20058 6316 22102
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6368 21888 6420 21894
rect 6368 21830 6420 21836
rect 6380 21486 6408 21830
rect 6460 21548 6512 21554
rect 6460 21490 6512 21496
rect 6368 21480 6420 21486
rect 6368 21422 6420 21428
rect 6472 20942 6500 21490
rect 6656 21146 6684 21966
rect 6840 21418 6868 22374
rect 6920 22092 6972 22098
rect 6920 22034 6972 22040
rect 6828 21412 6880 21418
rect 6828 21354 6880 21360
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 6656 21010 6684 21082
rect 6840 21078 6868 21354
rect 6828 21072 6880 21078
rect 6828 21014 6880 21020
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 6932 20942 6960 22034
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 7024 21418 7052 21490
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 6380 20398 6408 20878
rect 6932 20534 6960 20878
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6288 16998 6316 19450
rect 6380 19446 6408 20334
rect 6368 19440 6420 19446
rect 6368 19382 6420 19388
rect 6656 19378 6960 19394
rect 7024 19378 7052 20538
rect 7116 20262 7144 21286
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 7300 19718 7328 23734
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7392 22778 7420 23054
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7484 22094 7512 24806
rect 7760 24698 7788 24822
rect 8220 24818 8248 25298
rect 8392 25152 8444 25158
rect 8392 25094 8444 25100
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 7668 24670 7788 24698
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7576 24070 7604 24346
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7392 22066 7512 22094
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 6644 19372 6960 19378
rect 6696 19366 6960 19372
rect 6644 19314 6696 19320
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6840 19174 6868 19246
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6472 18766 6500 19110
rect 6840 18970 6868 19110
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6932 18630 6960 19366
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 7116 19242 7144 19654
rect 7300 19310 7328 19654
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7104 19236 7156 19242
rect 7104 19178 7156 19184
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6840 17610 6868 18566
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6840 17134 6868 17546
rect 7116 17542 7144 18634
rect 7208 18358 7236 18702
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6288 14618 6316 15370
rect 6564 15026 6592 15642
rect 6552 15020 6604 15026
rect 6380 14980 6552 15008
rect 6144 14572 6224 14600
rect 6276 14612 6328 14618
rect 6092 14554 6144 14560
rect 6276 14554 6328 14560
rect 5906 14512 5962 14521
rect 5827 14470 5906 14498
rect 6380 14498 6408 14980
rect 6552 14962 6604 14968
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 5632 14408 5684 14414
rect 5827 14396 5855 14470
rect 5906 14447 5908 14456
rect 5960 14447 5962 14456
rect 6196 14470 6408 14498
rect 5908 14418 5960 14424
rect 6196 14414 6224 14470
rect 6184 14408 6236 14414
rect 5827 14368 5856 14396
rect 5632 14350 5684 14356
rect 5644 14074 5672 14350
rect 5828 14090 5856 14368
rect 6184 14350 6236 14356
rect 5908 14340 5960 14346
rect 5960 14300 6040 14328
rect 5908 14282 5960 14288
rect 5828 14074 5948 14090
rect 6012 14074 6040 14300
rect 5632 14068 5684 14074
rect 5828 14068 5960 14074
rect 5828 14062 5908 14068
rect 5632 14010 5684 14016
rect 5908 14010 5960 14016
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 4896 14000 4948 14006
rect 4710 13968 4766 13977
rect 4896 13942 4948 13948
rect 5722 13968 5778 13977
rect 4766 13912 4844 13920
rect 4710 13903 4712 13912
rect 4764 13892 4844 13912
rect 4712 13874 4764 13880
rect 4816 13326 4844 13892
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4724 12850 4752 13262
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4724 11830 4752 12786
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 4724 11218 4752 11766
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4540 10254 4660 10282
rect 4540 10062 4568 10254
rect 4724 10130 4752 11154
rect 4908 11150 4936 13942
rect 5722 13906 5724 13912
rect 5776 13906 5778 13912
rect 5722 13903 5778 13906
rect 5724 13900 5776 13903
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5120 13628 5428 13648
rect 5120 13626 5126 13628
rect 5182 13626 5206 13628
rect 5262 13626 5286 13628
rect 5342 13626 5366 13628
rect 5422 13626 5428 13628
rect 5182 13574 5184 13626
rect 5364 13574 5366 13626
rect 5120 13572 5126 13574
rect 5182 13572 5206 13574
rect 5262 13572 5286 13574
rect 5342 13572 5366 13574
rect 5422 13572 5428 13574
rect 5120 13552 5428 13572
rect 5460 13433 5488 13738
rect 5446 13424 5502 13433
rect 5446 13359 5502 13368
rect 5814 13424 5870 13433
rect 5920 13394 5948 14010
rect 6564 13938 6592 14758
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6734 14512 6790 14521
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13530 6224 13670
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 5814 13359 5870 13368
rect 5908 13388 5960 13394
rect 5828 13326 5856 13359
rect 5908 13330 5960 13336
rect 6196 13326 6224 13466
rect 6656 13433 6684 14486
rect 6734 14447 6736 14456
rect 6788 14447 6790 14456
rect 6736 14418 6788 14424
rect 6642 13424 6698 13433
rect 6642 13359 6698 13368
rect 6656 13326 6684 13359
rect 6748 13326 6776 14418
rect 6840 14074 6868 16390
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6932 14600 6960 14962
rect 7012 14612 7064 14618
rect 6932 14572 7012 14600
rect 7012 14554 7064 14560
rect 7116 14482 7144 17478
rect 7300 15366 7328 19246
rect 7392 17252 7420 22066
rect 7576 21690 7604 24006
rect 7668 23662 7696 24670
rect 7852 24614 7880 24686
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8128 24342 8156 24550
rect 7840 24336 7892 24342
rect 7840 24278 7892 24284
rect 8116 24336 8168 24342
rect 8116 24278 8168 24284
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7668 23118 7696 23598
rect 7760 23322 7788 23666
rect 7852 23474 7880 24278
rect 8024 24200 8076 24206
rect 8220 24188 8248 24754
rect 8404 24274 8432 25094
rect 8484 24880 8536 24886
rect 8484 24822 8536 24828
rect 8392 24268 8444 24274
rect 8392 24210 8444 24216
rect 8024 24142 8076 24148
rect 8128 24160 8248 24188
rect 7932 24064 7984 24070
rect 7932 24006 7984 24012
rect 7944 23798 7972 24006
rect 8036 23866 8064 24142
rect 8024 23860 8076 23866
rect 8024 23802 8076 23808
rect 7932 23792 7984 23798
rect 7932 23734 7984 23740
rect 8022 23760 8078 23769
rect 8022 23695 8024 23704
rect 8076 23695 8078 23704
rect 8024 23666 8076 23672
rect 8024 23588 8076 23594
rect 8128 23576 8156 24160
rect 8392 24132 8444 24138
rect 8392 24074 8444 24080
rect 8404 23866 8432 24074
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8392 23860 8444 23866
rect 8392 23802 8444 23808
rect 8076 23548 8156 23576
rect 8024 23530 8076 23536
rect 7852 23446 7972 23474
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 7748 23180 7800 23186
rect 7748 23122 7800 23128
rect 7656 23112 7708 23118
rect 7656 23054 7708 23060
rect 7668 22234 7696 23054
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 7576 21570 7604 21626
rect 7484 21542 7604 21570
rect 7760 21554 7788 23122
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7656 21548 7708 21554
rect 7484 20942 7512 21542
rect 7656 21490 7708 21496
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7472 19236 7524 19242
rect 7472 19178 7524 19184
rect 7484 18698 7512 19178
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7392 17224 7512 17252
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7392 14618 7420 15846
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6920 13864 6972 13870
rect 6918 13832 6920 13841
rect 6972 13832 6974 13841
rect 6918 13767 6974 13776
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 13326 6960 13670
rect 7104 13524 7156 13530
rect 7208 13512 7236 14486
rect 7300 14346 7328 14554
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7156 13484 7236 13512
rect 7104 13466 7156 13472
rect 7012 13456 7064 13462
rect 7116 13433 7144 13466
rect 7012 13398 7064 13404
rect 7102 13424 7158 13433
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5120 12540 5428 12560
rect 5120 12538 5126 12540
rect 5182 12538 5206 12540
rect 5262 12538 5286 12540
rect 5342 12538 5366 12540
rect 5422 12538 5428 12540
rect 5182 12486 5184 12538
rect 5364 12486 5366 12538
rect 5120 12484 5126 12486
rect 5182 12484 5206 12486
rect 5262 12484 5286 12486
rect 5342 12484 5366 12486
rect 5422 12484 5428 12486
rect 5120 12464 5428 12484
rect 5120 11452 5428 11472
rect 5120 11450 5126 11452
rect 5182 11450 5206 11452
rect 5262 11450 5286 11452
rect 5342 11450 5366 11452
rect 5422 11450 5428 11452
rect 5182 11398 5184 11450
rect 5364 11398 5366 11450
rect 5120 11396 5126 11398
rect 5182 11396 5206 11398
rect 5262 11396 5286 11398
rect 5342 11396 5366 11398
rect 5422 11396 5428 11398
rect 5120 11376 5428 11396
rect 5460 11257 5488 12922
rect 5552 12850 5580 13126
rect 5644 12986 5672 13262
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5446 11248 5502 11257
rect 5446 11183 5502 11192
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4908 10674 4936 11086
rect 4988 10736 5040 10742
rect 4986 10704 4988 10713
rect 5040 10704 5042 10713
rect 4896 10668 4948 10674
rect 5460 10674 5488 11183
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5644 10742 5672 11018
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5736 10674 5764 10950
rect 5828 10810 5856 11018
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 6012 10713 6040 11494
rect 5998 10704 6054 10713
rect 4986 10639 5042 10648
rect 5448 10668 5500 10674
rect 4896 10610 4948 10616
rect 5448 10610 5500 10616
rect 5724 10668 5776 10674
rect 5998 10639 6054 10648
rect 5724 10610 5776 10616
rect 5120 10364 5428 10384
rect 5120 10362 5126 10364
rect 5182 10362 5206 10364
rect 5262 10362 5286 10364
rect 5342 10362 5366 10364
rect 5422 10362 5428 10364
rect 5182 10310 5184 10362
rect 5364 10310 5366 10362
rect 5120 10308 5126 10310
rect 5182 10308 5206 10310
rect 5262 10308 5286 10310
rect 5342 10308 5366 10310
rect 5422 10308 5428 10310
rect 5120 10288 5428 10308
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4540 9926 4568 9998
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4632 9874 4660 9930
rect 4632 9846 4752 9874
rect 4724 9586 4752 9846
rect 5552 9654 5580 9930
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 9722 5672 9862
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4724 9450 4752 9522
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4816 9382 4844 9522
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3804 7750 3832 7890
rect 4068 7880 4120 7886
rect 4172 7834 4200 8434
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4356 7954 4384 8230
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4120 7828 4200 7834
rect 4068 7822 4200 7828
rect 4080 7806 4200 7822
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 3620 6322 3648 7210
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3514 4856 3570 4865
rect 3514 4791 3570 4800
rect 3804 3466 3832 7686
rect 4068 6384 4120 6390
rect 4066 6352 4068 6361
rect 4120 6352 4122 6361
rect 4172 6322 4200 7806
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4356 7410 4384 7754
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4356 6866 4384 7346
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4066 6287 4122 6296
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4356 6186 4384 6802
rect 4540 6390 4568 9318
rect 5120 9276 5428 9296
rect 5120 9274 5126 9276
rect 5182 9274 5206 9276
rect 5262 9274 5286 9276
rect 5342 9274 5366 9276
rect 5422 9274 5428 9276
rect 5182 9222 5184 9274
rect 5364 9222 5366 9274
rect 5120 9220 5126 9222
rect 5182 9220 5206 9222
rect 5262 9220 5286 9222
rect 5342 9220 5366 9222
rect 5422 9220 5428 9222
rect 5120 9200 5428 9220
rect 5356 8492 5408 8498
rect 5460 8480 5488 9318
rect 5408 8452 5488 8480
rect 5356 8434 5408 8440
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5120 8188 5428 8208
rect 5120 8186 5126 8188
rect 5182 8186 5206 8188
rect 5262 8186 5286 8188
rect 5342 8186 5366 8188
rect 5422 8186 5428 8188
rect 5182 8134 5184 8186
rect 5364 8134 5366 8186
rect 5120 8132 5126 8134
rect 5182 8132 5206 8134
rect 5262 8132 5286 8134
rect 5342 8132 5366 8134
rect 5422 8132 5428 8134
rect 5120 8112 5428 8132
rect 5644 8090 5672 8366
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5736 7970 5764 10610
rect 6012 10606 6040 10639
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6104 8634 6132 10406
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5644 7942 5764 7970
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4724 7478 4752 7686
rect 4816 7546 4844 7822
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4356 5778 4384 6122
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 5234 4384 5714
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 3896 5030 3924 5170
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 4356 4842 4384 5170
rect 4816 5166 4844 7482
rect 5644 7206 5672 7942
rect 5920 7750 5948 8434
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 6012 7818 6040 8298
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 5908 7744 5960 7750
rect 5960 7692 6040 7698
rect 5908 7686 6040 7692
rect 5920 7670 6040 7686
rect 5920 7621 5948 7670
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5120 7100 5428 7120
rect 5120 7098 5126 7100
rect 5182 7098 5206 7100
rect 5262 7098 5286 7100
rect 5342 7098 5366 7100
rect 5422 7098 5428 7100
rect 5182 7046 5184 7098
rect 5364 7046 5366 7098
rect 5120 7044 5126 7046
rect 5182 7044 5206 7046
rect 5262 7044 5286 7046
rect 5342 7044 5366 7046
rect 5422 7044 5428 7046
rect 5120 7024 5428 7044
rect 5644 6866 5672 7142
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5552 6458 5580 6666
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5120 6012 5428 6032
rect 5120 6010 5126 6012
rect 5182 6010 5206 6012
rect 5262 6010 5286 6012
rect 5342 6010 5366 6012
rect 5422 6010 5428 6012
rect 5182 5958 5184 6010
rect 5364 5958 5366 6010
rect 5120 5956 5126 5958
rect 5182 5956 5206 5958
rect 5262 5956 5286 5958
rect 5342 5956 5366 5958
rect 5422 5956 5428 5958
rect 5120 5936 5428 5956
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4908 5234 4936 5510
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 5120 4924 5428 4944
rect 5120 4922 5126 4924
rect 5182 4922 5206 4924
rect 5262 4922 5286 4924
rect 5342 4922 5366 4924
rect 5422 4922 5428 4924
rect 5182 4870 5184 4922
rect 5364 4870 5366 4922
rect 5120 4868 5126 4870
rect 5182 4868 5206 4870
rect 5262 4868 5286 4870
rect 5342 4868 5366 4870
rect 5422 4868 5428 4870
rect 5120 4848 5428 4868
rect 4264 4826 4384 4842
rect 5460 4826 5488 5238
rect 4252 4820 4384 4826
rect 4304 4814 4384 4820
rect 4252 4762 4304 4768
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 3148 1352 3200 1358
rect 3148 1294 3200 1300
rect 570 0 626 800
rect 1674 0 1730 800
rect 2870 0 2926 800
rect 3160 785 3188 1294
rect 4080 800 4108 3674
rect 4356 3602 4384 4814
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4816 4282 4844 4490
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5000 4146 5028 4422
rect 5460 4146 5488 4762
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5552 4078 5580 5646
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5120 3836 5428 3856
rect 5120 3834 5126 3836
rect 5182 3834 5206 3836
rect 5262 3834 5286 3836
rect 5342 3834 5366 3836
rect 5422 3834 5428 3836
rect 5182 3782 5184 3834
rect 5364 3782 5366 3834
rect 5120 3780 5126 3782
rect 5182 3780 5206 3782
rect 5262 3780 5286 3782
rect 5342 3780 5366 3782
rect 5422 3780 5428 3782
rect 5120 3760 5428 3780
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4816 3194 4844 3402
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5460 3126 5488 3878
rect 5644 3738 5672 6802
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6338 5948 6598
rect 5828 6322 5948 6338
rect 5816 6316 5948 6322
rect 5868 6310 5948 6316
rect 5816 6258 5868 6264
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5736 5166 5764 5510
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5828 4826 5856 4966
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5736 3738 5764 4422
rect 5828 4282 5856 4762
rect 5920 4690 5948 6310
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 6012 4282 6040 7670
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5828 4026 5856 4218
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 5828 3998 5948 4026
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5448 3120 5500 3126
rect 5736 3074 5764 3674
rect 5448 3062 5500 3068
rect 5644 3058 5764 3074
rect 5828 3058 5856 3878
rect 5920 3126 5948 3998
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 6012 3194 6040 3402
rect 6104 3398 6132 4082
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 5632 3052 5764 3058
rect 5684 3046 5764 3052
rect 5816 3052 5868 3058
rect 5632 2994 5684 3000
rect 5816 2994 5868 3000
rect 5920 2922 5948 3062
rect 6104 2990 6132 3334
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 5120 2748 5428 2768
rect 5120 2746 5126 2748
rect 5182 2746 5206 2748
rect 5262 2746 5286 2748
rect 5342 2746 5366 2748
rect 5422 2746 5428 2748
rect 5182 2694 5184 2746
rect 5364 2694 5366 2746
rect 5120 2692 5126 2694
rect 5182 2692 5206 2694
rect 5262 2692 5286 2694
rect 5342 2692 5366 2694
rect 5422 2692 5428 2694
rect 5120 2672 5428 2692
rect 3146 776 3202 785
rect 3146 711 3202 720
rect 4066 0 4122 800
rect 5262 0 5318 800
rect 6196 762 6224 12922
rect 6472 12850 6500 13126
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6564 11762 6592 12174
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6840 11354 6868 12038
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6748 11150 6776 11222
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 9722 6776 11086
rect 6840 10674 6868 11290
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6932 10577 6960 11494
rect 6918 10568 6974 10577
rect 6918 10503 6974 10512
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6932 8922 6960 10503
rect 7024 9926 7052 13398
rect 7102 13359 7158 13368
rect 7116 13326 7144 13359
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7196 11824 7248 11830
rect 7196 11766 7248 11772
rect 7208 10810 7236 11766
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7300 10266 7328 13874
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7392 12986 7420 13330
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7024 9518 7052 9862
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7116 9042 7144 9454
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 6932 8894 7052 8922
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8566 6960 8774
rect 7024 8566 7052 8894
rect 7116 8634 7144 8978
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6380 6798 6408 8366
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6472 6866 6500 8026
rect 6656 7886 6684 8298
rect 6748 8090 6776 8366
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6932 7886 6960 8502
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7024 7886 7052 8026
rect 7116 7954 7144 8570
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7024 7732 7052 7822
rect 6932 7704 7052 7732
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6380 6390 6408 6734
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 6472 6254 6500 6802
rect 6748 6798 6776 7142
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 5030 6316 5510
rect 6380 5234 6408 6122
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 4622 6316 4966
rect 6564 4758 6592 5578
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6656 4826 6684 5170
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6288 4146 6316 4558
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6288 3194 6316 4082
rect 6748 4078 6776 6734
rect 6932 6730 6960 7704
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7024 6866 7052 7346
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7392 6746 7420 12922
rect 7484 10606 7512 17224
rect 7576 16998 7604 21354
rect 7668 21078 7696 21490
rect 7760 21146 7788 21490
rect 7852 21350 7880 22578
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7656 21072 7708 21078
rect 7656 21014 7708 21020
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7668 20602 7696 20878
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7944 20346 7972 23446
rect 8116 23316 8168 23322
rect 8116 23258 8168 23264
rect 8128 22234 8156 23258
rect 8220 23118 8248 23802
rect 8298 23760 8354 23769
rect 8298 23695 8354 23704
rect 8312 23186 8340 23695
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8312 23050 8340 23122
rect 8300 23044 8352 23050
rect 8300 22986 8352 22992
rect 8312 22778 8340 22986
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8404 22642 8432 23802
rect 8496 23662 8524 24822
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8772 24274 8800 24686
rect 8760 24268 8812 24274
rect 8760 24210 8812 24216
rect 8666 23760 8722 23769
rect 8666 23695 8668 23704
rect 8720 23695 8722 23704
rect 8760 23724 8812 23730
rect 8668 23666 8720 23672
rect 8760 23666 8812 23672
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 8496 23322 8524 23598
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8496 23100 8524 23258
rect 8772 23254 8800 23666
rect 8864 23610 8892 25638
rect 10416 25356 10468 25362
rect 10416 25298 10468 25304
rect 9220 25220 9272 25226
rect 9220 25162 9272 25168
rect 9232 24818 9260 25162
rect 9291 25052 9599 25072
rect 9291 25050 9297 25052
rect 9353 25050 9377 25052
rect 9433 25050 9457 25052
rect 9513 25050 9537 25052
rect 9593 25050 9599 25052
rect 9353 24998 9355 25050
rect 9535 24998 9537 25050
rect 9291 24996 9297 24998
rect 9353 24996 9377 24998
rect 9433 24996 9457 24998
rect 9513 24996 9537 24998
rect 9593 24996 9599 24998
rect 9291 24976 9599 24996
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 10428 24274 10456 25298
rect 10704 25294 10732 25638
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10968 24880 11020 24886
rect 10968 24822 11020 24828
rect 10980 24698 11008 24822
rect 11072 24818 11100 25842
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 10980 24670 11100 24698
rect 10508 24608 10560 24614
rect 10560 24568 10640 24596
rect 10508 24550 10560 24556
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 8944 24064 8996 24070
rect 8944 24006 8996 24012
rect 8956 23730 8984 24006
rect 9291 23964 9599 23984
rect 9291 23962 9297 23964
rect 9353 23962 9377 23964
rect 9433 23962 9457 23964
rect 9513 23962 9537 23964
rect 9593 23962 9599 23964
rect 9353 23910 9355 23962
rect 9535 23910 9537 23962
rect 9291 23908 9297 23910
rect 9353 23908 9377 23910
rect 9433 23908 9457 23910
rect 9513 23908 9537 23910
rect 9593 23908 9599 23910
rect 9291 23888 9599 23908
rect 10152 23866 10180 24074
rect 10612 24070 10640 24568
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 9772 23792 9824 23798
rect 9772 23734 9824 23740
rect 8944 23724 8996 23730
rect 9128 23724 9180 23730
rect 8944 23666 8996 23672
rect 9048 23684 9128 23712
rect 9048 23610 9076 23684
rect 9128 23666 9180 23672
rect 8864 23582 9076 23610
rect 8864 23526 8892 23582
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 8760 23248 8812 23254
rect 8760 23190 8812 23196
rect 8576 23112 8628 23118
rect 8496 23072 8576 23100
rect 8576 23054 8628 23060
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8760 22976 8812 22982
rect 8760 22918 8812 22924
rect 8588 22642 8616 22918
rect 8772 22642 8800 22918
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8208 22500 8260 22506
rect 8208 22442 8260 22448
rect 8116 22228 8168 22234
rect 8116 22170 8168 22176
rect 8220 21894 8248 22442
rect 8588 22030 8616 22578
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 8036 20942 8064 21422
rect 8220 21010 8248 21830
rect 8312 21418 8340 21966
rect 8484 21956 8536 21962
rect 8484 21898 8536 21904
rect 8300 21412 8352 21418
rect 8300 21354 8352 21360
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8024 20936 8076 20942
rect 8024 20878 8076 20884
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8300 20800 8352 20806
rect 8220 20748 8300 20754
rect 8220 20742 8352 20748
rect 8220 20726 8340 20742
rect 7944 20318 8064 20346
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 10713 7604 16934
rect 7668 14074 7696 18566
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 7760 18086 7788 18362
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7668 13394 7696 13806
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7760 13326 7788 18022
rect 7852 17678 7880 18294
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7852 17066 7880 17614
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7852 16590 7880 17002
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7852 16046 7880 16526
rect 8036 16522 8064 20318
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8128 18358 8156 19858
rect 8220 19514 8248 20726
rect 8300 20256 8352 20262
rect 8404 20244 8432 20878
rect 8352 20216 8432 20244
rect 8300 20198 8352 20204
rect 8312 19718 8340 20198
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8220 19378 8248 19450
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 8312 18086 8340 19110
rect 8496 18970 8524 21898
rect 8668 21888 8720 21894
rect 8668 21830 8720 21836
rect 8680 21486 8708 21830
rect 8956 21486 8984 23462
rect 9784 23118 9812 23734
rect 10140 23724 10192 23730
rect 10140 23666 10192 23672
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9876 23118 9904 23598
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 9220 23044 9272 23050
rect 9220 22986 9272 22992
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 9232 22642 9260 22986
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 9291 22876 9599 22896
rect 9291 22874 9297 22876
rect 9353 22874 9377 22876
rect 9433 22874 9457 22876
rect 9513 22874 9537 22876
rect 9593 22874 9599 22876
rect 9353 22822 9355 22874
rect 9535 22822 9537 22874
rect 9291 22820 9297 22822
rect 9353 22820 9377 22822
rect 9433 22820 9457 22822
rect 9513 22820 9537 22822
rect 9593 22820 9599 22822
rect 9291 22800 9599 22820
rect 9784 22642 9812 22918
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 8588 20602 8616 20946
rect 8680 20874 8708 21286
rect 8956 21146 8984 21422
rect 9140 21418 9168 22510
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9508 22234 9536 22374
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9680 22024 9732 22030
rect 9784 22012 9812 22374
rect 9956 22160 10008 22166
rect 9956 22102 10008 22108
rect 9864 22024 9916 22030
rect 9784 21984 9864 22012
rect 9680 21966 9732 21972
rect 9864 21966 9916 21972
rect 9291 21788 9599 21808
rect 9291 21786 9297 21788
rect 9353 21786 9377 21788
rect 9433 21786 9457 21788
rect 9513 21786 9537 21788
rect 9593 21786 9599 21788
rect 9353 21734 9355 21786
rect 9535 21734 9537 21786
rect 9291 21732 9297 21734
rect 9353 21732 9377 21734
rect 9433 21732 9457 21734
rect 9513 21732 9537 21734
rect 9593 21732 9599 21734
rect 9291 21712 9599 21732
rect 9692 21554 9720 21966
rect 9968 21894 9996 22102
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9876 21706 9904 21830
rect 10060 21706 10088 22986
rect 10152 22778 10180 23666
rect 10612 23526 10640 24006
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 10612 22574 10640 23462
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10140 22568 10192 22574
rect 10140 22510 10192 22516
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 10600 22568 10652 22574
rect 10600 22510 10652 22516
rect 10152 22234 10180 22510
rect 10336 22438 10364 22510
rect 10704 22506 10732 22578
rect 10692 22500 10744 22506
rect 10692 22442 10744 22448
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10416 22432 10468 22438
rect 10416 22374 10468 22380
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 10428 22030 10456 22374
rect 10704 22098 10732 22442
rect 10796 22098 10824 22918
rect 10692 22092 10744 22098
rect 10692 22034 10744 22040
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 9876 21678 10088 21706
rect 10796 21690 10824 22034
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9772 21480 9824 21486
rect 9876 21468 9904 21678
rect 9956 21548 10008 21554
rect 10060 21536 10088 21678
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10140 21548 10192 21554
rect 10060 21508 10140 21536
rect 9956 21490 10008 21496
rect 10140 21490 10192 21496
rect 9824 21440 9904 21468
rect 9772 21422 9824 21428
rect 9128 21412 9180 21418
rect 9128 21354 9180 21360
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 9784 21078 9812 21422
rect 9772 21072 9824 21078
rect 9772 21014 9824 21020
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 9291 20700 9599 20720
rect 9291 20698 9297 20700
rect 9353 20698 9377 20700
rect 9433 20698 9457 20700
rect 9513 20698 9537 20700
rect 9593 20698 9599 20700
rect 9353 20646 9355 20698
rect 9535 20646 9537 20698
rect 9291 20644 9297 20646
rect 9353 20644 9377 20646
rect 9433 20644 9457 20646
rect 9513 20644 9537 20646
rect 9593 20644 9599 20646
rect 9291 20624 9599 20644
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 9876 20466 9904 20946
rect 9968 20942 9996 21490
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 10152 20942 10180 21286
rect 10428 21078 10456 21286
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 9968 20602 9996 20878
rect 10796 20806 10824 21626
rect 10888 21486 10916 24210
rect 10968 23792 11020 23798
rect 10968 23734 11020 23740
rect 10980 23526 11008 23734
rect 11072 23730 11100 24670
rect 11164 24410 11192 25842
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 11348 24206 11376 24754
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11152 24132 11204 24138
rect 11152 24074 11204 24080
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 10888 20466 10916 20878
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10980 19854 11008 23462
rect 11072 20874 11100 23666
rect 11164 23526 11192 24074
rect 11256 23866 11284 24142
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 11624 23746 11652 25978
rect 11808 25430 11836 26318
rect 11796 25424 11848 25430
rect 11796 25366 11848 25372
rect 11704 25152 11756 25158
rect 11704 25094 11756 25100
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 11716 24818 11744 25094
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11888 24744 11940 24750
rect 11888 24686 11940 24692
rect 11900 23866 11928 24686
rect 11992 24410 12020 25094
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 11520 23724 11572 23730
rect 11624 23718 12020 23746
rect 11520 23666 11572 23672
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 11164 21690 11192 23462
rect 11532 23254 11560 23666
rect 11520 23248 11572 23254
rect 11520 23190 11572 23196
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11336 22976 11388 22982
rect 11336 22918 11388 22924
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11164 21418 11192 21626
rect 11152 21412 11204 21418
rect 11152 21354 11204 21360
rect 11152 21072 11204 21078
rect 11152 21014 11204 21020
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 11072 20058 11100 20810
rect 11164 20466 11192 21014
rect 11256 20466 11284 21966
rect 11348 21894 11376 22918
rect 11900 22642 11928 22986
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 11794 21992 11850 22001
rect 11612 21956 11664 21962
rect 11794 21927 11850 21936
rect 11612 21898 11664 21904
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11624 21690 11652 21898
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 11348 20602 11376 20742
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11164 20369 11192 20402
rect 11150 20360 11206 20369
rect 11150 20295 11206 20304
rect 11348 20262 11376 20538
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 9291 19612 9599 19632
rect 9291 19610 9297 19612
rect 9353 19610 9377 19612
rect 9433 19610 9457 19612
rect 9513 19610 9537 19612
rect 9593 19610 9599 19612
rect 9353 19558 9355 19610
rect 9535 19558 9537 19610
rect 9291 19556 9297 19558
rect 9353 19556 9377 19558
rect 9433 19556 9457 19558
rect 9513 19556 9537 19558
rect 9593 19556 9599 19558
rect 9291 19536 9599 19556
rect 11072 19378 11100 19994
rect 11520 19984 11572 19990
rect 11520 19926 11572 19932
rect 11336 19848 11388 19854
rect 11532 19825 11560 19926
rect 11336 19790 11388 19796
rect 11518 19816 11574 19825
rect 11152 19508 11204 19514
rect 11152 19450 11204 19456
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8404 18358 8432 18566
rect 8588 18426 8616 19314
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 9291 18524 9599 18544
rect 9291 18522 9297 18524
rect 9353 18522 9377 18524
rect 9433 18522 9457 18524
rect 9513 18522 9537 18524
rect 9593 18522 9599 18524
rect 9353 18470 9355 18522
rect 9535 18470 9537 18522
rect 9291 18468 9297 18470
rect 9353 18468 9377 18470
rect 9433 18468 9457 18470
rect 9513 18468 9537 18470
rect 9593 18468 9599 18470
rect 9291 18448 9599 18468
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8404 16522 8432 18294
rect 9291 17436 9599 17456
rect 9291 17434 9297 17436
rect 9353 17434 9377 17436
rect 9433 17434 9457 17436
rect 9513 17434 9537 17436
rect 9593 17434 9599 17436
rect 9353 17382 9355 17434
rect 9535 17382 9537 17434
rect 9291 17380 9297 17382
rect 9353 17380 9377 17382
rect 9433 17380 9457 17382
rect 9513 17380 9537 17382
rect 9593 17380 9599 17382
rect 9291 17360 9599 17380
rect 9692 17338 9720 18294
rect 10520 17814 10548 18634
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10704 17678 10732 18906
rect 11164 18766 11192 19450
rect 11242 19408 11298 19417
rect 11348 19378 11376 19790
rect 11518 19751 11574 19760
rect 11612 19780 11664 19786
rect 11242 19343 11298 19352
rect 11336 19372 11388 19378
rect 11256 19242 11284 19343
rect 11336 19314 11388 19320
rect 11244 19236 11296 19242
rect 11244 19178 11296 19184
rect 11532 18766 11560 19751
rect 11612 19722 11664 19728
rect 11624 19242 11652 19722
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11716 19378 11744 19654
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11612 19236 11664 19242
rect 11612 19178 11664 19184
rect 11624 18902 11652 19178
rect 11612 18896 11664 18902
rect 11612 18838 11664 18844
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 9876 17338 9904 17546
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9048 17202 9076 17274
rect 9692 17202 9720 17274
rect 10244 17202 10272 17478
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 8864 16794 8892 17138
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 9048 16590 9076 16934
rect 9324 16794 9352 17138
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 8392 16516 8444 16522
rect 8392 16458 8444 16464
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8312 16250 8340 16390
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7852 15638 7880 15982
rect 7840 15632 7892 15638
rect 7840 15574 7892 15580
rect 7852 15094 7880 15574
rect 8036 15502 8064 16118
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8128 15570 8156 16050
rect 8496 15706 8524 16458
rect 9291 16348 9599 16368
rect 9291 16346 9297 16348
rect 9353 16346 9377 16348
rect 9433 16346 9457 16348
rect 9513 16346 9537 16348
rect 9593 16346 9599 16348
rect 9353 16294 9355 16346
rect 9535 16294 9537 16346
rect 9291 16292 9297 16294
rect 9353 16292 9377 16294
rect 9433 16292 9457 16294
rect 9513 16292 9537 16294
rect 9593 16292 9599 16294
rect 9291 16272 9599 16292
rect 9968 16250 9996 17138
rect 10060 16998 10088 17138
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10152 16454 10180 16730
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9404 16176 9456 16182
rect 9968 16130 9996 16186
rect 9404 16118 9456 16124
rect 9324 15978 9352 16118
rect 9312 15972 9364 15978
rect 9312 15914 9364 15920
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7852 13870 7880 14418
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7944 13716 7972 15302
rect 8036 14822 8064 15438
rect 8496 15366 8524 15438
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 8036 14414 8064 14758
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8128 14414 8156 14554
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8128 14074 8156 14350
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 7852 13688 7972 13716
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11762 7788 12038
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7760 10742 7788 11698
rect 7748 10736 7800 10742
rect 7562 10704 7618 10713
rect 7748 10678 7800 10684
rect 7562 10639 7564 10648
rect 7616 10639 7618 10648
rect 7564 10610 7616 10616
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7576 6866 7604 10610
rect 7852 9761 7880 13688
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7838 9752 7894 9761
rect 7838 9687 7894 9696
rect 7944 9382 7972 12378
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8128 10266 8156 10610
rect 8220 10470 8248 14282
rect 8404 14006 8432 14554
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8312 12374 8340 13874
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8404 11762 8432 12242
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8300 11280 8352 11286
rect 8298 11248 8300 11257
rect 8352 11248 8354 11257
rect 8298 11183 8354 11192
rect 8312 11014 8340 11183
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8220 10062 8248 10406
rect 8208 10056 8260 10062
rect 8022 10024 8078 10033
rect 8208 9998 8260 10004
rect 8022 9959 8024 9968
rect 8076 9959 8078 9968
rect 8024 9930 8076 9936
rect 8206 9752 8262 9761
rect 8206 9687 8262 9696
rect 8220 9382 8248 9687
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 8036 8634 8064 8842
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7932 8560 7984 8566
rect 7932 8502 7984 8508
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7852 7886 7880 8026
rect 7944 7886 7972 8502
rect 8128 8090 8156 9318
rect 8312 8974 8340 10678
rect 8404 10062 8432 11698
rect 8496 11354 8524 12582
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8496 9518 8524 9998
rect 8588 9586 8616 14962
rect 8680 14618 8708 15098
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8772 14414 8800 15846
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 13938 8708 14214
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8680 13841 8708 13874
rect 8666 13832 8722 13841
rect 8666 13767 8722 13776
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8680 12918 8708 13466
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8680 12238 8708 12718
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8680 11082 8708 11698
rect 8772 11642 8800 14350
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 13938 8892 14214
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8864 13530 8892 13874
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8864 11762 8892 13194
rect 8956 12782 8984 13806
rect 9048 13462 9076 15642
rect 9416 15502 9444 16118
rect 9600 16114 9996 16130
rect 9588 16108 9996 16114
rect 9640 16102 9996 16108
rect 9588 16050 9640 16056
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9291 15260 9599 15280
rect 9291 15258 9297 15260
rect 9353 15258 9377 15260
rect 9433 15258 9457 15260
rect 9513 15258 9537 15260
rect 9593 15258 9599 15260
rect 9353 15206 9355 15258
rect 9535 15206 9537 15258
rect 9291 15204 9297 15206
rect 9353 15204 9377 15206
rect 9433 15204 9457 15206
rect 9513 15204 9537 15206
rect 9593 15204 9599 15206
rect 9291 15184 9599 15204
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9140 14822 9168 14962
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 9036 13320 9088 13326
rect 9140 13308 9168 14758
rect 9291 14172 9599 14192
rect 9291 14170 9297 14172
rect 9353 14170 9377 14172
rect 9433 14170 9457 14172
rect 9513 14170 9537 14172
rect 9593 14170 9599 14172
rect 9353 14118 9355 14170
rect 9535 14118 9537 14170
rect 9291 14116 9297 14118
rect 9353 14116 9377 14118
rect 9433 14116 9457 14118
rect 9513 14116 9537 14118
rect 9593 14116 9599 14118
rect 9291 14096 9599 14116
rect 9220 14000 9272 14006
rect 9680 14000 9732 14006
rect 9220 13942 9272 13948
rect 9586 13968 9642 13977
rect 9232 13462 9260 13942
rect 9680 13942 9732 13948
rect 9586 13903 9642 13912
rect 9600 13802 9628 13903
rect 9692 13841 9720 13942
rect 9678 13832 9734 13841
rect 9312 13796 9364 13802
rect 9588 13796 9640 13802
rect 9364 13756 9444 13784
rect 9312 13738 9364 13744
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9140 13280 9260 13308
rect 9416 13304 9444 13756
rect 9678 13767 9734 13776
rect 9588 13738 9640 13744
rect 9692 13326 9720 13767
rect 9680 13320 9732 13326
rect 9036 13262 9088 13268
rect 9048 12986 9076 13262
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 9140 12714 9168 13126
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 9048 12238 9076 12310
rect 9036 12232 9088 12238
rect 8956 12192 9036 12220
rect 8956 11898 8984 12192
rect 9036 12174 9088 12180
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8772 11614 8892 11642
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8680 10062 8708 10746
rect 8772 10130 8800 11290
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8864 9586 8892 11614
rect 8956 11218 8984 11698
rect 9048 11694 9076 12038
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8956 10674 8984 11154
rect 9048 11150 9076 11494
rect 9140 11234 9168 12650
rect 9232 12442 9260 13280
rect 9404 13298 9456 13304
rect 9680 13262 9732 13268
rect 9404 13240 9456 13246
rect 9291 13084 9599 13104
rect 9291 13082 9297 13084
rect 9353 13082 9377 13084
rect 9433 13082 9457 13084
rect 9513 13082 9537 13084
rect 9593 13082 9599 13084
rect 9353 13030 9355 13082
rect 9535 13030 9537 13082
rect 9291 13028 9297 13030
rect 9353 13028 9377 13030
rect 9433 13028 9457 13030
rect 9513 13028 9537 13030
rect 9593 13028 9599 13030
rect 9291 13008 9599 13028
rect 9678 13016 9734 13025
rect 9784 13002 9812 15370
rect 10152 15026 10180 16390
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10244 15094 10272 16050
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10336 15026 10364 15642
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9968 13734 9996 13874
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9968 13326 9996 13670
rect 10138 13424 10194 13433
rect 10138 13359 10194 13368
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9734 12974 9812 13002
rect 9678 12951 9680 12960
rect 9732 12951 9734 12960
rect 9680 12922 9732 12928
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9600 12238 9628 12378
rect 9784 12238 9812 12974
rect 9864 12912 9916 12918
rect 9968 12900 9996 13262
rect 10152 13258 10180 13359
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10322 13152 10378 13161
rect 9916 12872 9996 12900
rect 9864 12854 9916 12860
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9588 12232 9640 12238
rect 9772 12232 9824 12238
rect 9640 12180 9720 12186
rect 9588 12174 9720 12180
rect 9772 12174 9824 12180
rect 9232 11626 9260 12174
rect 9600 12158 9720 12174
rect 9291 11996 9599 12016
rect 9291 11994 9297 11996
rect 9353 11994 9377 11996
rect 9433 11994 9457 11996
rect 9513 11994 9537 11996
rect 9593 11994 9599 11996
rect 9353 11942 9355 11994
rect 9535 11942 9537 11994
rect 9291 11940 9297 11942
rect 9353 11940 9377 11942
rect 9433 11940 9457 11942
rect 9513 11940 9537 11942
rect 9593 11940 9599 11942
rect 9291 11920 9599 11940
rect 9692 11778 9720 12158
rect 9600 11750 9720 11778
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9232 11354 9260 11562
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9140 11206 9260 11234
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9034 10976 9090 10985
rect 9034 10911 9090 10920
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8496 8498 8524 8978
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8634 8616 8774
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8220 7954 8248 8366
rect 8300 8016 8352 8022
rect 8404 8004 8432 8366
rect 8352 7976 8432 8004
rect 8300 7958 8352 7964
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8312 7886 8340 7958
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7546 8340 7686
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 6920 6724 6972 6730
rect 7392 6718 7604 6746
rect 6920 6666 6972 6672
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4690 7512 4966
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7116 4146 7144 4422
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 7116 4010 7144 4082
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7484 3194 7512 4150
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7484 2514 7512 3130
rect 7576 2774 7604 6718
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6322 7788 6598
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7760 5642 7788 6258
rect 7944 6254 7972 7278
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7944 5846 7972 6190
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7944 5234 7972 5782
rect 8036 5302 8064 6054
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7840 5024 7892 5030
rect 7668 4984 7840 5012
rect 7668 4758 7696 4984
rect 7840 4966 7892 4972
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7760 4282 7788 4558
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7668 3738 7696 4014
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7760 3534 7788 4218
rect 7944 3602 7972 5170
rect 8036 4486 8064 5238
rect 8128 4622 8156 5306
rect 8220 5302 8248 5646
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8036 4146 8064 4422
rect 8220 4214 8248 4626
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8312 4078 8340 7142
rect 8404 6458 8432 7822
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8496 6390 8524 7686
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8404 4826 8432 5850
rect 8485 5704 8537 5710
rect 8485 5646 8537 5652
rect 8496 5370 8524 5646
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8496 4622 8524 5170
rect 8588 4690 8616 8570
rect 8680 8498 8708 9386
rect 8864 8974 8892 9522
rect 9048 9042 9076 10911
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9140 9926 9168 9998
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8498 8984 8842
rect 9048 8634 9076 8978
rect 9232 8906 9260 11206
rect 9600 11121 9628 11750
rect 9586 11112 9642 11121
rect 9586 11047 9642 11056
rect 9291 10908 9599 10928
rect 9291 10906 9297 10908
rect 9353 10906 9377 10908
rect 9433 10906 9457 10908
rect 9513 10906 9537 10908
rect 9593 10906 9599 10908
rect 9353 10854 9355 10906
rect 9535 10854 9537 10906
rect 9291 10852 9297 10854
rect 9353 10852 9377 10854
rect 9433 10852 9457 10854
rect 9513 10852 9537 10854
rect 9593 10852 9599 10854
rect 9291 10832 9599 10852
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9508 10062 9536 10678
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9692 10266 9720 10610
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9770 10024 9826 10033
rect 9680 9988 9732 9994
rect 9770 9959 9826 9968
rect 9680 9930 9732 9936
rect 9291 9820 9599 9840
rect 9291 9818 9297 9820
rect 9353 9818 9377 9820
rect 9433 9818 9457 9820
rect 9513 9818 9537 9820
rect 9593 9818 9599 9820
rect 9353 9766 9355 9818
rect 9535 9766 9537 9818
rect 9291 9764 9297 9766
rect 9353 9764 9377 9766
rect 9433 9764 9457 9766
rect 9513 9764 9537 9766
rect 9593 9764 9599 9766
rect 9291 9744 9599 9764
rect 9692 9722 9720 9930
rect 9784 9722 9812 9959
rect 9876 9926 9904 10066
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9291 8732 9599 8752
rect 9291 8730 9297 8732
rect 9353 8730 9377 8732
rect 9433 8730 9457 8732
rect 9513 8730 9537 8732
rect 9593 8730 9599 8732
rect 9353 8678 9355 8730
rect 9535 8678 9537 8730
rect 9291 8676 9297 8678
rect 9353 8676 9377 8678
rect 9433 8676 9457 8678
rect 9513 8676 9537 8678
rect 9593 8676 9599 8678
rect 9291 8656 9599 8676
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9048 7886 9076 8026
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9048 6662 9076 7482
rect 9140 7206 9168 7958
rect 9232 7886 9260 8298
rect 9876 8090 9904 9862
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9232 7410 9260 7686
rect 9291 7644 9599 7664
rect 9291 7642 9297 7644
rect 9353 7642 9377 7644
rect 9433 7642 9457 7644
rect 9513 7642 9537 7644
rect 9593 7642 9599 7644
rect 9353 7590 9355 7642
rect 9535 7590 9537 7642
rect 9291 7588 9297 7590
rect 9353 7588 9377 7590
rect 9433 7588 9457 7590
rect 9513 7588 9537 7590
rect 9593 7588 9599 7590
rect 9291 7568 9599 7588
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8680 4826 8708 5714
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8772 5370 8800 5646
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 9048 4146 9076 6598
rect 9291 6556 9599 6576
rect 9291 6554 9297 6556
rect 9353 6554 9377 6556
rect 9433 6554 9457 6556
rect 9513 6554 9537 6556
rect 9593 6554 9599 6556
rect 9353 6502 9355 6554
rect 9535 6502 9537 6554
rect 9291 6500 9297 6502
rect 9353 6500 9377 6502
rect 9433 6500 9457 6502
rect 9513 6500 9537 6502
rect 9593 6500 9599 6502
rect 9291 6480 9599 6500
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9232 5302 9260 6394
rect 9968 6254 9996 12872
rect 10060 12850 10088 13126
rect 10322 13087 10378 13096
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10152 12434 10180 12922
rect 10336 12646 10364 13087
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10428 12434 10456 16526
rect 10520 15706 10548 17546
rect 10796 17202 10824 18158
rect 10968 17740 11020 17746
rect 10888 17700 10968 17728
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10796 16794 10824 17138
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10888 15910 10916 17700
rect 10968 17682 11020 17688
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10600 15428 10652 15434
rect 10600 15370 10652 15376
rect 10612 15162 10640 15370
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10888 14958 10916 15846
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10612 12918 10640 13126
rect 10704 12986 10732 13262
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10060 12406 10180 12434
rect 10336 12406 10456 12434
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9291 5468 9599 5488
rect 9291 5466 9297 5468
rect 9353 5466 9377 5468
rect 9433 5466 9457 5468
rect 9513 5466 9537 5468
rect 9593 5466 9599 5468
rect 9353 5414 9355 5466
rect 9535 5414 9537 5466
rect 9291 5412 9297 5414
rect 9353 5412 9377 5414
rect 9433 5412 9457 5414
rect 9513 5412 9537 5414
rect 9593 5412 9599 5414
rect 9291 5392 9599 5412
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9232 4282 9260 4694
rect 9291 4380 9599 4400
rect 9291 4378 9297 4380
rect 9353 4378 9377 4380
rect 9433 4378 9457 4380
rect 9513 4378 9537 4380
rect 9593 4378 9599 4380
rect 9353 4326 9355 4378
rect 9535 4326 9537 4378
rect 9291 4324 9297 4326
rect 9353 4324 9377 4326
rect 9433 4324 9457 4326
rect 9513 4324 9537 4326
rect 9593 4324 9599 4326
rect 9291 4304 9599 4324
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8220 3602 8248 3946
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7576 2746 7696 2774
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 6380 870 6500 898
rect 6380 762 6408 870
rect 6472 800 6500 870
rect 7668 800 7696 2746
rect 7760 2446 7788 3470
rect 8220 2854 8248 3538
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8220 2650 8248 2790
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8312 2446 8340 3878
rect 8404 3670 8432 4082
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8496 3534 8524 3878
rect 10060 3738 10088 12406
rect 10230 11248 10286 11257
rect 10230 11183 10286 11192
rect 10244 11014 10272 11183
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10336 9586 10364 12406
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 10244 8430 10272 9386
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 6798 10180 7754
rect 10336 7342 10364 7822
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8588 2650 8616 2994
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8864 800 8892 3674
rect 9291 3292 9599 3312
rect 9291 3290 9297 3292
rect 9353 3290 9377 3292
rect 9433 3290 9457 3292
rect 9513 3290 9537 3292
rect 9593 3290 9599 3292
rect 9353 3238 9355 3290
rect 9535 3238 9537 3290
rect 9291 3236 9297 3238
rect 9353 3236 9377 3238
rect 9433 3236 9457 3238
rect 9513 3236 9537 3238
rect 9593 3236 9599 3238
rect 9291 3216 9599 3236
rect 10428 2774 10456 12038
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10612 11354 10640 11494
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10612 10198 10640 10950
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10796 9654 10824 14214
rect 10874 13424 10930 13433
rect 10874 13359 10876 13368
rect 10928 13359 10930 13368
rect 10876 13330 10928 13336
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12986 10916 13194
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 12102 10916 12242
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10612 7886 10640 8298
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10520 6798 10548 7278
rect 10704 6934 10732 9318
rect 10980 9110 11008 17070
rect 11164 15502 11192 18702
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11244 18352 11296 18358
rect 11244 18294 11296 18300
rect 11256 17202 11284 18294
rect 11348 17814 11376 18566
rect 11624 18290 11652 18838
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11532 17134 11560 17614
rect 11624 17542 11652 18226
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11716 16590 11744 19314
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11808 16522 11836 21927
rect 11900 21146 11928 22578
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 11992 20602 12020 23718
rect 12084 22001 12112 28750
rect 12438 28642 12494 29442
rect 12912 28750 13584 28778
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12360 26382 12388 26522
rect 12348 26376 12400 26382
rect 12348 26318 12400 26324
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 12360 25362 12388 26182
rect 12348 25356 12400 25362
rect 12348 25298 12400 25304
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 12164 24948 12216 24954
rect 12164 24890 12216 24896
rect 12176 24750 12204 24890
rect 12164 24744 12216 24750
rect 12164 24686 12216 24692
rect 12070 21992 12126 22001
rect 12070 21927 12126 21936
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11900 18290 11928 19178
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11992 17490 12020 18566
rect 12084 18290 12112 21830
rect 12176 21690 12204 24686
rect 12360 24682 12388 25094
rect 12348 24676 12400 24682
rect 12348 24618 12400 24624
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12268 23866 12296 24006
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12360 22438 12388 24142
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12268 21554 12296 21898
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12164 19712 12216 19718
rect 12164 19654 12216 19660
rect 12176 19378 12204 19654
rect 12268 19514 12296 19790
rect 12360 19786 12388 20538
rect 12348 19780 12400 19786
rect 12348 19722 12400 19728
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12346 19408 12402 19417
rect 12164 19372 12216 19378
rect 12346 19343 12402 19352
rect 12164 19314 12216 19320
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12176 18698 12204 19110
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12176 17678 12204 18022
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 11992 17462 12204 17490
rect 11796 16516 11848 16522
rect 11796 16458 11848 16464
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11072 14618 11100 15370
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11532 15026 11560 15302
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11532 14822 11560 14962
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11060 14612 11112 14618
rect 11532 14600 11560 14758
rect 11060 14554 11112 14560
rect 11440 14572 11560 14600
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11164 14074 11192 14418
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11164 13530 11192 14010
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11072 12238 11100 13398
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11164 12442 11192 13262
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11348 12714 11376 13126
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 11348 12306 11376 12650
rect 11440 12646 11468 14572
rect 11624 14414 11652 15574
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11532 12850 11560 13806
rect 11624 13326 11652 14010
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 13190 11652 13262
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11610 12880 11666 12889
rect 11520 12844 11572 12850
rect 11610 12815 11666 12824
rect 11520 12786 11572 12792
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11532 11694 11560 12786
rect 11624 12782 11652 12815
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11624 12238 11652 12378
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11612 12096 11664 12102
rect 11716 12050 11744 15438
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11900 14074 11928 14350
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11808 13530 11836 13874
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11796 13388 11848 13394
rect 11992 13376 12020 14418
rect 11848 13348 12020 13376
rect 11796 13330 11848 13336
rect 11808 13190 11836 13330
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11886 13152 11942 13161
rect 11886 13087 11942 13096
rect 11900 12850 11928 13087
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11888 12640 11940 12646
rect 12176 12594 12204 17462
rect 12360 16182 12388 19343
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 12452 15978 12480 28642
rect 12716 26308 12768 26314
rect 12716 26250 12768 26256
rect 12728 26042 12756 26250
rect 12716 26036 12768 26042
rect 12716 25978 12768 25984
rect 12624 25356 12676 25362
rect 12624 25298 12676 25304
rect 12636 24750 12664 25298
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12544 24410 12572 24550
rect 12820 24410 12848 25230
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12808 24404 12860 24410
rect 12808 24346 12860 24352
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12636 22982 12664 23598
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12912 22094 12940 28750
rect 13556 28642 13584 28750
rect 13634 28642 13690 29442
rect 14738 28642 14794 29442
rect 15934 28642 15990 29442
rect 17130 28642 17186 29442
rect 17972 28750 18276 28778
rect 13556 28614 13676 28642
rect 13462 26684 13770 26704
rect 13462 26682 13468 26684
rect 13524 26682 13548 26684
rect 13604 26682 13628 26684
rect 13684 26682 13708 26684
rect 13764 26682 13770 26684
rect 13524 26630 13526 26682
rect 13706 26630 13708 26682
rect 13462 26628 13468 26630
rect 13524 26628 13548 26630
rect 13604 26628 13628 26630
rect 13684 26628 13708 26630
rect 13764 26628 13770 26630
rect 13462 26608 13770 26628
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 14372 26376 14424 26382
rect 14424 26324 14504 26330
rect 14372 26318 14504 26324
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 13188 25498 13216 25842
rect 13462 25596 13770 25616
rect 13462 25594 13468 25596
rect 13524 25594 13548 25596
rect 13604 25594 13628 25596
rect 13684 25594 13708 25596
rect 13764 25594 13770 25596
rect 13524 25542 13526 25594
rect 13706 25542 13708 25594
rect 13462 25540 13468 25542
rect 13524 25540 13548 25542
rect 13604 25540 13628 25542
rect 13684 25540 13708 25542
rect 13764 25540 13770 25542
rect 13462 25520 13770 25540
rect 13176 25492 13228 25498
rect 13176 25434 13228 25440
rect 13832 25294 13860 26318
rect 14188 26308 14240 26314
rect 14384 26302 14504 26318
rect 14188 26250 14240 26256
rect 14200 25430 14228 26250
rect 14476 25702 14504 26302
rect 14556 26308 14608 26314
rect 14556 26250 14608 26256
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 14188 25424 14240 25430
rect 14188 25366 14240 25372
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 13188 24954 13216 25162
rect 13176 24948 13228 24954
rect 13176 24890 13228 24896
rect 14108 24818 14136 25230
rect 14384 24954 14412 25434
rect 14476 25362 14504 25638
rect 14464 25356 14516 25362
rect 14464 25298 14516 25304
rect 14464 25152 14516 25158
rect 14464 25094 14516 25100
rect 14372 24948 14424 24954
rect 14372 24890 14424 24896
rect 14280 24880 14332 24886
rect 14280 24822 14332 24828
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 13280 23866 13308 24754
rect 13372 24274 13400 24754
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 13462 24508 13770 24528
rect 13462 24506 13468 24508
rect 13524 24506 13548 24508
rect 13604 24506 13628 24508
rect 13684 24506 13708 24508
rect 13764 24506 13770 24508
rect 13524 24454 13526 24506
rect 13706 24454 13708 24506
rect 13462 24452 13468 24454
rect 13524 24452 13548 24454
rect 13604 24452 13628 24454
rect 13684 24452 13708 24454
rect 13764 24452 13770 24454
rect 13462 24432 13770 24452
rect 14016 24410 14044 24686
rect 14004 24404 14056 24410
rect 14004 24346 14056 24352
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 14188 24132 14240 24138
rect 14188 24074 14240 24080
rect 13268 23860 13320 23866
rect 13268 23802 13320 23808
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13280 23118 13308 23666
rect 13462 23420 13770 23440
rect 13462 23418 13468 23420
rect 13524 23418 13548 23420
rect 13604 23418 13628 23420
rect 13684 23418 13708 23420
rect 13764 23418 13770 23420
rect 13524 23366 13526 23418
rect 13706 23366 13708 23418
rect 13462 23364 13468 23366
rect 13524 23364 13548 23366
rect 13604 23364 13628 23366
rect 13684 23364 13708 23366
rect 13764 23364 13770 23366
rect 13462 23344 13770 23364
rect 14200 23322 14228 24074
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 12820 22066 12940 22094
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12636 19446 12664 19654
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12544 18630 12572 19246
rect 12636 18766 12664 19246
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12544 17270 12572 17818
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12636 16130 12664 17614
rect 12544 16114 12664 16130
rect 12532 16108 12664 16114
rect 12584 16102 12664 16108
rect 12532 16050 12584 16056
rect 12728 16046 12756 17682
rect 12716 16040 12768 16046
rect 12544 15988 12716 15994
rect 12544 15982 12768 15988
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12544 15966 12756 15982
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12360 15722 12388 15846
rect 12544 15722 12572 15966
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12360 15706 12572 15722
rect 12348 15700 12572 15706
rect 12400 15694 12572 15700
rect 12348 15642 12400 15648
rect 12440 15564 12492 15570
rect 12636 15552 12664 15846
rect 12492 15524 12664 15552
rect 12440 15506 12492 15512
rect 12256 15496 12308 15502
rect 12254 15464 12256 15473
rect 12308 15464 12310 15473
rect 12622 15464 12678 15473
rect 12254 15399 12310 15408
rect 12440 15428 12492 15434
rect 12622 15399 12678 15408
rect 12440 15370 12492 15376
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12268 13462 12296 14010
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12268 13274 12296 13398
rect 12268 13246 12388 13274
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12268 12646 12296 13126
rect 11888 12582 11940 12588
rect 11664 12044 11744 12050
rect 11612 12038 11744 12044
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11624 12022 11744 12038
rect 11808 11762 11836 12038
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11900 11234 11928 12582
rect 11992 12566 12204 12594
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 11992 11370 12020 12566
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12084 11762 12112 12174
rect 12268 12170 12296 12582
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11992 11342 12296 11370
rect 11900 11206 12112 11234
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11992 10470 12020 11086
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10888 8430 10916 8910
rect 10980 8566 11008 9046
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10520 5642 10548 6734
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10520 5234 10548 5578
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10520 4622 10548 5170
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10612 4826 10640 4966
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10520 3534 10548 4558
rect 10612 4282 10640 4762
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10796 3534 10824 8298
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 8090 11008 8230
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10980 7478 11008 8026
rect 11072 7886 11100 9114
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 11164 8634 11192 8842
rect 11624 8634 11652 8842
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11164 8537 11192 8570
rect 11150 8528 11206 8537
rect 11150 8463 11206 8472
rect 11808 8430 11836 8774
rect 11900 8566 11928 9318
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 11072 7410 11100 7822
rect 11624 7546 11652 8366
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11716 7410 11744 7958
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10888 5302 10916 5850
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10888 4690 10916 5238
rect 11164 5098 11192 5782
rect 11532 5710 11560 6258
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11440 5370 11468 5646
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10888 4214 10916 4626
rect 11532 4622 11560 5646
rect 11900 5642 11928 8502
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11624 5302 11652 5510
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 11532 4146 11560 4422
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11072 3534 11100 3878
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 10520 3058 10548 3470
rect 11256 3126 11284 3878
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11808 3058 11836 3878
rect 11992 3194 12020 10406
rect 12084 7342 12112 11206
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12176 7954 12204 9522
rect 12268 9382 12296 11342
rect 12360 11132 12388 13246
rect 12452 13025 12480 15370
rect 12532 13456 12584 13462
rect 12636 13433 12664 15399
rect 12532 13398 12584 13404
rect 12622 13424 12678 13433
rect 12438 13016 12494 13025
rect 12438 12951 12494 12960
rect 12452 12850 12480 12951
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12544 12730 12572 13398
rect 12622 13359 12624 13368
rect 12676 13359 12678 13368
rect 12624 13330 12676 13336
rect 12452 12714 12572 12730
rect 12440 12708 12572 12714
rect 12492 12702 12572 12708
rect 12440 12650 12492 12656
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12544 12238 12572 12582
rect 12636 12442 12664 13330
rect 12714 13288 12770 13297
rect 12714 13223 12770 13232
rect 12728 12714 12756 13223
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12636 11558 12664 12242
rect 12820 12170 12848 22066
rect 13096 21554 13124 22374
rect 13280 21570 13308 23054
rect 13360 22976 13412 22982
rect 13360 22918 13412 22924
rect 13372 22642 13400 22918
rect 14292 22778 14320 24822
rect 14476 24138 14504 25094
rect 14568 24818 14596 26250
rect 14648 25832 14700 25838
rect 14648 25774 14700 25780
rect 14660 25362 14688 25774
rect 14648 25356 14700 25362
rect 14648 25298 14700 25304
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14568 24410 14596 24550
rect 14556 24404 14608 24410
rect 14556 24346 14608 24352
rect 14464 24132 14516 24138
rect 14464 24074 14516 24080
rect 14464 23656 14516 23662
rect 14464 23598 14516 23604
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 14096 22636 14148 22642
rect 14096 22578 14148 22584
rect 13372 22234 13400 22578
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 13462 22332 13770 22352
rect 13462 22330 13468 22332
rect 13524 22330 13548 22332
rect 13604 22330 13628 22332
rect 13684 22330 13708 22332
rect 13764 22330 13770 22332
rect 13524 22278 13526 22330
rect 13706 22278 13708 22330
rect 13462 22276 13468 22278
rect 13524 22276 13548 22278
rect 13604 22276 13628 22278
rect 13684 22276 13708 22278
rect 13764 22276 13770 22278
rect 13462 22256 13770 22276
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13372 22030 13400 22170
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 13188 21542 13308 21570
rect 13832 21554 13860 22374
rect 13924 22166 13952 22510
rect 14108 22234 14136 22578
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 13912 22160 13964 22166
rect 13912 22102 13964 22108
rect 13820 21548 13872 21554
rect 12912 20369 12940 21490
rect 12898 20360 12954 20369
rect 12898 20295 12954 20304
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12912 19922 12940 20198
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12992 19848 13044 19854
rect 12990 19816 12992 19825
rect 13188 19836 13216 21542
rect 13820 21490 13872 21496
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13044 19816 13216 19836
rect 13046 19808 13216 19816
rect 12990 19751 13046 19760
rect 12900 18148 12952 18154
rect 12900 18090 12952 18096
rect 12912 17882 12940 18090
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12912 16114 12940 17818
rect 13096 17678 13124 18022
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13280 17762 13308 21422
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13462 21244 13770 21264
rect 13462 21242 13468 21244
rect 13524 21242 13548 21244
rect 13604 21242 13628 21244
rect 13684 21242 13708 21244
rect 13764 21242 13770 21244
rect 13524 21190 13526 21242
rect 13706 21190 13708 21242
rect 13462 21188 13468 21190
rect 13524 21188 13548 21190
rect 13604 21188 13628 21190
rect 13684 21188 13708 21190
rect 13764 21188 13770 21190
rect 13462 21168 13770 21188
rect 13462 20156 13770 20176
rect 13462 20154 13468 20156
rect 13524 20154 13548 20156
rect 13604 20154 13628 20156
rect 13684 20154 13708 20156
rect 13764 20154 13770 20156
rect 13524 20102 13526 20154
rect 13706 20102 13708 20154
rect 13462 20100 13468 20102
rect 13524 20100 13548 20102
rect 13604 20100 13628 20102
rect 13684 20100 13708 20102
rect 13764 20100 13770 20102
rect 13462 20080 13770 20100
rect 13832 19854 13860 21286
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13462 19068 13770 19088
rect 13462 19066 13468 19068
rect 13524 19066 13548 19068
rect 13604 19066 13628 19068
rect 13684 19066 13708 19068
rect 13764 19066 13770 19068
rect 13524 19014 13526 19066
rect 13706 19014 13708 19066
rect 13462 19012 13468 19014
rect 13524 19012 13548 19014
rect 13604 19012 13628 19014
rect 13684 19012 13708 19014
rect 13764 19012 13770 19014
rect 13462 18992 13770 19012
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13372 18290 13400 18702
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13464 18068 13492 18226
rect 13372 18040 13492 18068
rect 13372 17882 13400 18040
rect 13462 17980 13770 18000
rect 13462 17978 13468 17980
rect 13524 17978 13548 17980
rect 13604 17978 13628 17980
rect 13684 17978 13708 17980
rect 13764 17978 13770 17980
rect 13524 17926 13526 17978
rect 13706 17926 13708 17978
rect 13462 17924 13468 17926
rect 13524 17924 13548 17926
rect 13604 17924 13628 17926
rect 13684 17924 13708 17926
rect 13764 17924 13770 17926
rect 13462 17904 13770 17924
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 13096 16250 13124 16458
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 13188 16046 13216 17750
rect 13280 17734 13400 17762
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13280 17338 13308 17614
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 12992 15088 13044 15094
rect 12992 15030 13044 15036
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12912 14822 12940 14962
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12440 11144 12492 11150
rect 12360 11104 12440 11132
rect 12440 11086 12492 11092
rect 12808 11076 12860 11082
rect 12808 11018 12860 11024
rect 12820 10742 12848 11018
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12268 7886 12296 8910
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 6322 12204 7142
rect 12268 7002 12296 7822
rect 12360 7818 12388 8570
rect 12636 8412 12664 8910
rect 12714 8528 12770 8537
rect 12714 8463 12716 8472
rect 12768 8463 12770 8472
rect 12716 8434 12768 8440
rect 12452 8384 12664 8412
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12452 7426 12480 8384
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12544 7732 12572 8230
rect 12624 7744 12676 7750
rect 12544 7704 12624 7732
rect 12544 7546 12572 7704
rect 12624 7686 12676 7692
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12820 7478 12848 7686
rect 12808 7472 12860 7478
rect 12452 7410 12664 7426
rect 12808 7414 12860 7420
rect 12440 7404 12664 7410
rect 12492 7398 12664 7404
rect 12440 7346 12492 7352
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12268 6118 12296 6734
rect 12452 6458 12480 6802
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12268 5778 12296 6054
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12268 4690 12296 5714
rect 12544 5030 12572 7278
rect 12636 6934 12664 7398
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12084 4214 12112 4422
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 12176 4078 12204 4422
rect 12636 4146 12664 5238
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12360 3534 12388 3946
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12636 3194 12664 4082
rect 12728 3942 12756 4422
rect 12820 4146 12848 4966
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 10336 2746 10456 2774
rect 9291 2204 9599 2224
rect 9291 2202 9297 2204
rect 9353 2202 9377 2204
rect 9433 2202 9457 2204
rect 9513 2202 9537 2204
rect 9593 2202 9599 2204
rect 9353 2150 9355 2202
rect 9535 2150 9537 2202
rect 9291 2148 9297 2150
rect 9353 2148 9377 2150
rect 9433 2148 9457 2150
rect 9513 2148 9537 2150
rect 9593 2148 9599 2150
rect 9291 2128 9599 2148
rect 10060 870 10180 898
rect 10060 800 10088 870
rect 6196 734 6408 762
rect 6458 0 6514 800
rect 7654 0 7710 800
rect 8850 0 8906 800
rect 10046 0 10102 800
rect 10152 762 10180 870
rect 10336 762 10364 2746
rect 12452 800 12480 3130
rect 12912 1358 12940 14758
rect 13004 14074 13032 15030
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13096 13938 13124 14350
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13188 13462 13216 13874
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 13280 13326 13308 15506
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 12990 12880 13046 12889
rect 12990 12815 12992 12824
rect 13044 12815 13046 12824
rect 12992 12786 13044 12792
rect 13004 12238 13032 12786
rect 13096 12646 13124 13262
rect 13280 12782 13308 13262
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12992 11144 13044 11150
rect 13096 11132 13124 12582
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13188 11150 13216 11630
rect 13280 11286 13308 12038
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 13372 11268 13400 17734
rect 13832 17678 13860 18362
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13462 16892 13770 16912
rect 13462 16890 13468 16892
rect 13524 16890 13548 16892
rect 13604 16890 13628 16892
rect 13684 16890 13708 16892
rect 13764 16890 13770 16892
rect 13524 16838 13526 16890
rect 13706 16838 13708 16890
rect 13462 16836 13468 16838
rect 13524 16836 13548 16838
rect 13604 16836 13628 16838
rect 13684 16836 13708 16838
rect 13764 16836 13770 16838
rect 13462 16816 13770 16836
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13462 15804 13770 15824
rect 13462 15802 13468 15804
rect 13524 15802 13548 15804
rect 13604 15802 13628 15804
rect 13684 15802 13708 15804
rect 13764 15802 13770 15804
rect 13524 15750 13526 15802
rect 13706 15750 13708 15802
rect 13462 15748 13468 15750
rect 13524 15748 13548 15750
rect 13604 15748 13628 15750
rect 13684 15748 13708 15750
rect 13764 15748 13770 15750
rect 13462 15728 13770 15748
rect 13636 15496 13688 15502
rect 13634 15464 13636 15473
rect 13688 15464 13690 15473
rect 13634 15399 13690 15408
rect 13832 15026 13860 16118
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13462 14716 13770 14736
rect 13462 14714 13468 14716
rect 13524 14714 13548 14716
rect 13604 14714 13628 14716
rect 13684 14714 13708 14716
rect 13764 14714 13770 14716
rect 13524 14662 13526 14714
rect 13706 14662 13708 14714
rect 13462 14660 13468 14662
rect 13524 14660 13548 14662
rect 13604 14660 13628 14662
rect 13684 14660 13708 14662
rect 13764 14660 13770 14662
rect 13462 14640 13770 14660
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13462 13628 13770 13648
rect 13462 13626 13468 13628
rect 13524 13626 13548 13628
rect 13604 13626 13628 13628
rect 13684 13626 13708 13628
rect 13764 13626 13770 13628
rect 13524 13574 13526 13626
rect 13706 13574 13708 13626
rect 13462 13572 13468 13574
rect 13524 13572 13548 13574
rect 13604 13572 13628 13574
rect 13684 13572 13708 13574
rect 13764 13572 13770 13574
rect 13462 13552 13770 13572
rect 13544 13320 13596 13326
rect 13542 13288 13544 13297
rect 13596 13288 13598 13297
rect 13542 13223 13598 13232
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12850 13676 13126
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13462 12540 13770 12560
rect 13462 12538 13468 12540
rect 13524 12538 13548 12540
rect 13604 12538 13628 12540
rect 13684 12538 13708 12540
rect 13764 12538 13770 12540
rect 13524 12486 13526 12538
rect 13706 12486 13708 12538
rect 13462 12484 13468 12486
rect 13524 12484 13548 12486
rect 13604 12484 13628 12486
rect 13684 12484 13708 12486
rect 13764 12484 13770 12486
rect 13462 12464 13770 12484
rect 13462 11452 13770 11472
rect 13462 11450 13468 11452
rect 13524 11450 13548 11452
rect 13604 11450 13628 11452
rect 13684 11450 13708 11452
rect 13764 11450 13770 11452
rect 13524 11398 13526 11450
rect 13706 11398 13708 11450
rect 13462 11396 13468 11398
rect 13524 11396 13548 11398
rect 13604 11396 13628 11398
rect 13684 11396 13708 11398
rect 13764 11396 13770 11398
rect 13462 11376 13770 11396
rect 13452 11280 13504 11286
rect 13372 11240 13452 11268
rect 13280 11150 13308 11222
rect 13044 11104 13124 11132
rect 13176 11144 13228 11150
rect 12992 11086 13044 11092
rect 13176 11086 13228 11092
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13084 10464 13136 10470
rect 13004 10424 13084 10452
rect 13004 6746 13032 10424
rect 13084 10406 13136 10412
rect 13372 10266 13400 11240
rect 13452 11222 13504 11228
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13464 10538 13492 11086
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13462 10364 13770 10384
rect 13462 10362 13468 10364
rect 13524 10362 13548 10364
rect 13604 10362 13628 10364
rect 13684 10362 13708 10364
rect 13764 10362 13770 10364
rect 13524 10310 13526 10362
rect 13706 10310 13708 10362
rect 13462 10308 13468 10310
rect 13524 10308 13548 10310
rect 13604 10308 13628 10310
rect 13684 10308 13708 10310
rect 13764 10308 13770 10310
rect 13462 10288 13770 10308
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13372 9722 13400 10202
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13372 9586 13400 9658
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13372 9178 13400 9522
rect 13462 9276 13770 9296
rect 13462 9274 13468 9276
rect 13524 9274 13548 9276
rect 13604 9274 13628 9276
rect 13684 9274 13708 9276
rect 13764 9274 13770 9276
rect 13524 9222 13526 9274
rect 13706 9222 13708 9274
rect 13462 9220 13468 9222
rect 13524 9220 13548 9222
rect 13604 9220 13628 9222
rect 13684 9220 13708 9222
rect 13764 9220 13770 9222
rect 13462 9200 13770 9220
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13372 8974 13400 9114
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13096 6866 13124 8910
rect 13176 8832 13228 8838
rect 13360 8832 13412 8838
rect 13228 8792 13308 8820
rect 13176 8774 13228 8780
rect 13280 8430 13308 8792
rect 13360 8774 13412 8780
rect 13372 8634 13400 8774
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 7954 13308 8366
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13188 7002 13216 7686
rect 13280 7410 13308 7754
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13176 6792 13228 6798
rect 13004 6718 13124 6746
rect 13280 6780 13308 7346
rect 13228 6752 13308 6780
rect 13176 6734 13228 6740
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13004 5846 13032 6598
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13004 5234 13032 5646
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 12900 1352 12952 1358
rect 12900 1294 12952 1300
rect 10152 734 10364 762
rect 11242 0 11298 800
rect 12438 0 12494 800
rect 13096 762 13124 6718
rect 13372 4622 13400 8298
rect 13462 8188 13770 8208
rect 13462 8186 13468 8188
rect 13524 8186 13548 8188
rect 13604 8186 13628 8188
rect 13684 8186 13708 8188
rect 13764 8186 13770 8188
rect 13524 8134 13526 8186
rect 13706 8134 13708 8186
rect 13462 8132 13468 8134
rect 13524 8132 13548 8134
rect 13604 8132 13628 8134
rect 13684 8132 13708 8134
rect 13764 8132 13770 8134
rect 13462 8112 13770 8132
rect 13832 7954 13860 14554
rect 13924 10266 13952 22102
rect 14476 21894 14504 23598
rect 14660 23050 14688 25298
rect 14648 23044 14700 23050
rect 14648 22986 14700 22992
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 22574 14596 22918
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 14568 22098 14596 22510
rect 14556 22092 14608 22098
rect 14556 22034 14608 22040
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 14556 21888 14608 21894
rect 14556 21830 14608 21836
rect 14476 21078 14504 21830
rect 14568 21690 14596 21830
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 14464 21072 14516 21078
rect 14464 21014 14516 21020
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14476 20466 14504 20742
rect 14660 20534 14688 22986
rect 14752 21162 14780 28642
rect 15476 26308 15528 26314
rect 15476 26250 15528 26256
rect 15488 26042 15516 26250
rect 15476 26036 15528 26042
rect 15476 25978 15528 25984
rect 14924 25900 14976 25906
rect 14924 25842 14976 25848
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14844 24818 14872 25094
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14936 24682 14964 25842
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 14924 24676 14976 24682
rect 14924 24618 14976 24624
rect 15028 24410 15056 25230
rect 15108 25220 15160 25226
rect 15108 25162 15160 25168
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 15120 24206 15148 25162
rect 15384 24880 15436 24886
rect 15384 24822 15436 24828
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 15120 23798 15148 24142
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 15200 22636 15252 22642
rect 15200 22578 15252 22584
rect 14832 22568 14884 22574
rect 14832 22510 14884 22516
rect 14844 21690 14872 22510
rect 15212 22234 15240 22578
rect 15396 22506 15424 24822
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15580 24410 15608 24754
rect 15660 24744 15712 24750
rect 15660 24686 15712 24692
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15672 23526 15700 24686
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15384 22500 15436 22506
rect 15384 22442 15436 22448
rect 15200 22228 15252 22234
rect 15200 22170 15252 22176
rect 15212 22030 15240 22170
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15384 22024 15436 22030
rect 15384 21966 15436 21972
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 15028 21554 15056 21830
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 14752 21134 15056 21162
rect 14924 21072 14976 21078
rect 14924 21014 14976 21020
rect 14832 20936 14884 20942
rect 14832 20878 14884 20884
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14844 20058 14872 20878
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 14016 16250 14044 17206
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 14016 16046 14044 16186
rect 14108 16182 14136 19450
rect 14384 19446 14412 19790
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14752 18426 14780 19178
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14844 18426 14872 18566
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 14200 15552 14228 16050
rect 14108 15524 14228 15552
rect 14108 14414 14136 15524
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14200 14822 14228 15098
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14016 13734 14044 14214
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14016 11694 14044 13670
rect 14108 13462 14136 13942
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 14108 12986 14136 13398
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14200 11558 14228 14758
rect 14292 14618 14320 16934
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14384 15910 14412 16390
rect 14476 16114 14504 17750
rect 14740 17672 14792 17678
rect 14660 17632 14740 17660
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14568 16794 14596 17478
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14568 16658 14596 16730
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14292 14278 14320 14350
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14004 11552 14056 11558
rect 14002 11520 14004 11529
rect 14188 11552 14240 11558
rect 14056 11520 14058 11529
rect 14188 11494 14240 11500
rect 14002 11455 14058 11464
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14108 11082 14136 11222
rect 14292 11218 14320 13194
rect 14384 12434 14412 15846
rect 14476 15706 14504 16050
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14476 14482 14504 15642
rect 14568 14958 14596 16594
rect 14660 16046 14688 17632
rect 14740 17614 14792 17620
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14752 16114 14780 16390
rect 14844 16250 14872 16458
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14936 16130 14964 21014
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14844 16102 14964 16130
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14660 14521 14688 15982
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14646 14512 14702 14521
rect 14464 14476 14516 14482
rect 14646 14447 14648 14456
rect 14464 14418 14516 14424
rect 14700 14447 14702 14456
rect 14648 14418 14700 14424
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14476 13161 14504 13262
rect 14568 13258 14596 13670
rect 14660 13530 14688 14418
rect 14752 13938 14780 14826
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14752 13326 14780 13874
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14462 13152 14518 13161
rect 14462 13087 14518 13096
rect 14384 12406 14596 12434
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14016 10742 14044 11018
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13924 9722 13952 10202
rect 14108 10062 14136 11018
rect 14200 10130 14228 11086
rect 14476 10674 14504 11630
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14200 9586 14228 10066
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 13912 9444 13964 9450
rect 13912 9386 13964 9392
rect 13924 9110 13952 9386
rect 14016 9178 14044 9454
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13924 8566 13952 9046
rect 14384 9042 14412 9658
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14016 8634 14044 8978
rect 14476 8974 14504 9318
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 14016 8430 14044 8570
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13464 7528 13492 7890
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13544 7540 13596 7546
rect 13464 7500 13544 7528
rect 13464 7274 13492 7500
rect 13544 7482 13596 7488
rect 13924 7410 13952 7686
rect 14016 7546 14044 7754
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13462 7100 13770 7120
rect 13462 7098 13468 7100
rect 13524 7098 13548 7100
rect 13604 7098 13628 7100
rect 13684 7098 13708 7100
rect 13764 7098 13770 7100
rect 13524 7046 13526 7098
rect 13706 7046 13708 7098
rect 13462 7044 13468 7046
rect 13524 7044 13548 7046
rect 13604 7044 13628 7046
rect 13684 7044 13708 7046
rect 13764 7044 13770 7046
rect 13462 7024 13770 7044
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14200 6458 14228 6734
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13462 6012 13770 6032
rect 13462 6010 13468 6012
rect 13524 6010 13548 6012
rect 13604 6010 13628 6012
rect 13684 6010 13708 6012
rect 13764 6010 13770 6012
rect 13524 5958 13526 6010
rect 13706 5958 13708 6010
rect 13462 5956 13468 5958
rect 13524 5956 13548 5958
rect 13604 5956 13628 5958
rect 13684 5956 13708 5958
rect 13764 5956 13770 5958
rect 13462 5936 13770 5956
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13462 4924 13770 4944
rect 13462 4922 13468 4924
rect 13524 4922 13548 4924
rect 13604 4922 13628 4924
rect 13684 4922 13708 4924
rect 13764 4922 13770 4924
rect 13524 4870 13526 4922
rect 13706 4870 13708 4922
rect 13462 4868 13468 4870
rect 13524 4868 13548 4870
rect 13604 4868 13628 4870
rect 13684 4868 13708 4870
rect 13764 4868 13770 4870
rect 13462 4848 13770 4868
rect 13832 4622 13860 5034
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13832 4214 13860 4558
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13188 3194 13216 4082
rect 13462 3836 13770 3856
rect 13462 3834 13468 3836
rect 13524 3834 13548 3836
rect 13604 3834 13628 3836
rect 13684 3834 13708 3836
rect 13764 3834 13770 3836
rect 13524 3782 13526 3834
rect 13706 3782 13708 3834
rect 13462 3780 13468 3782
rect 13524 3780 13548 3782
rect 13604 3780 13628 3782
rect 13684 3780 13708 3782
rect 13764 3780 13770 3782
rect 13462 3760 13770 3780
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13280 3058 13308 3674
rect 13924 3126 13952 6190
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 14016 4214 14044 4762
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 14016 3738 14044 4150
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 14108 3670 14136 4422
rect 14292 4282 14320 4558
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 14292 3398 14320 4218
rect 14384 4146 14412 4490
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14476 3942 14504 4422
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14476 3534 14504 3878
rect 14568 3738 14596 12406
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14660 11082 14688 11494
rect 14844 11234 14872 16102
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14936 14414 14964 14758
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 15028 14278 15056 21134
rect 15212 20466 15240 21830
rect 15396 21622 15424 21966
rect 15476 21956 15528 21962
rect 15476 21898 15528 21904
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15488 21418 15516 21898
rect 15476 21412 15528 21418
rect 15476 21354 15528 21360
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 15304 20602 15332 20810
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15304 19514 15332 19722
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15120 18154 15148 18702
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15108 18148 15160 18154
rect 15108 18090 15160 18096
rect 15120 17610 15148 18090
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15304 16522 15332 18158
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15120 14618 15148 14962
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15212 14414 15240 15302
rect 15382 14512 15438 14521
rect 15382 14447 15384 14456
rect 15436 14447 15438 14456
rect 15384 14418 15436 14424
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15212 13954 15240 14010
rect 15212 13926 15332 13954
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14936 12646 14964 13126
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14936 12238 14964 12582
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15028 11694 15056 12786
rect 15106 12336 15162 12345
rect 15106 12271 15162 12280
rect 15120 12238 15148 12271
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15108 11280 15160 11286
rect 14844 11206 14964 11234
rect 15108 11222 15160 11228
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14660 10713 14688 11018
rect 14646 10704 14702 10713
rect 14646 10639 14702 10648
rect 14844 8566 14872 11018
rect 14936 9450 14964 11206
rect 15120 10674 15148 11222
rect 15212 11150 15240 11766
rect 15304 11286 15332 13926
rect 15488 12186 15516 21354
rect 15672 19922 15700 23462
rect 15844 22568 15896 22574
rect 15844 22510 15896 22516
rect 15856 21962 15884 22510
rect 15844 21956 15896 21962
rect 15844 21898 15896 21904
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15764 21690 15792 21830
rect 15752 21684 15804 21690
rect 15752 21626 15804 21632
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15856 19990 15884 20198
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15672 19310 15700 19858
rect 15660 19304 15712 19310
rect 15660 19246 15712 19252
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15580 18426 15608 18634
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15948 17882 15976 28642
rect 16396 26308 16448 26314
rect 16580 26308 16632 26314
rect 16448 26268 16528 26296
rect 16396 26250 16448 26256
rect 16500 25906 16528 26268
rect 16580 26250 16632 26256
rect 16672 26308 16724 26314
rect 16672 26250 16724 26256
rect 16488 25900 16540 25906
rect 16488 25842 16540 25848
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 16120 25764 16172 25770
rect 16120 25706 16172 25712
rect 16132 24818 16160 25706
rect 16408 25158 16436 25774
rect 16396 25152 16448 25158
rect 16396 25094 16448 25100
rect 16408 24818 16436 25094
rect 16500 24886 16528 25842
rect 16592 25702 16620 26250
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16592 25498 16620 25638
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 16488 24880 16540 24886
rect 16488 24822 16540 24828
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16580 24744 16632 24750
rect 16684 24732 16712 26250
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16776 24750 16804 25434
rect 16856 25220 16908 25226
rect 16856 25162 16908 25168
rect 16868 24954 16896 25162
rect 16856 24948 16908 24954
rect 16856 24890 16908 24896
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 16632 24704 16712 24732
rect 16580 24686 16632 24692
rect 16304 24608 16356 24614
rect 16684 24596 16712 24704
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 17052 24596 17080 24754
rect 16684 24568 17080 24596
rect 16304 24550 16356 24556
rect 16316 24274 16344 24550
rect 16304 24268 16356 24274
rect 16304 24210 16356 24216
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16028 24064 16080 24070
rect 16028 24006 16080 24012
rect 16040 23798 16068 24006
rect 16028 23792 16080 23798
rect 16028 23734 16080 23740
rect 16040 23254 16068 23734
rect 16408 23662 16436 24210
rect 17040 24132 17092 24138
rect 17040 24074 17092 24080
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16592 23322 16620 24006
rect 17052 23866 17080 24074
rect 17040 23860 17092 23866
rect 17040 23802 17092 23808
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16028 23248 16080 23254
rect 16028 23190 16080 23196
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 16132 22778 16160 22918
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 16132 22166 16160 22714
rect 16224 22234 16252 22918
rect 16684 22642 16712 23122
rect 16856 23044 16908 23050
rect 16856 22986 16908 22992
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16396 22432 16448 22438
rect 16396 22374 16448 22380
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 16120 22160 16172 22166
rect 16120 22102 16172 22108
rect 16408 22098 16436 22374
rect 16396 22092 16448 22098
rect 16396 22034 16448 22040
rect 16408 21418 16436 22034
rect 16396 21412 16448 21418
rect 16396 21354 16448 21360
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16500 20534 16528 20878
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16396 20392 16448 20398
rect 16396 20334 16448 20340
rect 16408 20058 16436 20334
rect 16500 20058 16528 20470
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19378 16068 19790
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 16592 19174 16620 19654
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15948 17338 15976 17818
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 15978 15884 16526
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15844 15972 15896 15978
rect 15844 15914 15896 15920
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15580 13938 15608 14350
rect 15672 14006 15700 14418
rect 15856 14414 15884 15914
rect 15948 15638 15976 16050
rect 16040 16046 16068 16458
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 16040 15706 16068 15982
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 15948 14550 15976 15574
rect 16040 14618 16068 15642
rect 16132 15162 16160 18566
rect 16408 18358 16436 18566
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 16592 18290 16620 18906
rect 16684 18630 16712 22578
rect 16868 22438 16896 22986
rect 16948 22568 17000 22574
rect 16948 22510 17000 22516
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 16764 22160 16816 22166
rect 16764 22102 16816 22108
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16408 16590 16436 18158
rect 16684 17134 16712 18362
rect 16776 17354 16804 22102
rect 16868 22098 16896 22374
rect 16960 22234 16988 22510
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 16856 22092 16908 22098
rect 17144 22094 17172 28642
rect 17632 27228 17940 27248
rect 17632 27226 17638 27228
rect 17694 27226 17718 27228
rect 17774 27226 17798 27228
rect 17854 27226 17878 27228
rect 17934 27226 17940 27228
rect 17694 27174 17696 27226
rect 17876 27174 17878 27226
rect 17632 27172 17638 27174
rect 17694 27172 17718 27174
rect 17774 27172 17798 27174
rect 17854 27172 17878 27174
rect 17934 27172 17940 27174
rect 17632 27152 17940 27172
rect 17632 26140 17940 26160
rect 17632 26138 17638 26140
rect 17694 26138 17718 26140
rect 17774 26138 17798 26140
rect 17854 26138 17878 26140
rect 17934 26138 17940 26140
rect 17694 26086 17696 26138
rect 17876 26086 17878 26138
rect 17632 26084 17638 26086
rect 17694 26084 17718 26086
rect 17774 26084 17798 26086
rect 17854 26084 17878 26086
rect 17934 26084 17940 26086
rect 17632 26064 17940 26084
rect 17632 25052 17940 25072
rect 17632 25050 17638 25052
rect 17694 25050 17718 25052
rect 17774 25050 17798 25052
rect 17854 25050 17878 25052
rect 17934 25050 17940 25052
rect 17694 24998 17696 25050
rect 17876 24998 17878 25050
rect 17632 24996 17638 24998
rect 17694 24996 17718 24998
rect 17774 24996 17798 24998
rect 17854 24996 17878 24998
rect 17934 24996 17940 24998
rect 17632 24976 17940 24996
rect 17632 23964 17940 23984
rect 17632 23962 17638 23964
rect 17694 23962 17718 23964
rect 17774 23962 17798 23964
rect 17854 23962 17878 23964
rect 17934 23962 17940 23964
rect 17694 23910 17696 23962
rect 17876 23910 17878 23962
rect 17632 23908 17638 23910
rect 17694 23908 17718 23910
rect 17774 23908 17798 23910
rect 17854 23908 17878 23910
rect 17934 23908 17940 23910
rect 17632 23888 17940 23908
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 17512 22778 17540 23666
rect 17632 22876 17940 22896
rect 17632 22874 17638 22876
rect 17694 22874 17718 22876
rect 17774 22874 17798 22876
rect 17854 22874 17878 22876
rect 17934 22874 17940 22876
rect 17694 22822 17696 22874
rect 17876 22822 17878 22874
rect 17632 22820 17638 22822
rect 17694 22820 17718 22822
rect 17774 22820 17798 22822
rect 17854 22820 17878 22822
rect 17934 22820 17940 22822
rect 17632 22800 17940 22820
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17408 22704 17460 22710
rect 17408 22646 17460 22652
rect 17776 22704 17828 22710
rect 17776 22646 17828 22652
rect 17420 22506 17448 22646
rect 17408 22500 17460 22506
rect 17408 22442 17460 22448
rect 17788 22438 17816 22646
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17144 22066 17264 22094
rect 16856 22034 16908 22040
rect 17040 21956 17092 21962
rect 17040 21898 17092 21904
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16960 19922 16988 20742
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16868 17882 16896 19722
rect 17052 18698 17080 21898
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 17144 18902 17172 21354
rect 17236 18970 17264 22066
rect 17632 21788 17940 21808
rect 17632 21786 17638 21788
rect 17694 21786 17718 21788
rect 17774 21786 17798 21788
rect 17854 21786 17878 21788
rect 17934 21786 17940 21788
rect 17694 21734 17696 21786
rect 17876 21734 17878 21786
rect 17632 21732 17638 21734
rect 17694 21732 17718 21734
rect 17774 21732 17798 21734
rect 17854 21732 17878 21734
rect 17934 21732 17940 21734
rect 17632 21712 17940 21732
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17696 21146 17724 21490
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 17632 20700 17940 20720
rect 17632 20698 17638 20700
rect 17694 20698 17718 20700
rect 17774 20698 17798 20700
rect 17854 20698 17878 20700
rect 17934 20698 17940 20700
rect 17694 20646 17696 20698
rect 17876 20646 17878 20698
rect 17632 20644 17638 20646
rect 17694 20644 17718 20646
rect 17774 20644 17798 20646
rect 17854 20644 17878 20646
rect 17934 20644 17940 20646
rect 17632 20624 17940 20644
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17040 18692 17092 18698
rect 17040 18634 17092 18640
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16960 18290 16988 18566
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16960 18086 16988 18226
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 16960 17746 16988 18022
rect 17144 17814 17172 18838
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17132 17808 17184 17814
rect 17132 17750 17184 17756
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 17144 17626 17172 17750
rect 17236 17678 17264 18566
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17052 17598 17172 17626
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17328 17626 17356 18226
rect 17420 18154 17448 19654
rect 17632 19612 17940 19632
rect 17632 19610 17638 19612
rect 17694 19610 17718 19612
rect 17774 19610 17798 19612
rect 17854 19610 17878 19612
rect 17934 19610 17940 19612
rect 17694 19558 17696 19610
rect 17876 19558 17878 19610
rect 17632 19556 17638 19558
rect 17694 19556 17718 19558
rect 17774 19556 17798 19558
rect 17854 19556 17878 19558
rect 17934 19556 17940 19558
rect 17632 19536 17940 19556
rect 17972 19242 18000 28750
rect 18248 28642 18276 28750
rect 18326 28642 18382 29442
rect 19522 28642 19578 29442
rect 20718 28642 20774 29442
rect 21914 28642 21970 29442
rect 23110 28642 23166 29442
rect 24306 28642 24362 29442
rect 25502 28642 25558 29442
rect 26698 28642 26754 29442
rect 18248 28614 18368 28642
rect 21928 27282 21956 28642
rect 21744 27254 21956 27282
rect 21744 25906 21772 27254
rect 21803 26684 22111 26704
rect 21803 26682 21809 26684
rect 21865 26682 21889 26684
rect 21945 26682 21969 26684
rect 22025 26682 22049 26684
rect 22105 26682 22111 26684
rect 21865 26630 21867 26682
rect 22047 26630 22049 26682
rect 21803 26628 21809 26630
rect 21865 26628 21889 26630
rect 21945 26628 21969 26630
rect 22025 26628 22049 26630
rect 22105 26628 22111 26630
rect 21803 26608 22111 26628
rect 23124 25906 23152 28642
rect 25516 25906 25544 28642
rect 26238 28520 26294 28529
rect 26238 28455 26240 28464
rect 26292 28455 26294 28464
rect 26240 28426 26292 28432
rect 21732 25900 21784 25906
rect 21732 25842 21784 25848
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 19248 25696 19300 25702
rect 19248 25638 19300 25644
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 18340 24206 18368 25230
rect 19260 24206 19288 25638
rect 21803 25596 22111 25616
rect 21803 25594 21809 25596
rect 21865 25594 21889 25596
rect 21945 25594 21969 25596
rect 22025 25594 22049 25596
rect 22105 25594 22111 25596
rect 21865 25542 21867 25594
rect 22047 25542 22049 25594
rect 21803 25540 21809 25542
rect 21865 25540 21889 25542
rect 21945 25540 21969 25542
rect 22025 25540 22049 25542
rect 22105 25540 22111 25542
rect 21803 25520 22111 25540
rect 25042 25392 25098 25401
rect 25042 25327 25044 25336
rect 25096 25327 25098 25336
rect 25044 25298 25096 25304
rect 21803 24508 22111 24528
rect 21803 24506 21809 24508
rect 21865 24506 21889 24508
rect 21945 24506 21969 24508
rect 22025 24506 22049 24508
rect 22105 24506 22111 24508
rect 21865 24454 21867 24506
rect 22047 24454 22049 24506
rect 21803 24452 21809 24454
rect 21865 24452 21889 24454
rect 21945 24452 21969 24454
rect 22025 24452 22049 24454
rect 22105 24452 22111 24454
rect 21803 24432 22111 24452
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 18604 24132 18656 24138
rect 18604 24074 18656 24080
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18524 23798 18552 24006
rect 18052 23792 18104 23798
rect 18052 23734 18104 23740
rect 18512 23792 18564 23798
rect 18512 23734 18564 23740
rect 18064 23050 18092 23734
rect 18524 23662 18552 23734
rect 18616 23730 18644 24074
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18892 23662 18920 24142
rect 18972 23860 19024 23866
rect 18972 23802 19024 23808
rect 18512 23656 18564 23662
rect 18512 23598 18564 23604
rect 18880 23656 18932 23662
rect 18880 23598 18932 23604
rect 18892 23254 18920 23598
rect 18512 23248 18564 23254
rect 18512 23190 18564 23196
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 18524 22438 18552 23190
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18708 22642 18736 23122
rect 18984 22642 19012 23802
rect 19156 23724 19208 23730
rect 19156 23666 19208 23672
rect 19168 22982 19196 23666
rect 19536 23526 19564 24142
rect 20444 24132 20496 24138
rect 20444 24074 20496 24080
rect 19616 24064 19668 24070
rect 19616 24006 19668 24012
rect 19248 23520 19300 23526
rect 19524 23520 19576 23526
rect 19300 23468 19380 23474
rect 19248 23462 19380 23468
rect 19524 23462 19576 23468
rect 19260 23446 19380 23462
rect 19352 23186 19380 23446
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18420 21412 18472 21418
rect 18420 21354 18472 21360
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 18064 20602 18092 20946
rect 18340 20942 18368 21286
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18052 19780 18104 19786
rect 18052 19722 18104 19728
rect 18064 19446 18092 19722
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 17960 19236 18012 19242
rect 17960 19178 18012 19184
rect 18248 18714 18276 20334
rect 18340 19378 18368 20878
rect 18432 20380 18460 21354
rect 18524 20942 18552 22374
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18524 20534 18552 20878
rect 18708 20806 18736 22578
rect 19352 22506 19380 22986
rect 19536 22574 19564 23462
rect 19628 22710 19656 24006
rect 20456 23730 20484 24074
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 21803 23420 22111 23440
rect 21803 23418 21809 23420
rect 21865 23418 21889 23420
rect 21945 23418 21969 23420
rect 22025 23418 22049 23420
rect 22105 23418 22111 23420
rect 21865 23366 21867 23418
rect 22047 23366 22049 23418
rect 21803 23364 21809 23366
rect 21865 23364 21889 23366
rect 21945 23364 21969 23366
rect 22025 23364 22049 23366
rect 22105 23364 22111 23366
rect 21803 23344 22111 23364
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 19708 22976 19760 22982
rect 19708 22918 19760 22924
rect 19720 22778 19748 22918
rect 19904 22778 19932 23054
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19892 22772 19944 22778
rect 19892 22714 19944 22720
rect 19616 22704 19668 22710
rect 19616 22646 19668 22652
rect 19708 22636 19760 22642
rect 19708 22578 19760 22584
rect 19524 22568 19576 22574
rect 19524 22510 19576 22516
rect 19720 22506 19748 22578
rect 18788 22500 18840 22506
rect 18788 22442 18840 22448
rect 19340 22500 19392 22506
rect 19340 22442 19392 22448
rect 19708 22500 19760 22506
rect 19708 22442 19760 22448
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18432 20352 18552 20380
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18432 20058 18460 20198
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18156 18686 18276 18714
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17512 18222 17540 18566
rect 17632 18524 17940 18544
rect 17632 18522 17638 18524
rect 17694 18522 17718 18524
rect 17774 18522 17798 18524
rect 17854 18522 17878 18524
rect 17934 18522 17940 18524
rect 17694 18470 17696 18522
rect 17876 18470 17878 18522
rect 17632 18468 17638 18470
rect 17694 18468 17718 18470
rect 17774 18468 17798 18470
rect 17854 18468 17878 18470
rect 17934 18468 17940 18470
rect 17632 18448 17940 18468
rect 18156 18290 18184 18686
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17408 18148 17460 18154
rect 17408 18090 17460 18096
rect 17328 17598 17448 17626
rect 16776 17326 16896 17354
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16408 16046 16436 16526
rect 16684 16046 16712 17070
rect 16776 16794 16804 17138
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16684 15026 16712 15982
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 14074 15884 14350
rect 15936 14340 15988 14346
rect 15988 14300 16068 14328
rect 15936 14282 15988 14288
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15580 13682 15608 13874
rect 15580 13654 15700 13682
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 12306 15608 12786
rect 15672 12345 15700 13654
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15752 12368 15804 12374
rect 15658 12336 15714 12345
rect 15568 12300 15620 12306
rect 15752 12310 15804 12316
rect 15658 12271 15714 12280
rect 15568 12242 15620 12248
rect 15384 12164 15436 12170
rect 15488 12158 15608 12186
rect 15384 12106 15436 12112
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15292 11144 15344 11150
rect 15396 11132 15424 12106
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15344 11104 15424 11132
rect 15292 11086 15344 11092
rect 15488 10674 15516 12038
rect 15580 10810 15608 12158
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15672 11354 15700 11698
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15764 11218 15792 12310
rect 15948 12238 15976 12854
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 15028 8906 15056 10542
rect 15120 10130 15148 10610
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15212 9926 15240 10542
rect 15488 10266 15516 10610
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15488 9586 15516 9862
rect 15580 9722 15608 10746
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 15028 8634 15056 8842
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 15028 7886 15056 8570
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14844 6322 14872 6598
rect 14936 6458 14964 6598
rect 15028 6458 15056 7822
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14660 5574 14688 6190
rect 15120 5710 15148 6326
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14752 3398 14780 3946
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14844 3194 14872 3470
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 14936 2922 14964 4422
rect 15120 4214 15148 4626
rect 15212 4622 15240 9046
rect 15304 8906 15332 9318
rect 15580 8906 15608 9658
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15844 8900 15896 8906
rect 15844 8842 15896 8848
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15396 5914 15424 6598
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15304 5166 15332 5510
rect 15488 5234 15516 6802
rect 15672 6798 15700 8774
rect 15856 8634 15884 8842
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15488 4758 15516 5170
rect 15580 5098 15608 6598
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15672 5778 15700 6054
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15764 5370 15792 6258
rect 15856 5710 15884 6666
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15568 5092 15620 5098
rect 15568 5034 15620 5040
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15764 4554 15792 5102
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15304 4214 15332 4422
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15120 4078 15148 4150
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 15028 2990 15056 3674
rect 15764 3126 15792 4490
rect 15856 3738 15884 5646
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 13462 2748 13770 2768
rect 13462 2746 13468 2748
rect 13524 2746 13548 2748
rect 13604 2746 13628 2748
rect 13684 2746 13708 2748
rect 13764 2746 13770 2748
rect 13524 2694 13526 2746
rect 13706 2694 13708 2746
rect 13462 2692 13468 2694
rect 13524 2692 13548 2694
rect 13604 2692 13628 2694
rect 13684 2692 13708 2694
rect 13764 2692 13770 2694
rect 13462 2672 13770 2692
rect 13556 870 13676 898
rect 13556 762 13584 870
rect 13648 800 13676 870
rect 14752 800 14780 2790
rect 15948 800 15976 11086
rect 16040 2854 16068 14300
rect 16408 11830 16436 14758
rect 16776 14618 16804 14962
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16500 14074 16528 14282
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16396 11824 16448 11830
rect 16396 11766 16448 11772
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 11150 16160 11494
rect 16592 11286 16620 12242
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 11762 16712 12038
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16580 11280 16632 11286
rect 16578 11248 16580 11257
rect 16632 11248 16634 11257
rect 16578 11183 16634 11192
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16488 11144 16540 11150
rect 16776 11132 16804 12310
rect 16868 11898 16896 17326
rect 17052 16794 17080 17598
rect 17132 17536 17184 17542
rect 17316 17536 17368 17542
rect 17184 17496 17264 17524
rect 17132 17478 17184 17484
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 17236 16726 17264 17496
rect 17316 17478 17368 17484
rect 17224 16720 17276 16726
rect 17224 16662 17276 16668
rect 17236 14074 17264 16662
rect 17328 16658 17356 17478
rect 17420 17202 17448 17598
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17420 16590 17448 17138
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17420 13870 17448 14214
rect 17512 13954 17540 18158
rect 18064 17882 18092 18226
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17632 17436 17940 17456
rect 17632 17434 17638 17436
rect 17694 17434 17718 17436
rect 17774 17434 17798 17436
rect 17854 17434 17878 17436
rect 17934 17434 17940 17436
rect 17694 17382 17696 17434
rect 17876 17382 17878 17434
rect 17632 17380 17638 17382
rect 17694 17380 17718 17382
rect 17774 17380 17798 17382
rect 17854 17380 17878 17382
rect 17934 17380 17940 17382
rect 17632 17360 17940 17380
rect 17972 16658 18000 17614
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 18064 16522 18092 17274
rect 18156 17134 18184 18226
rect 18248 17270 18276 18566
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18432 17542 18460 18226
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 17632 16348 17940 16368
rect 17632 16346 17638 16348
rect 17694 16346 17718 16348
rect 17774 16346 17798 16348
rect 17854 16346 17878 16348
rect 17934 16346 17940 16348
rect 17694 16294 17696 16346
rect 17876 16294 17878 16346
rect 17632 16292 17638 16294
rect 17694 16292 17718 16294
rect 17774 16292 17798 16294
rect 17854 16292 17878 16294
rect 17934 16292 17940 16294
rect 17632 16272 17940 16292
rect 17632 15260 17940 15280
rect 17632 15258 17638 15260
rect 17694 15258 17718 15260
rect 17774 15258 17798 15260
rect 17854 15258 17878 15260
rect 17934 15258 17940 15260
rect 17694 15206 17696 15258
rect 17876 15206 17878 15258
rect 17632 15204 17638 15206
rect 17694 15204 17718 15206
rect 17774 15204 17798 15206
rect 17854 15204 17878 15206
rect 17934 15204 17940 15206
rect 17632 15184 17940 15204
rect 18156 15162 18184 16662
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 18248 15434 18276 16594
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18340 15434 18368 16390
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18156 14958 18184 15098
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 17960 14408 18012 14414
rect 18156 14396 18184 14758
rect 18248 14414 18276 15370
rect 18340 14482 18368 15370
rect 18432 15314 18460 17478
rect 18524 17202 18552 20352
rect 18616 17882 18644 20402
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 18708 19514 18736 20334
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18524 16794 18552 17138
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18524 16658 18552 16730
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 18512 15360 18564 15366
rect 18432 15308 18512 15314
rect 18432 15302 18564 15308
rect 18432 15286 18552 15302
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18012 14368 18184 14396
rect 17960 14350 18012 14356
rect 17632 14172 17940 14192
rect 17632 14170 17638 14172
rect 17694 14170 17718 14172
rect 17774 14170 17798 14172
rect 17854 14170 17878 14172
rect 17934 14170 17940 14172
rect 17694 14118 17696 14170
rect 17876 14118 17878 14170
rect 17632 14116 17638 14118
rect 17694 14116 17718 14118
rect 17774 14116 17798 14118
rect 17854 14116 17878 14118
rect 17934 14116 17940 14118
rect 17632 14096 17940 14116
rect 18156 13954 18184 14368
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18340 14074 18368 14418
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 17512 13938 17632 13954
rect 17512 13932 17644 13938
rect 17512 13926 17592 13932
rect 18156 13926 18276 13954
rect 18432 13938 18460 15286
rect 18616 14346 18644 15370
rect 18708 14550 18736 15438
rect 18800 15162 18828 22442
rect 19720 22030 19748 22442
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18892 20262 18920 21422
rect 18972 20868 19024 20874
rect 18972 20810 19024 20816
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18892 19446 18920 20198
rect 18984 20058 19012 20810
rect 19168 20516 19196 21490
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19248 20528 19300 20534
rect 19168 20488 19248 20516
rect 19064 20460 19116 20466
rect 19168 20448 19196 20488
rect 19248 20470 19300 20476
rect 19116 20420 19196 20448
rect 19064 20402 19116 20408
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 19076 19378 19104 20402
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19444 19990 19472 20266
rect 19432 19984 19484 19990
rect 19432 19926 19484 19932
rect 19536 19802 19564 20742
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19798 20360 19854 20369
rect 19798 20295 19854 20304
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19628 20058 19656 20198
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19536 19774 19656 19802
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19536 19514 19564 19654
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19628 19446 19656 19774
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 19706 19408 19762 19417
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 19628 18766 19656 19382
rect 19706 19343 19708 19352
rect 19760 19343 19762 19352
rect 19708 19314 19760 19320
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19248 18148 19300 18154
rect 19248 18090 19300 18096
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 19076 17678 19104 18022
rect 19260 17746 19288 18090
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19168 17338 19196 17614
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19260 16794 19288 17682
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19628 17338 19656 17478
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19444 17134 19472 17206
rect 19812 17202 19840 20295
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19260 16250 19288 16730
rect 19340 16720 19392 16726
rect 19444 16708 19472 17070
rect 19536 16776 19564 17070
rect 19616 16788 19668 16794
rect 19536 16748 19616 16776
rect 19616 16730 19668 16736
rect 19392 16680 19472 16708
rect 19340 16662 19392 16668
rect 19444 16454 19472 16680
rect 19720 16658 19748 17138
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19536 16266 19564 16526
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19444 16238 19564 16266
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18604 14340 18656 14346
rect 18604 14282 18656 14288
rect 17592 13874 17644 13880
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16868 11218 16896 11834
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16540 11104 16804 11132
rect 16488 11086 16540 11092
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 3466 16160 7142
rect 16316 6866 16344 8434
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16316 6202 16344 6802
rect 16408 6730 16436 7890
rect 16500 7342 16528 8366
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16592 6866 16620 10950
rect 16684 9518 16712 11104
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16776 6798 16804 7414
rect 16868 7410 16896 11018
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16776 6458 16804 6598
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16316 6174 16436 6202
rect 16408 6118 16436 6174
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16316 5642 16344 6054
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16500 5642 16528 5850
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16500 5302 16528 5578
rect 16592 5370 16620 6258
rect 16960 5370 16988 11494
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17052 9178 17080 10746
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 17144 8634 17172 13126
rect 17236 12374 17264 13738
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17328 13326 17356 13670
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17512 13240 17540 13466
rect 17604 13394 17632 13874
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17696 13240 17724 13330
rect 18156 13326 18184 13670
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 17512 13212 17724 13240
rect 17512 12782 17540 13212
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17632 13084 17940 13104
rect 17632 13082 17638 13084
rect 17694 13082 17718 13084
rect 17774 13082 17798 13084
rect 17854 13082 17878 13084
rect 17934 13082 17940 13084
rect 17694 13030 17696 13082
rect 17876 13030 17878 13082
rect 17632 13028 17638 13030
rect 17694 13028 17718 13030
rect 17774 13028 17798 13030
rect 17854 13028 17878 13030
rect 17934 13028 17940 13030
rect 17632 13008 17940 13028
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 12374 17540 12718
rect 17224 12368 17276 12374
rect 17500 12368 17552 12374
rect 17276 12328 17356 12356
rect 17224 12310 17276 12316
rect 17328 11762 17356 12328
rect 17500 12310 17552 12316
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17512 11694 17540 12310
rect 17632 11996 17940 12016
rect 17632 11994 17638 11996
rect 17694 11994 17718 11996
rect 17774 11994 17798 11996
rect 17854 11994 17878 11996
rect 17934 11994 17940 11996
rect 17694 11942 17696 11994
rect 17876 11942 17878 11994
rect 17632 11940 17638 11942
rect 17694 11940 17718 11942
rect 17774 11940 17798 11942
rect 17854 11940 17878 11942
rect 17934 11940 17940 11942
rect 17632 11920 17940 11940
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17224 11552 17276 11558
rect 17222 11520 17224 11529
rect 17276 11520 17278 11529
rect 17222 11455 17278 11464
rect 17512 11286 17540 11630
rect 17500 11280 17552 11286
rect 17500 11222 17552 11228
rect 17512 10810 17540 11222
rect 17632 10908 17940 10928
rect 17632 10906 17638 10908
rect 17694 10906 17718 10908
rect 17774 10906 17798 10908
rect 17854 10906 17878 10908
rect 17934 10906 17940 10908
rect 17694 10854 17696 10906
rect 17876 10854 17878 10906
rect 17632 10852 17638 10854
rect 17694 10852 17718 10854
rect 17774 10852 17798 10854
rect 17854 10852 17878 10854
rect 17934 10852 17940 10854
rect 17632 10832 17940 10852
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17632 9820 17940 9840
rect 17632 9818 17638 9820
rect 17694 9818 17718 9820
rect 17774 9818 17798 9820
rect 17854 9818 17878 9820
rect 17934 9818 17940 9820
rect 17694 9766 17696 9818
rect 17876 9766 17878 9818
rect 17632 9764 17638 9766
rect 17694 9764 17718 9766
rect 17774 9764 17798 9766
rect 17854 9764 17878 9766
rect 17934 9764 17940 9766
rect 17632 9744 17940 9764
rect 17972 9654 18000 13126
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18156 11898 18184 12922
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17144 8090 17172 8366
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17236 8022 17264 9386
rect 17328 8090 17356 9522
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17420 7886 17448 8774
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17040 7812 17092 7818
rect 17040 7754 17092 7760
rect 17052 7342 17080 7754
rect 17420 7546 17448 7822
rect 17512 7818 17540 9318
rect 17972 9042 18000 9386
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17632 8732 17940 8752
rect 17632 8730 17638 8732
rect 17694 8730 17718 8732
rect 17774 8730 17798 8732
rect 17854 8730 17878 8732
rect 17934 8730 17940 8732
rect 17694 8678 17696 8730
rect 17876 8678 17878 8730
rect 17632 8676 17638 8678
rect 17694 8676 17718 8678
rect 17774 8676 17798 8678
rect 17854 8676 17878 8678
rect 17934 8676 17940 8678
rect 17632 8656 17940 8676
rect 17972 8616 18000 8978
rect 18064 8634 18092 9454
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17880 8588 18000 8616
rect 18052 8628 18104 8634
rect 17880 8430 17908 8588
rect 18052 8570 18104 8576
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17632 7644 17940 7664
rect 17632 7642 17638 7644
rect 17694 7642 17718 7644
rect 17774 7642 17798 7644
rect 17854 7642 17878 7644
rect 17934 7642 17940 7644
rect 17694 7590 17696 7642
rect 17876 7590 17878 7642
rect 17632 7588 17638 7590
rect 17694 7588 17718 7590
rect 17774 7588 17798 7590
rect 17854 7588 17878 7590
rect 17934 7588 17940 7590
rect 17632 7568 17940 7588
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17972 7410 18000 8434
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 18156 7206 18184 8774
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 17632 6556 17940 6576
rect 17632 6554 17638 6556
rect 17694 6554 17718 6556
rect 17774 6554 17798 6556
rect 17854 6554 17878 6556
rect 17934 6554 17940 6556
rect 17694 6502 17696 6554
rect 17876 6502 17878 6554
rect 17632 6500 17638 6502
rect 17694 6500 17718 6502
rect 17774 6500 17798 6502
rect 17854 6500 17878 6502
rect 17934 6500 17940 6502
rect 17632 6480 17940 6500
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17144 5574 17172 6190
rect 17328 5710 17356 6190
rect 17500 6180 17552 6186
rect 17500 6122 17552 6128
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17512 5642 17540 6122
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16500 4214 16528 5238
rect 16592 4690 16620 5306
rect 17144 5234 17172 5510
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16776 4758 16804 4966
rect 17236 4826 17264 5306
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16500 3942 16528 4150
rect 16592 4146 16620 4490
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16592 3670 16620 4082
rect 16776 3670 16804 4490
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17144 4146 17172 4422
rect 17420 4214 17448 5170
rect 17512 5030 17540 5578
rect 17632 5468 17940 5488
rect 17632 5466 17638 5468
rect 17694 5466 17718 5468
rect 17774 5466 17798 5468
rect 17854 5466 17878 5468
rect 17934 5466 17940 5468
rect 17694 5414 17696 5466
rect 17876 5414 17878 5466
rect 17632 5412 17638 5414
rect 17694 5412 17718 5414
rect 17774 5412 17798 5414
rect 17854 5412 17878 5414
rect 17934 5412 17940 5414
rect 17632 5392 17940 5412
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17696 4758 17724 5102
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 18064 4622 18092 4966
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17632 4380 17940 4400
rect 17632 4378 17638 4380
rect 17694 4378 17718 4380
rect 17774 4378 17798 4380
rect 17854 4378 17878 4380
rect 17934 4378 17940 4380
rect 17694 4326 17696 4378
rect 17876 4326 17878 4378
rect 17632 4324 17638 4326
rect 17694 4324 17718 4326
rect 17774 4324 17798 4326
rect 17854 4324 17878 4326
rect 17934 4324 17940 4326
rect 17632 4304 17940 4324
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 18248 4010 18276 13926
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18432 13394 18460 13874
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18800 12986 18828 15098
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18432 12374 18460 12786
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18340 11830 18368 12174
rect 18524 11898 18552 12174
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18340 11354 18368 11766
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18340 10742 18368 11290
rect 18420 11144 18472 11150
rect 18616 11132 18644 12174
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18800 11762 18828 12106
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18800 11218 18828 11698
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18892 11286 18920 11630
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18472 11104 18644 11132
rect 18420 11086 18472 11092
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18432 10538 18460 11086
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18340 7410 18368 7686
rect 18616 7546 18644 8434
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18432 5302 18460 5510
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 17144 800 17172 3946
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17328 3534 17356 3878
rect 18892 3738 18920 5102
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17632 3292 17940 3312
rect 17632 3290 17638 3292
rect 17694 3290 17718 3292
rect 17774 3290 17798 3292
rect 17854 3290 17878 3292
rect 17934 3290 17940 3292
rect 17694 3238 17696 3290
rect 17876 3238 17878 3290
rect 17632 3236 17638 3238
rect 17694 3236 17718 3238
rect 17774 3236 17798 3238
rect 17854 3236 17878 3238
rect 17934 3236 17940 3238
rect 17632 3216 17940 3236
rect 18984 2774 19012 15846
rect 19260 15706 19288 16186
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19260 15570 19288 15642
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19076 14074 19104 14894
rect 19444 14618 19472 16238
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19628 15162 19656 15302
rect 19616 15156 19668 15162
rect 19616 15098 19668 15104
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19536 14890 19564 14962
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19248 14340 19300 14346
rect 19248 14282 19300 14288
rect 19260 14074 19288 14282
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19444 13938 19472 14554
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19536 13920 19564 14826
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19628 14482 19656 14758
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19720 14346 19748 16594
rect 19812 16590 19840 16934
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19904 16454 19932 20402
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19996 15706 20024 22986
rect 20260 22976 20312 22982
rect 20260 22918 20312 22924
rect 20272 22234 20300 22918
rect 20364 22642 20392 23054
rect 22192 23044 22244 23050
rect 22192 22986 22244 22992
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 20352 22636 20404 22642
rect 20352 22578 20404 22584
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20180 20058 20208 20810
rect 20272 20806 20300 22170
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20548 20398 20576 20742
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20548 19718 20576 20334
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20456 18698 20484 19450
rect 20548 19174 20576 19654
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20628 18896 20680 18902
rect 20628 18838 20680 18844
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20640 18290 20668 18838
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20732 17082 20760 22578
rect 20904 22568 20956 22574
rect 20904 22510 20956 22516
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 20916 21622 20944 22510
rect 21100 22234 21128 22510
rect 22112 22420 22140 22918
rect 22204 22778 22232 22986
rect 23204 22976 23256 22982
rect 23204 22918 23256 22924
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 23216 22642 23244 22918
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 22112 22392 22232 22420
rect 21803 22332 22111 22352
rect 21803 22330 21809 22332
rect 21865 22330 21889 22332
rect 21945 22330 21969 22332
rect 22025 22330 22049 22332
rect 22105 22330 22111 22332
rect 21865 22278 21867 22330
rect 22047 22278 22049 22330
rect 21803 22276 21809 22278
rect 21865 22276 21889 22278
rect 21945 22276 21969 22278
rect 22025 22276 22049 22278
rect 22105 22276 22111 22278
rect 21803 22256 22111 22276
rect 21088 22228 21140 22234
rect 21088 22170 21140 22176
rect 22204 21622 22232 22392
rect 22296 22166 22324 22578
rect 22376 22432 22428 22438
rect 22376 22374 22428 22380
rect 22388 22234 22416 22374
rect 22376 22228 22428 22234
rect 22376 22170 22428 22176
rect 22284 22160 22336 22166
rect 22284 22102 22336 22108
rect 20904 21616 20956 21622
rect 20904 21558 20956 21564
rect 21732 21616 21784 21622
rect 21732 21558 21784 21564
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 22468 21616 22520 21622
rect 22468 21558 22520 21564
rect 21744 21010 21772 21558
rect 21803 21244 22111 21264
rect 21803 21242 21809 21244
rect 21865 21242 21889 21244
rect 21945 21242 21969 21244
rect 22025 21242 22049 21244
rect 22105 21242 22111 21244
rect 21865 21190 21867 21242
rect 22047 21190 22049 21242
rect 21803 21188 21809 21190
rect 21865 21188 21889 21190
rect 21945 21188 21969 21190
rect 22025 21188 22049 21190
rect 22105 21188 22111 21190
rect 21803 21168 22111 21188
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21468 20466 21496 20742
rect 21560 20534 21588 20742
rect 22388 20602 22416 20878
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22480 20534 22508 21558
rect 21548 20528 21600 20534
rect 21548 20470 21600 20476
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21560 19854 21588 20334
rect 21803 20156 22111 20176
rect 21803 20154 21809 20156
rect 21865 20154 21889 20156
rect 21945 20154 21969 20156
rect 22025 20154 22049 20156
rect 22105 20154 22111 20156
rect 21865 20102 21867 20154
rect 22047 20102 22049 20154
rect 21803 20100 21809 20102
rect 21865 20100 21889 20102
rect 21945 20100 21969 20102
rect 22025 20100 22049 20102
rect 22105 20100 22111 20102
rect 21803 20080 22111 20100
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 20824 18766 20852 19790
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 22468 19780 22520 19786
rect 22468 19722 22520 19728
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21192 19514 21220 19654
rect 21468 19514 21496 19722
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 22480 19446 22508 19722
rect 22468 19440 22520 19446
rect 22468 19382 22520 19388
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20824 18426 20852 18702
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20824 18154 20852 18362
rect 20916 18290 20944 19246
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20812 18148 20864 18154
rect 20812 18090 20864 18096
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20732 17054 20852 17082
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20732 16590 20760 16934
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20272 15706 20300 16390
rect 20824 16250 20852 17054
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20916 16182 20944 17274
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20640 15570 20760 15586
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20640 15564 20772 15570
rect 20640 15558 20720 15564
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20180 15162 20208 15438
rect 20548 15366 20576 15506
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19708 14340 19760 14346
rect 19708 14282 19760 14288
rect 19616 13932 19668 13938
rect 19536 13892 19616 13920
rect 19076 12850 19104 13874
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19352 12782 19380 13330
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 8974 19104 12038
rect 19352 11762 19380 12106
rect 19536 11898 19564 13892
rect 19616 13874 19668 13880
rect 19720 12306 19748 14282
rect 19996 14006 20024 15030
rect 20548 15026 20576 15302
rect 20640 15162 20668 15558
rect 20720 15506 20772 15512
rect 20916 15450 20944 16118
rect 21008 15978 21036 19314
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21284 19174 21312 19246
rect 22192 19236 22244 19242
rect 22192 19178 22244 19184
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 21100 18426 21128 18634
rect 21088 18420 21140 18426
rect 21088 18362 21140 18368
rect 21284 18358 21312 19110
rect 21803 19068 22111 19088
rect 21803 19066 21809 19068
rect 21865 19066 21889 19068
rect 21945 19066 21969 19068
rect 22025 19066 22049 19068
rect 22105 19066 22111 19068
rect 21865 19014 21867 19066
rect 22047 19014 22049 19066
rect 21803 19012 21809 19014
rect 21865 19012 21889 19014
rect 21945 19012 21969 19014
rect 22025 19012 22049 19014
rect 22105 19012 22111 19014
rect 21803 18992 22111 19012
rect 22204 18970 22232 19178
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21376 18426 21404 18566
rect 21744 18426 21772 18906
rect 22296 18426 22324 19110
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21732 18420 21784 18426
rect 21732 18362 21784 18368
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 21272 18352 21324 18358
rect 21272 18294 21324 18300
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 21803 17980 22111 18000
rect 21803 17978 21809 17980
rect 21865 17978 21889 17980
rect 21945 17978 21969 17980
rect 22025 17978 22049 17980
rect 22105 17978 22111 17980
rect 21865 17926 21867 17978
rect 22047 17926 22049 17978
rect 21803 17924 21809 17926
rect 21865 17924 21889 17926
rect 21945 17924 21969 17926
rect 22025 17924 22049 17926
rect 22105 17924 22111 17926
rect 21803 17904 22111 17924
rect 21548 17264 21600 17270
rect 21548 17206 21600 17212
rect 21560 16658 21588 17206
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 16250 21220 16390
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 20996 15972 21048 15978
rect 20996 15914 21048 15920
rect 21100 15706 21128 16050
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 20732 15422 20944 15450
rect 20996 15496 21048 15502
rect 21284 15450 21312 16186
rect 21468 15638 21496 16186
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21560 15570 21588 16594
rect 21744 16590 21772 16934
rect 21803 16892 22111 16912
rect 21803 16890 21809 16892
rect 21865 16890 21889 16892
rect 21945 16890 21969 16892
rect 22025 16890 22049 16892
rect 22105 16890 22111 16892
rect 21865 16838 21867 16890
rect 22047 16838 22049 16890
rect 21803 16836 21809 16838
rect 21865 16836 21889 16838
rect 21945 16836 21969 16838
rect 22025 16836 22049 16838
rect 22105 16836 22111 16838
rect 21803 16816 22111 16836
rect 22204 16674 22232 17138
rect 22112 16646 22232 16674
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 22112 16522 22140 16646
rect 22100 16516 22152 16522
rect 22100 16458 22152 16464
rect 22112 16130 22140 16458
rect 22572 16454 22600 18226
rect 22664 16454 22692 22578
rect 23020 22568 23072 22574
rect 23020 22510 23072 22516
rect 23032 22166 23060 22510
rect 23020 22160 23072 22166
rect 23020 22102 23072 22108
rect 23400 21554 23428 23054
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 21962 23520 22918
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 23664 22636 23716 22642
rect 23664 22578 23716 22584
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 24676 22636 24728 22642
rect 24676 22578 24728 22584
rect 23480 21956 23532 21962
rect 23480 21898 23532 21904
rect 23492 21622 23520 21898
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 22836 20936 22888 20942
rect 22836 20878 22888 20884
rect 22848 19922 22876 20878
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22756 19514 22784 19790
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22848 19310 22876 19858
rect 23308 19854 23336 21082
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 23216 18834 23244 19314
rect 23308 19174 23336 19790
rect 23584 19446 23612 21830
rect 23676 21350 23704 22578
rect 23848 22432 23900 22438
rect 23848 22374 23900 22380
rect 23860 22098 23888 22374
rect 23848 22092 23900 22098
rect 23848 22034 23900 22040
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23848 21888 23900 21894
rect 23848 21830 23900 21836
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 20942 23704 21286
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23492 18630 23520 19110
rect 23584 18698 23612 19382
rect 23676 18970 23704 20470
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23572 18692 23624 18698
rect 23572 18634 23624 18640
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23386 17776 23442 17785
rect 23386 17711 23442 17720
rect 23400 17678 23428 17711
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 23216 16658 23244 16934
rect 23204 16652 23256 16658
rect 23204 16594 23256 16600
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22848 16250 22876 16526
rect 22928 16516 22980 16522
rect 22928 16458 22980 16464
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22374 16144 22430 16153
rect 21640 16108 21692 16114
rect 22112 16102 22232 16130
rect 21640 16050 21692 16056
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 21048 15444 21312 15450
rect 20996 15438 21312 15444
rect 21008 15422 21312 15438
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20088 14074 20116 14350
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 20272 13920 20300 14418
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20456 13938 20484 14350
rect 20352 13932 20404 13938
rect 20272 13892 20352 13920
rect 20352 13874 20404 13880
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20364 13530 20392 13874
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20364 13190 20392 13330
rect 20456 13326 20484 13874
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19812 12306 19840 12718
rect 20364 12374 20392 13126
rect 20352 12368 20404 12374
rect 20352 12310 20404 12316
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19628 11898 19656 12038
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19720 11830 19748 12242
rect 19812 11880 19840 12242
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 19892 11892 19944 11898
rect 19812 11852 19892 11880
rect 19892 11834 19944 11840
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 20456 11762 20484 12106
rect 20548 11830 20576 14962
rect 20732 14958 20760 15422
rect 21284 15162 21312 15422
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20824 14550 20852 14962
rect 21100 14822 21128 14962
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21100 14618 21128 14758
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 20824 13938 20852 14214
rect 21192 13938 21220 14214
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20916 12986 20944 13126
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 20824 12374 20852 12786
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 20812 12368 20864 12374
rect 20812 12310 20864 12316
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20456 11354 20484 11698
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 19352 10810 19380 11222
rect 20548 11150 20576 11766
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20732 11558 20760 11698
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19628 10742 19656 11086
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 19352 8566 19380 8978
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19352 8090 19380 8502
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19536 7750 19564 8434
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19064 6724 19116 6730
rect 19064 6666 19116 6672
rect 19076 6458 19104 6666
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19076 6202 19104 6394
rect 19536 6390 19564 7346
rect 19720 6458 19748 10406
rect 20916 10062 20944 12038
rect 21008 11354 21036 12038
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19812 8566 19840 9454
rect 20074 9208 20130 9217
rect 20074 9143 20076 9152
rect 20128 9143 20130 9152
rect 20076 9114 20128 9120
rect 20258 9072 20314 9081
rect 20258 9007 20314 9016
rect 20272 8974 20300 9007
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19800 8560 19852 8566
rect 19800 8502 19852 8508
rect 19812 7750 19840 8502
rect 19996 8430 20024 8842
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20180 8498 20208 8774
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19904 7954 19932 8366
rect 19996 8090 20024 8366
rect 20180 8362 20208 8434
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19812 7546 19840 7686
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 20180 7274 20208 8298
rect 20272 7886 20300 8910
rect 20548 8566 20576 9862
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20640 8974 20668 9522
rect 20732 9382 20760 9998
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20536 8560 20588 8566
rect 20536 8502 20588 8508
rect 20824 8022 20852 9862
rect 21100 9654 21128 12582
rect 21192 11218 21220 13874
rect 21284 13326 21312 15098
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21376 13530 21404 13874
rect 21456 13796 21508 13802
rect 21456 13738 21508 13744
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21468 13394 21496 13738
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21284 12986 21312 13262
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21468 12306 21496 12718
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21180 11212 21232 11218
rect 21180 11154 21232 11160
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20916 9217 20944 9454
rect 20902 9208 20958 9217
rect 20902 9143 20958 9152
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 21008 8090 21036 8842
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19524 6384 19576 6390
rect 19524 6326 19576 6332
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19076 6174 19196 6202
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 19076 5846 19104 6054
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 19168 5710 19196 6174
rect 19156 5704 19208 5710
rect 19156 5646 19208 5652
rect 19260 5642 19288 6258
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19352 5914 19380 6190
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19628 5710 19656 6054
rect 19812 5710 19840 6326
rect 19996 5778 20024 7210
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 20272 5710 20300 7142
rect 20548 7002 20576 7346
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 21284 6882 21312 11494
rect 21376 11150 21404 12038
rect 21468 11694 21496 12242
rect 21560 11762 21588 13466
rect 21652 12986 21680 16050
rect 21803 15804 22111 15824
rect 21803 15802 21809 15804
rect 21865 15802 21889 15804
rect 21945 15802 21969 15804
rect 22025 15802 22049 15804
rect 22105 15802 22111 15804
rect 21865 15750 21867 15802
rect 22047 15750 22049 15802
rect 21803 15748 21809 15750
rect 21865 15748 21889 15750
rect 21945 15748 21969 15750
rect 22025 15748 22049 15750
rect 22105 15748 22111 15750
rect 21803 15728 22111 15748
rect 21803 14716 22111 14736
rect 21803 14714 21809 14716
rect 21865 14714 21889 14716
rect 21945 14714 21969 14716
rect 22025 14714 22049 14716
rect 22105 14714 22111 14716
rect 21865 14662 21867 14714
rect 22047 14662 22049 14714
rect 21803 14660 21809 14662
rect 21865 14660 21889 14662
rect 21945 14660 21969 14662
rect 22025 14660 22049 14662
rect 22105 14660 22111 14662
rect 21803 14640 22111 14660
rect 22204 13802 22232 16102
rect 22374 16079 22430 16088
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 21803 13628 22111 13648
rect 21803 13626 21809 13628
rect 21865 13626 21889 13628
rect 21945 13626 21969 13628
rect 22025 13626 22049 13628
rect 22105 13626 22111 13628
rect 21865 13574 21867 13626
rect 22047 13574 22049 13626
rect 21803 13572 21809 13574
rect 21865 13572 21889 13574
rect 21945 13572 21969 13574
rect 22025 13572 22049 13574
rect 22105 13572 22111 13574
rect 21803 13552 22111 13572
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21652 12866 21680 12922
rect 21652 12838 21772 12866
rect 21928 12850 21956 13262
rect 22008 13252 22060 13258
rect 22008 13194 22060 13200
rect 21640 12776 21692 12782
rect 21640 12718 21692 12724
rect 21652 12238 21680 12718
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21744 11830 21772 12838
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 22020 12782 22048 13194
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 21803 12540 22111 12560
rect 21803 12538 21809 12540
rect 21865 12538 21889 12540
rect 21945 12538 21969 12540
rect 22025 12538 22049 12540
rect 22105 12538 22111 12540
rect 21865 12486 21867 12538
rect 22047 12486 22049 12538
rect 21803 12484 21809 12486
rect 21865 12484 21889 12486
rect 21945 12484 21969 12486
rect 22025 12484 22049 12486
rect 22105 12484 22111 12486
rect 21803 12464 22111 12484
rect 22204 12356 22232 13738
rect 22388 12918 22416 16079
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22572 15570 22600 15982
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22664 15502 22692 15846
rect 22756 15706 22784 15982
rect 22940 15706 22968 16458
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 23032 16250 23060 16390
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23216 16046 23244 16594
rect 23664 16516 23716 16522
rect 23664 16458 23716 16464
rect 23204 16040 23256 16046
rect 23204 15982 23256 15988
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 23492 15570 23520 15982
rect 23676 15910 23704 16458
rect 23768 16454 23796 21830
rect 23860 21146 23888 21830
rect 23952 21146 23980 22578
rect 24400 22568 24452 22574
rect 24400 22510 24452 22516
rect 24032 21956 24084 21962
rect 24032 21898 24084 21904
rect 24044 21350 24072 21898
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24412 21146 24440 22510
rect 24688 22030 24716 22578
rect 24872 22234 24900 22714
rect 24860 22228 24912 22234
rect 24860 22170 24912 22176
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24688 21690 24716 21966
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 25056 21622 25084 21830
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 24400 21140 24452 21146
rect 24400 21082 24452 21088
rect 23860 20874 23888 21082
rect 24596 20942 24624 21286
rect 25044 21072 25096 21078
rect 25044 21014 25096 21020
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 23848 20868 23900 20874
rect 23848 20810 23900 20816
rect 24308 20460 24360 20466
rect 24308 20402 24360 20408
rect 24492 20460 24544 20466
rect 24492 20402 24544 20408
rect 24320 20330 24348 20402
rect 24308 20324 24360 20330
rect 24308 20266 24360 20272
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23860 19854 23888 20198
rect 24320 19990 24348 20266
rect 24308 19984 24360 19990
rect 24308 19926 24360 19932
rect 24504 19854 24532 20402
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24584 20256 24636 20262
rect 24584 20198 24636 20204
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 23860 19514 23888 19790
rect 23940 19780 23992 19786
rect 23940 19722 23992 19728
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 23952 18834 23980 19722
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 23940 18828 23992 18834
rect 23940 18770 23992 18776
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23860 16250 23888 18566
rect 24044 18222 24072 19246
rect 24228 18834 24256 19654
rect 24216 18828 24268 18834
rect 24216 18770 24268 18776
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24228 18426 24256 18566
rect 24216 18420 24268 18426
rect 24216 18362 24268 18368
rect 24596 18358 24624 20198
rect 24964 19854 24992 20334
rect 25056 19854 25084 21014
rect 25594 20768 25650 20777
rect 25594 20703 25650 20712
rect 25320 19984 25372 19990
rect 25320 19926 25372 19932
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 24964 19514 24992 19790
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 25240 18970 25268 19314
rect 25228 18964 25280 18970
rect 25228 18906 25280 18912
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 24584 18352 24636 18358
rect 24584 18294 24636 18300
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 23848 16244 23900 16250
rect 23848 16186 23900 16192
rect 24124 16176 24176 16182
rect 24124 16118 24176 16124
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23480 15564 23532 15570
rect 23480 15506 23532 15512
rect 23676 15502 23704 15846
rect 23768 15570 23796 15914
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23400 15162 23428 15302
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23768 15026 23796 15506
rect 24032 15496 24084 15502
rect 24032 15438 24084 15444
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23308 14550 23336 14962
rect 23676 14822 23704 14962
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23386 14648 23442 14657
rect 23386 14583 23442 14592
rect 23296 14544 23348 14550
rect 23296 14486 23348 14492
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 22468 13252 22520 13258
rect 22468 13194 22520 13200
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22480 12714 22508 13194
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22940 12918 22968 13126
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 22468 12708 22520 12714
rect 22468 12650 22520 12656
rect 22112 12328 22232 12356
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 21928 12170 21956 12242
rect 21916 12164 21968 12170
rect 21916 12106 21968 12112
rect 21928 11898 21956 12106
rect 22112 12102 22140 12328
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 22204 11694 22232 12038
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 21803 11452 22111 11472
rect 21803 11450 21809 11452
rect 21865 11450 21889 11452
rect 21945 11450 21969 11452
rect 22025 11450 22049 11452
rect 22105 11450 22111 11452
rect 21865 11398 21867 11450
rect 22047 11398 22049 11450
rect 21803 11396 21809 11398
rect 21865 11396 21889 11398
rect 21945 11396 21969 11398
rect 22025 11396 22049 11398
rect 22105 11396 22111 11398
rect 21803 11376 22111 11396
rect 22204 11354 22232 11630
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 22388 11286 22416 11630
rect 22480 11626 22508 12650
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22664 12434 22692 12582
rect 22572 12406 22692 12434
rect 22572 12238 22600 12406
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22848 12102 22876 12582
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22468 11620 22520 11626
rect 22468 11562 22520 11568
rect 22376 11280 22428 11286
rect 22376 11222 22428 11228
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 22836 11008 22888 11014
rect 22836 10950 22888 10956
rect 21803 10364 22111 10384
rect 21803 10362 21809 10364
rect 21865 10362 21889 10364
rect 21945 10362 21969 10364
rect 22025 10362 22049 10364
rect 22105 10362 22111 10364
rect 21865 10310 21867 10362
rect 22047 10310 22049 10362
rect 21803 10308 21809 10310
rect 21865 10308 21889 10310
rect 21945 10308 21969 10310
rect 22025 10308 22049 10310
rect 22105 10308 22111 10310
rect 21803 10288 22111 10308
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21468 9450 21496 10066
rect 22098 10024 22154 10033
rect 22098 9959 22100 9968
rect 22152 9959 22154 9968
rect 22652 9988 22704 9994
rect 22100 9930 22152 9936
rect 22652 9930 22704 9936
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 21732 9648 21784 9654
rect 21732 9590 21784 9596
rect 22192 9648 22244 9654
rect 22192 9590 22244 9596
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21376 9081 21404 9318
rect 21456 9172 21508 9178
rect 21560 9160 21588 9522
rect 21508 9132 21588 9160
rect 21456 9114 21508 9120
rect 21362 9072 21418 9081
rect 21362 9007 21418 9016
rect 21560 8634 21588 9132
rect 21744 8974 21772 9590
rect 21803 9276 22111 9296
rect 21803 9274 21809 9276
rect 21865 9274 21889 9276
rect 21945 9274 21969 9276
rect 22025 9274 22049 9276
rect 22105 9274 22111 9276
rect 21865 9222 21867 9274
rect 22047 9222 22049 9274
rect 21803 9220 21809 9222
rect 21865 9220 21889 9222
rect 21945 9220 21969 9222
rect 22025 9220 22049 9222
rect 22105 9220 22111 9222
rect 21803 9200 22111 9220
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21744 8566 21772 8910
rect 22020 8566 22048 8978
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 22204 8401 22232 9590
rect 22296 9110 22324 9862
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22664 8430 22692 9930
rect 22744 8900 22796 8906
rect 22744 8842 22796 8848
rect 22756 8498 22784 8842
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22652 8424 22704 8430
rect 22190 8392 22246 8401
rect 22652 8366 22704 8372
rect 22190 8327 22246 8336
rect 21803 8188 22111 8208
rect 21803 8186 21809 8188
rect 21865 8186 21889 8188
rect 21945 8186 21969 8188
rect 22025 8186 22049 8188
rect 22105 8186 22111 8188
rect 21865 8134 21867 8186
rect 22047 8134 22049 8186
rect 21803 8132 21809 8134
rect 21865 8132 21889 8134
rect 21945 8132 21969 8134
rect 22025 8132 22049 8134
rect 22105 8132 22111 8134
rect 21803 8112 22111 8132
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 21192 6854 21312 6882
rect 20364 6458 20392 6802
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20824 6458 20852 6598
rect 21192 6458 21220 6854
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21284 6390 21312 6734
rect 21272 6384 21324 6390
rect 21272 6326 21324 6332
rect 21284 5914 21312 6326
rect 21376 6254 21404 7278
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 21803 7100 22111 7120
rect 21803 7098 21809 7100
rect 21865 7098 21889 7100
rect 21945 7098 21969 7100
rect 22025 7098 22049 7100
rect 22105 7098 22111 7100
rect 21865 7046 21867 7098
rect 22047 7046 22049 7098
rect 21803 7044 21809 7046
rect 21865 7044 21889 7046
rect 21945 7044 21969 7046
rect 22025 7044 22049 7046
rect 22105 7044 22111 7046
rect 21803 7024 22111 7044
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21468 6322 21496 6734
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21560 6390 21588 6666
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19260 5030 19288 5578
rect 19812 5370 19840 5646
rect 19800 5364 19852 5370
rect 19800 5306 19852 5312
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 21652 3398 21680 6870
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22112 6100 22140 6258
rect 22112 6072 22232 6100
rect 21803 6012 22111 6032
rect 21803 6010 21809 6012
rect 21865 6010 21889 6012
rect 21945 6010 21969 6012
rect 22025 6010 22049 6012
rect 22105 6010 22111 6012
rect 21865 5958 21867 6010
rect 22047 5958 22049 6010
rect 21803 5956 21809 5958
rect 21865 5956 21889 5958
rect 21945 5956 21969 5958
rect 22025 5956 22049 5958
rect 22105 5956 22111 5958
rect 21803 5936 22111 5956
rect 22204 5914 22232 6072
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 22296 5846 22324 7142
rect 22572 6934 22600 7142
rect 22560 6928 22612 6934
rect 22560 6870 22612 6876
rect 22756 6866 22784 8434
rect 22848 7546 22876 10950
rect 23032 9602 23060 14418
rect 23204 14272 23256 14278
rect 23204 14214 23256 14220
rect 23216 13938 23244 14214
rect 23308 14074 23336 14486
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 23400 13462 23428 14583
rect 23676 14482 23704 14758
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23584 13938 23612 14350
rect 23756 14340 23808 14346
rect 23756 14282 23808 14288
rect 23664 14000 23716 14006
rect 23664 13942 23716 13948
rect 23572 13932 23624 13938
rect 23492 13892 23572 13920
rect 23388 13456 23440 13462
rect 23388 13398 23440 13404
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 23216 11150 23244 11494
rect 23296 11280 23348 11286
rect 23296 11222 23348 11228
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23112 10192 23164 10198
rect 23112 10134 23164 10140
rect 23124 9722 23152 10134
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23112 9716 23164 9722
rect 23112 9658 23164 9664
rect 23032 9574 23152 9602
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 22940 8974 22968 9318
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22940 8566 22968 8910
rect 22928 8560 22980 8566
rect 22928 8502 22980 8508
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22376 6724 22428 6730
rect 22376 6666 22428 6672
rect 22284 5840 22336 5846
rect 22284 5782 22336 5788
rect 22388 5778 22416 6666
rect 22756 6322 22784 6802
rect 23032 6798 23060 7686
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 22744 6316 22796 6322
rect 22744 6258 22796 6264
rect 22376 5772 22428 5778
rect 22376 5714 22428 5720
rect 21803 4924 22111 4944
rect 21803 4922 21809 4924
rect 21865 4922 21889 4924
rect 21945 4922 21969 4924
rect 22025 4922 22049 4924
rect 22105 4922 22111 4924
rect 21865 4870 21867 4922
rect 22047 4870 22049 4922
rect 21803 4868 21809 4870
rect 21865 4868 21889 4870
rect 21945 4868 21969 4870
rect 22025 4868 22049 4870
rect 22105 4868 22111 4870
rect 21803 4848 22111 4868
rect 22756 4214 22784 6258
rect 22744 4208 22796 4214
rect 22744 4150 22796 4156
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 21803 3836 22111 3856
rect 21803 3834 21809 3836
rect 21865 3834 21889 3836
rect 21945 3834 21969 3836
rect 22025 3834 22049 3836
rect 22105 3834 22111 3836
rect 21865 3782 21867 3834
rect 22047 3782 22049 3834
rect 21803 3780 21809 3782
rect 21865 3780 21889 3782
rect 21945 3780 21969 3782
rect 22025 3780 22049 3782
rect 22105 3780 22111 3782
rect 21803 3760 22111 3780
rect 22296 3738 22324 4082
rect 23124 4010 23152 9574
rect 23216 8974 23244 9862
rect 23308 9518 23336 11222
rect 23492 10810 23520 13892
rect 23572 13874 23624 13880
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 23584 12442 23612 13670
rect 23676 13530 23704 13942
rect 23768 13870 23796 14282
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23676 13326 23704 13466
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 23584 11898 23612 12378
rect 23676 12306 23704 13262
rect 23768 13190 23796 13806
rect 23860 13394 23888 13874
rect 23940 13796 23992 13802
rect 23940 13738 23992 13744
rect 23952 13394 23980 13738
rect 24044 13734 24072 15438
rect 24136 15026 24164 16118
rect 24228 15706 24256 17138
rect 24492 16992 24544 16998
rect 24492 16934 24544 16940
rect 24504 16658 24532 16934
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24320 15706 24348 16050
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 24596 15502 24624 16390
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24216 15428 24268 15434
rect 24216 15370 24268 15376
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 24136 13530 24164 14962
rect 24228 14482 24256 15370
rect 24216 14476 24268 14482
rect 24216 14418 24268 14424
rect 24308 14408 24360 14414
rect 24308 14350 24360 14356
rect 24320 13938 24348 14350
rect 24596 14074 24624 15438
rect 24688 15366 24716 16594
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24872 16250 24900 16390
rect 24964 16250 24992 16458
rect 25148 16454 25176 18634
rect 25332 18426 25360 19926
rect 25412 19440 25464 19446
rect 25412 19382 25464 19388
rect 25424 18766 25452 19382
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25320 18420 25372 18426
rect 25320 18362 25372 18368
rect 25412 17060 25464 17066
rect 25412 17002 25464 17008
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25424 16250 25452 17002
rect 25608 16794 25636 20703
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 25504 16040 25556 16046
rect 25504 15982 25556 15988
rect 25240 15706 25268 15982
rect 25228 15700 25280 15706
rect 25228 15642 25280 15648
rect 25516 15638 25544 15982
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 25504 15632 25556 15638
rect 25504 15574 25556 15580
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24688 14278 24716 15302
rect 24780 15094 24808 15574
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25424 15162 25452 15438
rect 25412 15156 25464 15162
rect 25412 15098 25464 15104
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24584 14068 24636 14074
rect 24584 14010 24636 14016
rect 24308 13932 24360 13938
rect 24308 13874 24360 13880
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23940 13388 23992 13394
rect 23940 13330 23992 13336
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23860 12850 23888 13330
rect 24136 12986 24164 13466
rect 24320 13258 24348 13874
rect 24308 13252 24360 13258
rect 24308 13194 24360 13200
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 24136 12850 24164 12922
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 24124 12708 24176 12714
rect 24124 12650 24176 12656
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23664 12300 23716 12306
rect 23664 12242 23716 12248
rect 23664 12096 23716 12102
rect 23664 12038 23716 12044
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23584 11150 23612 11834
rect 23676 11694 23704 12038
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23676 10742 23704 11630
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 23480 9580 23532 9586
rect 23480 9522 23532 9528
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23400 9042 23428 9454
rect 23492 9178 23520 9522
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23308 6662 23336 7822
rect 23400 7274 23428 8978
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23492 8430 23520 8774
rect 23676 8498 23704 9454
rect 23768 8974 23796 12582
rect 24136 12374 24164 12650
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 24136 12102 24164 12310
rect 24596 12238 24624 14010
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24124 12096 24176 12102
rect 24124 12038 24176 12044
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24412 11898 24440 12038
rect 24400 11892 24452 11898
rect 24400 11834 24452 11840
rect 24596 11830 24624 12174
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24308 11688 24360 11694
rect 24308 11630 24360 11636
rect 23848 11552 23900 11558
rect 23848 11494 23900 11500
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 23676 7886 23704 8230
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23860 7546 23888 11494
rect 24320 11218 24348 11630
rect 24688 11218 24716 14214
rect 24308 11212 24360 11218
rect 24308 11154 24360 11160
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 24688 10742 24716 11154
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24780 10810 24808 10950
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24676 10736 24728 10742
rect 24676 10678 24728 10684
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 25596 10056 25648 10062
rect 25596 9998 25648 10004
rect 24400 9988 24452 9994
rect 24400 9930 24452 9936
rect 24412 9654 24440 9930
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 24596 9382 24624 9998
rect 24964 9722 24992 9998
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 25608 9586 25636 9998
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23952 8090 23980 8434
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 23388 7268 23440 7274
rect 23388 7210 23440 7216
rect 23768 7002 23796 7278
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 24136 6458 24164 7346
rect 24320 6914 24348 7346
rect 24320 6886 24440 6914
rect 24412 6798 24440 6886
rect 24504 6866 24532 7346
rect 24872 7206 24900 8910
rect 25240 8634 25268 8910
rect 25608 8906 25636 9522
rect 25596 8900 25648 8906
rect 25596 8842 25648 8848
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 24872 6934 24900 7142
rect 24860 6928 24912 6934
rect 24860 6870 24912 6876
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24400 6792 24452 6798
rect 24400 6734 24452 6740
rect 24124 6452 24176 6458
rect 24124 6394 24176 6400
rect 24412 6322 24440 6734
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 23308 5710 23336 6054
rect 23584 5710 23612 6054
rect 23676 5846 23704 6258
rect 23664 5840 23716 5846
rect 23664 5782 23716 5788
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23112 4004 23164 4010
rect 23112 3946 23164 3952
rect 22374 3768 22430 3777
rect 22284 3732 22336 3738
rect 22374 3703 22430 3712
rect 22284 3674 22336 3680
rect 21732 3460 21784 3466
rect 21732 3402 21784 3408
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 18708 2746 19012 2774
rect 17632 2204 17940 2224
rect 17632 2202 17638 2204
rect 17694 2202 17718 2204
rect 17774 2202 17798 2204
rect 17854 2202 17878 2204
rect 17934 2202 17940 2204
rect 17694 2150 17696 2202
rect 17876 2150 17878 2202
rect 17632 2148 17638 2150
rect 17694 2148 17718 2150
rect 17774 2148 17798 2150
rect 17854 2148 17878 2150
rect 17934 2148 17940 2150
rect 17632 2128 17940 2148
rect 18340 870 18460 898
rect 18340 800 18368 870
rect 13096 734 13584 762
rect 13634 0 13690 800
rect 14738 0 14794 800
rect 15934 0 15990 800
rect 17130 0 17186 800
rect 18326 0 18382 800
rect 18432 762 18460 870
rect 18708 762 18736 2746
rect 19536 800 19564 2926
rect 21744 1714 21772 3402
rect 22388 3194 22416 3703
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22376 3188 22428 3194
rect 22376 3130 22428 3136
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 21803 2748 22111 2768
rect 21803 2746 21809 2748
rect 21865 2746 21889 2748
rect 21945 2746 21969 2748
rect 22025 2746 22049 2748
rect 22105 2746 22111 2748
rect 21865 2694 21867 2746
rect 22047 2694 22049 2746
rect 21803 2692 21809 2694
rect 21865 2692 21889 2694
rect 21945 2692 21969 2694
rect 22025 2692 22049 2694
rect 22105 2692 22111 2694
rect 21803 2672 22111 2692
rect 22204 2281 22232 3062
rect 22190 2272 22246 2281
rect 22190 2207 22246 2216
rect 21744 1686 21956 1714
rect 21928 800 21956 1686
rect 18432 734 18736 762
rect 19522 0 19578 800
rect 20718 0 20774 800
rect 21914 0 21970 800
rect 22664 785 22692 3334
rect 23124 800 23152 3470
rect 24320 800 24348 3470
rect 25516 800 25544 3470
rect 22650 776 22706 785
rect 22650 711 22706 720
rect 23110 0 23166 800
rect 24306 0 24362 800
rect 25502 0 25558 800
rect 26698 0 26754 800
<< via2 >>
rect 2134 24404 2190 24440
rect 2134 24384 2136 24404
rect 2136 24384 2188 24404
rect 2188 24384 2190 24404
rect 2134 23060 2136 23080
rect 2136 23060 2188 23080
rect 2188 23060 2190 23080
rect 2134 23024 2190 23060
rect 5126 26682 5182 26684
rect 5206 26682 5262 26684
rect 5286 26682 5342 26684
rect 5366 26682 5422 26684
rect 5126 26630 5172 26682
rect 5172 26630 5182 26682
rect 5206 26630 5236 26682
rect 5236 26630 5248 26682
rect 5248 26630 5262 26682
rect 5286 26630 5300 26682
rect 5300 26630 5312 26682
rect 5312 26630 5342 26682
rect 5366 26630 5376 26682
rect 5376 26630 5422 26682
rect 5126 26628 5182 26630
rect 5206 26628 5262 26630
rect 5286 26628 5342 26630
rect 5366 26628 5422 26630
rect 5126 25594 5182 25596
rect 5206 25594 5262 25596
rect 5286 25594 5342 25596
rect 5366 25594 5422 25596
rect 5126 25542 5172 25594
rect 5172 25542 5182 25594
rect 5206 25542 5236 25594
rect 5236 25542 5248 25594
rect 5248 25542 5262 25594
rect 5286 25542 5300 25594
rect 5300 25542 5312 25594
rect 5312 25542 5342 25594
rect 5366 25542 5376 25594
rect 5376 25542 5422 25594
rect 5126 25540 5182 25542
rect 5206 25540 5262 25542
rect 5286 25540 5342 25542
rect 5366 25540 5422 25542
rect 5126 24506 5182 24508
rect 5206 24506 5262 24508
rect 5286 24506 5342 24508
rect 5366 24506 5422 24508
rect 5126 24454 5172 24506
rect 5172 24454 5182 24506
rect 5206 24454 5236 24506
rect 5236 24454 5248 24506
rect 5248 24454 5262 24506
rect 5286 24454 5300 24506
rect 5300 24454 5312 24506
rect 5312 24454 5342 24506
rect 5366 24454 5376 24506
rect 5376 24454 5422 24506
rect 5126 24452 5182 24454
rect 5206 24452 5262 24454
rect 5286 24452 5342 24454
rect 5366 24452 5422 24454
rect 5126 23418 5182 23420
rect 5206 23418 5262 23420
rect 5286 23418 5342 23420
rect 5366 23418 5422 23420
rect 5126 23366 5172 23418
rect 5172 23366 5182 23418
rect 5206 23366 5236 23418
rect 5236 23366 5248 23418
rect 5248 23366 5262 23418
rect 5286 23366 5300 23418
rect 5300 23366 5312 23418
rect 5312 23366 5342 23418
rect 5366 23366 5376 23418
rect 5376 23366 5422 23418
rect 5126 23364 5182 23366
rect 5206 23364 5262 23366
rect 5286 23364 5342 23366
rect 5366 23364 5422 23366
rect 5126 22330 5182 22332
rect 5206 22330 5262 22332
rect 5286 22330 5342 22332
rect 5366 22330 5422 22332
rect 5126 22278 5172 22330
rect 5172 22278 5182 22330
rect 5206 22278 5236 22330
rect 5236 22278 5248 22330
rect 5248 22278 5262 22330
rect 5286 22278 5300 22330
rect 5300 22278 5312 22330
rect 5312 22278 5342 22330
rect 5366 22278 5376 22330
rect 5376 22278 5422 22330
rect 5126 22276 5182 22278
rect 5206 22276 5262 22278
rect 5286 22276 5342 22278
rect 5366 22276 5422 22278
rect 3422 14592 3478 14648
rect 4066 17448 4122 17504
rect 9297 27226 9353 27228
rect 9377 27226 9433 27228
rect 9457 27226 9513 27228
rect 9537 27226 9593 27228
rect 9297 27174 9343 27226
rect 9343 27174 9353 27226
rect 9377 27174 9407 27226
rect 9407 27174 9419 27226
rect 9419 27174 9433 27226
rect 9457 27174 9471 27226
rect 9471 27174 9483 27226
rect 9483 27174 9513 27226
rect 9537 27174 9547 27226
rect 9547 27174 9593 27226
rect 9297 27172 9353 27174
rect 9377 27172 9433 27174
rect 9457 27172 9513 27174
rect 9537 27172 9593 27174
rect 9297 26138 9353 26140
rect 9377 26138 9433 26140
rect 9457 26138 9513 26140
rect 9537 26138 9593 26140
rect 9297 26086 9343 26138
rect 9343 26086 9353 26138
rect 9377 26086 9407 26138
rect 9407 26086 9419 26138
rect 9419 26086 9433 26138
rect 9457 26086 9471 26138
rect 9471 26086 9483 26138
rect 9483 26086 9513 26138
rect 9537 26086 9547 26138
rect 9547 26086 9593 26138
rect 9297 26084 9353 26086
rect 9377 26084 9433 26086
rect 9457 26084 9513 26086
rect 9537 26084 9593 26086
rect 5998 21664 6054 21720
rect 5126 21242 5182 21244
rect 5206 21242 5262 21244
rect 5286 21242 5342 21244
rect 5366 21242 5422 21244
rect 5126 21190 5172 21242
rect 5172 21190 5182 21242
rect 5206 21190 5236 21242
rect 5236 21190 5248 21242
rect 5248 21190 5262 21242
rect 5286 21190 5300 21242
rect 5300 21190 5312 21242
rect 5312 21190 5342 21242
rect 5366 21190 5376 21242
rect 5376 21190 5422 21242
rect 5126 21188 5182 21190
rect 5206 21188 5262 21190
rect 5286 21188 5342 21190
rect 5366 21188 5422 21190
rect 5126 20154 5182 20156
rect 5206 20154 5262 20156
rect 5286 20154 5342 20156
rect 5366 20154 5422 20156
rect 5126 20102 5172 20154
rect 5172 20102 5182 20154
rect 5206 20102 5236 20154
rect 5236 20102 5248 20154
rect 5248 20102 5262 20154
rect 5286 20102 5300 20154
rect 5300 20102 5312 20154
rect 5312 20102 5342 20154
rect 5366 20102 5376 20154
rect 5376 20102 5422 20154
rect 5126 20100 5182 20102
rect 5206 20100 5262 20102
rect 5286 20100 5342 20102
rect 5366 20100 5422 20102
rect 5126 19066 5182 19068
rect 5206 19066 5262 19068
rect 5286 19066 5342 19068
rect 5366 19066 5422 19068
rect 5126 19014 5172 19066
rect 5172 19014 5182 19066
rect 5206 19014 5236 19066
rect 5236 19014 5248 19066
rect 5248 19014 5262 19066
rect 5286 19014 5300 19066
rect 5300 19014 5312 19066
rect 5312 19014 5342 19066
rect 5366 19014 5376 19066
rect 5376 19014 5422 19066
rect 5126 19012 5182 19014
rect 5206 19012 5262 19014
rect 5286 19012 5342 19014
rect 5366 19012 5422 19014
rect 5126 17978 5182 17980
rect 5206 17978 5262 17980
rect 5286 17978 5342 17980
rect 5366 17978 5422 17980
rect 5126 17926 5172 17978
rect 5172 17926 5182 17978
rect 5206 17926 5236 17978
rect 5236 17926 5248 17978
rect 5248 17926 5262 17978
rect 5286 17926 5300 17978
rect 5300 17926 5312 17978
rect 5312 17926 5342 17978
rect 5366 17926 5376 17978
rect 5376 17926 5422 17978
rect 5126 17924 5182 17926
rect 5206 17924 5262 17926
rect 5286 17924 5342 17926
rect 5366 17924 5422 17926
rect 4066 16088 4122 16144
rect 3054 9696 3110 9752
rect 2042 3440 2098 3496
rect 2778 2080 2834 2136
rect 3974 9036 4030 9072
rect 3974 9016 3976 9036
rect 3976 9016 4028 9036
rect 4028 9016 4030 9036
rect 5126 16890 5182 16892
rect 5206 16890 5262 16892
rect 5286 16890 5342 16892
rect 5366 16890 5422 16892
rect 5126 16838 5172 16890
rect 5172 16838 5182 16890
rect 5206 16838 5236 16890
rect 5236 16838 5248 16890
rect 5248 16838 5262 16890
rect 5286 16838 5300 16890
rect 5300 16838 5312 16890
rect 5312 16838 5342 16890
rect 5366 16838 5376 16890
rect 5376 16838 5422 16890
rect 5126 16836 5182 16838
rect 5206 16836 5262 16838
rect 5286 16836 5342 16838
rect 5366 16836 5422 16838
rect 5126 15802 5182 15804
rect 5206 15802 5262 15804
rect 5286 15802 5342 15804
rect 5366 15802 5422 15804
rect 5126 15750 5172 15802
rect 5172 15750 5182 15802
rect 5206 15750 5236 15802
rect 5236 15750 5248 15802
rect 5248 15750 5262 15802
rect 5286 15750 5300 15802
rect 5300 15750 5312 15802
rect 5312 15750 5342 15802
rect 5366 15750 5376 15802
rect 5376 15750 5422 15802
rect 5126 15748 5182 15750
rect 5206 15748 5262 15750
rect 5286 15748 5342 15750
rect 5366 15748 5422 15750
rect 4526 13812 4528 13832
rect 4528 13812 4580 13832
rect 4580 13812 4582 13832
rect 4526 13776 4582 13812
rect 5126 14714 5182 14716
rect 5206 14714 5262 14716
rect 5286 14714 5342 14716
rect 5366 14714 5422 14716
rect 5126 14662 5172 14714
rect 5172 14662 5182 14714
rect 5206 14662 5236 14714
rect 5236 14662 5248 14714
rect 5248 14662 5262 14714
rect 5286 14662 5300 14714
rect 5300 14662 5312 14714
rect 5312 14662 5342 14714
rect 5366 14662 5376 14714
rect 5376 14662 5422 14714
rect 5126 14660 5182 14662
rect 5206 14660 5262 14662
rect 5286 14660 5342 14662
rect 5366 14660 5422 14662
rect 5906 14476 5962 14512
rect 5906 14456 5908 14476
rect 5908 14456 5960 14476
rect 5960 14456 5962 14476
rect 4710 13932 4766 13968
rect 5722 13958 5778 13968
rect 4710 13912 4712 13932
rect 4712 13912 4764 13932
rect 4764 13912 4766 13932
rect 5722 13912 5724 13958
rect 5724 13912 5776 13958
rect 5776 13912 5778 13958
rect 5126 13626 5182 13628
rect 5206 13626 5262 13628
rect 5286 13626 5342 13628
rect 5366 13626 5422 13628
rect 5126 13574 5172 13626
rect 5172 13574 5182 13626
rect 5206 13574 5236 13626
rect 5236 13574 5248 13626
rect 5248 13574 5262 13626
rect 5286 13574 5300 13626
rect 5300 13574 5312 13626
rect 5312 13574 5342 13626
rect 5366 13574 5376 13626
rect 5376 13574 5422 13626
rect 5126 13572 5182 13574
rect 5206 13572 5262 13574
rect 5286 13572 5342 13574
rect 5366 13572 5422 13574
rect 5446 13368 5502 13424
rect 5814 13368 5870 13424
rect 6734 14476 6790 14512
rect 6734 14456 6736 14476
rect 6736 14456 6788 14476
rect 6788 14456 6790 14476
rect 6642 13368 6698 13424
rect 8022 23724 8078 23760
rect 8022 23704 8024 23724
rect 8024 23704 8076 23724
rect 8076 23704 8078 23724
rect 6918 13812 6920 13832
rect 6920 13812 6972 13832
rect 6972 13812 6974 13832
rect 6918 13776 6974 13812
rect 5126 12538 5182 12540
rect 5206 12538 5262 12540
rect 5286 12538 5342 12540
rect 5366 12538 5422 12540
rect 5126 12486 5172 12538
rect 5172 12486 5182 12538
rect 5206 12486 5236 12538
rect 5236 12486 5248 12538
rect 5248 12486 5262 12538
rect 5286 12486 5300 12538
rect 5300 12486 5312 12538
rect 5312 12486 5342 12538
rect 5366 12486 5376 12538
rect 5376 12486 5422 12538
rect 5126 12484 5182 12486
rect 5206 12484 5262 12486
rect 5286 12484 5342 12486
rect 5366 12484 5422 12486
rect 5126 11450 5182 11452
rect 5206 11450 5262 11452
rect 5286 11450 5342 11452
rect 5366 11450 5422 11452
rect 5126 11398 5172 11450
rect 5172 11398 5182 11450
rect 5206 11398 5236 11450
rect 5236 11398 5248 11450
rect 5248 11398 5262 11450
rect 5286 11398 5300 11450
rect 5300 11398 5312 11450
rect 5312 11398 5342 11450
rect 5366 11398 5376 11450
rect 5376 11398 5422 11450
rect 5126 11396 5182 11398
rect 5206 11396 5262 11398
rect 5286 11396 5342 11398
rect 5366 11396 5422 11398
rect 5446 11192 5502 11248
rect 4986 10684 4988 10704
rect 4988 10684 5040 10704
rect 5040 10684 5042 10704
rect 4986 10648 5042 10684
rect 5998 10648 6054 10704
rect 5126 10362 5182 10364
rect 5206 10362 5262 10364
rect 5286 10362 5342 10364
rect 5366 10362 5422 10364
rect 5126 10310 5172 10362
rect 5172 10310 5182 10362
rect 5206 10310 5236 10362
rect 5236 10310 5248 10362
rect 5248 10310 5262 10362
rect 5286 10310 5300 10362
rect 5300 10310 5312 10362
rect 5312 10310 5342 10362
rect 5366 10310 5376 10362
rect 5376 10310 5422 10362
rect 5126 10308 5182 10310
rect 5206 10308 5262 10310
rect 5286 10308 5342 10310
rect 5366 10308 5422 10310
rect 3514 4800 3570 4856
rect 4066 6332 4068 6352
rect 4068 6332 4120 6352
rect 4120 6332 4122 6352
rect 4066 6296 4122 6332
rect 5126 9274 5182 9276
rect 5206 9274 5262 9276
rect 5286 9274 5342 9276
rect 5366 9274 5422 9276
rect 5126 9222 5172 9274
rect 5172 9222 5182 9274
rect 5206 9222 5236 9274
rect 5236 9222 5248 9274
rect 5248 9222 5262 9274
rect 5286 9222 5300 9274
rect 5300 9222 5312 9274
rect 5312 9222 5342 9274
rect 5366 9222 5376 9274
rect 5376 9222 5422 9274
rect 5126 9220 5182 9222
rect 5206 9220 5262 9222
rect 5286 9220 5342 9222
rect 5366 9220 5422 9222
rect 5126 8186 5182 8188
rect 5206 8186 5262 8188
rect 5286 8186 5342 8188
rect 5366 8186 5422 8188
rect 5126 8134 5172 8186
rect 5172 8134 5182 8186
rect 5206 8134 5236 8186
rect 5236 8134 5248 8186
rect 5248 8134 5262 8186
rect 5286 8134 5300 8186
rect 5300 8134 5312 8186
rect 5312 8134 5342 8186
rect 5366 8134 5376 8186
rect 5376 8134 5422 8186
rect 5126 8132 5182 8134
rect 5206 8132 5262 8134
rect 5286 8132 5342 8134
rect 5366 8132 5422 8134
rect 5126 7098 5182 7100
rect 5206 7098 5262 7100
rect 5286 7098 5342 7100
rect 5366 7098 5422 7100
rect 5126 7046 5172 7098
rect 5172 7046 5182 7098
rect 5206 7046 5236 7098
rect 5236 7046 5248 7098
rect 5248 7046 5262 7098
rect 5286 7046 5300 7098
rect 5300 7046 5312 7098
rect 5312 7046 5342 7098
rect 5366 7046 5376 7098
rect 5376 7046 5422 7098
rect 5126 7044 5182 7046
rect 5206 7044 5262 7046
rect 5286 7044 5342 7046
rect 5366 7044 5422 7046
rect 5126 6010 5182 6012
rect 5206 6010 5262 6012
rect 5286 6010 5342 6012
rect 5366 6010 5422 6012
rect 5126 5958 5172 6010
rect 5172 5958 5182 6010
rect 5206 5958 5236 6010
rect 5236 5958 5248 6010
rect 5248 5958 5262 6010
rect 5286 5958 5300 6010
rect 5300 5958 5312 6010
rect 5312 5958 5342 6010
rect 5366 5958 5376 6010
rect 5376 5958 5422 6010
rect 5126 5956 5182 5958
rect 5206 5956 5262 5958
rect 5286 5956 5342 5958
rect 5366 5956 5422 5958
rect 5126 4922 5182 4924
rect 5206 4922 5262 4924
rect 5286 4922 5342 4924
rect 5366 4922 5422 4924
rect 5126 4870 5172 4922
rect 5172 4870 5182 4922
rect 5206 4870 5236 4922
rect 5236 4870 5248 4922
rect 5248 4870 5262 4922
rect 5286 4870 5300 4922
rect 5300 4870 5312 4922
rect 5312 4870 5342 4922
rect 5366 4870 5376 4922
rect 5376 4870 5422 4922
rect 5126 4868 5182 4870
rect 5206 4868 5262 4870
rect 5286 4868 5342 4870
rect 5366 4868 5422 4870
rect 5126 3834 5182 3836
rect 5206 3834 5262 3836
rect 5286 3834 5342 3836
rect 5366 3834 5422 3836
rect 5126 3782 5172 3834
rect 5172 3782 5182 3834
rect 5206 3782 5236 3834
rect 5236 3782 5248 3834
rect 5248 3782 5262 3834
rect 5286 3782 5300 3834
rect 5300 3782 5312 3834
rect 5312 3782 5342 3834
rect 5366 3782 5376 3834
rect 5376 3782 5422 3834
rect 5126 3780 5182 3782
rect 5206 3780 5262 3782
rect 5286 3780 5342 3782
rect 5366 3780 5422 3782
rect 5126 2746 5182 2748
rect 5206 2746 5262 2748
rect 5286 2746 5342 2748
rect 5366 2746 5422 2748
rect 5126 2694 5172 2746
rect 5172 2694 5182 2746
rect 5206 2694 5236 2746
rect 5236 2694 5248 2746
rect 5248 2694 5262 2746
rect 5286 2694 5300 2746
rect 5300 2694 5312 2746
rect 5312 2694 5342 2746
rect 5366 2694 5376 2746
rect 5376 2694 5422 2746
rect 5126 2692 5182 2694
rect 5206 2692 5262 2694
rect 5286 2692 5342 2694
rect 5366 2692 5422 2694
rect 3146 720 3202 776
rect 6918 10512 6974 10568
rect 7102 13368 7158 13424
rect 8298 23704 8354 23760
rect 8666 23724 8722 23760
rect 8666 23704 8668 23724
rect 8668 23704 8720 23724
rect 8720 23704 8722 23724
rect 9297 25050 9353 25052
rect 9377 25050 9433 25052
rect 9457 25050 9513 25052
rect 9537 25050 9593 25052
rect 9297 24998 9343 25050
rect 9343 24998 9353 25050
rect 9377 24998 9407 25050
rect 9407 24998 9419 25050
rect 9419 24998 9433 25050
rect 9457 24998 9471 25050
rect 9471 24998 9483 25050
rect 9483 24998 9513 25050
rect 9537 24998 9547 25050
rect 9547 24998 9593 25050
rect 9297 24996 9353 24998
rect 9377 24996 9433 24998
rect 9457 24996 9513 24998
rect 9537 24996 9593 24998
rect 9297 23962 9353 23964
rect 9377 23962 9433 23964
rect 9457 23962 9513 23964
rect 9537 23962 9593 23964
rect 9297 23910 9343 23962
rect 9343 23910 9353 23962
rect 9377 23910 9407 23962
rect 9407 23910 9419 23962
rect 9419 23910 9433 23962
rect 9457 23910 9471 23962
rect 9471 23910 9483 23962
rect 9483 23910 9513 23962
rect 9537 23910 9547 23962
rect 9547 23910 9593 23962
rect 9297 23908 9353 23910
rect 9377 23908 9433 23910
rect 9457 23908 9513 23910
rect 9537 23908 9593 23910
rect 9297 22874 9353 22876
rect 9377 22874 9433 22876
rect 9457 22874 9513 22876
rect 9537 22874 9593 22876
rect 9297 22822 9343 22874
rect 9343 22822 9353 22874
rect 9377 22822 9407 22874
rect 9407 22822 9419 22874
rect 9419 22822 9433 22874
rect 9457 22822 9471 22874
rect 9471 22822 9483 22874
rect 9483 22822 9513 22874
rect 9537 22822 9547 22874
rect 9547 22822 9593 22874
rect 9297 22820 9353 22822
rect 9377 22820 9433 22822
rect 9457 22820 9513 22822
rect 9537 22820 9593 22822
rect 9297 21786 9353 21788
rect 9377 21786 9433 21788
rect 9457 21786 9513 21788
rect 9537 21786 9593 21788
rect 9297 21734 9343 21786
rect 9343 21734 9353 21786
rect 9377 21734 9407 21786
rect 9407 21734 9419 21786
rect 9419 21734 9433 21786
rect 9457 21734 9471 21786
rect 9471 21734 9483 21786
rect 9483 21734 9513 21786
rect 9537 21734 9547 21786
rect 9547 21734 9593 21786
rect 9297 21732 9353 21734
rect 9377 21732 9433 21734
rect 9457 21732 9513 21734
rect 9537 21732 9593 21734
rect 9297 20698 9353 20700
rect 9377 20698 9433 20700
rect 9457 20698 9513 20700
rect 9537 20698 9593 20700
rect 9297 20646 9343 20698
rect 9343 20646 9353 20698
rect 9377 20646 9407 20698
rect 9407 20646 9419 20698
rect 9419 20646 9433 20698
rect 9457 20646 9471 20698
rect 9471 20646 9483 20698
rect 9483 20646 9513 20698
rect 9537 20646 9547 20698
rect 9547 20646 9593 20698
rect 9297 20644 9353 20646
rect 9377 20644 9433 20646
rect 9457 20644 9513 20646
rect 9537 20644 9593 20646
rect 11794 21936 11850 21992
rect 11150 20304 11206 20360
rect 9297 19610 9353 19612
rect 9377 19610 9433 19612
rect 9457 19610 9513 19612
rect 9537 19610 9593 19612
rect 9297 19558 9343 19610
rect 9343 19558 9353 19610
rect 9377 19558 9407 19610
rect 9407 19558 9419 19610
rect 9419 19558 9433 19610
rect 9457 19558 9471 19610
rect 9471 19558 9483 19610
rect 9483 19558 9513 19610
rect 9537 19558 9547 19610
rect 9547 19558 9593 19610
rect 9297 19556 9353 19558
rect 9377 19556 9433 19558
rect 9457 19556 9513 19558
rect 9537 19556 9593 19558
rect 9297 18522 9353 18524
rect 9377 18522 9433 18524
rect 9457 18522 9513 18524
rect 9537 18522 9593 18524
rect 9297 18470 9343 18522
rect 9343 18470 9353 18522
rect 9377 18470 9407 18522
rect 9407 18470 9419 18522
rect 9419 18470 9433 18522
rect 9457 18470 9471 18522
rect 9471 18470 9483 18522
rect 9483 18470 9513 18522
rect 9537 18470 9547 18522
rect 9547 18470 9593 18522
rect 9297 18468 9353 18470
rect 9377 18468 9433 18470
rect 9457 18468 9513 18470
rect 9537 18468 9593 18470
rect 9297 17434 9353 17436
rect 9377 17434 9433 17436
rect 9457 17434 9513 17436
rect 9537 17434 9593 17436
rect 9297 17382 9343 17434
rect 9343 17382 9353 17434
rect 9377 17382 9407 17434
rect 9407 17382 9419 17434
rect 9419 17382 9433 17434
rect 9457 17382 9471 17434
rect 9471 17382 9483 17434
rect 9483 17382 9513 17434
rect 9537 17382 9547 17434
rect 9547 17382 9593 17434
rect 9297 17380 9353 17382
rect 9377 17380 9433 17382
rect 9457 17380 9513 17382
rect 9537 17380 9593 17382
rect 11242 19352 11298 19408
rect 11518 19760 11574 19816
rect 9297 16346 9353 16348
rect 9377 16346 9433 16348
rect 9457 16346 9513 16348
rect 9537 16346 9593 16348
rect 9297 16294 9343 16346
rect 9343 16294 9353 16346
rect 9377 16294 9407 16346
rect 9407 16294 9419 16346
rect 9419 16294 9433 16346
rect 9457 16294 9471 16346
rect 9471 16294 9483 16346
rect 9483 16294 9513 16346
rect 9537 16294 9547 16346
rect 9547 16294 9593 16346
rect 9297 16292 9353 16294
rect 9377 16292 9433 16294
rect 9457 16292 9513 16294
rect 9537 16292 9593 16294
rect 7562 10668 7618 10704
rect 7562 10648 7564 10668
rect 7564 10648 7616 10668
rect 7616 10648 7618 10668
rect 7838 9696 7894 9752
rect 8298 11228 8300 11248
rect 8300 11228 8352 11248
rect 8352 11228 8354 11248
rect 8298 11192 8354 11228
rect 8022 9988 8078 10024
rect 8022 9968 8024 9988
rect 8024 9968 8076 9988
rect 8076 9968 8078 9988
rect 8206 9696 8262 9752
rect 8666 13776 8722 13832
rect 9297 15258 9353 15260
rect 9377 15258 9433 15260
rect 9457 15258 9513 15260
rect 9537 15258 9593 15260
rect 9297 15206 9343 15258
rect 9343 15206 9353 15258
rect 9377 15206 9407 15258
rect 9407 15206 9419 15258
rect 9419 15206 9433 15258
rect 9457 15206 9471 15258
rect 9471 15206 9483 15258
rect 9483 15206 9513 15258
rect 9537 15206 9547 15258
rect 9547 15206 9593 15258
rect 9297 15204 9353 15206
rect 9377 15204 9433 15206
rect 9457 15204 9513 15206
rect 9537 15204 9593 15206
rect 9297 14170 9353 14172
rect 9377 14170 9433 14172
rect 9457 14170 9513 14172
rect 9537 14170 9593 14172
rect 9297 14118 9343 14170
rect 9343 14118 9353 14170
rect 9377 14118 9407 14170
rect 9407 14118 9419 14170
rect 9419 14118 9433 14170
rect 9457 14118 9471 14170
rect 9471 14118 9483 14170
rect 9483 14118 9513 14170
rect 9537 14118 9547 14170
rect 9547 14118 9593 14170
rect 9297 14116 9353 14118
rect 9377 14116 9433 14118
rect 9457 14116 9513 14118
rect 9537 14116 9593 14118
rect 9586 13912 9642 13968
rect 9678 13776 9734 13832
rect 9297 13082 9353 13084
rect 9377 13082 9433 13084
rect 9457 13082 9513 13084
rect 9537 13082 9593 13084
rect 9297 13030 9343 13082
rect 9343 13030 9353 13082
rect 9377 13030 9407 13082
rect 9407 13030 9419 13082
rect 9419 13030 9433 13082
rect 9457 13030 9471 13082
rect 9471 13030 9483 13082
rect 9483 13030 9513 13082
rect 9537 13030 9547 13082
rect 9547 13030 9593 13082
rect 9297 13028 9353 13030
rect 9377 13028 9433 13030
rect 9457 13028 9513 13030
rect 9537 13028 9593 13030
rect 9678 12980 9734 13016
rect 10138 13368 10194 13424
rect 9678 12960 9680 12980
rect 9680 12960 9732 12980
rect 9732 12960 9734 12980
rect 9297 11994 9353 11996
rect 9377 11994 9433 11996
rect 9457 11994 9513 11996
rect 9537 11994 9593 11996
rect 9297 11942 9343 11994
rect 9343 11942 9353 11994
rect 9377 11942 9407 11994
rect 9407 11942 9419 11994
rect 9419 11942 9433 11994
rect 9457 11942 9471 11994
rect 9471 11942 9483 11994
rect 9483 11942 9513 11994
rect 9537 11942 9547 11994
rect 9547 11942 9593 11994
rect 9297 11940 9353 11942
rect 9377 11940 9433 11942
rect 9457 11940 9513 11942
rect 9537 11940 9593 11942
rect 9034 10920 9090 10976
rect 9586 11056 9642 11112
rect 9297 10906 9353 10908
rect 9377 10906 9433 10908
rect 9457 10906 9513 10908
rect 9537 10906 9593 10908
rect 9297 10854 9343 10906
rect 9343 10854 9353 10906
rect 9377 10854 9407 10906
rect 9407 10854 9419 10906
rect 9419 10854 9433 10906
rect 9457 10854 9471 10906
rect 9471 10854 9483 10906
rect 9483 10854 9513 10906
rect 9537 10854 9547 10906
rect 9547 10854 9593 10906
rect 9297 10852 9353 10854
rect 9377 10852 9433 10854
rect 9457 10852 9513 10854
rect 9537 10852 9593 10854
rect 9770 9968 9826 10024
rect 9297 9818 9353 9820
rect 9377 9818 9433 9820
rect 9457 9818 9513 9820
rect 9537 9818 9593 9820
rect 9297 9766 9343 9818
rect 9343 9766 9353 9818
rect 9377 9766 9407 9818
rect 9407 9766 9419 9818
rect 9419 9766 9433 9818
rect 9457 9766 9471 9818
rect 9471 9766 9483 9818
rect 9483 9766 9513 9818
rect 9537 9766 9547 9818
rect 9547 9766 9593 9818
rect 9297 9764 9353 9766
rect 9377 9764 9433 9766
rect 9457 9764 9513 9766
rect 9537 9764 9593 9766
rect 9297 8730 9353 8732
rect 9377 8730 9433 8732
rect 9457 8730 9513 8732
rect 9537 8730 9593 8732
rect 9297 8678 9343 8730
rect 9343 8678 9353 8730
rect 9377 8678 9407 8730
rect 9407 8678 9419 8730
rect 9419 8678 9433 8730
rect 9457 8678 9471 8730
rect 9471 8678 9483 8730
rect 9483 8678 9513 8730
rect 9537 8678 9547 8730
rect 9547 8678 9593 8730
rect 9297 8676 9353 8678
rect 9377 8676 9433 8678
rect 9457 8676 9513 8678
rect 9537 8676 9593 8678
rect 9297 7642 9353 7644
rect 9377 7642 9433 7644
rect 9457 7642 9513 7644
rect 9537 7642 9593 7644
rect 9297 7590 9343 7642
rect 9343 7590 9353 7642
rect 9377 7590 9407 7642
rect 9407 7590 9419 7642
rect 9419 7590 9433 7642
rect 9457 7590 9471 7642
rect 9471 7590 9483 7642
rect 9483 7590 9513 7642
rect 9537 7590 9547 7642
rect 9547 7590 9593 7642
rect 9297 7588 9353 7590
rect 9377 7588 9433 7590
rect 9457 7588 9513 7590
rect 9537 7588 9593 7590
rect 9297 6554 9353 6556
rect 9377 6554 9433 6556
rect 9457 6554 9513 6556
rect 9537 6554 9593 6556
rect 9297 6502 9343 6554
rect 9343 6502 9353 6554
rect 9377 6502 9407 6554
rect 9407 6502 9419 6554
rect 9419 6502 9433 6554
rect 9457 6502 9471 6554
rect 9471 6502 9483 6554
rect 9483 6502 9513 6554
rect 9537 6502 9547 6554
rect 9547 6502 9593 6554
rect 9297 6500 9353 6502
rect 9377 6500 9433 6502
rect 9457 6500 9513 6502
rect 9537 6500 9593 6502
rect 10322 13096 10378 13152
rect 9297 5466 9353 5468
rect 9377 5466 9433 5468
rect 9457 5466 9513 5468
rect 9537 5466 9593 5468
rect 9297 5414 9343 5466
rect 9343 5414 9353 5466
rect 9377 5414 9407 5466
rect 9407 5414 9419 5466
rect 9419 5414 9433 5466
rect 9457 5414 9471 5466
rect 9471 5414 9483 5466
rect 9483 5414 9513 5466
rect 9537 5414 9547 5466
rect 9547 5414 9593 5466
rect 9297 5412 9353 5414
rect 9377 5412 9433 5414
rect 9457 5412 9513 5414
rect 9537 5412 9593 5414
rect 9297 4378 9353 4380
rect 9377 4378 9433 4380
rect 9457 4378 9513 4380
rect 9537 4378 9593 4380
rect 9297 4326 9343 4378
rect 9343 4326 9353 4378
rect 9377 4326 9407 4378
rect 9407 4326 9419 4378
rect 9419 4326 9433 4378
rect 9457 4326 9471 4378
rect 9471 4326 9483 4378
rect 9483 4326 9513 4378
rect 9537 4326 9547 4378
rect 9547 4326 9593 4378
rect 9297 4324 9353 4326
rect 9377 4324 9433 4326
rect 9457 4324 9513 4326
rect 9537 4324 9593 4326
rect 10230 11192 10286 11248
rect 9297 3290 9353 3292
rect 9377 3290 9433 3292
rect 9457 3290 9513 3292
rect 9537 3290 9593 3292
rect 9297 3238 9343 3290
rect 9343 3238 9353 3290
rect 9377 3238 9407 3290
rect 9407 3238 9419 3290
rect 9419 3238 9433 3290
rect 9457 3238 9471 3290
rect 9471 3238 9483 3290
rect 9483 3238 9513 3290
rect 9537 3238 9547 3290
rect 9547 3238 9593 3290
rect 9297 3236 9353 3238
rect 9377 3236 9433 3238
rect 9457 3236 9513 3238
rect 9537 3236 9593 3238
rect 10874 13388 10930 13424
rect 10874 13368 10876 13388
rect 10876 13368 10928 13388
rect 10928 13368 10930 13388
rect 12070 21936 12126 21992
rect 12346 19352 12402 19408
rect 11610 12824 11666 12880
rect 11886 13096 11942 13152
rect 13468 26682 13524 26684
rect 13548 26682 13604 26684
rect 13628 26682 13684 26684
rect 13708 26682 13764 26684
rect 13468 26630 13514 26682
rect 13514 26630 13524 26682
rect 13548 26630 13578 26682
rect 13578 26630 13590 26682
rect 13590 26630 13604 26682
rect 13628 26630 13642 26682
rect 13642 26630 13654 26682
rect 13654 26630 13684 26682
rect 13708 26630 13718 26682
rect 13718 26630 13764 26682
rect 13468 26628 13524 26630
rect 13548 26628 13604 26630
rect 13628 26628 13684 26630
rect 13708 26628 13764 26630
rect 13468 25594 13524 25596
rect 13548 25594 13604 25596
rect 13628 25594 13684 25596
rect 13708 25594 13764 25596
rect 13468 25542 13514 25594
rect 13514 25542 13524 25594
rect 13548 25542 13578 25594
rect 13578 25542 13590 25594
rect 13590 25542 13604 25594
rect 13628 25542 13642 25594
rect 13642 25542 13654 25594
rect 13654 25542 13684 25594
rect 13708 25542 13718 25594
rect 13718 25542 13764 25594
rect 13468 25540 13524 25542
rect 13548 25540 13604 25542
rect 13628 25540 13684 25542
rect 13708 25540 13764 25542
rect 13468 24506 13524 24508
rect 13548 24506 13604 24508
rect 13628 24506 13684 24508
rect 13708 24506 13764 24508
rect 13468 24454 13514 24506
rect 13514 24454 13524 24506
rect 13548 24454 13578 24506
rect 13578 24454 13590 24506
rect 13590 24454 13604 24506
rect 13628 24454 13642 24506
rect 13642 24454 13654 24506
rect 13654 24454 13684 24506
rect 13708 24454 13718 24506
rect 13718 24454 13764 24506
rect 13468 24452 13524 24454
rect 13548 24452 13604 24454
rect 13628 24452 13684 24454
rect 13708 24452 13764 24454
rect 13468 23418 13524 23420
rect 13548 23418 13604 23420
rect 13628 23418 13684 23420
rect 13708 23418 13764 23420
rect 13468 23366 13514 23418
rect 13514 23366 13524 23418
rect 13548 23366 13578 23418
rect 13578 23366 13590 23418
rect 13590 23366 13604 23418
rect 13628 23366 13642 23418
rect 13642 23366 13654 23418
rect 13654 23366 13684 23418
rect 13708 23366 13718 23418
rect 13718 23366 13764 23418
rect 13468 23364 13524 23366
rect 13548 23364 13604 23366
rect 13628 23364 13684 23366
rect 13708 23364 13764 23366
rect 12254 15444 12256 15464
rect 12256 15444 12308 15464
rect 12308 15444 12310 15464
rect 12254 15408 12310 15444
rect 12622 15408 12678 15464
rect 11150 8472 11206 8528
rect 12438 12960 12494 13016
rect 12622 13388 12678 13424
rect 12622 13368 12624 13388
rect 12624 13368 12676 13388
rect 12676 13368 12678 13388
rect 12714 13232 12770 13288
rect 13468 22330 13524 22332
rect 13548 22330 13604 22332
rect 13628 22330 13684 22332
rect 13708 22330 13764 22332
rect 13468 22278 13514 22330
rect 13514 22278 13524 22330
rect 13548 22278 13578 22330
rect 13578 22278 13590 22330
rect 13590 22278 13604 22330
rect 13628 22278 13642 22330
rect 13642 22278 13654 22330
rect 13654 22278 13684 22330
rect 13708 22278 13718 22330
rect 13718 22278 13764 22330
rect 13468 22276 13524 22278
rect 13548 22276 13604 22278
rect 13628 22276 13684 22278
rect 13708 22276 13764 22278
rect 12898 20304 12954 20360
rect 12990 19796 12992 19816
rect 12992 19796 13044 19816
rect 13044 19796 13046 19816
rect 12990 19760 13046 19796
rect 13468 21242 13524 21244
rect 13548 21242 13604 21244
rect 13628 21242 13684 21244
rect 13708 21242 13764 21244
rect 13468 21190 13514 21242
rect 13514 21190 13524 21242
rect 13548 21190 13578 21242
rect 13578 21190 13590 21242
rect 13590 21190 13604 21242
rect 13628 21190 13642 21242
rect 13642 21190 13654 21242
rect 13654 21190 13684 21242
rect 13708 21190 13718 21242
rect 13718 21190 13764 21242
rect 13468 21188 13524 21190
rect 13548 21188 13604 21190
rect 13628 21188 13684 21190
rect 13708 21188 13764 21190
rect 13468 20154 13524 20156
rect 13548 20154 13604 20156
rect 13628 20154 13684 20156
rect 13708 20154 13764 20156
rect 13468 20102 13514 20154
rect 13514 20102 13524 20154
rect 13548 20102 13578 20154
rect 13578 20102 13590 20154
rect 13590 20102 13604 20154
rect 13628 20102 13642 20154
rect 13642 20102 13654 20154
rect 13654 20102 13684 20154
rect 13708 20102 13718 20154
rect 13718 20102 13764 20154
rect 13468 20100 13524 20102
rect 13548 20100 13604 20102
rect 13628 20100 13684 20102
rect 13708 20100 13764 20102
rect 13468 19066 13524 19068
rect 13548 19066 13604 19068
rect 13628 19066 13684 19068
rect 13708 19066 13764 19068
rect 13468 19014 13514 19066
rect 13514 19014 13524 19066
rect 13548 19014 13578 19066
rect 13578 19014 13590 19066
rect 13590 19014 13604 19066
rect 13628 19014 13642 19066
rect 13642 19014 13654 19066
rect 13654 19014 13684 19066
rect 13708 19014 13718 19066
rect 13718 19014 13764 19066
rect 13468 19012 13524 19014
rect 13548 19012 13604 19014
rect 13628 19012 13684 19014
rect 13708 19012 13764 19014
rect 13468 17978 13524 17980
rect 13548 17978 13604 17980
rect 13628 17978 13684 17980
rect 13708 17978 13764 17980
rect 13468 17926 13514 17978
rect 13514 17926 13524 17978
rect 13548 17926 13578 17978
rect 13578 17926 13590 17978
rect 13590 17926 13604 17978
rect 13628 17926 13642 17978
rect 13642 17926 13654 17978
rect 13654 17926 13684 17978
rect 13708 17926 13718 17978
rect 13718 17926 13764 17978
rect 13468 17924 13524 17926
rect 13548 17924 13604 17926
rect 13628 17924 13684 17926
rect 13708 17924 13764 17926
rect 12714 8492 12770 8528
rect 12714 8472 12716 8492
rect 12716 8472 12768 8492
rect 12768 8472 12770 8492
rect 9297 2202 9353 2204
rect 9377 2202 9433 2204
rect 9457 2202 9513 2204
rect 9537 2202 9593 2204
rect 9297 2150 9343 2202
rect 9343 2150 9353 2202
rect 9377 2150 9407 2202
rect 9407 2150 9419 2202
rect 9419 2150 9433 2202
rect 9457 2150 9471 2202
rect 9471 2150 9483 2202
rect 9483 2150 9513 2202
rect 9537 2150 9547 2202
rect 9547 2150 9593 2202
rect 9297 2148 9353 2150
rect 9377 2148 9433 2150
rect 9457 2148 9513 2150
rect 9537 2148 9593 2150
rect 12990 12844 13046 12880
rect 12990 12824 12992 12844
rect 12992 12824 13044 12844
rect 13044 12824 13046 12844
rect 13468 16890 13524 16892
rect 13548 16890 13604 16892
rect 13628 16890 13684 16892
rect 13708 16890 13764 16892
rect 13468 16838 13514 16890
rect 13514 16838 13524 16890
rect 13548 16838 13578 16890
rect 13578 16838 13590 16890
rect 13590 16838 13604 16890
rect 13628 16838 13642 16890
rect 13642 16838 13654 16890
rect 13654 16838 13684 16890
rect 13708 16838 13718 16890
rect 13718 16838 13764 16890
rect 13468 16836 13524 16838
rect 13548 16836 13604 16838
rect 13628 16836 13684 16838
rect 13708 16836 13764 16838
rect 13468 15802 13524 15804
rect 13548 15802 13604 15804
rect 13628 15802 13684 15804
rect 13708 15802 13764 15804
rect 13468 15750 13514 15802
rect 13514 15750 13524 15802
rect 13548 15750 13578 15802
rect 13578 15750 13590 15802
rect 13590 15750 13604 15802
rect 13628 15750 13642 15802
rect 13642 15750 13654 15802
rect 13654 15750 13684 15802
rect 13708 15750 13718 15802
rect 13718 15750 13764 15802
rect 13468 15748 13524 15750
rect 13548 15748 13604 15750
rect 13628 15748 13684 15750
rect 13708 15748 13764 15750
rect 13634 15444 13636 15464
rect 13636 15444 13688 15464
rect 13688 15444 13690 15464
rect 13634 15408 13690 15444
rect 13468 14714 13524 14716
rect 13548 14714 13604 14716
rect 13628 14714 13684 14716
rect 13708 14714 13764 14716
rect 13468 14662 13514 14714
rect 13514 14662 13524 14714
rect 13548 14662 13578 14714
rect 13578 14662 13590 14714
rect 13590 14662 13604 14714
rect 13628 14662 13642 14714
rect 13642 14662 13654 14714
rect 13654 14662 13684 14714
rect 13708 14662 13718 14714
rect 13718 14662 13764 14714
rect 13468 14660 13524 14662
rect 13548 14660 13604 14662
rect 13628 14660 13684 14662
rect 13708 14660 13764 14662
rect 13468 13626 13524 13628
rect 13548 13626 13604 13628
rect 13628 13626 13684 13628
rect 13708 13626 13764 13628
rect 13468 13574 13514 13626
rect 13514 13574 13524 13626
rect 13548 13574 13578 13626
rect 13578 13574 13590 13626
rect 13590 13574 13604 13626
rect 13628 13574 13642 13626
rect 13642 13574 13654 13626
rect 13654 13574 13684 13626
rect 13708 13574 13718 13626
rect 13718 13574 13764 13626
rect 13468 13572 13524 13574
rect 13548 13572 13604 13574
rect 13628 13572 13684 13574
rect 13708 13572 13764 13574
rect 13542 13268 13544 13288
rect 13544 13268 13596 13288
rect 13596 13268 13598 13288
rect 13542 13232 13598 13268
rect 13468 12538 13524 12540
rect 13548 12538 13604 12540
rect 13628 12538 13684 12540
rect 13708 12538 13764 12540
rect 13468 12486 13514 12538
rect 13514 12486 13524 12538
rect 13548 12486 13578 12538
rect 13578 12486 13590 12538
rect 13590 12486 13604 12538
rect 13628 12486 13642 12538
rect 13642 12486 13654 12538
rect 13654 12486 13684 12538
rect 13708 12486 13718 12538
rect 13718 12486 13764 12538
rect 13468 12484 13524 12486
rect 13548 12484 13604 12486
rect 13628 12484 13684 12486
rect 13708 12484 13764 12486
rect 13468 11450 13524 11452
rect 13548 11450 13604 11452
rect 13628 11450 13684 11452
rect 13708 11450 13764 11452
rect 13468 11398 13514 11450
rect 13514 11398 13524 11450
rect 13548 11398 13578 11450
rect 13578 11398 13590 11450
rect 13590 11398 13604 11450
rect 13628 11398 13642 11450
rect 13642 11398 13654 11450
rect 13654 11398 13684 11450
rect 13708 11398 13718 11450
rect 13718 11398 13764 11450
rect 13468 11396 13524 11398
rect 13548 11396 13604 11398
rect 13628 11396 13684 11398
rect 13708 11396 13764 11398
rect 13468 10362 13524 10364
rect 13548 10362 13604 10364
rect 13628 10362 13684 10364
rect 13708 10362 13764 10364
rect 13468 10310 13514 10362
rect 13514 10310 13524 10362
rect 13548 10310 13578 10362
rect 13578 10310 13590 10362
rect 13590 10310 13604 10362
rect 13628 10310 13642 10362
rect 13642 10310 13654 10362
rect 13654 10310 13684 10362
rect 13708 10310 13718 10362
rect 13718 10310 13764 10362
rect 13468 10308 13524 10310
rect 13548 10308 13604 10310
rect 13628 10308 13684 10310
rect 13708 10308 13764 10310
rect 13468 9274 13524 9276
rect 13548 9274 13604 9276
rect 13628 9274 13684 9276
rect 13708 9274 13764 9276
rect 13468 9222 13514 9274
rect 13514 9222 13524 9274
rect 13548 9222 13578 9274
rect 13578 9222 13590 9274
rect 13590 9222 13604 9274
rect 13628 9222 13642 9274
rect 13642 9222 13654 9274
rect 13654 9222 13684 9274
rect 13708 9222 13718 9274
rect 13718 9222 13764 9274
rect 13468 9220 13524 9222
rect 13548 9220 13604 9222
rect 13628 9220 13684 9222
rect 13708 9220 13764 9222
rect 13468 8186 13524 8188
rect 13548 8186 13604 8188
rect 13628 8186 13684 8188
rect 13708 8186 13764 8188
rect 13468 8134 13514 8186
rect 13514 8134 13524 8186
rect 13548 8134 13578 8186
rect 13578 8134 13590 8186
rect 13590 8134 13604 8186
rect 13628 8134 13642 8186
rect 13642 8134 13654 8186
rect 13654 8134 13684 8186
rect 13708 8134 13718 8186
rect 13718 8134 13764 8186
rect 13468 8132 13524 8134
rect 13548 8132 13604 8134
rect 13628 8132 13684 8134
rect 13708 8132 13764 8134
rect 14002 11500 14004 11520
rect 14004 11500 14056 11520
rect 14056 11500 14058 11520
rect 14002 11464 14058 11500
rect 14646 14476 14702 14512
rect 14646 14456 14648 14476
rect 14648 14456 14700 14476
rect 14700 14456 14702 14476
rect 14462 13096 14518 13152
rect 13468 7098 13524 7100
rect 13548 7098 13604 7100
rect 13628 7098 13684 7100
rect 13708 7098 13764 7100
rect 13468 7046 13514 7098
rect 13514 7046 13524 7098
rect 13548 7046 13578 7098
rect 13578 7046 13590 7098
rect 13590 7046 13604 7098
rect 13628 7046 13642 7098
rect 13642 7046 13654 7098
rect 13654 7046 13684 7098
rect 13708 7046 13718 7098
rect 13718 7046 13764 7098
rect 13468 7044 13524 7046
rect 13548 7044 13604 7046
rect 13628 7044 13684 7046
rect 13708 7044 13764 7046
rect 13468 6010 13524 6012
rect 13548 6010 13604 6012
rect 13628 6010 13684 6012
rect 13708 6010 13764 6012
rect 13468 5958 13514 6010
rect 13514 5958 13524 6010
rect 13548 5958 13578 6010
rect 13578 5958 13590 6010
rect 13590 5958 13604 6010
rect 13628 5958 13642 6010
rect 13642 5958 13654 6010
rect 13654 5958 13684 6010
rect 13708 5958 13718 6010
rect 13718 5958 13764 6010
rect 13468 5956 13524 5958
rect 13548 5956 13604 5958
rect 13628 5956 13684 5958
rect 13708 5956 13764 5958
rect 13468 4922 13524 4924
rect 13548 4922 13604 4924
rect 13628 4922 13684 4924
rect 13708 4922 13764 4924
rect 13468 4870 13514 4922
rect 13514 4870 13524 4922
rect 13548 4870 13578 4922
rect 13578 4870 13590 4922
rect 13590 4870 13604 4922
rect 13628 4870 13642 4922
rect 13642 4870 13654 4922
rect 13654 4870 13684 4922
rect 13708 4870 13718 4922
rect 13718 4870 13764 4922
rect 13468 4868 13524 4870
rect 13548 4868 13604 4870
rect 13628 4868 13684 4870
rect 13708 4868 13764 4870
rect 13468 3834 13524 3836
rect 13548 3834 13604 3836
rect 13628 3834 13684 3836
rect 13708 3834 13764 3836
rect 13468 3782 13514 3834
rect 13514 3782 13524 3834
rect 13548 3782 13578 3834
rect 13578 3782 13590 3834
rect 13590 3782 13604 3834
rect 13628 3782 13642 3834
rect 13642 3782 13654 3834
rect 13654 3782 13684 3834
rect 13708 3782 13718 3834
rect 13718 3782 13764 3834
rect 13468 3780 13524 3782
rect 13548 3780 13604 3782
rect 13628 3780 13684 3782
rect 13708 3780 13764 3782
rect 15382 14476 15438 14512
rect 15382 14456 15384 14476
rect 15384 14456 15436 14476
rect 15436 14456 15438 14476
rect 15106 12280 15162 12336
rect 14646 10648 14702 10704
rect 17638 27226 17694 27228
rect 17718 27226 17774 27228
rect 17798 27226 17854 27228
rect 17878 27226 17934 27228
rect 17638 27174 17684 27226
rect 17684 27174 17694 27226
rect 17718 27174 17748 27226
rect 17748 27174 17760 27226
rect 17760 27174 17774 27226
rect 17798 27174 17812 27226
rect 17812 27174 17824 27226
rect 17824 27174 17854 27226
rect 17878 27174 17888 27226
rect 17888 27174 17934 27226
rect 17638 27172 17694 27174
rect 17718 27172 17774 27174
rect 17798 27172 17854 27174
rect 17878 27172 17934 27174
rect 17638 26138 17694 26140
rect 17718 26138 17774 26140
rect 17798 26138 17854 26140
rect 17878 26138 17934 26140
rect 17638 26086 17684 26138
rect 17684 26086 17694 26138
rect 17718 26086 17748 26138
rect 17748 26086 17760 26138
rect 17760 26086 17774 26138
rect 17798 26086 17812 26138
rect 17812 26086 17824 26138
rect 17824 26086 17854 26138
rect 17878 26086 17888 26138
rect 17888 26086 17934 26138
rect 17638 26084 17694 26086
rect 17718 26084 17774 26086
rect 17798 26084 17854 26086
rect 17878 26084 17934 26086
rect 17638 25050 17694 25052
rect 17718 25050 17774 25052
rect 17798 25050 17854 25052
rect 17878 25050 17934 25052
rect 17638 24998 17684 25050
rect 17684 24998 17694 25050
rect 17718 24998 17748 25050
rect 17748 24998 17760 25050
rect 17760 24998 17774 25050
rect 17798 24998 17812 25050
rect 17812 24998 17824 25050
rect 17824 24998 17854 25050
rect 17878 24998 17888 25050
rect 17888 24998 17934 25050
rect 17638 24996 17694 24998
rect 17718 24996 17774 24998
rect 17798 24996 17854 24998
rect 17878 24996 17934 24998
rect 17638 23962 17694 23964
rect 17718 23962 17774 23964
rect 17798 23962 17854 23964
rect 17878 23962 17934 23964
rect 17638 23910 17684 23962
rect 17684 23910 17694 23962
rect 17718 23910 17748 23962
rect 17748 23910 17760 23962
rect 17760 23910 17774 23962
rect 17798 23910 17812 23962
rect 17812 23910 17824 23962
rect 17824 23910 17854 23962
rect 17878 23910 17888 23962
rect 17888 23910 17934 23962
rect 17638 23908 17694 23910
rect 17718 23908 17774 23910
rect 17798 23908 17854 23910
rect 17878 23908 17934 23910
rect 17638 22874 17694 22876
rect 17718 22874 17774 22876
rect 17798 22874 17854 22876
rect 17878 22874 17934 22876
rect 17638 22822 17684 22874
rect 17684 22822 17694 22874
rect 17718 22822 17748 22874
rect 17748 22822 17760 22874
rect 17760 22822 17774 22874
rect 17798 22822 17812 22874
rect 17812 22822 17824 22874
rect 17824 22822 17854 22874
rect 17878 22822 17888 22874
rect 17888 22822 17934 22874
rect 17638 22820 17694 22822
rect 17718 22820 17774 22822
rect 17798 22820 17854 22822
rect 17878 22820 17934 22822
rect 17638 21786 17694 21788
rect 17718 21786 17774 21788
rect 17798 21786 17854 21788
rect 17878 21786 17934 21788
rect 17638 21734 17684 21786
rect 17684 21734 17694 21786
rect 17718 21734 17748 21786
rect 17748 21734 17760 21786
rect 17760 21734 17774 21786
rect 17798 21734 17812 21786
rect 17812 21734 17824 21786
rect 17824 21734 17854 21786
rect 17878 21734 17888 21786
rect 17888 21734 17934 21786
rect 17638 21732 17694 21734
rect 17718 21732 17774 21734
rect 17798 21732 17854 21734
rect 17878 21732 17934 21734
rect 17638 20698 17694 20700
rect 17718 20698 17774 20700
rect 17798 20698 17854 20700
rect 17878 20698 17934 20700
rect 17638 20646 17684 20698
rect 17684 20646 17694 20698
rect 17718 20646 17748 20698
rect 17748 20646 17760 20698
rect 17760 20646 17774 20698
rect 17798 20646 17812 20698
rect 17812 20646 17824 20698
rect 17824 20646 17854 20698
rect 17878 20646 17888 20698
rect 17888 20646 17934 20698
rect 17638 20644 17694 20646
rect 17718 20644 17774 20646
rect 17798 20644 17854 20646
rect 17878 20644 17934 20646
rect 17638 19610 17694 19612
rect 17718 19610 17774 19612
rect 17798 19610 17854 19612
rect 17878 19610 17934 19612
rect 17638 19558 17684 19610
rect 17684 19558 17694 19610
rect 17718 19558 17748 19610
rect 17748 19558 17760 19610
rect 17760 19558 17774 19610
rect 17798 19558 17812 19610
rect 17812 19558 17824 19610
rect 17824 19558 17854 19610
rect 17878 19558 17888 19610
rect 17888 19558 17934 19610
rect 17638 19556 17694 19558
rect 17718 19556 17774 19558
rect 17798 19556 17854 19558
rect 17878 19556 17934 19558
rect 21809 26682 21865 26684
rect 21889 26682 21945 26684
rect 21969 26682 22025 26684
rect 22049 26682 22105 26684
rect 21809 26630 21855 26682
rect 21855 26630 21865 26682
rect 21889 26630 21919 26682
rect 21919 26630 21931 26682
rect 21931 26630 21945 26682
rect 21969 26630 21983 26682
rect 21983 26630 21995 26682
rect 21995 26630 22025 26682
rect 22049 26630 22059 26682
rect 22059 26630 22105 26682
rect 21809 26628 21865 26630
rect 21889 26628 21945 26630
rect 21969 26628 22025 26630
rect 22049 26628 22105 26630
rect 26238 28484 26294 28520
rect 26238 28464 26240 28484
rect 26240 28464 26292 28484
rect 26292 28464 26294 28484
rect 21809 25594 21865 25596
rect 21889 25594 21945 25596
rect 21969 25594 22025 25596
rect 22049 25594 22105 25596
rect 21809 25542 21855 25594
rect 21855 25542 21865 25594
rect 21889 25542 21919 25594
rect 21919 25542 21931 25594
rect 21931 25542 21945 25594
rect 21969 25542 21983 25594
rect 21983 25542 21995 25594
rect 21995 25542 22025 25594
rect 22049 25542 22059 25594
rect 22059 25542 22105 25594
rect 21809 25540 21865 25542
rect 21889 25540 21945 25542
rect 21969 25540 22025 25542
rect 22049 25540 22105 25542
rect 25042 25356 25098 25392
rect 25042 25336 25044 25356
rect 25044 25336 25096 25356
rect 25096 25336 25098 25356
rect 21809 24506 21865 24508
rect 21889 24506 21945 24508
rect 21969 24506 22025 24508
rect 22049 24506 22105 24508
rect 21809 24454 21855 24506
rect 21855 24454 21865 24506
rect 21889 24454 21919 24506
rect 21919 24454 21931 24506
rect 21931 24454 21945 24506
rect 21969 24454 21983 24506
rect 21983 24454 21995 24506
rect 21995 24454 22025 24506
rect 22049 24454 22059 24506
rect 22059 24454 22105 24506
rect 21809 24452 21865 24454
rect 21889 24452 21945 24454
rect 21969 24452 22025 24454
rect 22049 24452 22105 24454
rect 21809 23418 21865 23420
rect 21889 23418 21945 23420
rect 21969 23418 22025 23420
rect 22049 23418 22105 23420
rect 21809 23366 21855 23418
rect 21855 23366 21865 23418
rect 21889 23366 21919 23418
rect 21919 23366 21931 23418
rect 21931 23366 21945 23418
rect 21969 23366 21983 23418
rect 21983 23366 21995 23418
rect 21995 23366 22025 23418
rect 22049 23366 22059 23418
rect 22059 23366 22105 23418
rect 21809 23364 21865 23366
rect 21889 23364 21945 23366
rect 21969 23364 22025 23366
rect 22049 23364 22105 23366
rect 17638 18522 17694 18524
rect 17718 18522 17774 18524
rect 17798 18522 17854 18524
rect 17878 18522 17934 18524
rect 17638 18470 17684 18522
rect 17684 18470 17694 18522
rect 17718 18470 17748 18522
rect 17748 18470 17760 18522
rect 17760 18470 17774 18522
rect 17798 18470 17812 18522
rect 17812 18470 17824 18522
rect 17824 18470 17854 18522
rect 17878 18470 17888 18522
rect 17888 18470 17934 18522
rect 17638 18468 17694 18470
rect 17718 18468 17774 18470
rect 17798 18468 17854 18470
rect 17878 18468 17934 18470
rect 15658 12280 15714 12336
rect 13468 2746 13524 2748
rect 13548 2746 13604 2748
rect 13628 2746 13684 2748
rect 13708 2746 13764 2748
rect 13468 2694 13514 2746
rect 13514 2694 13524 2746
rect 13548 2694 13578 2746
rect 13578 2694 13590 2746
rect 13590 2694 13604 2746
rect 13628 2694 13642 2746
rect 13642 2694 13654 2746
rect 13654 2694 13684 2746
rect 13708 2694 13718 2746
rect 13718 2694 13764 2746
rect 13468 2692 13524 2694
rect 13548 2692 13604 2694
rect 13628 2692 13684 2694
rect 13708 2692 13764 2694
rect 16578 11228 16580 11248
rect 16580 11228 16632 11248
rect 16632 11228 16634 11248
rect 16578 11192 16634 11228
rect 17638 17434 17694 17436
rect 17718 17434 17774 17436
rect 17798 17434 17854 17436
rect 17878 17434 17934 17436
rect 17638 17382 17684 17434
rect 17684 17382 17694 17434
rect 17718 17382 17748 17434
rect 17748 17382 17760 17434
rect 17760 17382 17774 17434
rect 17798 17382 17812 17434
rect 17812 17382 17824 17434
rect 17824 17382 17854 17434
rect 17878 17382 17888 17434
rect 17888 17382 17934 17434
rect 17638 17380 17694 17382
rect 17718 17380 17774 17382
rect 17798 17380 17854 17382
rect 17878 17380 17934 17382
rect 17638 16346 17694 16348
rect 17718 16346 17774 16348
rect 17798 16346 17854 16348
rect 17878 16346 17934 16348
rect 17638 16294 17684 16346
rect 17684 16294 17694 16346
rect 17718 16294 17748 16346
rect 17748 16294 17760 16346
rect 17760 16294 17774 16346
rect 17798 16294 17812 16346
rect 17812 16294 17824 16346
rect 17824 16294 17854 16346
rect 17878 16294 17888 16346
rect 17888 16294 17934 16346
rect 17638 16292 17694 16294
rect 17718 16292 17774 16294
rect 17798 16292 17854 16294
rect 17878 16292 17934 16294
rect 17638 15258 17694 15260
rect 17718 15258 17774 15260
rect 17798 15258 17854 15260
rect 17878 15258 17934 15260
rect 17638 15206 17684 15258
rect 17684 15206 17694 15258
rect 17718 15206 17748 15258
rect 17748 15206 17760 15258
rect 17760 15206 17774 15258
rect 17798 15206 17812 15258
rect 17812 15206 17824 15258
rect 17824 15206 17854 15258
rect 17878 15206 17888 15258
rect 17888 15206 17934 15258
rect 17638 15204 17694 15206
rect 17718 15204 17774 15206
rect 17798 15204 17854 15206
rect 17878 15204 17934 15206
rect 17638 14170 17694 14172
rect 17718 14170 17774 14172
rect 17798 14170 17854 14172
rect 17878 14170 17934 14172
rect 17638 14118 17684 14170
rect 17684 14118 17694 14170
rect 17718 14118 17748 14170
rect 17748 14118 17760 14170
rect 17760 14118 17774 14170
rect 17798 14118 17812 14170
rect 17812 14118 17824 14170
rect 17824 14118 17854 14170
rect 17878 14118 17888 14170
rect 17888 14118 17934 14170
rect 17638 14116 17694 14118
rect 17718 14116 17774 14118
rect 17798 14116 17854 14118
rect 17878 14116 17934 14118
rect 19798 20304 19854 20360
rect 19706 19372 19762 19408
rect 19706 19352 19708 19372
rect 19708 19352 19760 19372
rect 19760 19352 19762 19372
rect 17638 13082 17694 13084
rect 17718 13082 17774 13084
rect 17798 13082 17854 13084
rect 17878 13082 17934 13084
rect 17638 13030 17684 13082
rect 17684 13030 17694 13082
rect 17718 13030 17748 13082
rect 17748 13030 17760 13082
rect 17760 13030 17774 13082
rect 17798 13030 17812 13082
rect 17812 13030 17824 13082
rect 17824 13030 17854 13082
rect 17878 13030 17888 13082
rect 17888 13030 17934 13082
rect 17638 13028 17694 13030
rect 17718 13028 17774 13030
rect 17798 13028 17854 13030
rect 17878 13028 17934 13030
rect 17638 11994 17694 11996
rect 17718 11994 17774 11996
rect 17798 11994 17854 11996
rect 17878 11994 17934 11996
rect 17638 11942 17684 11994
rect 17684 11942 17694 11994
rect 17718 11942 17748 11994
rect 17748 11942 17760 11994
rect 17760 11942 17774 11994
rect 17798 11942 17812 11994
rect 17812 11942 17824 11994
rect 17824 11942 17854 11994
rect 17878 11942 17888 11994
rect 17888 11942 17934 11994
rect 17638 11940 17694 11942
rect 17718 11940 17774 11942
rect 17798 11940 17854 11942
rect 17878 11940 17934 11942
rect 17222 11500 17224 11520
rect 17224 11500 17276 11520
rect 17276 11500 17278 11520
rect 17222 11464 17278 11500
rect 17638 10906 17694 10908
rect 17718 10906 17774 10908
rect 17798 10906 17854 10908
rect 17878 10906 17934 10908
rect 17638 10854 17684 10906
rect 17684 10854 17694 10906
rect 17718 10854 17748 10906
rect 17748 10854 17760 10906
rect 17760 10854 17774 10906
rect 17798 10854 17812 10906
rect 17812 10854 17824 10906
rect 17824 10854 17854 10906
rect 17878 10854 17888 10906
rect 17888 10854 17934 10906
rect 17638 10852 17694 10854
rect 17718 10852 17774 10854
rect 17798 10852 17854 10854
rect 17878 10852 17934 10854
rect 17638 9818 17694 9820
rect 17718 9818 17774 9820
rect 17798 9818 17854 9820
rect 17878 9818 17934 9820
rect 17638 9766 17684 9818
rect 17684 9766 17694 9818
rect 17718 9766 17748 9818
rect 17748 9766 17760 9818
rect 17760 9766 17774 9818
rect 17798 9766 17812 9818
rect 17812 9766 17824 9818
rect 17824 9766 17854 9818
rect 17878 9766 17888 9818
rect 17888 9766 17934 9818
rect 17638 9764 17694 9766
rect 17718 9764 17774 9766
rect 17798 9764 17854 9766
rect 17878 9764 17934 9766
rect 17638 8730 17694 8732
rect 17718 8730 17774 8732
rect 17798 8730 17854 8732
rect 17878 8730 17934 8732
rect 17638 8678 17684 8730
rect 17684 8678 17694 8730
rect 17718 8678 17748 8730
rect 17748 8678 17760 8730
rect 17760 8678 17774 8730
rect 17798 8678 17812 8730
rect 17812 8678 17824 8730
rect 17824 8678 17854 8730
rect 17878 8678 17888 8730
rect 17888 8678 17934 8730
rect 17638 8676 17694 8678
rect 17718 8676 17774 8678
rect 17798 8676 17854 8678
rect 17878 8676 17934 8678
rect 17638 7642 17694 7644
rect 17718 7642 17774 7644
rect 17798 7642 17854 7644
rect 17878 7642 17934 7644
rect 17638 7590 17684 7642
rect 17684 7590 17694 7642
rect 17718 7590 17748 7642
rect 17748 7590 17760 7642
rect 17760 7590 17774 7642
rect 17798 7590 17812 7642
rect 17812 7590 17824 7642
rect 17824 7590 17854 7642
rect 17878 7590 17888 7642
rect 17888 7590 17934 7642
rect 17638 7588 17694 7590
rect 17718 7588 17774 7590
rect 17798 7588 17854 7590
rect 17878 7588 17934 7590
rect 17638 6554 17694 6556
rect 17718 6554 17774 6556
rect 17798 6554 17854 6556
rect 17878 6554 17934 6556
rect 17638 6502 17684 6554
rect 17684 6502 17694 6554
rect 17718 6502 17748 6554
rect 17748 6502 17760 6554
rect 17760 6502 17774 6554
rect 17798 6502 17812 6554
rect 17812 6502 17824 6554
rect 17824 6502 17854 6554
rect 17878 6502 17888 6554
rect 17888 6502 17934 6554
rect 17638 6500 17694 6502
rect 17718 6500 17774 6502
rect 17798 6500 17854 6502
rect 17878 6500 17934 6502
rect 17638 5466 17694 5468
rect 17718 5466 17774 5468
rect 17798 5466 17854 5468
rect 17878 5466 17934 5468
rect 17638 5414 17684 5466
rect 17684 5414 17694 5466
rect 17718 5414 17748 5466
rect 17748 5414 17760 5466
rect 17760 5414 17774 5466
rect 17798 5414 17812 5466
rect 17812 5414 17824 5466
rect 17824 5414 17854 5466
rect 17878 5414 17888 5466
rect 17888 5414 17934 5466
rect 17638 5412 17694 5414
rect 17718 5412 17774 5414
rect 17798 5412 17854 5414
rect 17878 5412 17934 5414
rect 17638 4378 17694 4380
rect 17718 4378 17774 4380
rect 17798 4378 17854 4380
rect 17878 4378 17934 4380
rect 17638 4326 17684 4378
rect 17684 4326 17694 4378
rect 17718 4326 17748 4378
rect 17748 4326 17760 4378
rect 17760 4326 17774 4378
rect 17798 4326 17812 4378
rect 17812 4326 17824 4378
rect 17824 4326 17854 4378
rect 17878 4326 17888 4378
rect 17888 4326 17934 4378
rect 17638 4324 17694 4326
rect 17718 4324 17774 4326
rect 17798 4324 17854 4326
rect 17878 4324 17934 4326
rect 17638 3290 17694 3292
rect 17718 3290 17774 3292
rect 17798 3290 17854 3292
rect 17878 3290 17934 3292
rect 17638 3238 17684 3290
rect 17684 3238 17694 3290
rect 17718 3238 17748 3290
rect 17748 3238 17760 3290
rect 17760 3238 17774 3290
rect 17798 3238 17812 3290
rect 17812 3238 17824 3290
rect 17824 3238 17854 3290
rect 17878 3238 17888 3290
rect 17888 3238 17934 3290
rect 17638 3236 17694 3238
rect 17718 3236 17774 3238
rect 17798 3236 17854 3238
rect 17878 3236 17934 3238
rect 21809 22330 21865 22332
rect 21889 22330 21945 22332
rect 21969 22330 22025 22332
rect 22049 22330 22105 22332
rect 21809 22278 21855 22330
rect 21855 22278 21865 22330
rect 21889 22278 21919 22330
rect 21919 22278 21931 22330
rect 21931 22278 21945 22330
rect 21969 22278 21983 22330
rect 21983 22278 21995 22330
rect 21995 22278 22025 22330
rect 22049 22278 22059 22330
rect 22059 22278 22105 22330
rect 21809 22276 21865 22278
rect 21889 22276 21945 22278
rect 21969 22276 22025 22278
rect 22049 22276 22105 22278
rect 21809 21242 21865 21244
rect 21889 21242 21945 21244
rect 21969 21242 22025 21244
rect 22049 21242 22105 21244
rect 21809 21190 21855 21242
rect 21855 21190 21865 21242
rect 21889 21190 21919 21242
rect 21919 21190 21931 21242
rect 21931 21190 21945 21242
rect 21969 21190 21983 21242
rect 21983 21190 21995 21242
rect 21995 21190 22025 21242
rect 22049 21190 22059 21242
rect 22059 21190 22105 21242
rect 21809 21188 21865 21190
rect 21889 21188 21945 21190
rect 21969 21188 22025 21190
rect 22049 21188 22105 21190
rect 21809 20154 21865 20156
rect 21889 20154 21945 20156
rect 21969 20154 22025 20156
rect 22049 20154 22105 20156
rect 21809 20102 21855 20154
rect 21855 20102 21865 20154
rect 21889 20102 21919 20154
rect 21919 20102 21931 20154
rect 21931 20102 21945 20154
rect 21969 20102 21983 20154
rect 21983 20102 21995 20154
rect 21995 20102 22025 20154
rect 22049 20102 22059 20154
rect 22059 20102 22105 20154
rect 21809 20100 21865 20102
rect 21889 20100 21945 20102
rect 21969 20100 22025 20102
rect 22049 20100 22105 20102
rect 21809 19066 21865 19068
rect 21889 19066 21945 19068
rect 21969 19066 22025 19068
rect 22049 19066 22105 19068
rect 21809 19014 21855 19066
rect 21855 19014 21865 19066
rect 21889 19014 21919 19066
rect 21919 19014 21931 19066
rect 21931 19014 21945 19066
rect 21969 19014 21983 19066
rect 21983 19014 21995 19066
rect 21995 19014 22025 19066
rect 22049 19014 22059 19066
rect 22059 19014 22105 19066
rect 21809 19012 21865 19014
rect 21889 19012 21945 19014
rect 21969 19012 22025 19014
rect 22049 19012 22105 19014
rect 21809 17978 21865 17980
rect 21889 17978 21945 17980
rect 21969 17978 22025 17980
rect 22049 17978 22105 17980
rect 21809 17926 21855 17978
rect 21855 17926 21865 17978
rect 21889 17926 21919 17978
rect 21919 17926 21931 17978
rect 21931 17926 21945 17978
rect 21969 17926 21983 17978
rect 21983 17926 21995 17978
rect 21995 17926 22025 17978
rect 22049 17926 22059 17978
rect 22059 17926 22105 17978
rect 21809 17924 21865 17926
rect 21889 17924 21945 17926
rect 21969 17924 22025 17926
rect 22049 17924 22105 17926
rect 21809 16890 21865 16892
rect 21889 16890 21945 16892
rect 21969 16890 22025 16892
rect 22049 16890 22105 16892
rect 21809 16838 21855 16890
rect 21855 16838 21865 16890
rect 21889 16838 21919 16890
rect 21919 16838 21931 16890
rect 21931 16838 21945 16890
rect 21969 16838 21983 16890
rect 21983 16838 21995 16890
rect 21995 16838 22025 16890
rect 22049 16838 22059 16890
rect 22059 16838 22105 16890
rect 21809 16836 21865 16838
rect 21889 16836 21945 16838
rect 21969 16836 22025 16838
rect 22049 16836 22105 16838
rect 23386 17720 23442 17776
rect 20074 9172 20130 9208
rect 20074 9152 20076 9172
rect 20076 9152 20128 9172
rect 20128 9152 20130 9172
rect 20258 9016 20314 9072
rect 20902 9152 20958 9208
rect 21809 15802 21865 15804
rect 21889 15802 21945 15804
rect 21969 15802 22025 15804
rect 22049 15802 22105 15804
rect 21809 15750 21855 15802
rect 21855 15750 21865 15802
rect 21889 15750 21919 15802
rect 21919 15750 21931 15802
rect 21931 15750 21945 15802
rect 21969 15750 21983 15802
rect 21983 15750 21995 15802
rect 21995 15750 22025 15802
rect 22049 15750 22059 15802
rect 22059 15750 22105 15802
rect 21809 15748 21865 15750
rect 21889 15748 21945 15750
rect 21969 15748 22025 15750
rect 22049 15748 22105 15750
rect 21809 14714 21865 14716
rect 21889 14714 21945 14716
rect 21969 14714 22025 14716
rect 22049 14714 22105 14716
rect 21809 14662 21855 14714
rect 21855 14662 21865 14714
rect 21889 14662 21919 14714
rect 21919 14662 21931 14714
rect 21931 14662 21945 14714
rect 21969 14662 21983 14714
rect 21983 14662 21995 14714
rect 21995 14662 22025 14714
rect 22049 14662 22059 14714
rect 22059 14662 22105 14714
rect 21809 14660 21865 14662
rect 21889 14660 21945 14662
rect 21969 14660 22025 14662
rect 22049 14660 22105 14662
rect 22374 16088 22430 16144
rect 21809 13626 21865 13628
rect 21889 13626 21945 13628
rect 21969 13626 22025 13628
rect 22049 13626 22105 13628
rect 21809 13574 21855 13626
rect 21855 13574 21865 13626
rect 21889 13574 21919 13626
rect 21919 13574 21931 13626
rect 21931 13574 21945 13626
rect 21969 13574 21983 13626
rect 21983 13574 21995 13626
rect 21995 13574 22025 13626
rect 22049 13574 22059 13626
rect 22059 13574 22105 13626
rect 21809 13572 21865 13574
rect 21889 13572 21945 13574
rect 21969 13572 22025 13574
rect 22049 13572 22105 13574
rect 21809 12538 21865 12540
rect 21889 12538 21945 12540
rect 21969 12538 22025 12540
rect 22049 12538 22105 12540
rect 21809 12486 21855 12538
rect 21855 12486 21865 12538
rect 21889 12486 21919 12538
rect 21919 12486 21931 12538
rect 21931 12486 21945 12538
rect 21969 12486 21983 12538
rect 21983 12486 21995 12538
rect 21995 12486 22025 12538
rect 22049 12486 22059 12538
rect 22059 12486 22105 12538
rect 21809 12484 21865 12486
rect 21889 12484 21945 12486
rect 21969 12484 22025 12486
rect 22049 12484 22105 12486
rect 25594 20712 25650 20768
rect 23386 14592 23442 14648
rect 21809 11450 21865 11452
rect 21889 11450 21945 11452
rect 21969 11450 22025 11452
rect 22049 11450 22105 11452
rect 21809 11398 21855 11450
rect 21855 11398 21865 11450
rect 21889 11398 21919 11450
rect 21919 11398 21931 11450
rect 21931 11398 21945 11450
rect 21969 11398 21983 11450
rect 21983 11398 21995 11450
rect 21995 11398 22025 11450
rect 22049 11398 22059 11450
rect 22059 11398 22105 11450
rect 21809 11396 21865 11398
rect 21889 11396 21945 11398
rect 21969 11396 22025 11398
rect 22049 11396 22105 11398
rect 21809 10362 21865 10364
rect 21889 10362 21945 10364
rect 21969 10362 22025 10364
rect 22049 10362 22105 10364
rect 21809 10310 21855 10362
rect 21855 10310 21865 10362
rect 21889 10310 21919 10362
rect 21919 10310 21931 10362
rect 21931 10310 21945 10362
rect 21969 10310 21983 10362
rect 21983 10310 21995 10362
rect 21995 10310 22025 10362
rect 22049 10310 22059 10362
rect 22059 10310 22105 10362
rect 21809 10308 21865 10310
rect 21889 10308 21945 10310
rect 21969 10308 22025 10310
rect 22049 10308 22105 10310
rect 22098 9988 22154 10024
rect 22098 9968 22100 9988
rect 22100 9968 22152 9988
rect 22152 9968 22154 9988
rect 21362 9016 21418 9072
rect 21809 9274 21865 9276
rect 21889 9274 21945 9276
rect 21969 9274 22025 9276
rect 22049 9274 22105 9276
rect 21809 9222 21855 9274
rect 21855 9222 21865 9274
rect 21889 9222 21919 9274
rect 21919 9222 21931 9274
rect 21931 9222 21945 9274
rect 21969 9222 21983 9274
rect 21983 9222 21995 9274
rect 21995 9222 22025 9274
rect 22049 9222 22059 9274
rect 22059 9222 22105 9274
rect 21809 9220 21865 9222
rect 21889 9220 21945 9222
rect 21969 9220 22025 9222
rect 22049 9220 22105 9222
rect 22190 8336 22246 8392
rect 21809 8186 21865 8188
rect 21889 8186 21945 8188
rect 21969 8186 22025 8188
rect 22049 8186 22105 8188
rect 21809 8134 21855 8186
rect 21855 8134 21865 8186
rect 21889 8134 21919 8186
rect 21919 8134 21931 8186
rect 21931 8134 21945 8186
rect 21969 8134 21983 8186
rect 21983 8134 21995 8186
rect 21995 8134 22025 8186
rect 22049 8134 22059 8186
rect 22059 8134 22105 8186
rect 21809 8132 21865 8134
rect 21889 8132 21945 8134
rect 21969 8132 22025 8134
rect 22049 8132 22105 8134
rect 21809 7098 21865 7100
rect 21889 7098 21945 7100
rect 21969 7098 22025 7100
rect 22049 7098 22105 7100
rect 21809 7046 21855 7098
rect 21855 7046 21865 7098
rect 21889 7046 21919 7098
rect 21919 7046 21931 7098
rect 21931 7046 21945 7098
rect 21969 7046 21983 7098
rect 21983 7046 21995 7098
rect 21995 7046 22025 7098
rect 22049 7046 22059 7098
rect 22059 7046 22105 7098
rect 21809 7044 21865 7046
rect 21889 7044 21945 7046
rect 21969 7044 22025 7046
rect 22049 7044 22105 7046
rect 21809 6010 21865 6012
rect 21889 6010 21945 6012
rect 21969 6010 22025 6012
rect 22049 6010 22105 6012
rect 21809 5958 21855 6010
rect 21855 5958 21865 6010
rect 21889 5958 21919 6010
rect 21919 5958 21931 6010
rect 21931 5958 21945 6010
rect 21969 5958 21983 6010
rect 21983 5958 21995 6010
rect 21995 5958 22025 6010
rect 22049 5958 22059 6010
rect 22059 5958 22105 6010
rect 21809 5956 21865 5958
rect 21889 5956 21945 5958
rect 21969 5956 22025 5958
rect 22049 5956 22105 5958
rect 21809 4922 21865 4924
rect 21889 4922 21945 4924
rect 21969 4922 22025 4924
rect 22049 4922 22105 4924
rect 21809 4870 21855 4922
rect 21855 4870 21865 4922
rect 21889 4870 21919 4922
rect 21919 4870 21931 4922
rect 21931 4870 21945 4922
rect 21969 4870 21983 4922
rect 21983 4870 21995 4922
rect 21995 4870 22025 4922
rect 22049 4870 22059 4922
rect 22059 4870 22105 4922
rect 21809 4868 21865 4870
rect 21889 4868 21945 4870
rect 21969 4868 22025 4870
rect 22049 4868 22105 4870
rect 21809 3834 21865 3836
rect 21889 3834 21945 3836
rect 21969 3834 22025 3836
rect 22049 3834 22105 3836
rect 21809 3782 21855 3834
rect 21855 3782 21865 3834
rect 21889 3782 21919 3834
rect 21919 3782 21931 3834
rect 21931 3782 21945 3834
rect 21969 3782 21983 3834
rect 21983 3782 21995 3834
rect 21995 3782 22025 3834
rect 22049 3782 22059 3834
rect 22059 3782 22105 3834
rect 21809 3780 21865 3782
rect 21889 3780 21945 3782
rect 21969 3780 22025 3782
rect 22049 3780 22105 3782
rect 22374 3712 22430 3768
rect 17638 2202 17694 2204
rect 17718 2202 17774 2204
rect 17798 2202 17854 2204
rect 17878 2202 17934 2204
rect 17638 2150 17684 2202
rect 17684 2150 17694 2202
rect 17718 2150 17748 2202
rect 17748 2150 17760 2202
rect 17760 2150 17774 2202
rect 17798 2150 17812 2202
rect 17812 2150 17824 2202
rect 17824 2150 17854 2202
rect 17878 2150 17888 2202
rect 17888 2150 17934 2202
rect 17638 2148 17694 2150
rect 17718 2148 17774 2150
rect 17798 2148 17854 2150
rect 17878 2148 17934 2150
rect 21809 2746 21865 2748
rect 21889 2746 21945 2748
rect 21969 2746 22025 2748
rect 22049 2746 22105 2748
rect 21809 2694 21855 2746
rect 21855 2694 21865 2746
rect 21889 2694 21919 2746
rect 21919 2694 21931 2746
rect 21931 2694 21945 2746
rect 21969 2694 21983 2746
rect 21983 2694 21995 2746
rect 21995 2694 22025 2746
rect 22049 2694 22059 2746
rect 22059 2694 22105 2746
rect 21809 2692 21865 2694
rect 21889 2692 21945 2694
rect 21969 2692 22025 2694
rect 22049 2692 22105 2694
rect 22190 2216 22246 2272
rect 22650 720 22706 776
<< metal3 >>
rect 0 28568 800 28688
rect 26233 28522 26299 28525
rect 26498 28522 27298 28552
rect 26233 28520 27298 28522
rect 26233 28464 26238 28520
rect 26294 28464 27298 28520
rect 26233 28462 27298 28464
rect 26233 28459 26299 28462
rect 26498 28432 27298 28462
rect 0 27208 800 27328
rect 9285 27232 9605 27233
rect 9285 27168 9293 27232
rect 9357 27168 9373 27232
rect 9437 27168 9453 27232
rect 9517 27168 9533 27232
rect 9597 27168 9605 27232
rect 9285 27167 9605 27168
rect 17626 27232 17946 27233
rect 17626 27168 17634 27232
rect 17698 27168 17714 27232
rect 17778 27168 17794 27232
rect 17858 27168 17874 27232
rect 17938 27168 17946 27232
rect 17626 27167 17946 27168
rect 26498 26936 27298 27056
rect 5114 26688 5434 26689
rect 5114 26624 5122 26688
rect 5186 26624 5202 26688
rect 5266 26624 5282 26688
rect 5346 26624 5362 26688
rect 5426 26624 5434 26688
rect 5114 26623 5434 26624
rect 13456 26688 13776 26689
rect 13456 26624 13464 26688
rect 13528 26624 13544 26688
rect 13608 26624 13624 26688
rect 13688 26624 13704 26688
rect 13768 26624 13776 26688
rect 13456 26623 13776 26624
rect 21797 26688 22117 26689
rect 21797 26624 21805 26688
rect 21869 26624 21885 26688
rect 21949 26624 21965 26688
rect 22029 26624 22045 26688
rect 22109 26624 22117 26688
rect 21797 26623 22117 26624
rect 9285 26144 9605 26145
rect 9285 26080 9293 26144
rect 9357 26080 9373 26144
rect 9437 26080 9453 26144
rect 9517 26080 9533 26144
rect 9597 26080 9605 26144
rect 9285 26079 9605 26080
rect 17626 26144 17946 26145
rect 17626 26080 17634 26144
rect 17698 26080 17714 26144
rect 17778 26080 17794 26144
rect 17858 26080 17874 26144
rect 17938 26080 17946 26144
rect 17626 26079 17946 26080
rect 0 25848 800 25968
rect 5114 25600 5434 25601
rect 5114 25536 5122 25600
rect 5186 25536 5202 25600
rect 5266 25536 5282 25600
rect 5346 25536 5362 25600
rect 5426 25536 5434 25600
rect 5114 25535 5434 25536
rect 13456 25600 13776 25601
rect 13456 25536 13464 25600
rect 13528 25536 13544 25600
rect 13608 25536 13624 25600
rect 13688 25536 13704 25600
rect 13768 25536 13776 25600
rect 13456 25535 13776 25536
rect 21797 25600 22117 25601
rect 21797 25536 21805 25600
rect 21869 25536 21885 25600
rect 21949 25536 21965 25600
rect 22029 25536 22045 25600
rect 22109 25536 22117 25600
rect 21797 25535 22117 25536
rect 25037 25394 25103 25397
rect 26498 25394 27298 25424
rect 25037 25392 27298 25394
rect 25037 25336 25042 25392
rect 25098 25336 27298 25392
rect 25037 25334 27298 25336
rect 25037 25331 25103 25334
rect 26498 25304 27298 25334
rect 9285 25056 9605 25057
rect 9285 24992 9293 25056
rect 9357 24992 9373 25056
rect 9437 24992 9453 25056
rect 9517 24992 9533 25056
rect 9597 24992 9605 25056
rect 9285 24991 9605 24992
rect 17626 25056 17946 25057
rect 17626 24992 17634 25056
rect 17698 24992 17714 25056
rect 17778 24992 17794 25056
rect 17858 24992 17874 25056
rect 17938 24992 17946 25056
rect 17626 24991 17946 24992
rect 5114 24512 5434 24513
rect 0 24442 800 24472
rect 5114 24448 5122 24512
rect 5186 24448 5202 24512
rect 5266 24448 5282 24512
rect 5346 24448 5362 24512
rect 5426 24448 5434 24512
rect 5114 24447 5434 24448
rect 13456 24512 13776 24513
rect 13456 24448 13464 24512
rect 13528 24448 13544 24512
rect 13608 24448 13624 24512
rect 13688 24448 13704 24512
rect 13768 24448 13776 24512
rect 13456 24447 13776 24448
rect 21797 24512 22117 24513
rect 21797 24448 21805 24512
rect 21869 24448 21885 24512
rect 21949 24448 21965 24512
rect 22029 24448 22045 24512
rect 22109 24448 22117 24512
rect 21797 24447 22117 24448
rect 2129 24442 2195 24445
rect 0 24440 2195 24442
rect 0 24384 2134 24440
rect 2190 24384 2195 24440
rect 0 24382 2195 24384
rect 0 24352 800 24382
rect 2129 24379 2195 24382
rect 9285 23968 9605 23969
rect 9285 23904 9293 23968
rect 9357 23904 9373 23968
rect 9437 23904 9453 23968
rect 9517 23904 9533 23968
rect 9597 23904 9605 23968
rect 9285 23903 9605 23904
rect 17626 23968 17946 23969
rect 17626 23904 17634 23968
rect 17698 23904 17714 23968
rect 17778 23904 17794 23968
rect 17858 23904 17874 23968
rect 17938 23904 17946 23968
rect 17626 23903 17946 23904
rect 26498 23808 27298 23928
rect 8017 23762 8083 23765
rect 8293 23762 8359 23765
rect 8661 23762 8727 23765
rect 8017 23760 8727 23762
rect 8017 23704 8022 23760
rect 8078 23704 8298 23760
rect 8354 23704 8666 23760
rect 8722 23704 8727 23760
rect 8017 23702 8727 23704
rect 8017 23699 8083 23702
rect 8293 23699 8359 23702
rect 8661 23699 8727 23702
rect 5114 23424 5434 23425
rect 5114 23360 5122 23424
rect 5186 23360 5202 23424
rect 5266 23360 5282 23424
rect 5346 23360 5362 23424
rect 5426 23360 5434 23424
rect 5114 23359 5434 23360
rect 13456 23424 13776 23425
rect 13456 23360 13464 23424
rect 13528 23360 13544 23424
rect 13608 23360 13624 23424
rect 13688 23360 13704 23424
rect 13768 23360 13776 23424
rect 13456 23359 13776 23360
rect 21797 23424 22117 23425
rect 21797 23360 21805 23424
rect 21869 23360 21885 23424
rect 21949 23360 21965 23424
rect 22029 23360 22045 23424
rect 22109 23360 22117 23424
rect 21797 23359 22117 23360
rect 0 23082 800 23112
rect 2129 23082 2195 23085
rect 0 23080 2195 23082
rect 0 23024 2134 23080
rect 2190 23024 2195 23080
rect 0 23022 2195 23024
rect 0 22992 800 23022
rect 2129 23019 2195 23022
rect 9285 22880 9605 22881
rect 9285 22816 9293 22880
rect 9357 22816 9373 22880
rect 9437 22816 9453 22880
rect 9517 22816 9533 22880
rect 9597 22816 9605 22880
rect 9285 22815 9605 22816
rect 17626 22880 17946 22881
rect 17626 22816 17634 22880
rect 17698 22816 17714 22880
rect 17778 22816 17794 22880
rect 17858 22816 17874 22880
rect 17938 22816 17946 22880
rect 17626 22815 17946 22816
rect 5114 22336 5434 22337
rect 5114 22272 5122 22336
rect 5186 22272 5202 22336
rect 5266 22272 5282 22336
rect 5346 22272 5362 22336
rect 5426 22272 5434 22336
rect 5114 22271 5434 22272
rect 13456 22336 13776 22337
rect 13456 22272 13464 22336
rect 13528 22272 13544 22336
rect 13608 22272 13624 22336
rect 13688 22272 13704 22336
rect 13768 22272 13776 22336
rect 13456 22271 13776 22272
rect 21797 22336 22117 22337
rect 21797 22272 21805 22336
rect 21869 22272 21885 22336
rect 21949 22272 21965 22336
rect 22029 22272 22045 22336
rect 22109 22272 22117 22336
rect 26498 22312 27298 22432
rect 21797 22271 22117 22272
rect 11789 21994 11855 21997
rect 12065 21994 12131 21997
rect 11789 21992 12131 21994
rect 11789 21936 11794 21992
rect 11850 21936 12070 21992
rect 12126 21936 12131 21992
rect 11789 21934 12131 21936
rect 11789 21931 11855 21934
rect 12065 21931 12131 21934
rect 9285 21792 9605 21793
rect 0 21722 800 21752
rect 9285 21728 9293 21792
rect 9357 21728 9373 21792
rect 9437 21728 9453 21792
rect 9517 21728 9533 21792
rect 9597 21728 9605 21792
rect 9285 21727 9605 21728
rect 17626 21792 17946 21793
rect 17626 21728 17634 21792
rect 17698 21728 17714 21792
rect 17778 21728 17794 21792
rect 17858 21728 17874 21792
rect 17938 21728 17946 21792
rect 17626 21727 17946 21728
rect 5993 21722 6059 21725
rect 0 21720 6059 21722
rect 0 21664 5998 21720
rect 6054 21664 6059 21720
rect 0 21662 6059 21664
rect 0 21632 800 21662
rect 5993 21659 6059 21662
rect 5114 21248 5434 21249
rect 5114 21184 5122 21248
rect 5186 21184 5202 21248
rect 5266 21184 5282 21248
rect 5346 21184 5362 21248
rect 5426 21184 5434 21248
rect 5114 21183 5434 21184
rect 13456 21248 13776 21249
rect 13456 21184 13464 21248
rect 13528 21184 13544 21248
rect 13608 21184 13624 21248
rect 13688 21184 13704 21248
rect 13768 21184 13776 21248
rect 13456 21183 13776 21184
rect 21797 21248 22117 21249
rect 21797 21184 21805 21248
rect 21869 21184 21885 21248
rect 21949 21184 21965 21248
rect 22029 21184 22045 21248
rect 22109 21184 22117 21248
rect 21797 21183 22117 21184
rect 25589 20770 25655 20773
rect 26498 20770 27298 20800
rect 25589 20768 27298 20770
rect 25589 20712 25594 20768
rect 25650 20712 27298 20768
rect 25589 20710 27298 20712
rect 25589 20707 25655 20710
rect 9285 20704 9605 20705
rect 9285 20640 9293 20704
rect 9357 20640 9373 20704
rect 9437 20640 9453 20704
rect 9517 20640 9533 20704
rect 9597 20640 9605 20704
rect 9285 20639 9605 20640
rect 17626 20704 17946 20705
rect 17626 20640 17634 20704
rect 17698 20640 17714 20704
rect 17778 20640 17794 20704
rect 17858 20640 17874 20704
rect 17938 20640 17946 20704
rect 26498 20680 27298 20710
rect 17626 20639 17946 20640
rect 0 20272 800 20392
rect 11145 20362 11211 20365
rect 12893 20362 12959 20365
rect 19793 20362 19859 20365
rect 11145 20360 19859 20362
rect 11145 20304 11150 20360
rect 11206 20304 12898 20360
rect 12954 20304 19798 20360
rect 19854 20304 19859 20360
rect 11145 20302 19859 20304
rect 11145 20299 11211 20302
rect 12893 20299 12959 20302
rect 19793 20299 19859 20302
rect 5114 20160 5434 20161
rect 5114 20096 5122 20160
rect 5186 20096 5202 20160
rect 5266 20096 5282 20160
rect 5346 20096 5362 20160
rect 5426 20096 5434 20160
rect 5114 20095 5434 20096
rect 13456 20160 13776 20161
rect 13456 20096 13464 20160
rect 13528 20096 13544 20160
rect 13608 20096 13624 20160
rect 13688 20096 13704 20160
rect 13768 20096 13776 20160
rect 13456 20095 13776 20096
rect 21797 20160 22117 20161
rect 21797 20096 21805 20160
rect 21869 20096 21885 20160
rect 21949 20096 21965 20160
rect 22029 20096 22045 20160
rect 22109 20096 22117 20160
rect 21797 20095 22117 20096
rect 11513 19818 11579 19821
rect 12985 19818 13051 19821
rect 11513 19816 13051 19818
rect 11513 19760 11518 19816
rect 11574 19760 12990 19816
rect 13046 19760 13051 19816
rect 11513 19758 13051 19760
rect 11513 19755 11579 19758
rect 12985 19755 13051 19758
rect 9285 19616 9605 19617
rect 9285 19552 9293 19616
rect 9357 19552 9373 19616
rect 9437 19552 9453 19616
rect 9517 19552 9533 19616
rect 9597 19552 9605 19616
rect 9285 19551 9605 19552
rect 17626 19616 17946 19617
rect 17626 19552 17634 19616
rect 17698 19552 17714 19616
rect 17778 19552 17794 19616
rect 17858 19552 17874 19616
rect 17938 19552 17946 19616
rect 17626 19551 17946 19552
rect 11237 19410 11303 19413
rect 12341 19410 12407 19413
rect 19701 19410 19767 19413
rect 11237 19408 19767 19410
rect 11237 19352 11242 19408
rect 11298 19352 12346 19408
rect 12402 19352 19706 19408
rect 19762 19352 19767 19408
rect 11237 19350 19767 19352
rect 11237 19347 11303 19350
rect 12341 19347 12407 19350
rect 19701 19347 19767 19350
rect 26498 19184 27298 19304
rect 5114 19072 5434 19073
rect 5114 19008 5122 19072
rect 5186 19008 5202 19072
rect 5266 19008 5282 19072
rect 5346 19008 5362 19072
rect 5426 19008 5434 19072
rect 5114 19007 5434 19008
rect 13456 19072 13776 19073
rect 13456 19008 13464 19072
rect 13528 19008 13544 19072
rect 13608 19008 13624 19072
rect 13688 19008 13704 19072
rect 13768 19008 13776 19072
rect 13456 19007 13776 19008
rect 21797 19072 22117 19073
rect 21797 19008 21805 19072
rect 21869 19008 21885 19072
rect 21949 19008 21965 19072
rect 22029 19008 22045 19072
rect 22109 19008 22117 19072
rect 21797 19007 22117 19008
rect 0 18776 800 18896
rect 9285 18528 9605 18529
rect 9285 18464 9293 18528
rect 9357 18464 9373 18528
rect 9437 18464 9453 18528
rect 9517 18464 9533 18528
rect 9597 18464 9605 18528
rect 9285 18463 9605 18464
rect 17626 18528 17946 18529
rect 17626 18464 17634 18528
rect 17698 18464 17714 18528
rect 17778 18464 17794 18528
rect 17858 18464 17874 18528
rect 17938 18464 17946 18528
rect 17626 18463 17946 18464
rect 5114 17984 5434 17985
rect 5114 17920 5122 17984
rect 5186 17920 5202 17984
rect 5266 17920 5282 17984
rect 5346 17920 5362 17984
rect 5426 17920 5434 17984
rect 5114 17919 5434 17920
rect 13456 17984 13776 17985
rect 13456 17920 13464 17984
rect 13528 17920 13544 17984
rect 13608 17920 13624 17984
rect 13688 17920 13704 17984
rect 13768 17920 13776 17984
rect 13456 17919 13776 17920
rect 21797 17984 22117 17985
rect 21797 17920 21805 17984
rect 21869 17920 21885 17984
rect 21949 17920 21965 17984
rect 22029 17920 22045 17984
rect 22109 17920 22117 17984
rect 21797 17919 22117 17920
rect 23381 17778 23447 17781
rect 26498 17778 27298 17808
rect 23381 17776 27298 17778
rect 23381 17720 23386 17776
rect 23442 17720 27298 17776
rect 23381 17718 27298 17720
rect 23381 17715 23447 17718
rect 26498 17688 27298 17718
rect 0 17506 800 17536
rect 4061 17506 4127 17509
rect 0 17504 4127 17506
rect 0 17448 4066 17504
rect 4122 17448 4127 17504
rect 0 17446 4127 17448
rect 0 17416 800 17446
rect 4061 17443 4127 17446
rect 9285 17440 9605 17441
rect 9285 17376 9293 17440
rect 9357 17376 9373 17440
rect 9437 17376 9453 17440
rect 9517 17376 9533 17440
rect 9597 17376 9605 17440
rect 9285 17375 9605 17376
rect 17626 17440 17946 17441
rect 17626 17376 17634 17440
rect 17698 17376 17714 17440
rect 17778 17376 17794 17440
rect 17858 17376 17874 17440
rect 17938 17376 17946 17440
rect 17626 17375 17946 17376
rect 5114 16896 5434 16897
rect 5114 16832 5122 16896
rect 5186 16832 5202 16896
rect 5266 16832 5282 16896
rect 5346 16832 5362 16896
rect 5426 16832 5434 16896
rect 5114 16831 5434 16832
rect 13456 16896 13776 16897
rect 13456 16832 13464 16896
rect 13528 16832 13544 16896
rect 13608 16832 13624 16896
rect 13688 16832 13704 16896
rect 13768 16832 13776 16896
rect 13456 16831 13776 16832
rect 21797 16896 22117 16897
rect 21797 16832 21805 16896
rect 21869 16832 21885 16896
rect 21949 16832 21965 16896
rect 22029 16832 22045 16896
rect 22109 16832 22117 16896
rect 21797 16831 22117 16832
rect 9285 16352 9605 16353
rect 9285 16288 9293 16352
rect 9357 16288 9373 16352
rect 9437 16288 9453 16352
rect 9517 16288 9533 16352
rect 9597 16288 9605 16352
rect 9285 16287 9605 16288
rect 17626 16352 17946 16353
rect 17626 16288 17634 16352
rect 17698 16288 17714 16352
rect 17778 16288 17794 16352
rect 17858 16288 17874 16352
rect 17938 16288 17946 16352
rect 17626 16287 17946 16288
rect 0 16146 800 16176
rect 4061 16146 4127 16149
rect 0 16144 4127 16146
rect 0 16088 4066 16144
rect 4122 16088 4127 16144
rect 0 16086 4127 16088
rect 0 16056 800 16086
rect 4061 16083 4127 16086
rect 22369 16146 22435 16149
rect 26498 16146 27298 16176
rect 22369 16144 27298 16146
rect 22369 16088 22374 16144
rect 22430 16088 27298 16144
rect 22369 16086 27298 16088
rect 22369 16083 22435 16086
rect 26498 16056 27298 16086
rect 5114 15808 5434 15809
rect 5114 15744 5122 15808
rect 5186 15744 5202 15808
rect 5266 15744 5282 15808
rect 5346 15744 5362 15808
rect 5426 15744 5434 15808
rect 5114 15743 5434 15744
rect 13456 15808 13776 15809
rect 13456 15744 13464 15808
rect 13528 15744 13544 15808
rect 13608 15744 13624 15808
rect 13688 15744 13704 15808
rect 13768 15744 13776 15808
rect 13456 15743 13776 15744
rect 21797 15808 22117 15809
rect 21797 15744 21805 15808
rect 21869 15744 21885 15808
rect 21949 15744 21965 15808
rect 22029 15744 22045 15808
rect 22109 15744 22117 15808
rect 21797 15743 22117 15744
rect 12249 15466 12315 15469
rect 12617 15466 12683 15469
rect 13629 15466 13695 15469
rect 12249 15464 13695 15466
rect 12249 15408 12254 15464
rect 12310 15408 12622 15464
rect 12678 15408 13634 15464
rect 13690 15408 13695 15464
rect 12249 15406 13695 15408
rect 12249 15403 12315 15406
rect 12617 15403 12683 15406
rect 13629 15403 13695 15406
rect 9285 15264 9605 15265
rect 9285 15200 9293 15264
rect 9357 15200 9373 15264
rect 9437 15200 9453 15264
rect 9517 15200 9533 15264
rect 9597 15200 9605 15264
rect 9285 15199 9605 15200
rect 17626 15264 17946 15265
rect 17626 15200 17634 15264
rect 17698 15200 17714 15264
rect 17778 15200 17794 15264
rect 17858 15200 17874 15264
rect 17938 15200 17946 15264
rect 17626 15199 17946 15200
rect 5114 14720 5434 14721
rect 0 14650 800 14680
rect 5114 14656 5122 14720
rect 5186 14656 5202 14720
rect 5266 14656 5282 14720
rect 5346 14656 5362 14720
rect 5426 14656 5434 14720
rect 5114 14655 5434 14656
rect 13456 14720 13776 14721
rect 13456 14656 13464 14720
rect 13528 14656 13544 14720
rect 13608 14656 13624 14720
rect 13688 14656 13704 14720
rect 13768 14656 13776 14720
rect 13456 14655 13776 14656
rect 21797 14720 22117 14721
rect 21797 14656 21805 14720
rect 21869 14656 21885 14720
rect 21949 14656 21965 14720
rect 22029 14656 22045 14720
rect 22109 14656 22117 14720
rect 21797 14655 22117 14656
rect 3417 14650 3483 14653
rect 0 14648 3483 14650
rect 0 14592 3422 14648
rect 3478 14592 3483 14648
rect 0 14590 3483 14592
rect 0 14560 800 14590
rect 3417 14587 3483 14590
rect 23381 14650 23447 14653
rect 26498 14650 27298 14680
rect 23381 14648 27298 14650
rect 23381 14592 23386 14648
rect 23442 14592 27298 14648
rect 23381 14590 27298 14592
rect 23381 14587 23447 14590
rect 26498 14560 27298 14590
rect 5901 14514 5967 14517
rect 6729 14514 6795 14517
rect 5901 14512 6795 14514
rect 5901 14456 5906 14512
rect 5962 14456 6734 14512
rect 6790 14456 6795 14512
rect 5901 14454 6795 14456
rect 5901 14451 5967 14454
rect 6729 14451 6795 14454
rect 14641 14514 14707 14517
rect 15377 14514 15443 14517
rect 14641 14512 15443 14514
rect 14641 14456 14646 14512
rect 14702 14456 15382 14512
rect 15438 14456 15443 14512
rect 14641 14454 15443 14456
rect 14641 14451 14707 14454
rect 15377 14451 15443 14454
rect 9285 14176 9605 14177
rect 9285 14112 9293 14176
rect 9357 14112 9373 14176
rect 9437 14112 9453 14176
rect 9517 14112 9533 14176
rect 9597 14112 9605 14176
rect 9285 14111 9605 14112
rect 17626 14176 17946 14177
rect 17626 14112 17634 14176
rect 17698 14112 17714 14176
rect 17778 14112 17794 14176
rect 17858 14112 17874 14176
rect 17938 14112 17946 14176
rect 17626 14111 17946 14112
rect 4705 13970 4771 13973
rect 5717 13970 5783 13973
rect 9581 13970 9647 13973
rect 4705 13968 9647 13970
rect 4705 13912 4710 13968
rect 4766 13912 5722 13968
rect 5778 13912 9586 13968
rect 9642 13912 9647 13968
rect 4705 13910 9647 13912
rect 4705 13907 4771 13910
rect 5717 13907 5783 13910
rect 9581 13907 9647 13910
rect 4521 13834 4587 13837
rect 6913 13834 6979 13837
rect 4521 13832 6979 13834
rect 4521 13776 4526 13832
rect 4582 13776 6918 13832
rect 6974 13776 6979 13832
rect 4521 13774 6979 13776
rect 4521 13771 4587 13774
rect 6913 13771 6979 13774
rect 8661 13834 8727 13837
rect 9673 13834 9739 13837
rect 8661 13832 9739 13834
rect 8661 13776 8666 13832
rect 8722 13776 9678 13832
rect 9734 13776 9739 13832
rect 8661 13774 9739 13776
rect 8661 13771 8727 13774
rect 9673 13771 9739 13774
rect 5114 13632 5434 13633
rect 5114 13568 5122 13632
rect 5186 13568 5202 13632
rect 5266 13568 5282 13632
rect 5346 13568 5362 13632
rect 5426 13568 5434 13632
rect 5114 13567 5434 13568
rect 13456 13632 13776 13633
rect 13456 13568 13464 13632
rect 13528 13568 13544 13632
rect 13608 13568 13624 13632
rect 13688 13568 13704 13632
rect 13768 13568 13776 13632
rect 13456 13567 13776 13568
rect 21797 13632 22117 13633
rect 21797 13568 21805 13632
rect 21869 13568 21885 13632
rect 21949 13568 21965 13632
rect 22029 13568 22045 13632
rect 22109 13568 22117 13632
rect 21797 13567 22117 13568
rect 5441 13426 5507 13429
rect 5809 13426 5875 13429
rect 6637 13426 6703 13429
rect 5441 13424 6703 13426
rect 5441 13368 5446 13424
rect 5502 13368 5814 13424
rect 5870 13368 6642 13424
rect 6698 13368 6703 13424
rect 5441 13366 6703 13368
rect 5441 13363 5507 13366
rect 5809 13363 5875 13366
rect 6637 13363 6703 13366
rect 7097 13426 7163 13429
rect 10133 13426 10199 13429
rect 7097 13424 10199 13426
rect 7097 13368 7102 13424
rect 7158 13368 10138 13424
rect 10194 13368 10199 13424
rect 7097 13366 10199 13368
rect 7097 13363 7163 13366
rect 10133 13363 10199 13366
rect 10869 13426 10935 13429
rect 12617 13426 12683 13429
rect 10869 13424 12683 13426
rect 10869 13368 10874 13424
rect 10930 13368 12622 13424
rect 12678 13368 12683 13424
rect 10869 13366 12683 13368
rect 10869 13363 10935 13366
rect 12617 13363 12683 13366
rect 0 13290 800 13320
rect 12709 13290 12775 13293
rect 13537 13290 13603 13293
rect 0 13288 13603 13290
rect 0 13232 12714 13288
rect 12770 13232 13542 13288
rect 13598 13232 13603 13288
rect 0 13230 13603 13232
rect 0 13200 800 13230
rect 12709 13227 12775 13230
rect 13537 13227 13603 13230
rect 10317 13154 10383 13157
rect 11881 13154 11947 13157
rect 14457 13154 14523 13157
rect 10317 13152 14523 13154
rect 10317 13096 10322 13152
rect 10378 13096 11886 13152
rect 11942 13096 14462 13152
rect 14518 13096 14523 13152
rect 10317 13094 14523 13096
rect 10317 13091 10383 13094
rect 11881 13091 11947 13094
rect 14457 13091 14523 13094
rect 9285 13088 9605 13089
rect 9285 13024 9293 13088
rect 9357 13024 9373 13088
rect 9437 13024 9453 13088
rect 9517 13024 9533 13088
rect 9597 13024 9605 13088
rect 9285 13023 9605 13024
rect 17626 13088 17946 13089
rect 17626 13024 17634 13088
rect 17698 13024 17714 13088
rect 17778 13024 17794 13088
rect 17858 13024 17874 13088
rect 17938 13024 17946 13088
rect 17626 13023 17946 13024
rect 9673 13018 9739 13021
rect 12433 13018 12499 13021
rect 9673 13016 12499 13018
rect 9673 12960 9678 13016
rect 9734 12960 12438 13016
rect 12494 12960 12499 13016
rect 9673 12958 12499 12960
rect 9673 12955 9739 12958
rect 12433 12955 12499 12958
rect 26498 12928 27298 13048
rect 11605 12882 11671 12885
rect 12985 12882 13051 12885
rect 11605 12880 13051 12882
rect 11605 12824 11610 12880
rect 11666 12824 12990 12880
rect 13046 12824 13051 12880
rect 11605 12822 13051 12824
rect 11605 12819 11671 12822
rect 12985 12819 13051 12822
rect 5114 12544 5434 12545
rect 5114 12480 5122 12544
rect 5186 12480 5202 12544
rect 5266 12480 5282 12544
rect 5346 12480 5362 12544
rect 5426 12480 5434 12544
rect 5114 12479 5434 12480
rect 13456 12544 13776 12545
rect 13456 12480 13464 12544
rect 13528 12480 13544 12544
rect 13608 12480 13624 12544
rect 13688 12480 13704 12544
rect 13768 12480 13776 12544
rect 13456 12479 13776 12480
rect 21797 12544 22117 12545
rect 21797 12480 21805 12544
rect 21869 12480 21885 12544
rect 21949 12480 21965 12544
rect 22029 12480 22045 12544
rect 22109 12480 22117 12544
rect 21797 12479 22117 12480
rect 15101 12338 15167 12341
rect 15653 12338 15719 12341
rect 15101 12336 15719 12338
rect 15101 12280 15106 12336
rect 15162 12280 15658 12336
rect 15714 12280 15719 12336
rect 15101 12278 15719 12280
rect 15101 12275 15167 12278
rect 15653 12275 15719 12278
rect 9285 12000 9605 12001
rect 0 11840 800 11960
rect 9285 11936 9293 12000
rect 9357 11936 9373 12000
rect 9437 11936 9453 12000
rect 9517 11936 9533 12000
rect 9597 11936 9605 12000
rect 9285 11935 9605 11936
rect 17626 12000 17946 12001
rect 17626 11936 17634 12000
rect 17698 11936 17714 12000
rect 17778 11936 17794 12000
rect 17858 11936 17874 12000
rect 17938 11936 17946 12000
rect 17626 11935 17946 11936
rect 13997 11522 14063 11525
rect 17217 11522 17283 11525
rect 13997 11520 17283 11522
rect 13997 11464 14002 11520
rect 14058 11464 17222 11520
rect 17278 11464 17283 11520
rect 13997 11462 17283 11464
rect 13997 11459 14063 11462
rect 17217 11459 17283 11462
rect 5114 11456 5434 11457
rect 5114 11392 5122 11456
rect 5186 11392 5202 11456
rect 5266 11392 5282 11456
rect 5346 11392 5362 11456
rect 5426 11392 5434 11456
rect 5114 11391 5434 11392
rect 13456 11456 13776 11457
rect 13456 11392 13464 11456
rect 13528 11392 13544 11456
rect 13608 11392 13624 11456
rect 13688 11392 13704 11456
rect 13768 11392 13776 11456
rect 13456 11391 13776 11392
rect 21797 11456 22117 11457
rect 21797 11392 21805 11456
rect 21869 11392 21885 11456
rect 21949 11392 21965 11456
rect 22029 11392 22045 11456
rect 22109 11392 22117 11456
rect 26498 11432 27298 11552
rect 21797 11391 22117 11392
rect 5441 11250 5507 11253
rect 8293 11250 8359 11253
rect 5441 11248 8359 11250
rect 5441 11192 5446 11248
rect 5502 11192 8298 11248
rect 8354 11192 8359 11248
rect 5441 11190 8359 11192
rect 5441 11187 5507 11190
rect 8293 11187 8359 11190
rect 10225 11250 10291 11253
rect 16573 11250 16639 11253
rect 10225 11248 16639 11250
rect 10225 11192 10230 11248
rect 10286 11192 16578 11248
rect 16634 11192 16639 11248
rect 10225 11190 16639 11192
rect 10225 11187 10291 11190
rect 16573 11187 16639 11190
rect 9581 11114 9647 11117
rect 9078 11112 9647 11114
rect 9078 11056 9586 11112
rect 9642 11056 9647 11112
rect 9078 11054 9647 11056
rect 9078 10981 9138 11054
rect 9581 11051 9647 11054
rect 9029 10976 9138 10981
rect 9029 10920 9034 10976
rect 9090 10920 9138 10976
rect 9029 10918 9138 10920
rect 9029 10915 9095 10918
rect 9285 10912 9605 10913
rect 9285 10848 9293 10912
rect 9357 10848 9373 10912
rect 9437 10848 9453 10912
rect 9517 10848 9533 10912
rect 9597 10848 9605 10912
rect 9285 10847 9605 10848
rect 17626 10912 17946 10913
rect 17626 10848 17634 10912
rect 17698 10848 17714 10912
rect 17778 10848 17794 10912
rect 17858 10848 17874 10912
rect 17938 10848 17946 10912
rect 17626 10847 17946 10848
rect 4981 10706 5047 10709
rect 5993 10706 6059 10709
rect 4981 10704 6059 10706
rect 4981 10648 4986 10704
rect 5042 10648 5998 10704
rect 6054 10648 6059 10704
rect 4981 10646 6059 10648
rect 4981 10643 5047 10646
rect 5993 10643 6059 10646
rect 7557 10706 7623 10709
rect 14641 10706 14707 10709
rect 7557 10704 14707 10706
rect 7557 10648 7562 10704
rect 7618 10648 14646 10704
rect 14702 10648 14707 10704
rect 7557 10646 14707 10648
rect 7557 10643 7623 10646
rect 14641 10643 14707 10646
rect 0 10570 800 10600
rect 6913 10570 6979 10573
rect 0 10568 6979 10570
rect 0 10512 6918 10568
rect 6974 10512 6979 10568
rect 0 10510 6979 10512
rect 0 10480 800 10510
rect 6913 10507 6979 10510
rect 5114 10368 5434 10369
rect 5114 10304 5122 10368
rect 5186 10304 5202 10368
rect 5266 10304 5282 10368
rect 5346 10304 5362 10368
rect 5426 10304 5434 10368
rect 5114 10303 5434 10304
rect 13456 10368 13776 10369
rect 13456 10304 13464 10368
rect 13528 10304 13544 10368
rect 13608 10304 13624 10368
rect 13688 10304 13704 10368
rect 13768 10304 13776 10368
rect 13456 10303 13776 10304
rect 21797 10368 22117 10369
rect 21797 10304 21805 10368
rect 21869 10304 21885 10368
rect 21949 10304 21965 10368
rect 22029 10304 22045 10368
rect 22109 10304 22117 10368
rect 21797 10303 22117 10304
rect 8017 10026 8083 10029
rect 9765 10026 9831 10029
rect 8017 10024 9831 10026
rect 8017 9968 8022 10024
rect 8078 9968 9770 10024
rect 9826 9968 9831 10024
rect 8017 9966 9831 9968
rect 8017 9963 8083 9966
rect 9765 9963 9831 9966
rect 22093 10026 22159 10029
rect 26498 10026 27298 10056
rect 22093 10024 27298 10026
rect 22093 9968 22098 10024
rect 22154 9968 27298 10024
rect 22093 9966 27298 9968
rect 22093 9963 22159 9966
rect 26498 9936 27298 9966
rect 9285 9824 9605 9825
rect 9285 9760 9293 9824
rect 9357 9760 9373 9824
rect 9437 9760 9453 9824
rect 9517 9760 9533 9824
rect 9597 9760 9605 9824
rect 9285 9759 9605 9760
rect 17626 9824 17946 9825
rect 17626 9760 17634 9824
rect 17698 9760 17714 9824
rect 17778 9760 17794 9824
rect 17858 9760 17874 9824
rect 17938 9760 17946 9824
rect 17626 9759 17946 9760
rect 3049 9754 3115 9757
rect 7833 9754 7899 9757
rect 8201 9754 8267 9757
rect 3049 9752 8267 9754
rect 3049 9696 3054 9752
rect 3110 9696 7838 9752
rect 7894 9696 8206 9752
rect 8262 9696 8267 9752
rect 3049 9694 8267 9696
rect 3049 9691 3115 9694
rect 7833 9691 7899 9694
rect 8201 9691 8267 9694
rect 5114 9280 5434 9281
rect 5114 9216 5122 9280
rect 5186 9216 5202 9280
rect 5266 9216 5282 9280
rect 5346 9216 5362 9280
rect 5426 9216 5434 9280
rect 5114 9215 5434 9216
rect 13456 9280 13776 9281
rect 13456 9216 13464 9280
rect 13528 9216 13544 9280
rect 13608 9216 13624 9280
rect 13688 9216 13704 9280
rect 13768 9216 13776 9280
rect 13456 9215 13776 9216
rect 21797 9280 22117 9281
rect 21797 9216 21805 9280
rect 21869 9216 21885 9280
rect 21949 9216 21965 9280
rect 22029 9216 22045 9280
rect 22109 9216 22117 9280
rect 21797 9215 22117 9216
rect 20069 9210 20135 9213
rect 20897 9210 20963 9213
rect 20069 9208 20963 9210
rect 20069 9152 20074 9208
rect 20130 9152 20902 9208
rect 20958 9152 20963 9208
rect 20069 9150 20963 9152
rect 20069 9147 20135 9150
rect 20897 9147 20963 9150
rect 0 9074 800 9104
rect 3969 9074 4035 9077
rect 0 9072 4035 9074
rect 0 9016 3974 9072
rect 4030 9016 4035 9072
rect 0 9014 4035 9016
rect 0 8984 800 9014
rect 3969 9011 4035 9014
rect 20253 9074 20319 9077
rect 21357 9074 21423 9077
rect 20253 9072 21423 9074
rect 20253 9016 20258 9072
rect 20314 9016 21362 9072
rect 21418 9016 21423 9072
rect 20253 9014 21423 9016
rect 20253 9011 20319 9014
rect 21357 9011 21423 9014
rect 9285 8736 9605 8737
rect 9285 8672 9293 8736
rect 9357 8672 9373 8736
rect 9437 8672 9453 8736
rect 9517 8672 9533 8736
rect 9597 8672 9605 8736
rect 9285 8671 9605 8672
rect 17626 8736 17946 8737
rect 17626 8672 17634 8736
rect 17698 8672 17714 8736
rect 17778 8672 17794 8736
rect 17858 8672 17874 8736
rect 17938 8672 17946 8736
rect 17626 8671 17946 8672
rect 11145 8530 11211 8533
rect 12709 8530 12775 8533
rect 11145 8528 12775 8530
rect 11145 8472 11150 8528
rect 11206 8472 12714 8528
rect 12770 8472 12775 8528
rect 11145 8470 12775 8472
rect 11145 8467 11211 8470
rect 12709 8467 12775 8470
rect 22185 8394 22251 8397
rect 26498 8394 27298 8424
rect 22185 8392 27298 8394
rect 22185 8336 22190 8392
rect 22246 8336 27298 8392
rect 22185 8334 27298 8336
rect 22185 8331 22251 8334
rect 26498 8304 27298 8334
rect 5114 8192 5434 8193
rect 5114 8128 5122 8192
rect 5186 8128 5202 8192
rect 5266 8128 5282 8192
rect 5346 8128 5362 8192
rect 5426 8128 5434 8192
rect 5114 8127 5434 8128
rect 13456 8192 13776 8193
rect 13456 8128 13464 8192
rect 13528 8128 13544 8192
rect 13608 8128 13624 8192
rect 13688 8128 13704 8192
rect 13768 8128 13776 8192
rect 13456 8127 13776 8128
rect 21797 8192 22117 8193
rect 21797 8128 21805 8192
rect 21869 8128 21885 8192
rect 21949 8128 21965 8192
rect 22029 8128 22045 8192
rect 22109 8128 22117 8192
rect 21797 8127 22117 8128
rect 0 7624 800 7744
rect 9285 7648 9605 7649
rect 9285 7584 9293 7648
rect 9357 7584 9373 7648
rect 9437 7584 9453 7648
rect 9517 7584 9533 7648
rect 9597 7584 9605 7648
rect 9285 7583 9605 7584
rect 17626 7648 17946 7649
rect 17626 7584 17634 7648
rect 17698 7584 17714 7648
rect 17778 7584 17794 7648
rect 17858 7584 17874 7648
rect 17938 7584 17946 7648
rect 17626 7583 17946 7584
rect 5114 7104 5434 7105
rect 5114 7040 5122 7104
rect 5186 7040 5202 7104
rect 5266 7040 5282 7104
rect 5346 7040 5362 7104
rect 5426 7040 5434 7104
rect 5114 7039 5434 7040
rect 13456 7104 13776 7105
rect 13456 7040 13464 7104
rect 13528 7040 13544 7104
rect 13608 7040 13624 7104
rect 13688 7040 13704 7104
rect 13768 7040 13776 7104
rect 13456 7039 13776 7040
rect 21797 7104 22117 7105
rect 21797 7040 21805 7104
rect 21869 7040 21885 7104
rect 21949 7040 21965 7104
rect 22029 7040 22045 7104
rect 22109 7040 22117 7104
rect 21797 7039 22117 7040
rect 26498 6808 27298 6928
rect 9285 6560 9605 6561
rect 9285 6496 9293 6560
rect 9357 6496 9373 6560
rect 9437 6496 9453 6560
rect 9517 6496 9533 6560
rect 9597 6496 9605 6560
rect 9285 6495 9605 6496
rect 17626 6560 17946 6561
rect 17626 6496 17634 6560
rect 17698 6496 17714 6560
rect 17778 6496 17794 6560
rect 17858 6496 17874 6560
rect 17938 6496 17946 6560
rect 17626 6495 17946 6496
rect 0 6354 800 6384
rect 4061 6354 4127 6357
rect 0 6352 4127 6354
rect 0 6296 4066 6352
rect 4122 6296 4127 6352
rect 0 6294 4127 6296
rect 0 6264 800 6294
rect 4061 6291 4127 6294
rect 5114 6016 5434 6017
rect 5114 5952 5122 6016
rect 5186 5952 5202 6016
rect 5266 5952 5282 6016
rect 5346 5952 5362 6016
rect 5426 5952 5434 6016
rect 5114 5951 5434 5952
rect 13456 6016 13776 6017
rect 13456 5952 13464 6016
rect 13528 5952 13544 6016
rect 13608 5952 13624 6016
rect 13688 5952 13704 6016
rect 13768 5952 13776 6016
rect 13456 5951 13776 5952
rect 21797 6016 22117 6017
rect 21797 5952 21805 6016
rect 21869 5952 21885 6016
rect 21949 5952 21965 6016
rect 22029 5952 22045 6016
rect 22109 5952 22117 6016
rect 21797 5951 22117 5952
rect 9285 5472 9605 5473
rect 9285 5408 9293 5472
rect 9357 5408 9373 5472
rect 9437 5408 9453 5472
rect 9517 5408 9533 5472
rect 9597 5408 9605 5472
rect 9285 5407 9605 5408
rect 17626 5472 17946 5473
rect 17626 5408 17634 5472
rect 17698 5408 17714 5472
rect 17778 5408 17794 5472
rect 17858 5408 17874 5472
rect 17938 5408 17946 5472
rect 17626 5407 17946 5408
rect 26498 5312 27298 5432
rect 5114 4928 5434 4929
rect 0 4858 800 4888
rect 5114 4864 5122 4928
rect 5186 4864 5202 4928
rect 5266 4864 5282 4928
rect 5346 4864 5362 4928
rect 5426 4864 5434 4928
rect 5114 4863 5434 4864
rect 13456 4928 13776 4929
rect 13456 4864 13464 4928
rect 13528 4864 13544 4928
rect 13608 4864 13624 4928
rect 13688 4864 13704 4928
rect 13768 4864 13776 4928
rect 13456 4863 13776 4864
rect 21797 4928 22117 4929
rect 21797 4864 21805 4928
rect 21869 4864 21885 4928
rect 21949 4864 21965 4928
rect 22029 4864 22045 4928
rect 22109 4864 22117 4928
rect 21797 4863 22117 4864
rect 3509 4858 3575 4861
rect 0 4856 3575 4858
rect 0 4800 3514 4856
rect 3570 4800 3575 4856
rect 0 4798 3575 4800
rect 0 4768 800 4798
rect 3509 4795 3575 4798
rect 9285 4384 9605 4385
rect 9285 4320 9293 4384
rect 9357 4320 9373 4384
rect 9437 4320 9453 4384
rect 9517 4320 9533 4384
rect 9597 4320 9605 4384
rect 9285 4319 9605 4320
rect 17626 4384 17946 4385
rect 17626 4320 17634 4384
rect 17698 4320 17714 4384
rect 17778 4320 17794 4384
rect 17858 4320 17874 4384
rect 17938 4320 17946 4384
rect 17626 4319 17946 4320
rect 5114 3840 5434 3841
rect 5114 3776 5122 3840
rect 5186 3776 5202 3840
rect 5266 3776 5282 3840
rect 5346 3776 5362 3840
rect 5426 3776 5434 3840
rect 5114 3775 5434 3776
rect 13456 3840 13776 3841
rect 13456 3776 13464 3840
rect 13528 3776 13544 3840
rect 13608 3776 13624 3840
rect 13688 3776 13704 3840
rect 13768 3776 13776 3840
rect 13456 3775 13776 3776
rect 21797 3840 22117 3841
rect 21797 3776 21805 3840
rect 21869 3776 21885 3840
rect 21949 3776 21965 3840
rect 22029 3776 22045 3840
rect 22109 3776 22117 3840
rect 21797 3775 22117 3776
rect 22369 3770 22435 3773
rect 26498 3770 27298 3800
rect 22369 3768 27298 3770
rect 22369 3712 22374 3768
rect 22430 3712 27298 3768
rect 22369 3710 27298 3712
rect 22369 3707 22435 3710
rect 26498 3680 27298 3710
rect 0 3498 800 3528
rect 2037 3498 2103 3501
rect 0 3496 2103 3498
rect 0 3440 2042 3496
rect 2098 3440 2103 3496
rect 0 3438 2103 3440
rect 0 3408 800 3438
rect 2037 3435 2103 3438
rect 9285 3296 9605 3297
rect 9285 3232 9293 3296
rect 9357 3232 9373 3296
rect 9437 3232 9453 3296
rect 9517 3232 9533 3296
rect 9597 3232 9605 3296
rect 9285 3231 9605 3232
rect 17626 3296 17946 3297
rect 17626 3232 17634 3296
rect 17698 3232 17714 3296
rect 17778 3232 17794 3296
rect 17858 3232 17874 3296
rect 17938 3232 17946 3296
rect 17626 3231 17946 3232
rect 5114 2752 5434 2753
rect 5114 2688 5122 2752
rect 5186 2688 5202 2752
rect 5266 2688 5282 2752
rect 5346 2688 5362 2752
rect 5426 2688 5434 2752
rect 5114 2687 5434 2688
rect 13456 2752 13776 2753
rect 13456 2688 13464 2752
rect 13528 2688 13544 2752
rect 13608 2688 13624 2752
rect 13688 2688 13704 2752
rect 13768 2688 13776 2752
rect 13456 2687 13776 2688
rect 21797 2752 22117 2753
rect 21797 2688 21805 2752
rect 21869 2688 21885 2752
rect 21949 2688 21965 2752
rect 22029 2688 22045 2752
rect 22109 2688 22117 2752
rect 21797 2687 22117 2688
rect 22185 2274 22251 2277
rect 26498 2274 27298 2304
rect 22185 2272 27298 2274
rect 22185 2216 22190 2272
rect 22246 2216 27298 2272
rect 22185 2214 27298 2216
rect 22185 2211 22251 2214
rect 9285 2208 9605 2209
rect 0 2138 800 2168
rect 9285 2144 9293 2208
rect 9357 2144 9373 2208
rect 9437 2144 9453 2208
rect 9517 2144 9533 2208
rect 9597 2144 9605 2208
rect 9285 2143 9605 2144
rect 17626 2208 17946 2209
rect 17626 2144 17634 2208
rect 17698 2144 17714 2208
rect 17778 2144 17794 2208
rect 17858 2144 17874 2208
rect 17938 2144 17946 2208
rect 26498 2184 27298 2214
rect 17626 2143 17946 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 0 2048 800 2078
rect 2773 2075 2839 2078
rect 0 778 800 808
rect 3141 778 3207 781
rect 0 776 3207 778
rect 0 720 3146 776
rect 3202 720 3207 776
rect 0 718 3207 720
rect 0 688 800 718
rect 3141 715 3207 718
rect 22645 778 22711 781
rect 26498 778 27298 808
rect 22645 776 27298 778
rect 22645 720 22650 776
rect 22706 720 27298 776
rect 22645 718 27298 720
rect 22645 715 22711 718
rect 26498 688 27298 718
<< via3 >>
rect 9293 27228 9357 27232
rect 9293 27172 9297 27228
rect 9297 27172 9353 27228
rect 9353 27172 9357 27228
rect 9293 27168 9357 27172
rect 9373 27228 9437 27232
rect 9373 27172 9377 27228
rect 9377 27172 9433 27228
rect 9433 27172 9437 27228
rect 9373 27168 9437 27172
rect 9453 27228 9517 27232
rect 9453 27172 9457 27228
rect 9457 27172 9513 27228
rect 9513 27172 9517 27228
rect 9453 27168 9517 27172
rect 9533 27228 9597 27232
rect 9533 27172 9537 27228
rect 9537 27172 9593 27228
rect 9593 27172 9597 27228
rect 9533 27168 9597 27172
rect 17634 27228 17698 27232
rect 17634 27172 17638 27228
rect 17638 27172 17694 27228
rect 17694 27172 17698 27228
rect 17634 27168 17698 27172
rect 17714 27228 17778 27232
rect 17714 27172 17718 27228
rect 17718 27172 17774 27228
rect 17774 27172 17778 27228
rect 17714 27168 17778 27172
rect 17794 27228 17858 27232
rect 17794 27172 17798 27228
rect 17798 27172 17854 27228
rect 17854 27172 17858 27228
rect 17794 27168 17858 27172
rect 17874 27228 17938 27232
rect 17874 27172 17878 27228
rect 17878 27172 17934 27228
rect 17934 27172 17938 27228
rect 17874 27168 17938 27172
rect 5122 26684 5186 26688
rect 5122 26628 5126 26684
rect 5126 26628 5182 26684
rect 5182 26628 5186 26684
rect 5122 26624 5186 26628
rect 5202 26684 5266 26688
rect 5202 26628 5206 26684
rect 5206 26628 5262 26684
rect 5262 26628 5266 26684
rect 5202 26624 5266 26628
rect 5282 26684 5346 26688
rect 5282 26628 5286 26684
rect 5286 26628 5342 26684
rect 5342 26628 5346 26684
rect 5282 26624 5346 26628
rect 5362 26684 5426 26688
rect 5362 26628 5366 26684
rect 5366 26628 5422 26684
rect 5422 26628 5426 26684
rect 5362 26624 5426 26628
rect 13464 26684 13528 26688
rect 13464 26628 13468 26684
rect 13468 26628 13524 26684
rect 13524 26628 13528 26684
rect 13464 26624 13528 26628
rect 13544 26684 13608 26688
rect 13544 26628 13548 26684
rect 13548 26628 13604 26684
rect 13604 26628 13608 26684
rect 13544 26624 13608 26628
rect 13624 26684 13688 26688
rect 13624 26628 13628 26684
rect 13628 26628 13684 26684
rect 13684 26628 13688 26684
rect 13624 26624 13688 26628
rect 13704 26684 13768 26688
rect 13704 26628 13708 26684
rect 13708 26628 13764 26684
rect 13764 26628 13768 26684
rect 13704 26624 13768 26628
rect 21805 26684 21869 26688
rect 21805 26628 21809 26684
rect 21809 26628 21865 26684
rect 21865 26628 21869 26684
rect 21805 26624 21869 26628
rect 21885 26684 21949 26688
rect 21885 26628 21889 26684
rect 21889 26628 21945 26684
rect 21945 26628 21949 26684
rect 21885 26624 21949 26628
rect 21965 26684 22029 26688
rect 21965 26628 21969 26684
rect 21969 26628 22025 26684
rect 22025 26628 22029 26684
rect 21965 26624 22029 26628
rect 22045 26684 22109 26688
rect 22045 26628 22049 26684
rect 22049 26628 22105 26684
rect 22105 26628 22109 26684
rect 22045 26624 22109 26628
rect 9293 26140 9357 26144
rect 9293 26084 9297 26140
rect 9297 26084 9353 26140
rect 9353 26084 9357 26140
rect 9293 26080 9357 26084
rect 9373 26140 9437 26144
rect 9373 26084 9377 26140
rect 9377 26084 9433 26140
rect 9433 26084 9437 26140
rect 9373 26080 9437 26084
rect 9453 26140 9517 26144
rect 9453 26084 9457 26140
rect 9457 26084 9513 26140
rect 9513 26084 9517 26140
rect 9453 26080 9517 26084
rect 9533 26140 9597 26144
rect 9533 26084 9537 26140
rect 9537 26084 9593 26140
rect 9593 26084 9597 26140
rect 9533 26080 9597 26084
rect 17634 26140 17698 26144
rect 17634 26084 17638 26140
rect 17638 26084 17694 26140
rect 17694 26084 17698 26140
rect 17634 26080 17698 26084
rect 17714 26140 17778 26144
rect 17714 26084 17718 26140
rect 17718 26084 17774 26140
rect 17774 26084 17778 26140
rect 17714 26080 17778 26084
rect 17794 26140 17858 26144
rect 17794 26084 17798 26140
rect 17798 26084 17854 26140
rect 17854 26084 17858 26140
rect 17794 26080 17858 26084
rect 17874 26140 17938 26144
rect 17874 26084 17878 26140
rect 17878 26084 17934 26140
rect 17934 26084 17938 26140
rect 17874 26080 17938 26084
rect 5122 25596 5186 25600
rect 5122 25540 5126 25596
rect 5126 25540 5182 25596
rect 5182 25540 5186 25596
rect 5122 25536 5186 25540
rect 5202 25596 5266 25600
rect 5202 25540 5206 25596
rect 5206 25540 5262 25596
rect 5262 25540 5266 25596
rect 5202 25536 5266 25540
rect 5282 25596 5346 25600
rect 5282 25540 5286 25596
rect 5286 25540 5342 25596
rect 5342 25540 5346 25596
rect 5282 25536 5346 25540
rect 5362 25596 5426 25600
rect 5362 25540 5366 25596
rect 5366 25540 5422 25596
rect 5422 25540 5426 25596
rect 5362 25536 5426 25540
rect 13464 25596 13528 25600
rect 13464 25540 13468 25596
rect 13468 25540 13524 25596
rect 13524 25540 13528 25596
rect 13464 25536 13528 25540
rect 13544 25596 13608 25600
rect 13544 25540 13548 25596
rect 13548 25540 13604 25596
rect 13604 25540 13608 25596
rect 13544 25536 13608 25540
rect 13624 25596 13688 25600
rect 13624 25540 13628 25596
rect 13628 25540 13684 25596
rect 13684 25540 13688 25596
rect 13624 25536 13688 25540
rect 13704 25596 13768 25600
rect 13704 25540 13708 25596
rect 13708 25540 13764 25596
rect 13764 25540 13768 25596
rect 13704 25536 13768 25540
rect 21805 25596 21869 25600
rect 21805 25540 21809 25596
rect 21809 25540 21865 25596
rect 21865 25540 21869 25596
rect 21805 25536 21869 25540
rect 21885 25596 21949 25600
rect 21885 25540 21889 25596
rect 21889 25540 21945 25596
rect 21945 25540 21949 25596
rect 21885 25536 21949 25540
rect 21965 25596 22029 25600
rect 21965 25540 21969 25596
rect 21969 25540 22025 25596
rect 22025 25540 22029 25596
rect 21965 25536 22029 25540
rect 22045 25596 22109 25600
rect 22045 25540 22049 25596
rect 22049 25540 22105 25596
rect 22105 25540 22109 25596
rect 22045 25536 22109 25540
rect 9293 25052 9357 25056
rect 9293 24996 9297 25052
rect 9297 24996 9353 25052
rect 9353 24996 9357 25052
rect 9293 24992 9357 24996
rect 9373 25052 9437 25056
rect 9373 24996 9377 25052
rect 9377 24996 9433 25052
rect 9433 24996 9437 25052
rect 9373 24992 9437 24996
rect 9453 25052 9517 25056
rect 9453 24996 9457 25052
rect 9457 24996 9513 25052
rect 9513 24996 9517 25052
rect 9453 24992 9517 24996
rect 9533 25052 9597 25056
rect 9533 24996 9537 25052
rect 9537 24996 9593 25052
rect 9593 24996 9597 25052
rect 9533 24992 9597 24996
rect 17634 25052 17698 25056
rect 17634 24996 17638 25052
rect 17638 24996 17694 25052
rect 17694 24996 17698 25052
rect 17634 24992 17698 24996
rect 17714 25052 17778 25056
rect 17714 24996 17718 25052
rect 17718 24996 17774 25052
rect 17774 24996 17778 25052
rect 17714 24992 17778 24996
rect 17794 25052 17858 25056
rect 17794 24996 17798 25052
rect 17798 24996 17854 25052
rect 17854 24996 17858 25052
rect 17794 24992 17858 24996
rect 17874 25052 17938 25056
rect 17874 24996 17878 25052
rect 17878 24996 17934 25052
rect 17934 24996 17938 25052
rect 17874 24992 17938 24996
rect 5122 24508 5186 24512
rect 5122 24452 5126 24508
rect 5126 24452 5182 24508
rect 5182 24452 5186 24508
rect 5122 24448 5186 24452
rect 5202 24508 5266 24512
rect 5202 24452 5206 24508
rect 5206 24452 5262 24508
rect 5262 24452 5266 24508
rect 5202 24448 5266 24452
rect 5282 24508 5346 24512
rect 5282 24452 5286 24508
rect 5286 24452 5342 24508
rect 5342 24452 5346 24508
rect 5282 24448 5346 24452
rect 5362 24508 5426 24512
rect 5362 24452 5366 24508
rect 5366 24452 5422 24508
rect 5422 24452 5426 24508
rect 5362 24448 5426 24452
rect 13464 24508 13528 24512
rect 13464 24452 13468 24508
rect 13468 24452 13524 24508
rect 13524 24452 13528 24508
rect 13464 24448 13528 24452
rect 13544 24508 13608 24512
rect 13544 24452 13548 24508
rect 13548 24452 13604 24508
rect 13604 24452 13608 24508
rect 13544 24448 13608 24452
rect 13624 24508 13688 24512
rect 13624 24452 13628 24508
rect 13628 24452 13684 24508
rect 13684 24452 13688 24508
rect 13624 24448 13688 24452
rect 13704 24508 13768 24512
rect 13704 24452 13708 24508
rect 13708 24452 13764 24508
rect 13764 24452 13768 24508
rect 13704 24448 13768 24452
rect 21805 24508 21869 24512
rect 21805 24452 21809 24508
rect 21809 24452 21865 24508
rect 21865 24452 21869 24508
rect 21805 24448 21869 24452
rect 21885 24508 21949 24512
rect 21885 24452 21889 24508
rect 21889 24452 21945 24508
rect 21945 24452 21949 24508
rect 21885 24448 21949 24452
rect 21965 24508 22029 24512
rect 21965 24452 21969 24508
rect 21969 24452 22025 24508
rect 22025 24452 22029 24508
rect 21965 24448 22029 24452
rect 22045 24508 22109 24512
rect 22045 24452 22049 24508
rect 22049 24452 22105 24508
rect 22105 24452 22109 24508
rect 22045 24448 22109 24452
rect 9293 23964 9357 23968
rect 9293 23908 9297 23964
rect 9297 23908 9353 23964
rect 9353 23908 9357 23964
rect 9293 23904 9357 23908
rect 9373 23964 9437 23968
rect 9373 23908 9377 23964
rect 9377 23908 9433 23964
rect 9433 23908 9437 23964
rect 9373 23904 9437 23908
rect 9453 23964 9517 23968
rect 9453 23908 9457 23964
rect 9457 23908 9513 23964
rect 9513 23908 9517 23964
rect 9453 23904 9517 23908
rect 9533 23964 9597 23968
rect 9533 23908 9537 23964
rect 9537 23908 9593 23964
rect 9593 23908 9597 23964
rect 9533 23904 9597 23908
rect 17634 23964 17698 23968
rect 17634 23908 17638 23964
rect 17638 23908 17694 23964
rect 17694 23908 17698 23964
rect 17634 23904 17698 23908
rect 17714 23964 17778 23968
rect 17714 23908 17718 23964
rect 17718 23908 17774 23964
rect 17774 23908 17778 23964
rect 17714 23904 17778 23908
rect 17794 23964 17858 23968
rect 17794 23908 17798 23964
rect 17798 23908 17854 23964
rect 17854 23908 17858 23964
rect 17794 23904 17858 23908
rect 17874 23964 17938 23968
rect 17874 23908 17878 23964
rect 17878 23908 17934 23964
rect 17934 23908 17938 23964
rect 17874 23904 17938 23908
rect 5122 23420 5186 23424
rect 5122 23364 5126 23420
rect 5126 23364 5182 23420
rect 5182 23364 5186 23420
rect 5122 23360 5186 23364
rect 5202 23420 5266 23424
rect 5202 23364 5206 23420
rect 5206 23364 5262 23420
rect 5262 23364 5266 23420
rect 5202 23360 5266 23364
rect 5282 23420 5346 23424
rect 5282 23364 5286 23420
rect 5286 23364 5342 23420
rect 5342 23364 5346 23420
rect 5282 23360 5346 23364
rect 5362 23420 5426 23424
rect 5362 23364 5366 23420
rect 5366 23364 5422 23420
rect 5422 23364 5426 23420
rect 5362 23360 5426 23364
rect 13464 23420 13528 23424
rect 13464 23364 13468 23420
rect 13468 23364 13524 23420
rect 13524 23364 13528 23420
rect 13464 23360 13528 23364
rect 13544 23420 13608 23424
rect 13544 23364 13548 23420
rect 13548 23364 13604 23420
rect 13604 23364 13608 23420
rect 13544 23360 13608 23364
rect 13624 23420 13688 23424
rect 13624 23364 13628 23420
rect 13628 23364 13684 23420
rect 13684 23364 13688 23420
rect 13624 23360 13688 23364
rect 13704 23420 13768 23424
rect 13704 23364 13708 23420
rect 13708 23364 13764 23420
rect 13764 23364 13768 23420
rect 13704 23360 13768 23364
rect 21805 23420 21869 23424
rect 21805 23364 21809 23420
rect 21809 23364 21865 23420
rect 21865 23364 21869 23420
rect 21805 23360 21869 23364
rect 21885 23420 21949 23424
rect 21885 23364 21889 23420
rect 21889 23364 21945 23420
rect 21945 23364 21949 23420
rect 21885 23360 21949 23364
rect 21965 23420 22029 23424
rect 21965 23364 21969 23420
rect 21969 23364 22025 23420
rect 22025 23364 22029 23420
rect 21965 23360 22029 23364
rect 22045 23420 22109 23424
rect 22045 23364 22049 23420
rect 22049 23364 22105 23420
rect 22105 23364 22109 23420
rect 22045 23360 22109 23364
rect 9293 22876 9357 22880
rect 9293 22820 9297 22876
rect 9297 22820 9353 22876
rect 9353 22820 9357 22876
rect 9293 22816 9357 22820
rect 9373 22876 9437 22880
rect 9373 22820 9377 22876
rect 9377 22820 9433 22876
rect 9433 22820 9437 22876
rect 9373 22816 9437 22820
rect 9453 22876 9517 22880
rect 9453 22820 9457 22876
rect 9457 22820 9513 22876
rect 9513 22820 9517 22876
rect 9453 22816 9517 22820
rect 9533 22876 9597 22880
rect 9533 22820 9537 22876
rect 9537 22820 9593 22876
rect 9593 22820 9597 22876
rect 9533 22816 9597 22820
rect 17634 22876 17698 22880
rect 17634 22820 17638 22876
rect 17638 22820 17694 22876
rect 17694 22820 17698 22876
rect 17634 22816 17698 22820
rect 17714 22876 17778 22880
rect 17714 22820 17718 22876
rect 17718 22820 17774 22876
rect 17774 22820 17778 22876
rect 17714 22816 17778 22820
rect 17794 22876 17858 22880
rect 17794 22820 17798 22876
rect 17798 22820 17854 22876
rect 17854 22820 17858 22876
rect 17794 22816 17858 22820
rect 17874 22876 17938 22880
rect 17874 22820 17878 22876
rect 17878 22820 17934 22876
rect 17934 22820 17938 22876
rect 17874 22816 17938 22820
rect 5122 22332 5186 22336
rect 5122 22276 5126 22332
rect 5126 22276 5182 22332
rect 5182 22276 5186 22332
rect 5122 22272 5186 22276
rect 5202 22332 5266 22336
rect 5202 22276 5206 22332
rect 5206 22276 5262 22332
rect 5262 22276 5266 22332
rect 5202 22272 5266 22276
rect 5282 22332 5346 22336
rect 5282 22276 5286 22332
rect 5286 22276 5342 22332
rect 5342 22276 5346 22332
rect 5282 22272 5346 22276
rect 5362 22332 5426 22336
rect 5362 22276 5366 22332
rect 5366 22276 5422 22332
rect 5422 22276 5426 22332
rect 5362 22272 5426 22276
rect 13464 22332 13528 22336
rect 13464 22276 13468 22332
rect 13468 22276 13524 22332
rect 13524 22276 13528 22332
rect 13464 22272 13528 22276
rect 13544 22332 13608 22336
rect 13544 22276 13548 22332
rect 13548 22276 13604 22332
rect 13604 22276 13608 22332
rect 13544 22272 13608 22276
rect 13624 22332 13688 22336
rect 13624 22276 13628 22332
rect 13628 22276 13684 22332
rect 13684 22276 13688 22332
rect 13624 22272 13688 22276
rect 13704 22332 13768 22336
rect 13704 22276 13708 22332
rect 13708 22276 13764 22332
rect 13764 22276 13768 22332
rect 13704 22272 13768 22276
rect 21805 22332 21869 22336
rect 21805 22276 21809 22332
rect 21809 22276 21865 22332
rect 21865 22276 21869 22332
rect 21805 22272 21869 22276
rect 21885 22332 21949 22336
rect 21885 22276 21889 22332
rect 21889 22276 21945 22332
rect 21945 22276 21949 22332
rect 21885 22272 21949 22276
rect 21965 22332 22029 22336
rect 21965 22276 21969 22332
rect 21969 22276 22025 22332
rect 22025 22276 22029 22332
rect 21965 22272 22029 22276
rect 22045 22332 22109 22336
rect 22045 22276 22049 22332
rect 22049 22276 22105 22332
rect 22105 22276 22109 22332
rect 22045 22272 22109 22276
rect 9293 21788 9357 21792
rect 9293 21732 9297 21788
rect 9297 21732 9353 21788
rect 9353 21732 9357 21788
rect 9293 21728 9357 21732
rect 9373 21788 9437 21792
rect 9373 21732 9377 21788
rect 9377 21732 9433 21788
rect 9433 21732 9437 21788
rect 9373 21728 9437 21732
rect 9453 21788 9517 21792
rect 9453 21732 9457 21788
rect 9457 21732 9513 21788
rect 9513 21732 9517 21788
rect 9453 21728 9517 21732
rect 9533 21788 9597 21792
rect 9533 21732 9537 21788
rect 9537 21732 9593 21788
rect 9593 21732 9597 21788
rect 9533 21728 9597 21732
rect 17634 21788 17698 21792
rect 17634 21732 17638 21788
rect 17638 21732 17694 21788
rect 17694 21732 17698 21788
rect 17634 21728 17698 21732
rect 17714 21788 17778 21792
rect 17714 21732 17718 21788
rect 17718 21732 17774 21788
rect 17774 21732 17778 21788
rect 17714 21728 17778 21732
rect 17794 21788 17858 21792
rect 17794 21732 17798 21788
rect 17798 21732 17854 21788
rect 17854 21732 17858 21788
rect 17794 21728 17858 21732
rect 17874 21788 17938 21792
rect 17874 21732 17878 21788
rect 17878 21732 17934 21788
rect 17934 21732 17938 21788
rect 17874 21728 17938 21732
rect 5122 21244 5186 21248
rect 5122 21188 5126 21244
rect 5126 21188 5182 21244
rect 5182 21188 5186 21244
rect 5122 21184 5186 21188
rect 5202 21244 5266 21248
rect 5202 21188 5206 21244
rect 5206 21188 5262 21244
rect 5262 21188 5266 21244
rect 5202 21184 5266 21188
rect 5282 21244 5346 21248
rect 5282 21188 5286 21244
rect 5286 21188 5342 21244
rect 5342 21188 5346 21244
rect 5282 21184 5346 21188
rect 5362 21244 5426 21248
rect 5362 21188 5366 21244
rect 5366 21188 5422 21244
rect 5422 21188 5426 21244
rect 5362 21184 5426 21188
rect 13464 21244 13528 21248
rect 13464 21188 13468 21244
rect 13468 21188 13524 21244
rect 13524 21188 13528 21244
rect 13464 21184 13528 21188
rect 13544 21244 13608 21248
rect 13544 21188 13548 21244
rect 13548 21188 13604 21244
rect 13604 21188 13608 21244
rect 13544 21184 13608 21188
rect 13624 21244 13688 21248
rect 13624 21188 13628 21244
rect 13628 21188 13684 21244
rect 13684 21188 13688 21244
rect 13624 21184 13688 21188
rect 13704 21244 13768 21248
rect 13704 21188 13708 21244
rect 13708 21188 13764 21244
rect 13764 21188 13768 21244
rect 13704 21184 13768 21188
rect 21805 21244 21869 21248
rect 21805 21188 21809 21244
rect 21809 21188 21865 21244
rect 21865 21188 21869 21244
rect 21805 21184 21869 21188
rect 21885 21244 21949 21248
rect 21885 21188 21889 21244
rect 21889 21188 21945 21244
rect 21945 21188 21949 21244
rect 21885 21184 21949 21188
rect 21965 21244 22029 21248
rect 21965 21188 21969 21244
rect 21969 21188 22025 21244
rect 22025 21188 22029 21244
rect 21965 21184 22029 21188
rect 22045 21244 22109 21248
rect 22045 21188 22049 21244
rect 22049 21188 22105 21244
rect 22105 21188 22109 21244
rect 22045 21184 22109 21188
rect 9293 20700 9357 20704
rect 9293 20644 9297 20700
rect 9297 20644 9353 20700
rect 9353 20644 9357 20700
rect 9293 20640 9357 20644
rect 9373 20700 9437 20704
rect 9373 20644 9377 20700
rect 9377 20644 9433 20700
rect 9433 20644 9437 20700
rect 9373 20640 9437 20644
rect 9453 20700 9517 20704
rect 9453 20644 9457 20700
rect 9457 20644 9513 20700
rect 9513 20644 9517 20700
rect 9453 20640 9517 20644
rect 9533 20700 9597 20704
rect 9533 20644 9537 20700
rect 9537 20644 9593 20700
rect 9593 20644 9597 20700
rect 9533 20640 9597 20644
rect 17634 20700 17698 20704
rect 17634 20644 17638 20700
rect 17638 20644 17694 20700
rect 17694 20644 17698 20700
rect 17634 20640 17698 20644
rect 17714 20700 17778 20704
rect 17714 20644 17718 20700
rect 17718 20644 17774 20700
rect 17774 20644 17778 20700
rect 17714 20640 17778 20644
rect 17794 20700 17858 20704
rect 17794 20644 17798 20700
rect 17798 20644 17854 20700
rect 17854 20644 17858 20700
rect 17794 20640 17858 20644
rect 17874 20700 17938 20704
rect 17874 20644 17878 20700
rect 17878 20644 17934 20700
rect 17934 20644 17938 20700
rect 17874 20640 17938 20644
rect 5122 20156 5186 20160
rect 5122 20100 5126 20156
rect 5126 20100 5182 20156
rect 5182 20100 5186 20156
rect 5122 20096 5186 20100
rect 5202 20156 5266 20160
rect 5202 20100 5206 20156
rect 5206 20100 5262 20156
rect 5262 20100 5266 20156
rect 5202 20096 5266 20100
rect 5282 20156 5346 20160
rect 5282 20100 5286 20156
rect 5286 20100 5342 20156
rect 5342 20100 5346 20156
rect 5282 20096 5346 20100
rect 5362 20156 5426 20160
rect 5362 20100 5366 20156
rect 5366 20100 5422 20156
rect 5422 20100 5426 20156
rect 5362 20096 5426 20100
rect 13464 20156 13528 20160
rect 13464 20100 13468 20156
rect 13468 20100 13524 20156
rect 13524 20100 13528 20156
rect 13464 20096 13528 20100
rect 13544 20156 13608 20160
rect 13544 20100 13548 20156
rect 13548 20100 13604 20156
rect 13604 20100 13608 20156
rect 13544 20096 13608 20100
rect 13624 20156 13688 20160
rect 13624 20100 13628 20156
rect 13628 20100 13684 20156
rect 13684 20100 13688 20156
rect 13624 20096 13688 20100
rect 13704 20156 13768 20160
rect 13704 20100 13708 20156
rect 13708 20100 13764 20156
rect 13764 20100 13768 20156
rect 13704 20096 13768 20100
rect 21805 20156 21869 20160
rect 21805 20100 21809 20156
rect 21809 20100 21865 20156
rect 21865 20100 21869 20156
rect 21805 20096 21869 20100
rect 21885 20156 21949 20160
rect 21885 20100 21889 20156
rect 21889 20100 21945 20156
rect 21945 20100 21949 20156
rect 21885 20096 21949 20100
rect 21965 20156 22029 20160
rect 21965 20100 21969 20156
rect 21969 20100 22025 20156
rect 22025 20100 22029 20156
rect 21965 20096 22029 20100
rect 22045 20156 22109 20160
rect 22045 20100 22049 20156
rect 22049 20100 22105 20156
rect 22105 20100 22109 20156
rect 22045 20096 22109 20100
rect 9293 19612 9357 19616
rect 9293 19556 9297 19612
rect 9297 19556 9353 19612
rect 9353 19556 9357 19612
rect 9293 19552 9357 19556
rect 9373 19612 9437 19616
rect 9373 19556 9377 19612
rect 9377 19556 9433 19612
rect 9433 19556 9437 19612
rect 9373 19552 9437 19556
rect 9453 19612 9517 19616
rect 9453 19556 9457 19612
rect 9457 19556 9513 19612
rect 9513 19556 9517 19612
rect 9453 19552 9517 19556
rect 9533 19612 9597 19616
rect 9533 19556 9537 19612
rect 9537 19556 9593 19612
rect 9593 19556 9597 19612
rect 9533 19552 9597 19556
rect 17634 19612 17698 19616
rect 17634 19556 17638 19612
rect 17638 19556 17694 19612
rect 17694 19556 17698 19612
rect 17634 19552 17698 19556
rect 17714 19612 17778 19616
rect 17714 19556 17718 19612
rect 17718 19556 17774 19612
rect 17774 19556 17778 19612
rect 17714 19552 17778 19556
rect 17794 19612 17858 19616
rect 17794 19556 17798 19612
rect 17798 19556 17854 19612
rect 17854 19556 17858 19612
rect 17794 19552 17858 19556
rect 17874 19612 17938 19616
rect 17874 19556 17878 19612
rect 17878 19556 17934 19612
rect 17934 19556 17938 19612
rect 17874 19552 17938 19556
rect 5122 19068 5186 19072
rect 5122 19012 5126 19068
rect 5126 19012 5182 19068
rect 5182 19012 5186 19068
rect 5122 19008 5186 19012
rect 5202 19068 5266 19072
rect 5202 19012 5206 19068
rect 5206 19012 5262 19068
rect 5262 19012 5266 19068
rect 5202 19008 5266 19012
rect 5282 19068 5346 19072
rect 5282 19012 5286 19068
rect 5286 19012 5342 19068
rect 5342 19012 5346 19068
rect 5282 19008 5346 19012
rect 5362 19068 5426 19072
rect 5362 19012 5366 19068
rect 5366 19012 5422 19068
rect 5422 19012 5426 19068
rect 5362 19008 5426 19012
rect 13464 19068 13528 19072
rect 13464 19012 13468 19068
rect 13468 19012 13524 19068
rect 13524 19012 13528 19068
rect 13464 19008 13528 19012
rect 13544 19068 13608 19072
rect 13544 19012 13548 19068
rect 13548 19012 13604 19068
rect 13604 19012 13608 19068
rect 13544 19008 13608 19012
rect 13624 19068 13688 19072
rect 13624 19012 13628 19068
rect 13628 19012 13684 19068
rect 13684 19012 13688 19068
rect 13624 19008 13688 19012
rect 13704 19068 13768 19072
rect 13704 19012 13708 19068
rect 13708 19012 13764 19068
rect 13764 19012 13768 19068
rect 13704 19008 13768 19012
rect 21805 19068 21869 19072
rect 21805 19012 21809 19068
rect 21809 19012 21865 19068
rect 21865 19012 21869 19068
rect 21805 19008 21869 19012
rect 21885 19068 21949 19072
rect 21885 19012 21889 19068
rect 21889 19012 21945 19068
rect 21945 19012 21949 19068
rect 21885 19008 21949 19012
rect 21965 19068 22029 19072
rect 21965 19012 21969 19068
rect 21969 19012 22025 19068
rect 22025 19012 22029 19068
rect 21965 19008 22029 19012
rect 22045 19068 22109 19072
rect 22045 19012 22049 19068
rect 22049 19012 22105 19068
rect 22105 19012 22109 19068
rect 22045 19008 22109 19012
rect 9293 18524 9357 18528
rect 9293 18468 9297 18524
rect 9297 18468 9353 18524
rect 9353 18468 9357 18524
rect 9293 18464 9357 18468
rect 9373 18524 9437 18528
rect 9373 18468 9377 18524
rect 9377 18468 9433 18524
rect 9433 18468 9437 18524
rect 9373 18464 9437 18468
rect 9453 18524 9517 18528
rect 9453 18468 9457 18524
rect 9457 18468 9513 18524
rect 9513 18468 9517 18524
rect 9453 18464 9517 18468
rect 9533 18524 9597 18528
rect 9533 18468 9537 18524
rect 9537 18468 9593 18524
rect 9593 18468 9597 18524
rect 9533 18464 9597 18468
rect 17634 18524 17698 18528
rect 17634 18468 17638 18524
rect 17638 18468 17694 18524
rect 17694 18468 17698 18524
rect 17634 18464 17698 18468
rect 17714 18524 17778 18528
rect 17714 18468 17718 18524
rect 17718 18468 17774 18524
rect 17774 18468 17778 18524
rect 17714 18464 17778 18468
rect 17794 18524 17858 18528
rect 17794 18468 17798 18524
rect 17798 18468 17854 18524
rect 17854 18468 17858 18524
rect 17794 18464 17858 18468
rect 17874 18524 17938 18528
rect 17874 18468 17878 18524
rect 17878 18468 17934 18524
rect 17934 18468 17938 18524
rect 17874 18464 17938 18468
rect 5122 17980 5186 17984
rect 5122 17924 5126 17980
rect 5126 17924 5182 17980
rect 5182 17924 5186 17980
rect 5122 17920 5186 17924
rect 5202 17980 5266 17984
rect 5202 17924 5206 17980
rect 5206 17924 5262 17980
rect 5262 17924 5266 17980
rect 5202 17920 5266 17924
rect 5282 17980 5346 17984
rect 5282 17924 5286 17980
rect 5286 17924 5342 17980
rect 5342 17924 5346 17980
rect 5282 17920 5346 17924
rect 5362 17980 5426 17984
rect 5362 17924 5366 17980
rect 5366 17924 5422 17980
rect 5422 17924 5426 17980
rect 5362 17920 5426 17924
rect 13464 17980 13528 17984
rect 13464 17924 13468 17980
rect 13468 17924 13524 17980
rect 13524 17924 13528 17980
rect 13464 17920 13528 17924
rect 13544 17980 13608 17984
rect 13544 17924 13548 17980
rect 13548 17924 13604 17980
rect 13604 17924 13608 17980
rect 13544 17920 13608 17924
rect 13624 17980 13688 17984
rect 13624 17924 13628 17980
rect 13628 17924 13684 17980
rect 13684 17924 13688 17980
rect 13624 17920 13688 17924
rect 13704 17980 13768 17984
rect 13704 17924 13708 17980
rect 13708 17924 13764 17980
rect 13764 17924 13768 17980
rect 13704 17920 13768 17924
rect 21805 17980 21869 17984
rect 21805 17924 21809 17980
rect 21809 17924 21865 17980
rect 21865 17924 21869 17980
rect 21805 17920 21869 17924
rect 21885 17980 21949 17984
rect 21885 17924 21889 17980
rect 21889 17924 21945 17980
rect 21945 17924 21949 17980
rect 21885 17920 21949 17924
rect 21965 17980 22029 17984
rect 21965 17924 21969 17980
rect 21969 17924 22025 17980
rect 22025 17924 22029 17980
rect 21965 17920 22029 17924
rect 22045 17980 22109 17984
rect 22045 17924 22049 17980
rect 22049 17924 22105 17980
rect 22105 17924 22109 17980
rect 22045 17920 22109 17924
rect 9293 17436 9357 17440
rect 9293 17380 9297 17436
rect 9297 17380 9353 17436
rect 9353 17380 9357 17436
rect 9293 17376 9357 17380
rect 9373 17436 9437 17440
rect 9373 17380 9377 17436
rect 9377 17380 9433 17436
rect 9433 17380 9437 17436
rect 9373 17376 9437 17380
rect 9453 17436 9517 17440
rect 9453 17380 9457 17436
rect 9457 17380 9513 17436
rect 9513 17380 9517 17436
rect 9453 17376 9517 17380
rect 9533 17436 9597 17440
rect 9533 17380 9537 17436
rect 9537 17380 9593 17436
rect 9593 17380 9597 17436
rect 9533 17376 9597 17380
rect 17634 17436 17698 17440
rect 17634 17380 17638 17436
rect 17638 17380 17694 17436
rect 17694 17380 17698 17436
rect 17634 17376 17698 17380
rect 17714 17436 17778 17440
rect 17714 17380 17718 17436
rect 17718 17380 17774 17436
rect 17774 17380 17778 17436
rect 17714 17376 17778 17380
rect 17794 17436 17858 17440
rect 17794 17380 17798 17436
rect 17798 17380 17854 17436
rect 17854 17380 17858 17436
rect 17794 17376 17858 17380
rect 17874 17436 17938 17440
rect 17874 17380 17878 17436
rect 17878 17380 17934 17436
rect 17934 17380 17938 17436
rect 17874 17376 17938 17380
rect 5122 16892 5186 16896
rect 5122 16836 5126 16892
rect 5126 16836 5182 16892
rect 5182 16836 5186 16892
rect 5122 16832 5186 16836
rect 5202 16892 5266 16896
rect 5202 16836 5206 16892
rect 5206 16836 5262 16892
rect 5262 16836 5266 16892
rect 5202 16832 5266 16836
rect 5282 16892 5346 16896
rect 5282 16836 5286 16892
rect 5286 16836 5342 16892
rect 5342 16836 5346 16892
rect 5282 16832 5346 16836
rect 5362 16892 5426 16896
rect 5362 16836 5366 16892
rect 5366 16836 5422 16892
rect 5422 16836 5426 16892
rect 5362 16832 5426 16836
rect 13464 16892 13528 16896
rect 13464 16836 13468 16892
rect 13468 16836 13524 16892
rect 13524 16836 13528 16892
rect 13464 16832 13528 16836
rect 13544 16892 13608 16896
rect 13544 16836 13548 16892
rect 13548 16836 13604 16892
rect 13604 16836 13608 16892
rect 13544 16832 13608 16836
rect 13624 16892 13688 16896
rect 13624 16836 13628 16892
rect 13628 16836 13684 16892
rect 13684 16836 13688 16892
rect 13624 16832 13688 16836
rect 13704 16892 13768 16896
rect 13704 16836 13708 16892
rect 13708 16836 13764 16892
rect 13764 16836 13768 16892
rect 13704 16832 13768 16836
rect 21805 16892 21869 16896
rect 21805 16836 21809 16892
rect 21809 16836 21865 16892
rect 21865 16836 21869 16892
rect 21805 16832 21869 16836
rect 21885 16892 21949 16896
rect 21885 16836 21889 16892
rect 21889 16836 21945 16892
rect 21945 16836 21949 16892
rect 21885 16832 21949 16836
rect 21965 16892 22029 16896
rect 21965 16836 21969 16892
rect 21969 16836 22025 16892
rect 22025 16836 22029 16892
rect 21965 16832 22029 16836
rect 22045 16892 22109 16896
rect 22045 16836 22049 16892
rect 22049 16836 22105 16892
rect 22105 16836 22109 16892
rect 22045 16832 22109 16836
rect 9293 16348 9357 16352
rect 9293 16292 9297 16348
rect 9297 16292 9353 16348
rect 9353 16292 9357 16348
rect 9293 16288 9357 16292
rect 9373 16348 9437 16352
rect 9373 16292 9377 16348
rect 9377 16292 9433 16348
rect 9433 16292 9437 16348
rect 9373 16288 9437 16292
rect 9453 16348 9517 16352
rect 9453 16292 9457 16348
rect 9457 16292 9513 16348
rect 9513 16292 9517 16348
rect 9453 16288 9517 16292
rect 9533 16348 9597 16352
rect 9533 16292 9537 16348
rect 9537 16292 9593 16348
rect 9593 16292 9597 16348
rect 9533 16288 9597 16292
rect 17634 16348 17698 16352
rect 17634 16292 17638 16348
rect 17638 16292 17694 16348
rect 17694 16292 17698 16348
rect 17634 16288 17698 16292
rect 17714 16348 17778 16352
rect 17714 16292 17718 16348
rect 17718 16292 17774 16348
rect 17774 16292 17778 16348
rect 17714 16288 17778 16292
rect 17794 16348 17858 16352
rect 17794 16292 17798 16348
rect 17798 16292 17854 16348
rect 17854 16292 17858 16348
rect 17794 16288 17858 16292
rect 17874 16348 17938 16352
rect 17874 16292 17878 16348
rect 17878 16292 17934 16348
rect 17934 16292 17938 16348
rect 17874 16288 17938 16292
rect 5122 15804 5186 15808
rect 5122 15748 5126 15804
rect 5126 15748 5182 15804
rect 5182 15748 5186 15804
rect 5122 15744 5186 15748
rect 5202 15804 5266 15808
rect 5202 15748 5206 15804
rect 5206 15748 5262 15804
rect 5262 15748 5266 15804
rect 5202 15744 5266 15748
rect 5282 15804 5346 15808
rect 5282 15748 5286 15804
rect 5286 15748 5342 15804
rect 5342 15748 5346 15804
rect 5282 15744 5346 15748
rect 5362 15804 5426 15808
rect 5362 15748 5366 15804
rect 5366 15748 5422 15804
rect 5422 15748 5426 15804
rect 5362 15744 5426 15748
rect 13464 15804 13528 15808
rect 13464 15748 13468 15804
rect 13468 15748 13524 15804
rect 13524 15748 13528 15804
rect 13464 15744 13528 15748
rect 13544 15804 13608 15808
rect 13544 15748 13548 15804
rect 13548 15748 13604 15804
rect 13604 15748 13608 15804
rect 13544 15744 13608 15748
rect 13624 15804 13688 15808
rect 13624 15748 13628 15804
rect 13628 15748 13684 15804
rect 13684 15748 13688 15804
rect 13624 15744 13688 15748
rect 13704 15804 13768 15808
rect 13704 15748 13708 15804
rect 13708 15748 13764 15804
rect 13764 15748 13768 15804
rect 13704 15744 13768 15748
rect 21805 15804 21869 15808
rect 21805 15748 21809 15804
rect 21809 15748 21865 15804
rect 21865 15748 21869 15804
rect 21805 15744 21869 15748
rect 21885 15804 21949 15808
rect 21885 15748 21889 15804
rect 21889 15748 21945 15804
rect 21945 15748 21949 15804
rect 21885 15744 21949 15748
rect 21965 15804 22029 15808
rect 21965 15748 21969 15804
rect 21969 15748 22025 15804
rect 22025 15748 22029 15804
rect 21965 15744 22029 15748
rect 22045 15804 22109 15808
rect 22045 15748 22049 15804
rect 22049 15748 22105 15804
rect 22105 15748 22109 15804
rect 22045 15744 22109 15748
rect 9293 15260 9357 15264
rect 9293 15204 9297 15260
rect 9297 15204 9353 15260
rect 9353 15204 9357 15260
rect 9293 15200 9357 15204
rect 9373 15260 9437 15264
rect 9373 15204 9377 15260
rect 9377 15204 9433 15260
rect 9433 15204 9437 15260
rect 9373 15200 9437 15204
rect 9453 15260 9517 15264
rect 9453 15204 9457 15260
rect 9457 15204 9513 15260
rect 9513 15204 9517 15260
rect 9453 15200 9517 15204
rect 9533 15260 9597 15264
rect 9533 15204 9537 15260
rect 9537 15204 9593 15260
rect 9593 15204 9597 15260
rect 9533 15200 9597 15204
rect 17634 15260 17698 15264
rect 17634 15204 17638 15260
rect 17638 15204 17694 15260
rect 17694 15204 17698 15260
rect 17634 15200 17698 15204
rect 17714 15260 17778 15264
rect 17714 15204 17718 15260
rect 17718 15204 17774 15260
rect 17774 15204 17778 15260
rect 17714 15200 17778 15204
rect 17794 15260 17858 15264
rect 17794 15204 17798 15260
rect 17798 15204 17854 15260
rect 17854 15204 17858 15260
rect 17794 15200 17858 15204
rect 17874 15260 17938 15264
rect 17874 15204 17878 15260
rect 17878 15204 17934 15260
rect 17934 15204 17938 15260
rect 17874 15200 17938 15204
rect 5122 14716 5186 14720
rect 5122 14660 5126 14716
rect 5126 14660 5182 14716
rect 5182 14660 5186 14716
rect 5122 14656 5186 14660
rect 5202 14716 5266 14720
rect 5202 14660 5206 14716
rect 5206 14660 5262 14716
rect 5262 14660 5266 14716
rect 5202 14656 5266 14660
rect 5282 14716 5346 14720
rect 5282 14660 5286 14716
rect 5286 14660 5342 14716
rect 5342 14660 5346 14716
rect 5282 14656 5346 14660
rect 5362 14716 5426 14720
rect 5362 14660 5366 14716
rect 5366 14660 5422 14716
rect 5422 14660 5426 14716
rect 5362 14656 5426 14660
rect 13464 14716 13528 14720
rect 13464 14660 13468 14716
rect 13468 14660 13524 14716
rect 13524 14660 13528 14716
rect 13464 14656 13528 14660
rect 13544 14716 13608 14720
rect 13544 14660 13548 14716
rect 13548 14660 13604 14716
rect 13604 14660 13608 14716
rect 13544 14656 13608 14660
rect 13624 14716 13688 14720
rect 13624 14660 13628 14716
rect 13628 14660 13684 14716
rect 13684 14660 13688 14716
rect 13624 14656 13688 14660
rect 13704 14716 13768 14720
rect 13704 14660 13708 14716
rect 13708 14660 13764 14716
rect 13764 14660 13768 14716
rect 13704 14656 13768 14660
rect 21805 14716 21869 14720
rect 21805 14660 21809 14716
rect 21809 14660 21865 14716
rect 21865 14660 21869 14716
rect 21805 14656 21869 14660
rect 21885 14716 21949 14720
rect 21885 14660 21889 14716
rect 21889 14660 21945 14716
rect 21945 14660 21949 14716
rect 21885 14656 21949 14660
rect 21965 14716 22029 14720
rect 21965 14660 21969 14716
rect 21969 14660 22025 14716
rect 22025 14660 22029 14716
rect 21965 14656 22029 14660
rect 22045 14716 22109 14720
rect 22045 14660 22049 14716
rect 22049 14660 22105 14716
rect 22105 14660 22109 14716
rect 22045 14656 22109 14660
rect 9293 14172 9357 14176
rect 9293 14116 9297 14172
rect 9297 14116 9353 14172
rect 9353 14116 9357 14172
rect 9293 14112 9357 14116
rect 9373 14172 9437 14176
rect 9373 14116 9377 14172
rect 9377 14116 9433 14172
rect 9433 14116 9437 14172
rect 9373 14112 9437 14116
rect 9453 14172 9517 14176
rect 9453 14116 9457 14172
rect 9457 14116 9513 14172
rect 9513 14116 9517 14172
rect 9453 14112 9517 14116
rect 9533 14172 9597 14176
rect 9533 14116 9537 14172
rect 9537 14116 9593 14172
rect 9593 14116 9597 14172
rect 9533 14112 9597 14116
rect 17634 14172 17698 14176
rect 17634 14116 17638 14172
rect 17638 14116 17694 14172
rect 17694 14116 17698 14172
rect 17634 14112 17698 14116
rect 17714 14172 17778 14176
rect 17714 14116 17718 14172
rect 17718 14116 17774 14172
rect 17774 14116 17778 14172
rect 17714 14112 17778 14116
rect 17794 14172 17858 14176
rect 17794 14116 17798 14172
rect 17798 14116 17854 14172
rect 17854 14116 17858 14172
rect 17794 14112 17858 14116
rect 17874 14172 17938 14176
rect 17874 14116 17878 14172
rect 17878 14116 17934 14172
rect 17934 14116 17938 14172
rect 17874 14112 17938 14116
rect 5122 13628 5186 13632
rect 5122 13572 5126 13628
rect 5126 13572 5182 13628
rect 5182 13572 5186 13628
rect 5122 13568 5186 13572
rect 5202 13628 5266 13632
rect 5202 13572 5206 13628
rect 5206 13572 5262 13628
rect 5262 13572 5266 13628
rect 5202 13568 5266 13572
rect 5282 13628 5346 13632
rect 5282 13572 5286 13628
rect 5286 13572 5342 13628
rect 5342 13572 5346 13628
rect 5282 13568 5346 13572
rect 5362 13628 5426 13632
rect 5362 13572 5366 13628
rect 5366 13572 5422 13628
rect 5422 13572 5426 13628
rect 5362 13568 5426 13572
rect 13464 13628 13528 13632
rect 13464 13572 13468 13628
rect 13468 13572 13524 13628
rect 13524 13572 13528 13628
rect 13464 13568 13528 13572
rect 13544 13628 13608 13632
rect 13544 13572 13548 13628
rect 13548 13572 13604 13628
rect 13604 13572 13608 13628
rect 13544 13568 13608 13572
rect 13624 13628 13688 13632
rect 13624 13572 13628 13628
rect 13628 13572 13684 13628
rect 13684 13572 13688 13628
rect 13624 13568 13688 13572
rect 13704 13628 13768 13632
rect 13704 13572 13708 13628
rect 13708 13572 13764 13628
rect 13764 13572 13768 13628
rect 13704 13568 13768 13572
rect 21805 13628 21869 13632
rect 21805 13572 21809 13628
rect 21809 13572 21865 13628
rect 21865 13572 21869 13628
rect 21805 13568 21869 13572
rect 21885 13628 21949 13632
rect 21885 13572 21889 13628
rect 21889 13572 21945 13628
rect 21945 13572 21949 13628
rect 21885 13568 21949 13572
rect 21965 13628 22029 13632
rect 21965 13572 21969 13628
rect 21969 13572 22025 13628
rect 22025 13572 22029 13628
rect 21965 13568 22029 13572
rect 22045 13628 22109 13632
rect 22045 13572 22049 13628
rect 22049 13572 22105 13628
rect 22105 13572 22109 13628
rect 22045 13568 22109 13572
rect 9293 13084 9357 13088
rect 9293 13028 9297 13084
rect 9297 13028 9353 13084
rect 9353 13028 9357 13084
rect 9293 13024 9357 13028
rect 9373 13084 9437 13088
rect 9373 13028 9377 13084
rect 9377 13028 9433 13084
rect 9433 13028 9437 13084
rect 9373 13024 9437 13028
rect 9453 13084 9517 13088
rect 9453 13028 9457 13084
rect 9457 13028 9513 13084
rect 9513 13028 9517 13084
rect 9453 13024 9517 13028
rect 9533 13084 9597 13088
rect 9533 13028 9537 13084
rect 9537 13028 9593 13084
rect 9593 13028 9597 13084
rect 9533 13024 9597 13028
rect 17634 13084 17698 13088
rect 17634 13028 17638 13084
rect 17638 13028 17694 13084
rect 17694 13028 17698 13084
rect 17634 13024 17698 13028
rect 17714 13084 17778 13088
rect 17714 13028 17718 13084
rect 17718 13028 17774 13084
rect 17774 13028 17778 13084
rect 17714 13024 17778 13028
rect 17794 13084 17858 13088
rect 17794 13028 17798 13084
rect 17798 13028 17854 13084
rect 17854 13028 17858 13084
rect 17794 13024 17858 13028
rect 17874 13084 17938 13088
rect 17874 13028 17878 13084
rect 17878 13028 17934 13084
rect 17934 13028 17938 13084
rect 17874 13024 17938 13028
rect 5122 12540 5186 12544
rect 5122 12484 5126 12540
rect 5126 12484 5182 12540
rect 5182 12484 5186 12540
rect 5122 12480 5186 12484
rect 5202 12540 5266 12544
rect 5202 12484 5206 12540
rect 5206 12484 5262 12540
rect 5262 12484 5266 12540
rect 5202 12480 5266 12484
rect 5282 12540 5346 12544
rect 5282 12484 5286 12540
rect 5286 12484 5342 12540
rect 5342 12484 5346 12540
rect 5282 12480 5346 12484
rect 5362 12540 5426 12544
rect 5362 12484 5366 12540
rect 5366 12484 5422 12540
rect 5422 12484 5426 12540
rect 5362 12480 5426 12484
rect 13464 12540 13528 12544
rect 13464 12484 13468 12540
rect 13468 12484 13524 12540
rect 13524 12484 13528 12540
rect 13464 12480 13528 12484
rect 13544 12540 13608 12544
rect 13544 12484 13548 12540
rect 13548 12484 13604 12540
rect 13604 12484 13608 12540
rect 13544 12480 13608 12484
rect 13624 12540 13688 12544
rect 13624 12484 13628 12540
rect 13628 12484 13684 12540
rect 13684 12484 13688 12540
rect 13624 12480 13688 12484
rect 13704 12540 13768 12544
rect 13704 12484 13708 12540
rect 13708 12484 13764 12540
rect 13764 12484 13768 12540
rect 13704 12480 13768 12484
rect 21805 12540 21869 12544
rect 21805 12484 21809 12540
rect 21809 12484 21865 12540
rect 21865 12484 21869 12540
rect 21805 12480 21869 12484
rect 21885 12540 21949 12544
rect 21885 12484 21889 12540
rect 21889 12484 21945 12540
rect 21945 12484 21949 12540
rect 21885 12480 21949 12484
rect 21965 12540 22029 12544
rect 21965 12484 21969 12540
rect 21969 12484 22025 12540
rect 22025 12484 22029 12540
rect 21965 12480 22029 12484
rect 22045 12540 22109 12544
rect 22045 12484 22049 12540
rect 22049 12484 22105 12540
rect 22105 12484 22109 12540
rect 22045 12480 22109 12484
rect 9293 11996 9357 12000
rect 9293 11940 9297 11996
rect 9297 11940 9353 11996
rect 9353 11940 9357 11996
rect 9293 11936 9357 11940
rect 9373 11996 9437 12000
rect 9373 11940 9377 11996
rect 9377 11940 9433 11996
rect 9433 11940 9437 11996
rect 9373 11936 9437 11940
rect 9453 11996 9517 12000
rect 9453 11940 9457 11996
rect 9457 11940 9513 11996
rect 9513 11940 9517 11996
rect 9453 11936 9517 11940
rect 9533 11996 9597 12000
rect 9533 11940 9537 11996
rect 9537 11940 9593 11996
rect 9593 11940 9597 11996
rect 9533 11936 9597 11940
rect 17634 11996 17698 12000
rect 17634 11940 17638 11996
rect 17638 11940 17694 11996
rect 17694 11940 17698 11996
rect 17634 11936 17698 11940
rect 17714 11996 17778 12000
rect 17714 11940 17718 11996
rect 17718 11940 17774 11996
rect 17774 11940 17778 11996
rect 17714 11936 17778 11940
rect 17794 11996 17858 12000
rect 17794 11940 17798 11996
rect 17798 11940 17854 11996
rect 17854 11940 17858 11996
rect 17794 11936 17858 11940
rect 17874 11996 17938 12000
rect 17874 11940 17878 11996
rect 17878 11940 17934 11996
rect 17934 11940 17938 11996
rect 17874 11936 17938 11940
rect 5122 11452 5186 11456
rect 5122 11396 5126 11452
rect 5126 11396 5182 11452
rect 5182 11396 5186 11452
rect 5122 11392 5186 11396
rect 5202 11452 5266 11456
rect 5202 11396 5206 11452
rect 5206 11396 5262 11452
rect 5262 11396 5266 11452
rect 5202 11392 5266 11396
rect 5282 11452 5346 11456
rect 5282 11396 5286 11452
rect 5286 11396 5342 11452
rect 5342 11396 5346 11452
rect 5282 11392 5346 11396
rect 5362 11452 5426 11456
rect 5362 11396 5366 11452
rect 5366 11396 5422 11452
rect 5422 11396 5426 11452
rect 5362 11392 5426 11396
rect 13464 11452 13528 11456
rect 13464 11396 13468 11452
rect 13468 11396 13524 11452
rect 13524 11396 13528 11452
rect 13464 11392 13528 11396
rect 13544 11452 13608 11456
rect 13544 11396 13548 11452
rect 13548 11396 13604 11452
rect 13604 11396 13608 11452
rect 13544 11392 13608 11396
rect 13624 11452 13688 11456
rect 13624 11396 13628 11452
rect 13628 11396 13684 11452
rect 13684 11396 13688 11452
rect 13624 11392 13688 11396
rect 13704 11452 13768 11456
rect 13704 11396 13708 11452
rect 13708 11396 13764 11452
rect 13764 11396 13768 11452
rect 13704 11392 13768 11396
rect 21805 11452 21869 11456
rect 21805 11396 21809 11452
rect 21809 11396 21865 11452
rect 21865 11396 21869 11452
rect 21805 11392 21869 11396
rect 21885 11452 21949 11456
rect 21885 11396 21889 11452
rect 21889 11396 21945 11452
rect 21945 11396 21949 11452
rect 21885 11392 21949 11396
rect 21965 11452 22029 11456
rect 21965 11396 21969 11452
rect 21969 11396 22025 11452
rect 22025 11396 22029 11452
rect 21965 11392 22029 11396
rect 22045 11452 22109 11456
rect 22045 11396 22049 11452
rect 22049 11396 22105 11452
rect 22105 11396 22109 11452
rect 22045 11392 22109 11396
rect 9293 10908 9357 10912
rect 9293 10852 9297 10908
rect 9297 10852 9353 10908
rect 9353 10852 9357 10908
rect 9293 10848 9357 10852
rect 9373 10908 9437 10912
rect 9373 10852 9377 10908
rect 9377 10852 9433 10908
rect 9433 10852 9437 10908
rect 9373 10848 9437 10852
rect 9453 10908 9517 10912
rect 9453 10852 9457 10908
rect 9457 10852 9513 10908
rect 9513 10852 9517 10908
rect 9453 10848 9517 10852
rect 9533 10908 9597 10912
rect 9533 10852 9537 10908
rect 9537 10852 9593 10908
rect 9593 10852 9597 10908
rect 9533 10848 9597 10852
rect 17634 10908 17698 10912
rect 17634 10852 17638 10908
rect 17638 10852 17694 10908
rect 17694 10852 17698 10908
rect 17634 10848 17698 10852
rect 17714 10908 17778 10912
rect 17714 10852 17718 10908
rect 17718 10852 17774 10908
rect 17774 10852 17778 10908
rect 17714 10848 17778 10852
rect 17794 10908 17858 10912
rect 17794 10852 17798 10908
rect 17798 10852 17854 10908
rect 17854 10852 17858 10908
rect 17794 10848 17858 10852
rect 17874 10908 17938 10912
rect 17874 10852 17878 10908
rect 17878 10852 17934 10908
rect 17934 10852 17938 10908
rect 17874 10848 17938 10852
rect 5122 10364 5186 10368
rect 5122 10308 5126 10364
rect 5126 10308 5182 10364
rect 5182 10308 5186 10364
rect 5122 10304 5186 10308
rect 5202 10364 5266 10368
rect 5202 10308 5206 10364
rect 5206 10308 5262 10364
rect 5262 10308 5266 10364
rect 5202 10304 5266 10308
rect 5282 10364 5346 10368
rect 5282 10308 5286 10364
rect 5286 10308 5342 10364
rect 5342 10308 5346 10364
rect 5282 10304 5346 10308
rect 5362 10364 5426 10368
rect 5362 10308 5366 10364
rect 5366 10308 5422 10364
rect 5422 10308 5426 10364
rect 5362 10304 5426 10308
rect 13464 10364 13528 10368
rect 13464 10308 13468 10364
rect 13468 10308 13524 10364
rect 13524 10308 13528 10364
rect 13464 10304 13528 10308
rect 13544 10364 13608 10368
rect 13544 10308 13548 10364
rect 13548 10308 13604 10364
rect 13604 10308 13608 10364
rect 13544 10304 13608 10308
rect 13624 10364 13688 10368
rect 13624 10308 13628 10364
rect 13628 10308 13684 10364
rect 13684 10308 13688 10364
rect 13624 10304 13688 10308
rect 13704 10364 13768 10368
rect 13704 10308 13708 10364
rect 13708 10308 13764 10364
rect 13764 10308 13768 10364
rect 13704 10304 13768 10308
rect 21805 10364 21869 10368
rect 21805 10308 21809 10364
rect 21809 10308 21865 10364
rect 21865 10308 21869 10364
rect 21805 10304 21869 10308
rect 21885 10364 21949 10368
rect 21885 10308 21889 10364
rect 21889 10308 21945 10364
rect 21945 10308 21949 10364
rect 21885 10304 21949 10308
rect 21965 10364 22029 10368
rect 21965 10308 21969 10364
rect 21969 10308 22025 10364
rect 22025 10308 22029 10364
rect 21965 10304 22029 10308
rect 22045 10364 22109 10368
rect 22045 10308 22049 10364
rect 22049 10308 22105 10364
rect 22105 10308 22109 10364
rect 22045 10304 22109 10308
rect 9293 9820 9357 9824
rect 9293 9764 9297 9820
rect 9297 9764 9353 9820
rect 9353 9764 9357 9820
rect 9293 9760 9357 9764
rect 9373 9820 9437 9824
rect 9373 9764 9377 9820
rect 9377 9764 9433 9820
rect 9433 9764 9437 9820
rect 9373 9760 9437 9764
rect 9453 9820 9517 9824
rect 9453 9764 9457 9820
rect 9457 9764 9513 9820
rect 9513 9764 9517 9820
rect 9453 9760 9517 9764
rect 9533 9820 9597 9824
rect 9533 9764 9537 9820
rect 9537 9764 9593 9820
rect 9593 9764 9597 9820
rect 9533 9760 9597 9764
rect 17634 9820 17698 9824
rect 17634 9764 17638 9820
rect 17638 9764 17694 9820
rect 17694 9764 17698 9820
rect 17634 9760 17698 9764
rect 17714 9820 17778 9824
rect 17714 9764 17718 9820
rect 17718 9764 17774 9820
rect 17774 9764 17778 9820
rect 17714 9760 17778 9764
rect 17794 9820 17858 9824
rect 17794 9764 17798 9820
rect 17798 9764 17854 9820
rect 17854 9764 17858 9820
rect 17794 9760 17858 9764
rect 17874 9820 17938 9824
rect 17874 9764 17878 9820
rect 17878 9764 17934 9820
rect 17934 9764 17938 9820
rect 17874 9760 17938 9764
rect 5122 9276 5186 9280
rect 5122 9220 5126 9276
rect 5126 9220 5182 9276
rect 5182 9220 5186 9276
rect 5122 9216 5186 9220
rect 5202 9276 5266 9280
rect 5202 9220 5206 9276
rect 5206 9220 5262 9276
rect 5262 9220 5266 9276
rect 5202 9216 5266 9220
rect 5282 9276 5346 9280
rect 5282 9220 5286 9276
rect 5286 9220 5342 9276
rect 5342 9220 5346 9276
rect 5282 9216 5346 9220
rect 5362 9276 5426 9280
rect 5362 9220 5366 9276
rect 5366 9220 5422 9276
rect 5422 9220 5426 9276
rect 5362 9216 5426 9220
rect 13464 9276 13528 9280
rect 13464 9220 13468 9276
rect 13468 9220 13524 9276
rect 13524 9220 13528 9276
rect 13464 9216 13528 9220
rect 13544 9276 13608 9280
rect 13544 9220 13548 9276
rect 13548 9220 13604 9276
rect 13604 9220 13608 9276
rect 13544 9216 13608 9220
rect 13624 9276 13688 9280
rect 13624 9220 13628 9276
rect 13628 9220 13684 9276
rect 13684 9220 13688 9276
rect 13624 9216 13688 9220
rect 13704 9276 13768 9280
rect 13704 9220 13708 9276
rect 13708 9220 13764 9276
rect 13764 9220 13768 9276
rect 13704 9216 13768 9220
rect 21805 9276 21869 9280
rect 21805 9220 21809 9276
rect 21809 9220 21865 9276
rect 21865 9220 21869 9276
rect 21805 9216 21869 9220
rect 21885 9276 21949 9280
rect 21885 9220 21889 9276
rect 21889 9220 21945 9276
rect 21945 9220 21949 9276
rect 21885 9216 21949 9220
rect 21965 9276 22029 9280
rect 21965 9220 21969 9276
rect 21969 9220 22025 9276
rect 22025 9220 22029 9276
rect 21965 9216 22029 9220
rect 22045 9276 22109 9280
rect 22045 9220 22049 9276
rect 22049 9220 22105 9276
rect 22105 9220 22109 9276
rect 22045 9216 22109 9220
rect 9293 8732 9357 8736
rect 9293 8676 9297 8732
rect 9297 8676 9353 8732
rect 9353 8676 9357 8732
rect 9293 8672 9357 8676
rect 9373 8732 9437 8736
rect 9373 8676 9377 8732
rect 9377 8676 9433 8732
rect 9433 8676 9437 8732
rect 9373 8672 9437 8676
rect 9453 8732 9517 8736
rect 9453 8676 9457 8732
rect 9457 8676 9513 8732
rect 9513 8676 9517 8732
rect 9453 8672 9517 8676
rect 9533 8732 9597 8736
rect 9533 8676 9537 8732
rect 9537 8676 9593 8732
rect 9593 8676 9597 8732
rect 9533 8672 9597 8676
rect 17634 8732 17698 8736
rect 17634 8676 17638 8732
rect 17638 8676 17694 8732
rect 17694 8676 17698 8732
rect 17634 8672 17698 8676
rect 17714 8732 17778 8736
rect 17714 8676 17718 8732
rect 17718 8676 17774 8732
rect 17774 8676 17778 8732
rect 17714 8672 17778 8676
rect 17794 8732 17858 8736
rect 17794 8676 17798 8732
rect 17798 8676 17854 8732
rect 17854 8676 17858 8732
rect 17794 8672 17858 8676
rect 17874 8732 17938 8736
rect 17874 8676 17878 8732
rect 17878 8676 17934 8732
rect 17934 8676 17938 8732
rect 17874 8672 17938 8676
rect 5122 8188 5186 8192
rect 5122 8132 5126 8188
rect 5126 8132 5182 8188
rect 5182 8132 5186 8188
rect 5122 8128 5186 8132
rect 5202 8188 5266 8192
rect 5202 8132 5206 8188
rect 5206 8132 5262 8188
rect 5262 8132 5266 8188
rect 5202 8128 5266 8132
rect 5282 8188 5346 8192
rect 5282 8132 5286 8188
rect 5286 8132 5342 8188
rect 5342 8132 5346 8188
rect 5282 8128 5346 8132
rect 5362 8188 5426 8192
rect 5362 8132 5366 8188
rect 5366 8132 5422 8188
rect 5422 8132 5426 8188
rect 5362 8128 5426 8132
rect 13464 8188 13528 8192
rect 13464 8132 13468 8188
rect 13468 8132 13524 8188
rect 13524 8132 13528 8188
rect 13464 8128 13528 8132
rect 13544 8188 13608 8192
rect 13544 8132 13548 8188
rect 13548 8132 13604 8188
rect 13604 8132 13608 8188
rect 13544 8128 13608 8132
rect 13624 8188 13688 8192
rect 13624 8132 13628 8188
rect 13628 8132 13684 8188
rect 13684 8132 13688 8188
rect 13624 8128 13688 8132
rect 13704 8188 13768 8192
rect 13704 8132 13708 8188
rect 13708 8132 13764 8188
rect 13764 8132 13768 8188
rect 13704 8128 13768 8132
rect 21805 8188 21869 8192
rect 21805 8132 21809 8188
rect 21809 8132 21865 8188
rect 21865 8132 21869 8188
rect 21805 8128 21869 8132
rect 21885 8188 21949 8192
rect 21885 8132 21889 8188
rect 21889 8132 21945 8188
rect 21945 8132 21949 8188
rect 21885 8128 21949 8132
rect 21965 8188 22029 8192
rect 21965 8132 21969 8188
rect 21969 8132 22025 8188
rect 22025 8132 22029 8188
rect 21965 8128 22029 8132
rect 22045 8188 22109 8192
rect 22045 8132 22049 8188
rect 22049 8132 22105 8188
rect 22105 8132 22109 8188
rect 22045 8128 22109 8132
rect 9293 7644 9357 7648
rect 9293 7588 9297 7644
rect 9297 7588 9353 7644
rect 9353 7588 9357 7644
rect 9293 7584 9357 7588
rect 9373 7644 9437 7648
rect 9373 7588 9377 7644
rect 9377 7588 9433 7644
rect 9433 7588 9437 7644
rect 9373 7584 9437 7588
rect 9453 7644 9517 7648
rect 9453 7588 9457 7644
rect 9457 7588 9513 7644
rect 9513 7588 9517 7644
rect 9453 7584 9517 7588
rect 9533 7644 9597 7648
rect 9533 7588 9537 7644
rect 9537 7588 9593 7644
rect 9593 7588 9597 7644
rect 9533 7584 9597 7588
rect 17634 7644 17698 7648
rect 17634 7588 17638 7644
rect 17638 7588 17694 7644
rect 17694 7588 17698 7644
rect 17634 7584 17698 7588
rect 17714 7644 17778 7648
rect 17714 7588 17718 7644
rect 17718 7588 17774 7644
rect 17774 7588 17778 7644
rect 17714 7584 17778 7588
rect 17794 7644 17858 7648
rect 17794 7588 17798 7644
rect 17798 7588 17854 7644
rect 17854 7588 17858 7644
rect 17794 7584 17858 7588
rect 17874 7644 17938 7648
rect 17874 7588 17878 7644
rect 17878 7588 17934 7644
rect 17934 7588 17938 7644
rect 17874 7584 17938 7588
rect 5122 7100 5186 7104
rect 5122 7044 5126 7100
rect 5126 7044 5182 7100
rect 5182 7044 5186 7100
rect 5122 7040 5186 7044
rect 5202 7100 5266 7104
rect 5202 7044 5206 7100
rect 5206 7044 5262 7100
rect 5262 7044 5266 7100
rect 5202 7040 5266 7044
rect 5282 7100 5346 7104
rect 5282 7044 5286 7100
rect 5286 7044 5342 7100
rect 5342 7044 5346 7100
rect 5282 7040 5346 7044
rect 5362 7100 5426 7104
rect 5362 7044 5366 7100
rect 5366 7044 5422 7100
rect 5422 7044 5426 7100
rect 5362 7040 5426 7044
rect 13464 7100 13528 7104
rect 13464 7044 13468 7100
rect 13468 7044 13524 7100
rect 13524 7044 13528 7100
rect 13464 7040 13528 7044
rect 13544 7100 13608 7104
rect 13544 7044 13548 7100
rect 13548 7044 13604 7100
rect 13604 7044 13608 7100
rect 13544 7040 13608 7044
rect 13624 7100 13688 7104
rect 13624 7044 13628 7100
rect 13628 7044 13684 7100
rect 13684 7044 13688 7100
rect 13624 7040 13688 7044
rect 13704 7100 13768 7104
rect 13704 7044 13708 7100
rect 13708 7044 13764 7100
rect 13764 7044 13768 7100
rect 13704 7040 13768 7044
rect 21805 7100 21869 7104
rect 21805 7044 21809 7100
rect 21809 7044 21865 7100
rect 21865 7044 21869 7100
rect 21805 7040 21869 7044
rect 21885 7100 21949 7104
rect 21885 7044 21889 7100
rect 21889 7044 21945 7100
rect 21945 7044 21949 7100
rect 21885 7040 21949 7044
rect 21965 7100 22029 7104
rect 21965 7044 21969 7100
rect 21969 7044 22025 7100
rect 22025 7044 22029 7100
rect 21965 7040 22029 7044
rect 22045 7100 22109 7104
rect 22045 7044 22049 7100
rect 22049 7044 22105 7100
rect 22105 7044 22109 7100
rect 22045 7040 22109 7044
rect 9293 6556 9357 6560
rect 9293 6500 9297 6556
rect 9297 6500 9353 6556
rect 9353 6500 9357 6556
rect 9293 6496 9357 6500
rect 9373 6556 9437 6560
rect 9373 6500 9377 6556
rect 9377 6500 9433 6556
rect 9433 6500 9437 6556
rect 9373 6496 9437 6500
rect 9453 6556 9517 6560
rect 9453 6500 9457 6556
rect 9457 6500 9513 6556
rect 9513 6500 9517 6556
rect 9453 6496 9517 6500
rect 9533 6556 9597 6560
rect 9533 6500 9537 6556
rect 9537 6500 9593 6556
rect 9593 6500 9597 6556
rect 9533 6496 9597 6500
rect 17634 6556 17698 6560
rect 17634 6500 17638 6556
rect 17638 6500 17694 6556
rect 17694 6500 17698 6556
rect 17634 6496 17698 6500
rect 17714 6556 17778 6560
rect 17714 6500 17718 6556
rect 17718 6500 17774 6556
rect 17774 6500 17778 6556
rect 17714 6496 17778 6500
rect 17794 6556 17858 6560
rect 17794 6500 17798 6556
rect 17798 6500 17854 6556
rect 17854 6500 17858 6556
rect 17794 6496 17858 6500
rect 17874 6556 17938 6560
rect 17874 6500 17878 6556
rect 17878 6500 17934 6556
rect 17934 6500 17938 6556
rect 17874 6496 17938 6500
rect 5122 6012 5186 6016
rect 5122 5956 5126 6012
rect 5126 5956 5182 6012
rect 5182 5956 5186 6012
rect 5122 5952 5186 5956
rect 5202 6012 5266 6016
rect 5202 5956 5206 6012
rect 5206 5956 5262 6012
rect 5262 5956 5266 6012
rect 5202 5952 5266 5956
rect 5282 6012 5346 6016
rect 5282 5956 5286 6012
rect 5286 5956 5342 6012
rect 5342 5956 5346 6012
rect 5282 5952 5346 5956
rect 5362 6012 5426 6016
rect 5362 5956 5366 6012
rect 5366 5956 5422 6012
rect 5422 5956 5426 6012
rect 5362 5952 5426 5956
rect 13464 6012 13528 6016
rect 13464 5956 13468 6012
rect 13468 5956 13524 6012
rect 13524 5956 13528 6012
rect 13464 5952 13528 5956
rect 13544 6012 13608 6016
rect 13544 5956 13548 6012
rect 13548 5956 13604 6012
rect 13604 5956 13608 6012
rect 13544 5952 13608 5956
rect 13624 6012 13688 6016
rect 13624 5956 13628 6012
rect 13628 5956 13684 6012
rect 13684 5956 13688 6012
rect 13624 5952 13688 5956
rect 13704 6012 13768 6016
rect 13704 5956 13708 6012
rect 13708 5956 13764 6012
rect 13764 5956 13768 6012
rect 13704 5952 13768 5956
rect 21805 6012 21869 6016
rect 21805 5956 21809 6012
rect 21809 5956 21865 6012
rect 21865 5956 21869 6012
rect 21805 5952 21869 5956
rect 21885 6012 21949 6016
rect 21885 5956 21889 6012
rect 21889 5956 21945 6012
rect 21945 5956 21949 6012
rect 21885 5952 21949 5956
rect 21965 6012 22029 6016
rect 21965 5956 21969 6012
rect 21969 5956 22025 6012
rect 22025 5956 22029 6012
rect 21965 5952 22029 5956
rect 22045 6012 22109 6016
rect 22045 5956 22049 6012
rect 22049 5956 22105 6012
rect 22105 5956 22109 6012
rect 22045 5952 22109 5956
rect 9293 5468 9357 5472
rect 9293 5412 9297 5468
rect 9297 5412 9353 5468
rect 9353 5412 9357 5468
rect 9293 5408 9357 5412
rect 9373 5468 9437 5472
rect 9373 5412 9377 5468
rect 9377 5412 9433 5468
rect 9433 5412 9437 5468
rect 9373 5408 9437 5412
rect 9453 5468 9517 5472
rect 9453 5412 9457 5468
rect 9457 5412 9513 5468
rect 9513 5412 9517 5468
rect 9453 5408 9517 5412
rect 9533 5468 9597 5472
rect 9533 5412 9537 5468
rect 9537 5412 9593 5468
rect 9593 5412 9597 5468
rect 9533 5408 9597 5412
rect 17634 5468 17698 5472
rect 17634 5412 17638 5468
rect 17638 5412 17694 5468
rect 17694 5412 17698 5468
rect 17634 5408 17698 5412
rect 17714 5468 17778 5472
rect 17714 5412 17718 5468
rect 17718 5412 17774 5468
rect 17774 5412 17778 5468
rect 17714 5408 17778 5412
rect 17794 5468 17858 5472
rect 17794 5412 17798 5468
rect 17798 5412 17854 5468
rect 17854 5412 17858 5468
rect 17794 5408 17858 5412
rect 17874 5468 17938 5472
rect 17874 5412 17878 5468
rect 17878 5412 17934 5468
rect 17934 5412 17938 5468
rect 17874 5408 17938 5412
rect 5122 4924 5186 4928
rect 5122 4868 5126 4924
rect 5126 4868 5182 4924
rect 5182 4868 5186 4924
rect 5122 4864 5186 4868
rect 5202 4924 5266 4928
rect 5202 4868 5206 4924
rect 5206 4868 5262 4924
rect 5262 4868 5266 4924
rect 5202 4864 5266 4868
rect 5282 4924 5346 4928
rect 5282 4868 5286 4924
rect 5286 4868 5342 4924
rect 5342 4868 5346 4924
rect 5282 4864 5346 4868
rect 5362 4924 5426 4928
rect 5362 4868 5366 4924
rect 5366 4868 5422 4924
rect 5422 4868 5426 4924
rect 5362 4864 5426 4868
rect 13464 4924 13528 4928
rect 13464 4868 13468 4924
rect 13468 4868 13524 4924
rect 13524 4868 13528 4924
rect 13464 4864 13528 4868
rect 13544 4924 13608 4928
rect 13544 4868 13548 4924
rect 13548 4868 13604 4924
rect 13604 4868 13608 4924
rect 13544 4864 13608 4868
rect 13624 4924 13688 4928
rect 13624 4868 13628 4924
rect 13628 4868 13684 4924
rect 13684 4868 13688 4924
rect 13624 4864 13688 4868
rect 13704 4924 13768 4928
rect 13704 4868 13708 4924
rect 13708 4868 13764 4924
rect 13764 4868 13768 4924
rect 13704 4864 13768 4868
rect 21805 4924 21869 4928
rect 21805 4868 21809 4924
rect 21809 4868 21865 4924
rect 21865 4868 21869 4924
rect 21805 4864 21869 4868
rect 21885 4924 21949 4928
rect 21885 4868 21889 4924
rect 21889 4868 21945 4924
rect 21945 4868 21949 4924
rect 21885 4864 21949 4868
rect 21965 4924 22029 4928
rect 21965 4868 21969 4924
rect 21969 4868 22025 4924
rect 22025 4868 22029 4924
rect 21965 4864 22029 4868
rect 22045 4924 22109 4928
rect 22045 4868 22049 4924
rect 22049 4868 22105 4924
rect 22105 4868 22109 4924
rect 22045 4864 22109 4868
rect 9293 4380 9357 4384
rect 9293 4324 9297 4380
rect 9297 4324 9353 4380
rect 9353 4324 9357 4380
rect 9293 4320 9357 4324
rect 9373 4380 9437 4384
rect 9373 4324 9377 4380
rect 9377 4324 9433 4380
rect 9433 4324 9437 4380
rect 9373 4320 9437 4324
rect 9453 4380 9517 4384
rect 9453 4324 9457 4380
rect 9457 4324 9513 4380
rect 9513 4324 9517 4380
rect 9453 4320 9517 4324
rect 9533 4380 9597 4384
rect 9533 4324 9537 4380
rect 9537 4324 9593 4380
rect 9593 4324 9597 4380
rect 9533 4320 9597 4324
rect 17634 4380 17698 4384
rect 17634 4324 17638 4380
rect 17638 4324 17694 4380
rect 17694 4324 17698 4380
rect 17634 4320 17698 4324
rect 17714 4380 17778 4384
rect 17714 4324 17718 4380
rect 17718 4324 17774 4380
rect 17774 4324 17778 4380
rect 17714 4320 17778 4324
rect 17794 4380 17858 4384
rect 17794 4324 17798 4380
rect 17798 4324 17854 4380
rect 17854 4324 17858 4380
rect 17794 4320 17858 4324
rect 17874 4380 17938 4384
rect 17874 4324 17878 4380
rect 17878 4324 17934 4380
rect 17934 4324 17938 4380
rect 17874 4320 17938 4324
rect 5122 3836 5186 3840
rect 5122 3780 5126 3836
rect 5126 3780 5182 3836
rect 5182 3780 5186 3836
rect 5122 3776 5186 3780
rect 5202 3836 5266 3840
rect 5202 3780 5206 3836
rect 5206 3780 5262 3836
rect 5262 3780 5266 3836
rect 5202 3776 5266 3780
rect 5282 3836 5346 3840
rect 5282 3780 5286 3836
rect 5286 3780 5342 3836
rect 5342 3780 5346 3836
rect 5282 3776 5346 3780
rect 5362 3836 5426 3840
rect 5362 3780 5366 3836
rect 5366 3780 5422 3836
rect 5422 3780 5426 3836
rect 5362 3776 5426 3780
rect 13464 3836 13528 3840
rect 13464 3780 13468 3836
rect 13468 3780 13524 3836
rect 13524 3780 13528 3836
rect 13464 3776 13528 3780
rect 13544 3836 13608 3840
rect 13544 3780 13548 3836
rect 13548 3780 13604 3836
rect 13604 3780 13608 3836
rect 13544 3776 13608 3780
rect 13624 3836 13688 3840
rect 13624 3780 13628 3836
rect 13628 3780 13684 3836
rect 13684 3780 13688 3836
rect 13624 3776 13688 3780
rect 13704 3836 13768 3840
rect 13704 3780 13708 3836
rect 13708 3780 13764 3836
rect 13764 3780 13768 3836
rect 13704 3776 13768 3780
rect 21805 3836 21869 3840
rect 21805 3780 21809 3836
rect 21809 3780 21865 3836
rect 21865 3780 21869 3836
rect 21805 3776 21869 3780
rect 21885 3836 21949 3840
rect 21885 3780 21889 3836
rect 21889 3780 21945 3836
rect 21945 3780 21949 3836
rect 21885 3776 21949 3780
rect 21965 3836 22029 3840
rect 21965 3780 21969 3836
rect 21969 3780 22025 3836
rect 22025 3780 22029 3836
rect 21965 3776 22029 3780
rect 22045 3836 22109 3840
rect 22045 3780 22049 3836
rect 22049 3780 22105 3836
rect 22105 3780 22109 3836
rect 22045 3776 22109 3780
rect 9293 3292 9357 3296
rect 9293 3236 9297 3292
rect 9297 3236 9353 3292
rect 9353 3236 9357 3292
rect 9293 3232 9357 3236
rect 9373 3292 9437 3296
rect 9373 3236 9377 3292
rect 9377 3236 9433 3292
rect 9433 3236 9437 3292
rect 9373 3232 9437 3236
rect 9453 3292 9517 3296
rect 9453 3236 9457 3292
rect 9457 3236 9513 3292
rect 9513 3236 9517 3292
rect 9453 3232 9517 3236
rect 9533 3292 9597 3296
rect 9533 3236 9537 3292
rect 9537 3236 9593 3292
rect 9593 3236 9597 3292
rect 9533 3232 9597 3236
rect 17634 3292 17698 3296
rect 17634 3236 17638 3292
rect 17638 3236 17694 3292
rect 17694 3236 17698 3292
rect 17634 3232 17698 3236
rect 17714 3292 17778 3296
rect 17714 3236 17718 3292
rect 17718 3236 17774 3292
rect 17774 3236 17778 3292
rect 17714 3232 17778 3236
rect 17794 3292 17858 3296
rect 17794 3236 17798 3292
rect 17798 3236 17854 3292
rect 17854 3236 17858 3292
rect 17794 3232 17858 3236
rect 17874 3292 17938 3296
rect 17874 3236 17878 3292
rect 17878 3236 17934 3292
rect 17934 3236 17938 3292
rect 17874 3232 17938 3236
rect 5122 2748 5186 2752
rect 5122 2692 5126 2748
rect 5126 2692 5182 2748
rect 5182 2692 5186 2748
rect 5122 2688 5186 2692
rect 5202 2748 5266 2752
rect 5202 2692 5206 2748
rect 5206 2692 5262 2748
rect 5262 2692 5266 2748
rect 5202 2688 5266 2692
rect 5282 2748 5346 2752
rect 5282 2692 5286 2748
rect 5286 2692 5342 2748
rect 5342 2692 5346 2748
rect 5282 2688 5346 2692
rect 5362 2748 5426 2752
rect 5362 2692 5366 2748
rect 5366 2692 5422 2748
rect 5422 2692 5426 2748
rect 5362 2688 5426 2692
rect 13464 2748 13528 2752
rect 13464 2692 13468 2748
rect 13468 2692 13524 2748
rect 13524 2692 13528 2748
rect 13464 2688 13528 2692
rect 13544 2748 13608 2752
rect 13544 2692 13548 2748
rect 13548 2692 13604 2748
rect 13604 2692 13608 2748
rect 13544 2688 13608 2692
rect 13624 2748 13688 2752
rect 13624 2692 13628 2748
rect 13628 2692 13684 2748
rect 13684 2692 13688 2748
rect 13624 2688 13688 2692
rect 13704 2748 13768 2752
rect 13704 2692 13708 2748
rect 13708 2692 13764 2748
rect 13764 2692 13768 2748
rect 13704 2688 13768 2692
rect 21805 2748 21869 2752
rect 21805 2692 21809 2748
rect 21809 2692 21865 2748
rect 21865 2692 21869 2748
rect 21805 2688 21869 2692
rect 21885 2748 21949 2752
rect 21885 2692 21889 2748
rect 21889 2692 21945 2748
rect 21945 2692 21949 2748
rect 21885 2688 21949 2692
rect 21965 2748 22029 2752
rect 21965 2692 21969 2748
rect 21969 2692 22025 2748
rect 22025 2692 22029 2748
rect 21965 2688 22029 2692
rect 22045 2748 22109 2752
rect 22045 2692 22049 2748
rect 22049 2692 22105 2748
rect 22105 2692 22109 2748
rect 22045 2688 22109 2692
rect 9293 2204 9357 2208
rect 9293 2148 9297 2204
rect 9297 2148 9353 2204
rect 9353 2148 9357 2204
rect 9293 2144 9357 2148
rect 9373 2204 9437 2208
rect 9373 2148 9377 2204
rect 9377 2148 9433 2204
rect 9433 2148 9437 2204
rect 9373 2144 9437 2148
rect 9453 2204 9517 2208
rect 9453 2148 9457 2204
rect 9457 2148 9513 2204
rect 9513 2148 9517 2204
rect 9453 2144 9517 2148
rect 9533 2204 9597 2208
rect 9533 2148 9537 2204
rect 9537 2148 9593 2204
rect 9593 2148 9597 2204
rect 9533 2144 9597 2148
rect 17634 2204 17698 2208
rect 17634 2148 17638 2204
rect 17638 2148 17694 2204
rect 17694 2148 17698 2204
rect 17634 2144 17698 2148
rect 17714 2204 17778 2208
rect 17714 2148 17718 2204
rect 17718 2148 17774 2204
rect 17774 2148 17778 2204
rect 17714 2144 17778 2148
rect 17794 2204 17858 2208
rect 17794 2148 17798 2204
rect 17798 2148 17854 2204
rect 17854 2148 17858 2204
rect 17794 2144 17858 2148
rect 17874 2204 17938 2208
rect 17874 2148 17878 2204
rect 17878 2148 17934 2204
rect 17934 2148 17938 2204
rect 17874 2144 17938 2148
<< metal4 >>
rect 5114 26688 5435 27248
rect 5114 26624 5122 26688
rect 5186 26624 5202 26688
rect 5266 26624 5282 26688
rect 5346 26624 5362 26688
rect 5426 26624 5435 26688
rect 5114 25600 5435 26624
rect 5114 25536 5122 25600
rect 5186 25536 5202 25600
rect 5266 25536 5282 25600
rect 5346 25536 5362 25600
rect 5426 25536 5435 25600
rect 5114 24512 5435 25536
rect 5114 24448 5122 24512
rect 5186 24448 5202 24512
rect 5266 24448 5282 24512
rect 5346 24448 5362 24512
rect 5426 24448 5435 24512
rect 5114 23424 5435 24448
rect 5114 23360 5122 23424
rect 5186 23360 5202 23424
rect 5266 23360 5282 23424
rect 5346 23360 5362 23424
rect 5426 23360 5435 23424
rect 5114 22336 5435 23360
rect 5114 22272 5122 22336
rect 5186 22272 5202 22336
rect 5266 22272 5282 22336
rect 5346 22272 5362 22336
rect 5426 22272 5435 22336
rect 5114 21248 5435 22272
rect 5114 21184 5122 21248
rect 5186 21184 5202 21248
rect 5266 21184 5282 21248
rect 5346 21184 5362 21248
rect 5426 21184 5435 21248
rect 5114 20160 5435 21184
rect 5114 20096 5122 20160
rect 5186 20096 5202 20160
rect 5266 20096 5282 20160
rect 5346 20096 5362 20160
rect 5426 20096 5435 20160
rect 5114 19072 5435 20096
rect 5114 19008 5122 19072
rect 5186 19008 5202 19072
rect 5266 19008 5282 19072
rect 5346 19008 5362 19072
rect 5426 19008 5435 19072
rect 5114 17984 5435 19008
rect 5114 17920 5122 17984
rect 5186 17920 5202 17984
rect 5266 17920 5282 17984
rect 5346 17920 5362 17984
rect 5426 17920 5435 17984
rect 5114 16896 5435 17920
rect 5114 16832 5122 16896
rect 5186 16832 5202 16896
rect 5266 16832 5282 16896
rect 5346 16832 5362 16896
rect 5426 16832 5435 16896
rect 5114 15808 5435 16832
rect 5114 15744 5122 15808
rect 5186 15744 5202 15808
rect 5266 15744 5282 15808
rect 5346 15744 5362 15808
rect 5426 15744 5435 15808
rect 5114 14720 5435 15744
rect 5114 14656 5122 14720
rect 5186 14656 5202 14720
rect 5266 14656 5282 14720
rect 5346 14656 5362 14720
rect 5426 14656 5435 14720
rect 5114 13632 5435 14656
rect 5114 13568 5122 13632
rect 5186 13568 5202 13632
rect 5266 13568 5282 13632
rect 5346 13568 5362 13632
rect 5426 13568 5435 13632
rect 5114 12544 5435 13568
rect 5114 12480 5122 12544
rect 5186 12480 5202 12544
rect 5266 12480 5282 12544
rect 5346 12480 5362 12544
rect 5426 12480 5435 12544
rect 5114 11456 5435 12480
rect 5114 11392 5122 11456
rect 5186 11392 5202 11456
rect 5266 11392 5282 11456
rect 5346 11392 5362 11456
rect 5426 11392 5435 11456
rect 5114 10368 5435 11392
rect 5114 10304 5122 10368
rect 5186 10304 5202 10368
rect 5266 10304 5282 10368
rect 5346 10304 5362 10368
rect 5426 10304 5435 10368
rect 5114 9280 5435 10304
rect 5114 9216 5122 9280
rect 5186 9216 5202 9280
rect 5266 9216 5282 9280
rect 5346 9216 5362 9280
rect 5426 9216 5435 9280
rect 5114 8192 5435 9216
rect 5114 8128 5122 8192
rect 5186 8128 5202 8192
rect 5266 8128 5282 8192
rect 5346 8128 5362 8192
rect 5426 8128 5435 8192
rect 5114 7104 5435 8128
rect 5114 7040 5122 7104
rect 5186 7040 5202 7104
rect 5266 7040 5282 7104
rect 5346 7040 5362 7104
rect 5426 7040 5435 7104
rect 5114 6016 5435 7040
rect 5114 5952 5122 6016
rect 5186 5952 5202 6016
rect 5266 5952 5282 6016
rect 5346 5952 5362 6016
rect 5426 5952 5435 6016
rect 5114 4928 5435 5952
rect 5114 4864 5122 4928
rect 5186 4864 5202 4928
rect 5266 4864 5282 4928
rect 5346 4864 5362 4928
rect 5426 4864 5435 4928
rect 5114 3840 5435 4864
rect 5114 3776 5122 3840
rect 5186 3776 5202 3840
rect 5266 3776 5282 3840
rect 5346 3776 5362 3840
rect 5426 3776 5435 3840
rect 5114 2752 5435 3776
rect 5114 2688 5122 2752
rect 5186 2688 5202 2752
rect 5266 2688 5282 2752
rect 5346 2688 5362 2752
rect 5426 2688 5435 2752
rect 5114 2128 5435 2688
rect 9285 27232 9605 27248
rect 9285 27168 9293 27232
rect 9357 27168 9373 27232
rect 9437 27168 9453 27232
rect 9517 27168 9533 27232
rect 9597 27168 9605 27232
rect 9285 26144 9605 27168
rect 9285 26080 9293 26144
rect 9357 26080 9373 26144
rect 9437 26080 9453 26144
rect 9517 26080 9533 26144
rect 9597 26080 9605 26144
rect 9285 25056 9605 26080
rect 9285 24992 9293 25056
rect 9357 24992 9373 25056
rect 9437 24992 9453 25056
rect 9517 24992 9533 25056
rect 9597 24992 9605 25056
rect 9285 23968 9605 24992
rect 9285 23904 9293 23968
rect 9357 23904 9373 23968
rect 9437 23904 9453 23968
rect 9517 23904 9533 23968
rect 9597 23904 9605 23968
rect 9285 22880 9605 23904
rect 9285 22816 9293 22880
rect 9357 22816 9373 22880
rect 9437 22816 9453 22880
rect 9517 22816 9533 22880
rect 9597 22816 9605 22880
rect 9285 21792 9605 22816
rect 9285 21728 9293 21792
rect 9357 21728 9373 21792
rect 9437 21728 9453 21792
rect 9517 21728 9533 21792
rect 9597 21728 9605 21792
rect 9285 20704 9605 21728
rect 9285 20640 9293 20704
rect 9357 20640 9373 20704
rect 9437 20640 9453 20704
rect 9517 20640 9533 20704
rect 9597 20640 9605 20704
rect 9285 19616 9605 20640
rect 9285 19552 9293 19616
rect 9357 19552 9373 19616
rect 9437 19552 9453 19616
rect 9517 19552 9533 19616
rect 9597 19552 9605 19616
rect 9285 18528 9605 19552
rect 9285 18464 9293 18528
rect 9357 18464 9373 18528
rect 9437 18464 9453 18528
rect 9517 18464 9533 18528
rect 9597 18464 9605 18528
rect 9285 17440 9605 18464
rect 9285 17376 9293 17440
rect 9357 17376 9373 17440
rect 9437 17376 9453 17440
rect 9517 17376 9533 17440
rect 9597 17376 9605 17440
rect 9285 16352 9605 17376
rect 9285 16288 9293 16352
rect 9357 16288 9373 16352
rect 9437 16288 9453 16352
rect 9517 16288 9533 16352
rect 9597 16288 9605 16352
rect 9285 15264 9605 16288
rect 9285 15200 9293 15264
rect 9357 15200 9373 15264
rect 9437 15200 9453 15264
rect 9517 15200 9533 15264
rect 9597 15200 9605 15264
rect 9285 14176 9605 15200
rect 9285 14112 9293 14176
rect 9357 14112 9373 14176
rect 9437 14112 9453 14176
rect 9517 14112 9533 14176
rect 9597 14112 9605 14176
rect 9285 13088 9605 14112
rect 9285 13024 9293 13088
rect 9357 13024 9373 13088
rect 9437 13024 9453 13088
rect 9517 13024 9533 13088
rect 9597 13024 9605 13088
rect 9285 12000 9605 13024
rect 9285 11936 9293 12000
rect 9357 11936 9373 12000
rect 9437 11936 9453 12000
rect 9517 11936 9533 12000
rect 9597 11936 9605 12000
rect 9285 10912 9605 11936
rect 9285 10848 9293 10912
rect 9357 10848 9373 10912
rect 9437 10848 9453 10912
rect 9517 10848 9533 10912
rect 9597 10848 9605 10912
rect 9285 9824 9605 10848
rect 9285 9760 9293 9824
rect 9357 9760 9373 9824
rect 9437 9760 9453 9824
rect 9517 9760 9533 9824
rect 9597 9760 9605 9824
rect 9285 8736 9605 9760
rect 9285 8672 9293 8736
rect 9357 8672 9373 8736
rect 9437 8672 9453 8736
rect 9517 8672 9533 8736
rect 9597 8672 9605 8736
rect 9285 7648 9605 8672
rect 9285 7584 9293 7648
rect 9357 7584 9373 7648
rect 9437 7584 9453 7648
rect 9517 7584 9533 7648
rect 9597 7584 9605 7648
rect 9285 6560 9605 7584
rect 9285 6496 9293 6560
rect 9357 6496 9373 6560
rect 9437 6496 9453 6560
rect 9517 6496 9533 6560
rect 9597 6496 9605 6560
rect 9285 5472 9605 6496
rect 9285 5408 9293 5472
rect 9357 5408 9373 5472
rect 9437 5408 9453 5472
rect 9517 5408 9533 5472
rect 9597 5408 9605 5472
rect 9285 4384 9605 5408
rect 9285 4320 9293 4384
rect 9357 4320 9373 4384
rect 9437 4320 9453 4384
rect 9517 4320 9533 4384
rect 9597 4320 9605 4384
rect 9285 3296 9605 4320
rect 9285 3232 9293 3296
rect 9357 3232 9373 3296
rect 9437 3232 9453 3296
rect 9517 3232 9533 3296
rect 9597 3232 9605 3296
rect 9285 2208 9605 3232
rect 9285 2144 9293 2208
rect 9357 2144 9373 2208
rect 9437 2144 9453 2208
rect 9517 2144 9533 2208
rect 9597 2144 9605 2208
rect 9285 2128 9605 2144
rect 13456 26688 13776 27248
rect 13456 26624 13464 26688
rect 13528 26624 13544 26688
rect 13608 26624 13624 26688
rect 13688 26624 13704 26688
rect 13768 26624 13776 26688
rect 13456 25600 13776 26624
rect 13456 25536 13464 25600
rect 13528 25536 13544 25600
rect 13608 25536 13624 25600
rect 13688 25536 13704 25600
rect 13768 25536 13776 25600
rect 13456 24512 13776 25536
rect 13456 24448 13464 24512
rect 13528 24448 13544 24512
rect 13608 24448 13624 24512
rect 13688 24448 13704 24512
rect 13768 24448 13776 24512
rect 13456 23424 13776 24448
rect 13456 23360 13464 23424
rect 13528 23360 13544 23424
rect 13608 23360 13624 23424
rect 13688 23360 13704 23424
rect 13768 23360 13776 23424
rect 13456 22336 13776 23360
rect 13456 22272 13464 22336
rect 13528 22272 13544 22336
rect 13608 22272 13624 22336
rect 13688 22272 13704 22336
rect 13768 22272 13776 22336
rect 13456 21248 13776 22272
rect 13456 21184 13464 21248
rect 13528 21184 13544 21248
rect 13608 21184 13624 21248
rect 13688 21184 13704 21248
rect 13768 21184 13776 21248
rect 13456 20160 13776 21184
rect 13456 20096 13464 20160
rect 13528 20096 13544 20160
rect 13608 20096 13624 20160
rect 13688 20096 13704 20160
rect 13768 20096 13776 20160
rect 13456 19072 13776 20096
rect 13456 19008 13464 19072
rect 13528 19008 13544 19072
rect 13608 19008 13624 19072
rect 13688 19008 13704 19072
rect 13768 19008 13776 19072
rect 13456 17984 13776 19008
rect 13456 17920 13464 17984
rect 13528 17920 13544 17984
rect 13608 17920 13624 17984
rect 13688 17920 13704 17984
rect 13768 17920 13776 17984
rect 13456 16896 13776 17920
rect 13456 16832 13464 16896
rect 13528 16832 13544 16896
rect 13608 16832 13624 16896
rect 13688 16832 13704 16896
rect 13768 16832 13776 16896
rect 13456 15808 13776 16832
rect 13456 15744 13464 15808
rect 13528 15744 13544 15808
rect 13608 15744 13624 15808
rect 13688 15744 13704 15808
rect 13768 15744 13776 15808
rect 13456 14720 13776 15744
rect 13456 14656 13464 14720
rect 13528 14656 13544 14720
rect 13608 14656 13624 14720
rect 13688 14656 13704 14720
rect 13768 14656 13776 14720
rect 13456 13632 13776 14656
rect 13456 13568 13464 13632
rect 13528 13568 13544 13632
rect 13608 13568 13624 13632
rect 13688 13568 13704 13632
rect 13768 13568 13776 13632
rect 13456 12544 13776 13568
rect 13456 12480 13464 12544
rect 13528 12480 13544 12544
rect 13608 12480 13624 12544
rect 13688 12480 13704 12544
rect 13768 12480 13776 12544
rect 13456 11456 13776 12480
rect 13456 11392 13464 11456
rect 13528 11392 13544 11456
rect 13608 11392 13624 11456
rect 13688 11392 13704 11456
rect 13768 11392 13776 11456
rect 13456 10368 13776 11392
rect 13456 10304 13464 10368
rect 13528 10304 13544 10368
rect 13608 10304 13624 10368
rect 13688 10304 13704 10368
rect 13768 10304 13776 10368
rect 13456 9280 13776 10304
rect 13456 9216 13464 9280
rect 13528 9216 13544 9280
rect 13608 9216 13624 9280
rect 13688 9216 13704 9280
rect 13768 9216 13776 9280
rect 13456 8192 13776 9216
rect 13456 8128 13464 8192
rect 13528 8128 13544 8192
rect 13608 8128 13624 8192
rect 13688 8128 13704 8192
rect 13768 8128 13776 8192
rect 13456 7104 13776 8128
rect 13456 7040 13464 7104
rect 13528 7040 13544 7104
rect 13608 7040 13624 7104
rect 13688 7040 13704 7104
rect 13768 7040 13776 7104
rect 13456 6016 13776 7040
rect 13456 5952 13464 6016
rect 13528 5952 13544 6016
rect 13608 5952 13624 6016
rect 13688 5952 13704 6016
rect 13768 5952 13776 6016
rect 13456 4928 13776 5952
rect 13456 4864 13464 4928
rect 13528 4864 13544 4928
rect 13608 4864 13624 4928
rect 13688 4864 13704 4928
rect 13768 4864 13776 4928
rect 13456 3840 13776 4864
rect 13456 3776 13464 3840
rect 13528 3776 13544 3840
rect 13608 3776 13624 3840
rect 13688 3776 13704 3840
rect 13768 3776 13776 3840
rect 13456 2752 13776 3776
rect 13456 2688 13464 2752
rect 13528 2688 13544 2752
rect 13608 2688 13624 2752
rect 13688 2688 13704 2752
rect 13768 2688 13776 2752
rect 13456 2128 13776 2688
rect 17626 27232 17946 27248
rect 17626 27168 17634 27232
rect 17698 27168 17714 27232
rect 17778 27168 17794 27232
rect 17858 27168 17874 27232
rect 17938 27168 17946 27232
rect 17626 26144 17946 27168
rect 17626 26080 17634 26144
rect 17698 26080 17714 26144
rect 17778 26080 17794 26144
rect 17858 26080 17874 26144
rect 17938 26080 17946 26144
rect 17626 25056 17946 26080
rect 17626 24992 17634 25056
rect 17698 24992 17714 25056
rect 17778 24992 17794 25056
rect 17858 24992 17874 25056
rect 17938 24992 17946 25056
rect 17626 23968 17946 24992
rect 17626 23904 17634 23968
rect 17698 23904 17714 23968
rect 17778 23904 17794 23968
rect 17858 23904 17874 23968
rect 17938 23904 17946 23968
rect 17626 22880 17946 23904
rect 17626 22816 17634 22880
rect 17698 22816 17714 22880
rect 17778 22816 17794 22880
rect 17858 22816 17874 22880
rect 17938 22816 17946 22880
rect 17626 21792 17946 22816
rect 17626 21728 17634 21792
rect 17698 21728 17714 21792
rect 17778 21728 17794 21792
rect 17858 21728 17874 21792
rect 17938 21728 17946 21792
rect 17626 20704 17946 21728
rect 17626 20640 17634 20704
rect 17698 20640 17714 20704
rect 17778 20640 17794 20704
rect 17858 20640 17874 20704
rect 17938 20640 17946 20704
rect 17626 19616 17946 20640
rect 17626 19552 17634 19616
rect 17698 19552 17714 19616
rect 17778 19552 17794 19616
rect 17858 19552 17874 19616
rect 17938 19552 17946 19616
rect 17626 18528 17946 19552
rect 17626 18464 17634 18528
rect 17698 18464 17714 18528
rect 17778 18464 17794 18528
rect 17858 18464 17874 18528
rect 17938 18464 17946 18528
rect 17626 17440 17946 18464
rect 17626 17376 17634 17440
rect 17698 17376 17714 17440
rect 17778 17376 17794 17440
rect 17858 17376 17874 17440
rect 17938 17376 17946 17440
rect 17626 16352 17946 17376
rect 17626 16288 17634 16352
rect 17698 16288 17714 16352
rect 17778 16288 17794 16352
rect 17858 16288 17874 16352
rect 17938 16288 17946 16352
rect 17626 15264 17946 16288
rect 17626 15200 17634 15264
rect 17698 15200 17714 15264
rect 17778 15200 17794 15264
rect 17858 15200 17874 15264
rect 17938 15200 17946 15264
rect 17626 14176 17946 15200
rect 17626 14112 17634 14176
rect 17698 14112 17714 14176
rect 17778 14112 17794 14176
rect 17858 14112 17874 14176
rect 17938 14112 17946 14176
rect 17626 13088 17946 14112
rect 17626 13024 17634 13088
rect 17698 13024 17714 13088
rect 17778 13024 17794 13088
rect 17858 13024 17874 13088
rect 17938 13024 17946 13088
rect 17626 12000 17946 13024
rect 17626 11936 17634 12000
rect 17698 11936 17714 12000
rect 17778 11936 17794 12000
rect 17858 11936 17874 12000
rect 17938 11936 17946 12000
rect 17626 10912 17946 11936
rect 17626 10848 17634 10912
rect 17698 10848 17714 10912
rect 17778 10848 17794 10912
rect 17858 10848 17874 10912
rect 17938 10848 17946 10912
rect 17626 9824 17946 10848
rect 17626 9760 17634 9824
rect 17698 9760 17714 9824
rect 17778 9760 17794 9824
rect 17858 9760 17874 9824
rect 17938 9760 17946 9824
rect 17626 8736 17946 9760
rect 17626 8672 17634 8736
rect 17698 8672 17714 8736
rect 17778 8672 17794 8736
rect 17858 8672 17874 8736
rect 17938 8672 17946 8736
rect 17626 7648 17946 8672
rect 17626 7584 17634 7648
rect 17698 7584 17714 7648
rect 17778 7584 17794 7648
rect 17858 7584 17874 7648
rect 17938 7584 17946 7648
rect 17626 6560 17946 7584
rect 17626 6496 17634 6560
rect 17698 6496 17714 6560
rect 17778 6496 17794 6560
rect 17858 6496 17874 6560
rect 17938 6496 17946 6560
rect 17626 5472 17946 6496
rect 17626 5408 17634 5472
rect 17698 5408 17714 5472
rect 17778 5408 17794 5472
rect 17858 5408 17874 5472
rect 17938 5408 17946 5472
rect 17626 4384 17946 5408
rect 17626 4320 17634 4384
rect 17698 4320 17714 4384
rect 17778 4320 17794 4384
rect 17858 4320 17874 4384
rect 17938 4320 17946 4384
rect 17626 3296 17946 4320
rect 17626 3232 17634 3296
rect 17698 3232 17714 3296
rect 17778 3232 17794 3296
rect 17858 3232 17874 3296
rect 17938 3232 17946 3296
rect 17626 2208 17946 3232
rect 17626 2144 17634 2208
rect 17698 2144 17714 2208
rect 17778 2144 17794 2208
rect 17858 2144 17874 2208
rect 17938 2144 17946 2208
rect 17626 2128 17946 2144
rect 21797 26688 22117 27248
rect 21797 26624 21805 26688
rect 21869 26624 21885 26688
rect 21949 26624 21965 26688
rect 22029 26624 22045 26688
rect 22109 26624 22117 26688
rect 21797 25600 22117 26624
rect 21797 25536 21805 25600
rect 21869 25536 21885 25600
rect 21949 25536 21965 25600
rect 22029 25536 22045 25600
rect 22109 25536 22117 25600
rect 21797 24512 22117 25536
rect 21797 24448 21805 24512
rect 21869 24448 21885 24512
rect 21949 24448 21965 24512
rect 22029 24448 22045 24512
rect 22109 24448 22117 24512
rect 21797 23424 22117 24448
rect 21797 23360 21805 23424
rect 21869 23360 21885 23424
rect 21949 23360 21965 23424
rect 22029 23360 22045 23424
rect 22109 23360 22117 23424
rect 21797 22336 22117 23360
rect 21797 22272 21805 22336
rect 21869 22272 21885 22336
rect 21949 22272 21965 22336
rect 22029 22272 22045 22336
rect 22109 22272 22117 22336
rect 21797 21248 22117 22272
rect 21797 21184 21805 21248
rect 21869 21184 21885 21248
rect 21949 21184 21965 21248
rect 22029 21184 22045 21248
rect 22109 21184 22117 21248
rect 21797 20160 22117 21184
rect 21797 20096 21805 20160
rect 21869 20096 21885 20160
rect 21949 20096 21965 20160
rect 22029 20096 22045 20160
rect 22109 20096 22117 20160
rect 21797 19072 22117 20096
rect 21797 19008 21805 19072
rect 21869 19008 21885 19072
rect 21949 19008 21965 19072
rect 22029 19008 22045 19072
rect 22109 19008 22117 19072
rect 21797 17984 22117 19008
rect 21797 17920 21805 17984
rect 21869 17920 21885 17984
rect 21949 17920 21965 17984
rect 22029 17920 22045 17984
rect 22109 17920 22117 17984
rect 21797 16896 22117 17920
rect 21797 16832 21805 16896
rect 21869 16832 21885 16896
rect 21949 16832 21965 16896
rect 22029 16832 22045 16896
rect 22109 16832 22117 16896
rect 21797 15808 22117 16832
rect 21797 15744 21805 15808
rect 21869 15744 21885 15808
rect 21949 15744 21965 15808
rect 22029 15744 22045 15808
rect 22109 15744 22117 15808
rect 21797 14720 22117 15744
rect 21797 14656 21805 14720
rect 21869 14656 21885 14720
rect 21949 14656 21965 14720
rect 22029 14656 22045 14720
rect 22109 14656 22117 14720
rect 21797 13632 22117 14656
rect 21797 13568 21805 13632
rect 21869 13568 21885 13632
rect 21949 13568 21965 13632
rect 22029 13568 22045 13632
rect 22109 13568 22117 13632
rect 21797 12544 22117 13568
rect 21797 12480 21805 12544
rect 21869 12480 21885 12544
rect 21949 12480 21965 12544
rect 22029 12480 22045 12544
rect 22109 12480 22117 12544
rect 21797 11456 22117 12480
rect 21797 11392 21805 11456
rect 21869 11392 21885 11456
rect 21949 11392 21965 11456
rect 22029 11392 22045 11456
rect 22109 11392 22117 11456
rect 21797 10368 22117 11392
rect 21797 10304 21805 10368
rect 21869 10304 21885 10368
rect 21949 10304 21965 10368
rect 22029 10304 22045 10368
rect 22109 10304 22117 10368
rect 21797 9280 22117 10304
rect 21797 9216 21805 9280
rect 21869 9216 21885 9280
rect 21949 9216 21965 9280
rect 22029 9216 22045 9280
rect 22109 9216 22117 9280
rect 21797 8192 22117 9216
rect 21797 8128 21805 8192
rect 21869 8128 21885 8192
rect 21949 8128 21965 8192
rect 22029 8128 22045 8192
rect 22109 8128 22117 8192
rect 21797 7104 22117 8128
rect 21797 7040 21805 7104
rect 21869 7040 21885 7104
rect 21949 7040 21965 7104
rect 22029 7040 22045 7104
rect 22109 7040 22117 7104
rect 21797 6016 22117 7040
rect 21797 5952 21805 6016
rect 21869 5952 21885 6016
rect 21949 5952 21965 6016
rect 22029 5952 22045 6016
rect 22109 5952 22117 6016
rect 21797 4928 22117 5952
rect 21797 4864 21805 4928
rect 21869 4864 21885 4928
rect 21949 4864 21965 4928
rect 22029 4864 22045 4928
rect 22109 4864 22117 4928
rect 21797 3840 22117 4864
rect 21797 3776 21805 3840
rect 21869 3776 21885 3840
rect 21949 3776 21965 3840
rect 22029 3776 22045 3840
rect 22109 3776 22117 3840
rect 21797 2752 22117 3776
rect 21797 2688 21805 2752
rect 21869 2688 21885 2752
rect 21949 2688 21965 2752
rect 22029 2688 22045 2752
rect 22109 2688 22117 2752
rect 21797 2128 22117 2688
use sky130_fd_sc_hd__decap_12  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1639504043
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1639504043
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1639504043
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1639504043
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1639504043
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1639504043
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1639504043
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1003_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 4692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__S $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1639504043
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1639504043
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1639504043
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 6532 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1639504043
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1639504043
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1002_
timestamp 1639504043
transform -1 0 6164 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73
timestamp 1639504043
transform 1 0 7820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_67
timestamp 1639504043
transform 1 0 7268 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1001_
timestamp 1639504043
transform -1 0 8648 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 8924 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1639504043
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1639504043
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_85
timestamp 1639504043
transform 1 0 8924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_97
timestamp 1639504043
transform 1 0 10028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1639504043
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1639504043
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1639504043
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1639504043
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1639504043
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1639504043
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1639504043
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1333_
timestamp 1639504043
transform 1 0 11500 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1639504043
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1639504043
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_133
timestamp 1639504043
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_145
timestamp 1639504043
transform 1 0 14444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1639504043
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0911_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 13064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1639504043
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1639504043
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_155
timestamp 1639504043
transform 1 0 15364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_2  _0907_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 15364 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1639504043
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1639504043
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1639504043
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1639504043
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1639504043
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1639504043
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1639504043
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1639504043
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1639504043
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1639504043
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1639504043
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1639504043
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1639504043
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1639504043
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1639504043
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1639504043
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1639504043
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1639504043
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1639504043
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1639504043
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1639504043
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1639504043
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1639504043
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1639504043
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1639504043
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_261
timestamp 1639504043
transform 1 0 25116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1639504043
transform -1 0 26128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1639504043
transform -1 0 26128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1639504043
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A
timestamp 1639504043
transform -1 0 2576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_16
timestamp 1639504043
transform 1 0 2576 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1639504043
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_9
timestamp 1639504043
transform 1 0 1932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1639504043
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1639504043
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_35
timestamp 1639504043
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1639504043
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1296_
timestamp 1639504043
transform 1 0 4416 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1297_
timestamp 1639504043
transform -1 0 7544 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__S
timestamp 1639504043
transform 1 0 7544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1639504043
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _1000_
timestamp 1639504043
transform -1 0 8832 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1639504043
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1299_
timestamp 1639504043
transform -1 0 10488 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1303_
timestamp 1639504043
transform 1 0 10488 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_1  _0913_
timestamp 1639504043
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1334_
timestamp 1639504043
transform 1 0 12328 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1639504043
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1639504043
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0908_
timestamp 1639504043
transform 1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1336_
timestamp 1639504043
transform 1 0 15088 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_2_186
timestamp 1639504043
transform 1 0 18216 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1339_
timestamp 1639504043
transform -1 0 18216 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1639504043
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1639504043
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1639504043
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A
timestamp 1639504043
transform 1 0 21620 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1639504043
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1639504043
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _0989_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 22264 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B
timestamp 1639504043
transform -1 0 22724 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_235
timestamp 1639504043
transform 1 0 22724 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_240
timestamp 1639504043
transform 1 0 23184 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0990_
timestamp 1639504043
transform -1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 22908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_256
timestamp 1639504043
transform 1 0 24656 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_261
timestamp 1639504043
transform 1 0 25116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1639504043
transform -1 0 26128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1639504043
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1162_
timestamp 1639504043
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1164_
timestamp 1639504043
transform 1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1639504043
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1639504043
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1639504043
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1639504043
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_2  _1004_
timestamp 1639504043
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1639504043
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1205_
timestamp 1639504043
transform 1 0 5428 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A1
timestamp 1639504043
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_71
timestamp 1639504043
transform 1 0 7636 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0996_
timestamp 1639504043
transform -1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0999_
timestamp 1639504043
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1258_
timestamp 1639504043
transform 1 0 8004 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__S
timestamp 1639504043
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__S
timestamp 1639504043
transform 1 0 9844 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_97
timestamp 1639504043
transform 1 0 10028 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0912_
timestamp 1639504043
transform -1 0 10764 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1255_
timestamp 1639504043
transform 1 0 8832 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_116
timestamp 1639504043
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1639504043
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0910_
timestamp 1639504043
transform 1 0 10764 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0915_
timestamp 1639504043
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1132_
timestamp 1639504043
transform 1 0 12052 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_127
timestamp 1639504043
transform 1 0 12788 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1134_
timestamp 1639504043
transform 1 0 14444 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1335_
timestamp 1639504043
transform 1 0 12880 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_3_158
timestamp 1639504043
transform 1 0 15640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1133_
timestamp 1639504043
transform 1 0 15180 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1138_
timestamp 1639504043
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1639504043
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_177
timestamp 1639504043
transform 1 0 17388 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1639504043
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0902_
timestamp 1639504043
transform 1 0 17112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1137_
timestamp 1639504043
transform 1 0 16652 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_3_189
timestamp 1639504043
transform 1 0 18492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_201
timestamp 1639504043
transform 1 0 19596 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_213
timestamp 1639504043
transform 1 0 20700 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_221
timestamp 1639504043
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1639504043
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1639504043
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1304_
timestamp 1639504043
transform 1 0 21988 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_3_244
timestamp 1639504043
transform 1 0 23552 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_256
timestamp 1639504043
transform 1 0 24656 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_268
timestamp 1639504043
transform 1 0 25760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1639504043
transform -1 0 26128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_14
timestamp 1639504043
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1639504043
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp 1639504043
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1639504043
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1168_
timestamp 1639504043
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1639504043
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1639504043
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1639504043
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1295_
timestamp 1639504043
transform 1 0 3864 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__o22a_2  _0995_
timestamp 1639504043
transform -1 0 6992 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1182_
timestamp 1639504043
transform 1 0 5428 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0993_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 6992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0998_
timestamp 1639504043
transform 1 0 7268 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1257_
timestamp 1639504043
transform -1 0 8832 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__S
timestamp 1639504043
transform 1 0 10488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1639504043
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0914_
timestamp 1639504043
transform 1 0 10672 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1300_
timestamp 1639504043
transform -1 0 10488 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1220_
timestamp 1639504043
transform 1 0 12144 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1224_
timestamp 1639504043
transform 1 0 11316 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1639504043
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1639504043
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1232_
timestamp 1639504043
transform 1 0 12972 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_147
timestamp 1639504043
transform 1 0 14628 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_158
timestamp 1639504043
transform 1 0 15640 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_166
timestamp 1639504043
transform 1 0 16376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__and2b_2  _0901_
timestamp 1639504043
transform 1 0 15732 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1228_
timestamp 1639504043
transform 1 0 14812 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_181
timestamp 1639504043
transform 1 0 17756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _0732_
timestamp 1639504043
transform 1 0 16560 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1143_
timestamp 1639504043
transform -1 0 17756 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1639504043
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1639504043
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1639504043
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1639504043
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1639504043
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1639504043
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1639504043
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1639504043
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1639504043
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_265
timestamp 1639504043
transform 1 0 25484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1639504043
transform -1 0 26128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1639504043
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1639504043
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1639504043
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1639504043
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1294_
timestamp 1639504043
transform -1 0 4232 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _1005_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 4968 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__S
timestamp 1639504043
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1639504043
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0992_
timestamp 1639504043
transform -1 0 6072 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1206_
timestamp 1639504043
transform 1 0 4968 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1302_
timestamp 1639504043
transform 1 0 6348 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1301_
timestamp 1639504043
transform 1 0 7912 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__S
timestamp 1639504043
transform 1 0 10304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_102
timestamp 1639504043
transform 1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1234_
timestamp 1639504043
transform 1 0 9476 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1639504043
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0916_
timestamp 1639504043
transform 1 0 10764 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1332_
timestamp 1639504043
transform 1 0 11500 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1639504043
transform 1 0 13524 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _0733_
timestamp 1639504043
transform 1 0 13064 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_5_147
timestamp 1639504043
transform 1 0 14628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_160
timestamp 1639504043
transform 1 0 15824 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__and2b_2  _0903_
timestamp 1639504043
transform 1 0 15180 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1141_
timestamp 1639504043
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 1639504043
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_186
timestamp 1639504043
transform 1 0 18216 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1639504043
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _0735_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 17572 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1175_
timestamp 1639504043
transform 1 0 16744 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_192
timestamp 1639504043
transform 1 0 18768 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1340_
timestamp 1639504043
transform 1 0 18860 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_5_210
timestamp 1639504043
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1639504043
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1639504043
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1639504043
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1639504043
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1639504043
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_261
timestamp 1639504043
transform 1 0 25116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1639504043
transform -1 0 26128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1639504043
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1639504043
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1639504043
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1639504043
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1639504043
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 2484 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 2484 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1355_
timestamp 1639504043
transform -1 0 3036 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__a21boi_2  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 3956 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0856_
timestamp 1639504043
transform 1 0 3956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1639504043
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1639504043
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_21
timestamp 1639504043
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B1
timestamp 1639504043
transform -1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _0771_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 4876 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_38
timestamp 1639504043
transform 1 0 4600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1639504043
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1639504043
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__B1
timestamp 1639504043
transform -1 0 4876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1639504043
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__S
timestamp 1639504043
transform 1 0 5796 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_48
timestamp 1639504043
transform 1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1639504043
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1639504043
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1639504043
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1639504043
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0994_
timestamp 1639504043
transform -1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 6072 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1639504043
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_73
timestamp 1639504043
transform 1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 1639504043
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _0997_
timestamp 1639504043
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1392_
timestamp 1639504043
transform 1 0 8004 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_6_103
timestamp 1639504043
transform 1 0 10580 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1639504043
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_91
timestamp 1639504043
transform 1 0 9476 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1639504043
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_92
timestamp 1639504043
transform 1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1639504043
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_clk
timestamp 1639504043
transform 1 0 9108 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1639504043
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_111
timestamp 1639504043
transform 1 0 11316 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1639504043
transform 1 0 12512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_121
timestamp 1639504043
transform 1 0 12236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1639504043
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0917_
timestamp 1639504043
transform 1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0991_
timestamp 1639504043
transform -1 0 12236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1229_
timestamp 1639504043
transform 1 0 11684 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_132
timestamp 1639504043
transform 1 0 13248 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1639504043
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_133
timestamp 1639504043
transform 1 0 13340 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1639504043
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0905_
timestamp 1639504043
transform -1 0 14720 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0909_
timestamp 1639504043
transform -1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1639504043
transform 1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_150
timestamp 1639504043
transform 1 0 14904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0900_
timestamp 1639504043
transform -1 0 14904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0904_
timestamp 1639504043
transform -1 0 16560 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1140_
timestamp 1639504043
transform 1 0 15088 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1337_
timestamp 1639504043
transform 1 0 14720 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1338_
timestamp 1639504043
transform 1 0 15824 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1639504043
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_177
timestamp 1639504043
transform 1 0 17388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1639504043
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0899_
timestamp 1639504043
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1139_
timestamp 1639504043
transform 1 0 17388 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1142_
timestamp 1639504043
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_189
timestamp 1639504043
transform 1 0 18492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1639504043
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0736_
timestamp 1639504043
transform 1 0 19872 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0891_
timestamp 1639504043
transform 1 0 18768 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0898_
timestamp 1639504043
transform -1 0 19136 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1144_
timestamp 1639504043
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1178_
timestamp 1639504043
transform 1 0 19044 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1341_
timestamp 1639504043
transform 1 0 19964 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_6_222
timestamp 1639504043
transform 1 0 21528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1639504043
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_225
timestamp 1639504043
transform 1 0 21804 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1639504043
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0737_
timestamp 1639504043
transform 1 0 21160 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _0894_
timestamp 1639504043
transform 1 0 21896 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0895_
timestamp 1639504043
transform 1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1172_
timestamp 1639504043
transform 1 0 20332 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1342_
timestamp 1639504043
transform 1 0 22172 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_6_233
timestamp 1639504043
transform 1 0 22540 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_246
timestamp 1639504043
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0738_
timestamp 1639504043
transform 1 0 23276 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1146_
timestamp 1639504043
transform -1 0 24472 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1639504043
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp 1639504043
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_254
timestamp 1639504043
transform 1 0 24472 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_266
timestamp 1639504043
transform 1 0 25576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1639504043
transform -1 0 26128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1639504043
transform -1 0 26128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1639504043
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1639504043
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1639504043
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1639504043
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1639504043
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1639504043
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1639504043
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1387_
timestamp 1639504043
transform 1 0 4508 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__o221a_2  _0768_
timestamp 1639504043
transform 1 0 6072 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_A
timestamp 1639504043
transform 1 0 8004 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_63
timestamp 1639504043
transform 1 0 6900 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1639504043
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1639504043
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clk
timestamp 1639504043
transform -1 0 8004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_102
timestamp 1639504043
transform 1 0 10488 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1639504043
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1391_
timestamp 1639504043
transform -1 0 10488 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_8_114
timestamp 1639504043
transform 1 0 11592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_118
timestamp 1639504043
transform 1 0 11960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_122
timestamp 1639504043
transform 1 0 12328 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1639504043
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__A0
timestamp 1639504043
transform 1 0 13524 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_128
timestamp 1639504043
transform 1 0 12880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1639504043
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_141
timestamp 1639504043
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1639504043
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0881_
timestamp 1639504043
transform -1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1639504043
transform 1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0906_
timestamp 1639504043
transform 1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1181_
timestamp 1639504043
transform 1 0 15732 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1223_
timestamp 1639504043
transform 1 0 14904 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_172
timestamp 1639504043
transform 1 0 16928 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1639504043
transform 1 0 18032 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_clk
timestamp 1639504043
transform -1 0 16928 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp 1639504043
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_203
timestamp 1639504043
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1639504043
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0896_
timestamp 1639504043
transform 1 0 19872 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_8_211
timestamp 1639504043
transform 1 0 20516 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_221
timestamp 1639504043
transform 1 0 21436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_227
timestamp 1639504043
transform 1 0 21988 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0892_
timestamp 1639504043
transform 1 0 22080 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1145_
timestamp 1639504043
transform 1 0 20700 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1343_
timestamp 1639504043
transform 1 0 22724 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_8_261
timestamp 1639504043
transform 1 0 25116 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1639504043
transform -1 0 26128 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1639504043
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1147_
timestamp 1639504043
transform -1 0 25116 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1639504043
transform 1 0 1840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1639504043
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1639504043
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1639504043
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0871_
timestamp 1639504043
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0872_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 2484 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_9_28
timestamp 1639504043
transform 1 0 3680 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_34
timestamp 1639504043
transform 1 0 4232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0855_
timestamp 1639504043
transform 1 0 3220 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1386_
timestamp 1639504043
transform 1 0 4324 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__B1
timestamp 1639504043
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1639504043
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1639504043
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1389_
timestamp 1639504043
transform -1 0 7912 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_9_74
timestamp 1639504043
transform 1 0 7912 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1390_
timestamp 1639504043
transform -1 0 9844 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_9_95
timestamp 1639504043
transform 1 0 9844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_107
timestamp 1639504043
transform 1 0 10948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_118
timestamp 1639504043
transform 1 0 11960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1639504043
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1639504043
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _0730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 11960 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1236_
timestamp 1639504043
transform 1 0 12052 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A2
timestamp 1639504043
transform 1 0 13524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__S
timestamp 1639504043
transform 1 0 14168 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_131
timestamp 1639504043
transform 1 0 13156 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_144
timestamp 1639504043
transform 1 0 14352 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0728_
timestamp 1639504043
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0874_
timestamp 1639504043
transform 1 0 13248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0919_
timestamp 1639504043
transform 1 0 13708 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_9_156
timestamp 1639504043
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_A
timestamp 1639504043
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1639504043
transform 1 0 17848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1639504043
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0745_
timestamp 1639504043
transform -1 0 18400 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _0879_
timestamp 1639504043
transform 1 0 17204 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clk
timestamp 1639504043
transform 1 0 16836 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_191
timestamp 1639504043
transform 1 0 18676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_201
timestamp 1639504043
transform 1 0 19596 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_205
timestamp 1639504043
transform 1 0 19964 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0880_
timestamp 1639504043
transform 1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0882_
timestamp 1639504043
transform 1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_clk
timestamp 1639504043
transform 1 0 19228 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_212
timestamp 1639504043
transform 1 0 20608 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1639504043
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1639504043
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0897_
timestamp 1639504043
transform -1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_231
timestamp 1639504043
transform 1 0 22356 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_250
timestamp 1639504043
transform 1 0 24104 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1281_
timestamp 1639504043
transform 1 0 22448 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1287_
timestamp 1639504043
transform 1 0 23276 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_256
timestamp 1639504043
transform 1 0 24656 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_268
timestamp 1639504043
transform 1 0 25760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1639504043
transform -1 0 26128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0739_
timestamp 1639504043
transform 1 0 24196 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1639504043
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1639504043
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1351_
timestamp 1639504043
transform 1 0 1564 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B1
timestamp 1639504043
transform 1 0 3864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1639504043
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1639504043
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1639504043
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0772_
timestamp 1639504043
transform 1 0 4048 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1639504043
transform -1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1388_
timestamp 1639504043
transform -1 0 6440 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_1  _0766_
timestamp 1639504043
transform -1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0767_
timestamp 1639504043
transform -1 0 6992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1639504043
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _0763_
timestamp 1639504043
transform 1 0 7820 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0764_
timestamp 1639504043
transform 1 0 6992 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B1
timestamp 1639504043
transform 1 0 9752 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_96
timestamp 1639504043
transform 1 0 9936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1639504043
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0765_
timestamp 1639504043
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1394_
timestamp 1639504043
transform 1 0 10304 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_2  _0851_
timestamp 1639504043
transform 1 0 11868 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _0873_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 13156 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B1
timestamp 1639504043
transform 1 0 13156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1639504043
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _0918_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 13340 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1331_
timestamp 1639504043
transform -1 0 15640 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_10_158
timestamp 1639504043
transform 1 0 15640 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _1155_
timestamp 1639504043
transform 1 0 16192 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _0877_
timestamp 1639504043
transform 1 0 16836 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1349_
timestamp 1639504043
transform 1 0 17480 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1639504043
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_208
timestamp 1639504043
transform 1 0 20240 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1639504043
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0744_
timestamp 1639504043
transform -1 0 19780 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1152_
timestamp 1639504043
transform -1 0 20240 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_10_220
timestamp 1639504043
transform 1 0 21344 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_2  _0885_
timestamp 1639504043
transform 1 0 20424 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0886_
timestamp 1639504043
transform -1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_232
timestamp 1639504043
transform 1 0 22448 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_238
timestamp 1639504043
transform 1 0 23000 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_242
timestamp 1639504043
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1639504043
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0890_
timestamp 1639504043
transform 1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0893_
timestamp 1639504043
transform -1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1639504043
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1639504043
transform 1 0 25484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1639504043
transform -1 0 26128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1639504043
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1639504043
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1639504043
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _0869_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 2484 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_11_31
timestamp 1639504043
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0852_
timestamp 1639504043
transform -1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0853_
timestamp 1639504043
transform 1 0 3128 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B1
timestamp 1639504043
transform -1 0 6256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_43
timestamp 1639504043
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1639504043
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_61
timestamp 1639504043
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1639504043
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1639504043
transform 1 0 6808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0770_
timestamp 1639504043
transform 1 0 5244 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B1
timestamp 1639504043
transform 1 0 7636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B1
timestamp 1639504043
transform 1 0 7084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_70
timestamp 1639504043
transform 1 0 7544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_73
timestamp 1639504043
transform 1 0 7820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0759_
timestamp 1639504043
transform 1 0 7268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0760_
timestamp 1639504043
transform -1 0 9016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0761_
timestamp 1639504043
transform -1 0 8740 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B1
timestamp 1639504043
transform -1 0 9200 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_88
timestamp 1639504043
transform 1 0 9200 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_96
timestamp 1639504043
transform 1 0 9936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _0756_
timestamp 1639504043
transform 1 0 10212 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1639504043
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1639504043
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1639504043
transform 1 0 11040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0731_
timestamp 1639504043
transform 1 0 12420 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_2  _0749_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 11500 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__S
timestamp 1639504043
transform 1 0 13892 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__S
timestamp 1639504043
transform 1 0 14076 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_138
timestamp 1639504043
transform 1 0 13800 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_143
timestamp 1639504043
transform 1 0 14260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1231_
timestamp 1639504043
transform -1 0 13800 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1639504043
transform 1 0 15180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_157
timestamp 1639504043
transform 1 0 15548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0875_
timestamp 1639504043
transform -1 0 16560 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0876_
timestamp 1639504043
transform 1 0 15640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_clk
timestamp 1639504043
transform 1 0 14812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1639504043
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0746_
timestamp 1639504043
transform -1 0 17756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1284_
timestamp 1639504043
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1348_
timestamp 1639504043
transform -1 0 19320 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_11_206
timestamp 1639504043
transform 1 0 20056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1154_
timestamp 1639504043
transform 1 0 19320 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1347_
timestamp 1639504043
transform 1 0 20148 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1639504043
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0742_
timestamp 1639504043
transform -1 0 22264 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_11_230
timestamp 1639504043
transform 1 0 22264 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_245
timestamp 1639504043
transform 1 0 23644 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__and2b_2  _0889_
timestamp 1639504043
transform 1 0 23000 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1344_
timestamp 1639504043
transform 1 0 23828 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_11_264
timestamp 1639504043
transform 1 0 25392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_268
timestamp 1639504043
transform 1 0 25760 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1639504043
transform -1 0 26128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1639504043
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1639504043
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1352_
timestamp 1639504043
transform 1 0 1656 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1639504043
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1639504043
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_36
timestamp 1639504043
transform 1 0 4416 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1639504043
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _0726_
timestamp 1639504043
transform 1 0 3772 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_12_48
timestamp 1639504043
transform 1 0 5520 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_60
timestamp 1639504043
transform 1 0 6624 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_66
timestamp 1639504043
transform 1 0 7176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1393_
timestamp 1639504043
transform 1 0 7268 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_12_100
timestamp 1639504043
transform 1 0 10304 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_90
timestamp 1639504043
transform 1 0 9384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_94
timestamp 1639504043
transform 1 0 9752 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1639504043
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0754_
timestamp 1639504043
transform 1 0 9844 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0757_
timestamp 1639504043
transform -1 0 9384 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1396_
timestamp 1639504043
transform -1 0 12052 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2
timestamp 1639504043
transform 1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__B1
timestamp 1639504043
transform 1 0 12604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_122
timestamp 1639504043
transform 1 0 12328 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0748_
timestamp 1639504043
transform -1 0 12328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A2
timestamp 1639504043
transform 1 0 13524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__S
timestamp 1639504043
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_137
timestamp 1639504043
transform 1 0 13708 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1639504043
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1136_
timestamp 1639504043
transform -1 0 13524 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1227_
timestamp 1639504043
transform -1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_12_159
timestamp 1639504043
transform 1 0 15732 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_165
timestamp 1639504043
transform 1 0 16284 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1222_
timestamp 1639504043
transform -1 0 15732 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1350_
timestamp 1639504043
transform 1 0 16376 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1639504043
transform 1 0 17940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1264_
timestamp 1639504043
transform 1 0 18124 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1639504043
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1639504043
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1151_
timestamp 1639504043
transform 1 0 19964 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1153_
timestamp 1639504043
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1346_
timestamp 1639504043
transform 1 0 20700 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_12_238
timestamp 1639504043
transform 1 0 23000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0888_
timestamp 1639504043
transform 1 0 23184 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1150_
timestamp 1639504043
transform 1 0 22264 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1275_
timestamp 1639504043
transform 1 0 23460 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_266
timestamp 1639504043
transform 1 0 25576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1639504043
transform -1 0 26128 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1639504043
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0740_
timestamp 1639504043
transform 1 0 25116 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1148_
timestamp 1639504043
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1639504043
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1639504043
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1639504043
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1639504043
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1639504043
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_2  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 2300 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _0868_
timestamp 1639504043
transform 1 0 2576 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0870_
timestamp 1639504043
transform 1 0 1932 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1639504043
transform -1 0 3680 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1639504043
transform -1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0860_
timestamp 1639504043
transform -1 0 3772 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _0725_
timestamp 1639504043
transform 1 0 3956 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1639504043
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_29
timestamp 1639504043
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B1
timestamp 1639504043
transform -1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _0724_
timestamp 1639504043
transform 1 0 4692 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B1
timestamp 1639504043
transform 1 0 4508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1397_
timestamp 1639504043
transform 1 0 4784 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A1
timestamp 1639504043
transform 1 0 5520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1639504043
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1639504043
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1639504043
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1398_
timestamp 1639504043
transform 1 0 6348 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B1
timestamp 1639504043
transform -1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1639504043
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1639504043
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1639504043
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0715_
timestamp 1639504043
transform -1 0 8740 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0722_
timestamp 1639504043
transform -1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0762_
timestamp 1639504043
transform -1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B1
timestamp 1639504043
transform -1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 1639504043
transform 1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1639504043
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_96
timestamp 1639504043
transform 1 0 9936 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1639504043
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0677_
timestamp 1639504043
transform 1 0 9660 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0716_
timestamp 1639504043
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0755_
timestamp 1639504043
transform -1 0 10580 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__C1
timestamp 1639504043
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1639504043
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1639504043
transform 1 0 11684 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_108
timestamp 1639504043
transform 1 0 11040 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_120
timestamp 1639504043
transform 1 0 12144 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1639504043
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1639504043
transform 1 0 13248 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_132
timestamp 1639504043
transform 1 0 13248 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_127
timestamp 1639504043
transform 1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1639504043
transform 1 0 13064 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1226_
timestamp 1639504043
transform 1 0 14168 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1033_
timestamp 1639504043
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1032_
timestamp 1639504043
transform -1 0 14812 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1639504043
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_135
timestamp 1639504043
transform 1 0 13524 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__S
timestamp 1639504043
transform 1 0 13800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__S
timestamp 1639504043
transform 1 0 13984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A2
timestamp 1639504043
transform 1 0 13524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1639504043
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_149
timestamp 1639504043
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_155
timestamp 1639504043
transform 1 0 15364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1039_
timestamp 1639504043
transform 1 0 14904 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1221_
timestamp 1639504043
transform 1 0 14996 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1639504043
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1639504043
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_167
timestamp 1639504043
transform 1 0 16468 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_179
timestamp 1639504043
transform 1 0 17572 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1639504043
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0878_
timestamp 1639504043
transform 1 0 17296 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1272_
timestamp 1639504043
transform 1 0 17572 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_188
timestamp 1639504043
transform 1 0 18400 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_200
timestamp 1639504043
transform 1 0 19504 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1639504043
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1639504043
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1639504043
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1639504043
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0883_
timestamp 1639504043
transform 1 0 19780 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1639504043
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1639504043
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_223
timestamp 1639504043
transform 1 0 21620 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1639504043
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0743_
timestamp 1639504043
transform -1 0 21712 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0884_
timestamp 1639504043
transform -1 0 20792 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1251_
timestamp 1639504043
transform 1 0 20424 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1278_
timestamp 1639504043
transform 1 0 20792 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_233
timestamp 1639504043
transform 1 0 22540 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_235
timestamp 1639504043
transform 1 0 22724 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_243
timestamp 1639504043
transform 1 0 23460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _0887_
timestamp 1639504043
transform 1 0 22816 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1290_
timestamp 1639504043
transform 1 0 22816 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1345_
timestamp 1639504043
transform 1 0 23644 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_13_267
timestamp 1639504043
transform 1 0 25668 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1639504043
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_261
timestamp 1639504043
transform 1 0 25116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1639504043
transform -1 0 26128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1639504043
transform -1 0 26128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1639504043
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0741_
timestamp 1639504043
transform -1 0 25668 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1149_
timestamp 1639504043
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1639504043
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1639504043
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1639504043
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1354_
timestamp 1639504043
transform 1 0 1840 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__o221a_2  _0723_
timestamp 1639504043
transform 1 0 4324 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _0862_
timestamp 1639504043
transform -1 0 4048 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1639504043
transform 1 0 4048 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B1
timestamp 1639504043
transform 1 0 5980 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1639504043
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_60
timestamp 1639504043
transform 1 0 6624 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1639504043
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0717_
timestamp 1639504043
transform -1 0 6624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0719_
timestamp 1639504043
transform -1 0 5980 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_A
timestamp 1639504043
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_64
timestamp 1639504043
transform 1 0 6992 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1639504043
transform 1 0 7636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1402_
timestamp 1639504043
transform 1 0 7820 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clk
timestamp 1639504043
transform -1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1401_
timestamp 1639504043
transform 1 0 9384 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1639504043
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1639504043
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1639504043
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1639504043
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1639504043
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1374_
timestamp 1639504043
transform -1 0 13524 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1375_
timestamp 1639504043
transform -1 0 15088 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1639504043
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_2  _1040_
timestamp 1639504043
transform -1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1041_
timestamp 1639504043
transform -1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__S
timestamp 1639504043
transform 1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1639504043
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1639504043
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_174
timestamp 1639504043
transform 1 0 17112 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_186
timestamp 1639504043
transform 1 0 18216 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1639504043
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__S
timestamp 1639504043
transform 1 0 18768 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_203
timestamp 1639504043
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1177_
timestamp 1639504043
transform -1 0 19780 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1639504043
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1639504043
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1639504043
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1639504043
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__S
timestamp 1639504043
transform 1 0 23276 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1639504043
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1288_
timestamp 1639504043
transform -1 0 24288 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_252
timestamp 1639504043
transform 1 0 24288 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_264
timestamp 1639504043
transform 1 0 25392 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_268
timestamp 1639504043
transform 1 0 25760 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1639504043
transform -1 0 26128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1639504043
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1639504043
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1353_
timestamp 1639504043
transform -1 0 3220 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1639504043
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_31
timestamp 1639504043
transform 1 0 3956 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_39
timestamp 1639504043
transform 1 0 4692 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1639504043
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _0867_
timestamp 1639504043
transform -1 0 3680 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__B1
timestamp 1639504043
transform -1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_44
timestamp 1639504043
transform 1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1399_
timestamp 1639504043
transform 1 0 5336 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_16_80
timestamp 1639504043
transform 1 0 8464 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0710_
timestamp 1639504043
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1400_
timestamp 1639504043
transform 1 0 6900 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_16_102
timestamp 1639504043
transform 1 0 10488 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1639504043
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1403_
timestamp 1639504043
transform 1 0 8924 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_16_114
timestamp 1639504043
transform 1 0 11592 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _0798_
timestamp 1639504043
transform -1 0 12972 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B
timestamp 1639504043
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1639504043
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0797_
timestamp 1639504043
transform 1 0 12972 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _1031_
timestamp 1639504043
transform 1 0 14076 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__S
timestamp 1639504043
transform 1 0 16100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_150
timestamp 1639504043
transform 1 0 14904 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_160
timestamp 1639504043
transform 1 0 15824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0794_
timestamp 1639504043
transform 1 0 14996 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1179_
timestamp 1639504043
transform -1 0 17112 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clk
timestamp 1639504043
transform 1 0 14536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_183
timestamp 1639504043
transform 1 0 17940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _1058_
timestamp 1639504043
transform 1 0 18308 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1180_
timestamp 1639504043
transform 1 0 17112 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__S
timestamp 1639504043
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_193
timestamp 1639504043
transform 1 0 18860 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1639504043
transform 1 0 20056 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1639504043
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1176_
timestamp 1639504043
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__S
timestamp 1639504043
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__S
timestamp 1639504043
transform 1 0 20792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_227
timestamp 1639504043
transform 1 0 21988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1276_
timestamp 1639504043
transform 1 0 20976 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__S
timestamp 1639504043
transform 1 0 22632 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__S
timestamp 1639504043
transform 1 0 23644 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__S
timestamp 1639504043
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_233
timestamp 1639504043
transform 1 0 22540 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_247
timestamp 1639504043
transform 1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1280_
timestamp 1639504043
transform 1 0 22816 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_262
timestamp 1639504043
transform 1 0 25208 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_268
timestamp 1639504043
transform 1 0 25760 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1639504043
transform -1 0 26128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1639504043
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1289_
timestamp 1639504043
transform 1 0 24380 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_11
timestamp 1639504043
transform 1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1639504043
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1639504043
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_2  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 2392 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B1
timestamp 1639504043
transform -1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1639504043
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_37
timestamp 1639504043
transform 1 0 4508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1639504043
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp 1639504043
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_60
timestamp 1639504043
transform 1 0 6624 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1639504043
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0718_
timestamp 1639504043
transform -1 0 6624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_clk
timestamp 1639504043
transform -1 0 5520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B1
timestamp 1639504043
transform 1 0 7728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_83
timestamp 1639504043
transform 1 0 8740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _0714_
timestamp 1639504043
transform 1 0 7912 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1404_
timestamp 1639504043
transform 1 0 9292 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_clk
timestamp 1639504043
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1639504043
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1639504043
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1405_
timestamp 1639504043
transform 1 0 11500 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_A
timestamp 1639504043
transform 1 0 14352 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_130
timestamp 1639504043
transform 1 0 13064 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1639504043
transform 1 0 14168 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_146
timestamp 1639504043
transform 1 0 14536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_150
timestamp 1639504043
transform 1 0 14904 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1377_
timestamp 1639504043
transform 1 0 14996 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1639504043
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1047_
timestamp 1639504043
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1173_
timestamp 1639504043
transform 1 0 17756 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1174_
timestamp 1639504043
transform 1 0 16928 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1052_
timestamp 1639504043
transform 1 0 18584 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1059_
timestamp 1639504043
transform 1 0 19872 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1262_
timestamp 1639504043
transform -1 0 19872 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__S
timestamp 1639504043
transform 1 0 20608 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_211
timestamp 1639504043
transform 1 0 20516 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1639504043
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1639504043
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1170_
timestamp 1639504043
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1171_
timestamp 1639504043
transform 1 0 20792 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__S
timestamp 1639504043
transform 1 0 22724 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_234
timestamp 1639504043
transform 1 0 22632 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1279_
timestamp 1639504043
transform 1 0 22908 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1286_
timestamp 1639504043
transform 1 0 23736 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_255
timestamp 1639504043
transform 1 0 24564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_267
timestamp 1639504043
transform 1 0 25668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1639504043
transform -1 0 26128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1639504043
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1639504043
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1639504043
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1639504043
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1639504043
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1639504043
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1639504043
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_53
timestamp 1639504043
transform 1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_61
timestamp 1639504043
transform 1 0 6716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1639504043
transform 1 0 7176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_78
timestamp 1639504043
transform 1 0 8280 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1639504043
transform 1 0 6900 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0713_
timestamp 1639504043
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B1
timestamp 1639504043
transform 1 0 10304 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_102
timestamp 1639504043
transform 1 0 10488 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1639504043
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0706_
timestamp 1639504043
transform -1 0 10304 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0711_
timestamp 1639504043
transform -1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0712_
timestamp 1639504043
transform -1 0 9752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__B1
timestamp 1639504043
transform -1 0 11040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1639504043
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1639504043
transform 1 0 12236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_125
timestamp 1639504043
transform 1 0 12604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0709_
timestamp 1639504043
transform 1 0 11040 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0775_
timestamp 1639504043
transform -1 0 12604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_132
timestamp 1639504043
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 1639504043
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1639504043
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0792_
timestamp 1639504043
transform 1 0 12696 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0793_
timestamp 1639504043
transform 1 0 12972 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_149
timestamp 1639504043
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_159
timestamp 1639504043
transform 1 0 15732 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0796_
timestamp 1639504043
transform 1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _1046_
timestamp 1639504043
transform -1 0 16744 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__S
timestamp 1639504043
transform 1 0 17572 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__S
timestamp 1639504043
transform 1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_177
timestamp 1639504043
transform 1 0 17388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_181
timestamp 1639504043
transform 1 0 17756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1045_
timestamp 1639504043
transform 1 0 16744 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1053_
timestamp 1639504043
transform 1 0 17940 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__S
timestamp 1639504043
transform 1 0 18860 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1639504043
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_206
timestamp 1639504043
transform 1 0 20056 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1639504043
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1639504043
transform 1 0 18584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1066_
timestamp 1639504043
transform -1 0 20884 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1263_
timestamp 1639504043
transform 1 0 19228 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__S
timestamp 1639504043
transform 1 0 22172 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1065_
timestamp 1639504043
transform 1 0 21712 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1277_
timestamp 1639504043
transform 1 0 20884 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__S
timestamp 1639504043
transform 1 0 23644 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__S
timestamp 1639504043
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1639504043
transform 1 0 22356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_236
timestamp 1639504043
transform 1 0 22816 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_244
timestamp 1639504043
transform 1 0 23552 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_247
timestamp 1639504043
transform 1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1075_
timestamp 1639504043
transform 1 0 22540 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_262
timestamp 1639504043
transform 1 0 25208 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_268
timestamp 1639504043
transform 1 0 25760 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1639504043
transform -1 0 26128 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1639504043
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1285_
timestamp 1639504043
transform 1 0 24380 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1639504043
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1639504043
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1639504043
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1639504043
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1639504043
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1365_
timestamp 1639504043
transform -1 0 3036 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1367_
timestamp 1639504043
transform 1 0 1840 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1235_
timestamp 1639504043
transform 1 0 3404 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1233_
timestamp 1639504043
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1639504043
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1639504043
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1639504043
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0812_
timestamp 1639504043
transform -1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_41
timestamp 1639504043
transform 1 0 4876 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_38
timestamp 1639504043
transform 1 0 4600 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_34
timestamp 1639504043
transform 1 0 4232 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1370_
timestamp 1639504043
transform 1 0 4692 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1639504043
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0806_
timestamp 1639504043
transform -1 0 7084 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0807_
timestamp 1639504043
transform -1 0 6256 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1371_
timestamp 1639504043
transform 1 0 6348 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_19_74
timestamp 1639504043
transform 1 0 7912 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_82
timestamp 1639504043
transform 1 0 8648 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_74
timestamp 1639504043
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1639504043
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1225_
timestamp 1639504043
transform 1 0 7084 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _0773_
timestamp 1639504043
transform 1 0 9660 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0696_
timestamp 1639504043
transform 1 0 9476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _0692_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 9660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0691_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 9016 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1639504043
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A
timestamp 1639504043
transform -1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _0801_
timestamp 1639504043
transform -1 0 11316 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_101
timestamp 1639504043
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_94
timestamp 1639504043
transform 1 0 9752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A1
timestamp 1639504043
transform 1 0 10212 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1372_
timestamp 1639504043
transform -1 0 11408 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_19_116
timestamp 1639504043
transform 1 0 11776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1639504043
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0703_
timestamp 1639504043
transform 1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0704_
timestamp 1639504043
transform 1 0 12144 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0707_
timestamp 1639504043
transform 1 0 11316 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0708_
timestamp 1639504043
transform 1 0 12144 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1639504043
transform -1 0 12696 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0777_
timestamp 1639504043
transform -1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B1
timestamp 1639504043
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1639504043
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_145
timestamp 1639504043
transform 1 0 14444 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1639504043
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0695_
timestamp 1639504043
transform 1 0 14444 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0799_
timestamp 1639504043
transform 1 0 12972 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1373_
timestamp 1639504043
transform -1 0 14444 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_clk
timestamp 1639504043
transform -1 0 14444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_151
timestamp 1639504043
transform 1 0 14996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_163
timestamp 1639504043
transform 1 0 16100 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0795_
timestamp 1639504043
transform 1 0 14720 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1376_
timestamp 1639504043
transform 1 0 14996 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__S
timestamp 1639504043
transform 1 0 17756 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__S
timestamp 1639504043
transform 1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1639504043
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_183
timestamp 1639504043
transform 1 0 17940 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_171
timestamp 1639504043
transform 1 0 16836 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1639504043
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1639504043
transform -1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1271_
timestamp 1639504043
transform 1 0 17940 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1283_
timestamp 1639504043
transform 1 0 17112 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__S
timestamp 1639504043
transform 1 0 20240 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__S
timestamp 1639504043
transform 1 0 19044 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_189
timestamp 1639504043
transform 1 0 18492 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_197
timestamp 1639504043
transform 1 0 19228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1639504043
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1639504043
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_205
timestamp 1639504043
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1639504043
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1250_
timestamp 1639504043
transform 1 0 20516 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1249_
timestamp 1639504043
transform -1 0 21252 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__S
timestamp 1639504043
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__or4_2  _1102_
timestamp 1639504043
transform -1 0 21988 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1074_
timestamp 1639504043
transform -1 0 22816 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1073_
timestamp 1639504043
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1072_
timestamp 1639504043
transform 1 0 21988 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1067_
timestamp 1639504043
transform 1 0 21344 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1639504043
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1639504043
transform 1 0 21252 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1639504043
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__S
timestamp 1639504043
transform 1 0 22816 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_232
timestamp 1639504043
transform 1 0 22448 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_236
timestamp 1639504043
transform 1 0 22816 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1639504043
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_2  _1082_
timestamp 1639504043
transform 1 0 23460 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1088_
timestamp 1639504043
transform 1 0 22908 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1273_
timestamp 1639504043
transform 1 0 23828 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1274_
timestamp 1639504043
transform -1 0 23828 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_256
timestamp 1639504043
transform 1 0 24656 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_268
timestamp 1639504043
transform 1 0 25760 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_263
timestamp 1639504043
transform 1 0 25300 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1639504043
transform -1 0 26128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1639504043
transform -1 0 26128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1639504043
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1639504043
transform 1 0 25024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1089_
timestamp 1639504043
transform -1 0 25024 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_21_15
timestamp 1639504043
transform 1 0 2484 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1639504043
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1639504043
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0813_
timestamp 1639504043
transform -1 0 3588 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_27
timestamp 1639504043
transform 1 0 3588 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1639504043
transform -1 0 4784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0811_
timestamp 1639504043
transform -1 0 5060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1200_
timestamp 1639504043
transform 1 0 3680 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_46
timestamp 1639504043
transform 1 0 5336 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1639504043
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0800_
timestamp 1639504043
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0804_
timestamp 1639504043
transform 1 0 5060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0805_
timestamp 1639504043
transform 1 0 5704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0809_
timestamp 1639504043
transform -1 0 5704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1199_
timestamp 1639504043
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1639504043
transform -1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__B
timestamp 1639504043
transform -1 0 8372 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_79
timestamp 1639504043
transform 1 0 8372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1639504043
transform 1 0 8648 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1256_
timestamp 1639504043
transform 1 0 7176 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1639504043
transform 1 0 9844 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A
timestamp 1639504043
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A
timestamp 1639504043
transform 1 0 10028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_101
timestamp 1639504043
transform 1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0693_
timestamp 1639504043
transform -1 0 9384 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0802_
timestamp 1639504043
transform -1 0 9844 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B1
timestamp 1639504043
transform 1 0 11132 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1639504043
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1639504043
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1407_
timestamp 1639504043
transform 1 0 11500 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1406_
timestamp 1639504043
transform 1 0 13064 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_21_150
timestamp 1639504043
transform 1 0 14904 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0788_
timestamp 1639504043
transform 1 0 14628 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1409_
timestamp 1639504043
transform 1 0 14996 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__S
timestamp 1639504043
transform -1 0 17296 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__S
timestamp 1639504043
transform -1 0 17112 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_169
timestamp 1639504043
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1639504043
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1270_
timestamp 1639504043
transform 1 0 18124 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1282_
timestamp 1639504043
transform 1 0 17296 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1639504043
transform 1 0 19412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _1056_
timestamp 1639504043
transform -1 0 19412 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1108_
timestamp 1639504043
transform -1 0 20608 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1114_
timestamp 1639504043
transform -1 0 20148 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1639504043
transform 1 0 20608 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1639504043
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1639504043
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1639504043
transform 1 0 20792 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1101_
timestamp 1639504043
transform 1 0 21068 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1103_
timestamp 1639504043
transform -1 0 22448 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_21_232
timestamp 1639504043
transform 1 0 22448 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1081_
timestamp 1639504043
transform -1 0 24288 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1095_
timestamp 1639504043
transform -1 0 23828 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_21_255
timestamp 1639504043
transform 1 0 24564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_267
timestamp 1639504043
transform 1 0 25668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1639504043
transform -1 0 26128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1639504043
transform 1 0 24288 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1639504043
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1639504043
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1639504043
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0815_
timestamp 1639504043
transform -1 0 3404 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1639504043
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1639504043
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1366_
timestamp 1639504043
transform 1 0 3772 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_22_46
timestamp 1639504043
transform 1 0 5336 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0808_
timestamp 1639504043
transform 1 0 6440 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0810_
timestamp 1639504043
transform 1 0 5612 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1639504043
transform 1 0 8096 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__or3_2  _0689_
timestamp 1639504043
transform -1 0 8832 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1230_
timestamp 1639504043
transform 1 0 7268 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__C
timestamp 1639504043
transform -1 0 9844 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_95
timestamp 1639504043
transform 1 0 9844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1639504043
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_2  _0688_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__B1
timestamp 1639504043
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1639504043
transform 1 0 10948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 1639504043
transform 1 0 11316 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0705_
timestamp 1639504043
transform 1 0 11592 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1408_
timestamp 1639504043
transform 1 0 12420 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1639504043
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1639504043
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0701_
timestamp 1639504043
transform 1 0 14168 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0702_
timestamp 1639504043
transform 1 0 14996 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0790_
timestamp 1639504043
transform 1 0 15824 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B1
timestamp 1639504043
transform -1 0 16836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_171
timestamp 1639504043
transform 1 0 16836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_183
timestamp 1639504043
transform 1 0 17940 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1121_
timestamp 1639504043
transform -1 0 18768 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1639504043
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1639504043
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1639504043
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1109_
timestamp 1639504043
transform -1 0 20700 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1115_
timestamp 1639504043
transform -1 0 20056 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_22_213
timestamp 1639504043
transform 1 0 20700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_225
timestamp 1639504043
transform 1 0 21804 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_237
timestamp 1639504043
transform 1 0 22908 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_246
timestamp 1639504043
transform 1 0 23736 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1086_
timestamp 1639504043
transform 1 0 23828 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1094_
timestamp 1639504043
transform -1 0 23736 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_22_256
timestamp 1639504043
transform 1 0 24656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_268
timestamp 1639504043
transform 1 0 25760 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1639504043
transform -1 0 26128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1639504043
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1639504043
transform 1 0 24380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1639504043
transform 1 0 1380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1639504043
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1364_
timestamp 1639504043
transform -1 0 3036 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1639504043
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _0814_
timestamp 1639504043
transform 1 0 3404 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1269_
timestamp 1639504043
transform 1 0 4232 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A1
timestamp 1639504043
transform 1 0 6440 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A0
timestamp 1639504043
transform 1 0 5060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1639504043
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1639504043
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1639504043
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1639504043
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1369_
timestamp 1639504043
transform 1 0 6624 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B
timestamp 1639504043
transform 1 0 8740 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_77
timestamp 1639504043
transform 1 0 8188 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_88
timestamp 1639504043
transform 1 0 9200 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0769_
timestamp 1639504043
transform 1 0 8924 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0779_
timestamp 1639504043
transform 1 0 9936 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A1
timestamp 1639504043
transform 1 0 10764 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1639504043
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1639504043
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1639504043
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_125
timestamp 1639504043
transform 1 0 12604 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1639504043
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1639504043
transform 1 0 12696 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 12880 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _0787_
timestamp 1639504043
transform -1 0 14996 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1410_
timestamp 1639504043
transform 1 0 14996 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__S
timestamp 1639504043
transform 1 0 18216 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1639504043
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1379_
timestamp 1639504043
transform 1 0 16652 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__S
timestamp 1639504043
transform 1 0 19964 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_197
timestamp 1639504043
transform 1 0 19228 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_203
timestamp 1639504043
transform 1 0 19780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__and2_2  _1063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform -1 0 20700 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1639504043
transform 1 0 19504 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1186_
timestamp 1639504043
transform -1 0 19228 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A
timestamp 1639504043
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1639504043
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1639504043
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1639504043
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1639504043
transform 1 0 21160 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1112_
timestamp 1639504043
transform -1 0 21160 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A
timestamp 1639504043
transform 1 0 23644 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_237
timestamp 1639504043
transform 1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_247
timestamp 1639504043
transform 1 0 23828 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1092_
timestamp 1639504043
transform 1 0 23920 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1099_
timestamp 1639504043
transform -1 0 23644 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A
timestamp 1639504043
transform -1 0 24656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__S
timestamp 1639504043
transform 1 0 24656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_258
timestamp 1639504043
transform 1 0 24840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_266
timestamp 1639504043
transform 1 0 25576 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1639504043
transform -1 0 26128 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_15
timestamp 1639504043
transform 1 0 2484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1639504043
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1639504043
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0817_
timestamp 1639504043
transform -1 0 3588 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__C1
timestamp 1639504043
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1639504043
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_31
timestamp 1639504043
transform 1 0 3956 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1639504043
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_43
timestamp 1639504043
transform 1 0 5060 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1368_
timestamp 1639504043
transform 1 0 5612 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A
timestamp 1639504043
transform 1 0 8004 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A1
timestamp 1639504043
transform 1 0 7268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_66
timestamp 1639504043
transform 1 0 7176 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_69
timestamp 1639504043
transform 1 0 7452 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1639504043
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _0753_
timestamp 1639504043
transform -1 0 8648 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1639504043
transform 1 0 9660 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1639504043
transform 1 0 10028 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1639504043
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _0752_
timestamp 1639504043
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1385_
timestamp 1639504043
transform 1 0 10120 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_24_118
timestamp 1639504043
transform 1 0 11960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_125
timestamp 1639504043
transform 1 0 12604 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0699_
timestamp 1639504043
transform 1 0 11684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0776_
timestamp 1639504043
transform -1 0 12328 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0778_
timestamp 1639504043
transform -1 0 12604 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1639504043
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1639504043
transform 1 0 14352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1639504043
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0697_
timestamp 1639504043
transform 1 0 13340 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0784_
timestamp 1639504043
transform 1 0 13616 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0785_
timestamp 1639504043
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B1
timestamp 1639504043
transform -1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_148
timestamp 1639504043
transform 1 0 14720 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_151
timestamp 1639504043
transform 1 0 14996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_163
timestamp 1639504043
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_175
timestamp 1639504043
transform 1 0 17204 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_183
timestamp 1639504043
transform 1 0 17940 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1120_
timestamp 1639504043
transform -1 0 18676 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__S
timestamp 1639504043
transform -1 0 19136 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_206
timestamp 1639504043
transform 1 0 20056 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1639504043
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1064_
timestamp 1639504043
transform 1 0 20148 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1122_
timestamp 1639504043
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1187_
timestamp 1639504043
transform -1 0 20056 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__S
timestamp 1639504043
transform 1 0 22080 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1252_
timestamp 1639504043
transform 1 0 20424 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1259_
timestamp 1639504043
transform 1 0 21252 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__S
timestamp 1639504043
transform 1 0 22448 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__S
timestamp 1639504043
transform 1 0 22264 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1071_
timestamp 1639504043
transform 1 0 22632 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1079_
timestamp 1639504043
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1237_
timestamp 1639504043
transform 1 0 22908 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__S
timestamp 1639504043
transform -1 0 25668 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_267
timestamp 1639504043
transform 1 0 25668 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1639504043
transform -1 0 26128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1639504043
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1093_
timestamp 1639504043
transform -1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1240_
timestamp 1639504043
transform 1 0 24380 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1639504043
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1639504043
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1639504043
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0671_
timestamp 1639504043
transform -1 0 3680 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_28
timestamp 1639504043
transform 1 0 3680 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_40
timestamp 1639504043
transform 1 0 4784 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1639504043
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1639504043
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1639504043
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1639504043
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1395_
timestamp 1639504043
transform 1 0 7820 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1639504043
transform -1 0 10120 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_102
timestamp 1639504043
transform 1 0 10488 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_98
timestamp 1639504043
transform 1 0 10120 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1639504043
transform -1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0721_
timestamp 1639504043
transform -1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1639504043
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0780_
timestamp 1639504043
transform 1 0 10212 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1639504043
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1639504043
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_121
timestamp 1639504043
transform 1 0 12236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1639504043
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0783_
timestamp 1639504043
transform 1 0 12420 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__B1
timestamp 1639504043
transform -1 0 14168 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A1
timestamp 1639504043
transform 1 0 13248 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_134
timestamp 1639504043
transform 1 0 13432 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _0700_
timestamp 1639504043
transform 1 0 14168 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_25_151
timestamp 1639504043
transform 1 0 14996 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_157
timestamp 1639504043
transform 1 0 15548 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0789_
timestamp 1639504043
transform 1 0 15640 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1639504043
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_186
timestamp 1639504043
transform 1 0 18216 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1639504043
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1380_
timestamp 1639504043
transform 1 0 16652 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__S
timestamp 1639504043
transform 1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__S
timestamp 1639504043
transform 1 0 19596 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_198
timestamp 1639504043
transform 1 0 19320 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1260_
timestamp 1639504043
transform -1 0 20792 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1639504043
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_225
timestamp 1639504043
transform 1 0 21804 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1639504043
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1070_
timestamp 1639504043
transform 1 0 21896 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1244_
timestamp 1639504043
transform 1 0 20792 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1196_
timestamp 1639504043
transform -1 0 24932 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1241_
timestamp 1639504043
transform -1 0 24104 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1265_
timestamp 1639504043
transform -1 0 23276 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_268
timestamp 1639504043
transform 1 0 25760 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1639504043
transform -1 0 26128 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1246_
timestamp 1639504043
transform 1 0 24932 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1639504043
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1639504043
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1639504043
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1639504043
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1639504043
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1420_
timestamp 1639504043
transform 1 0 1840 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1421_
timestamp 1639504043
transform 1 0 2116 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_27_25
timestamp 1639504043
transform 1 0 3404 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1639504043
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0673_
timestamp 1639504043
transform -1 0 4600 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1419_
timestamp 1639504043
transform 1 0 3496 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1423_
timestamp 1639504043
transform 1 0 4600 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A
timestamp 1639504043
transform 1 0 6808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_55
timestamp 1639504043
transform 1 0 6164 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1639504043
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1639504043
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1639504043
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0674_
timestamp 1639504043
transform -1 0 6164 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0675_
timestamp 1639504043
transform -1 0 5888 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clk
timestamp 1639504043
transform -1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A2
timestamp 1639504043
transform 1 0 8096 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_A
timestamp 1639504043
transform 1 0 6992 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_67
timestamp 1639504043
transform 1 0 7268 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_66
timestamp 1639504043
transform 1 0 7176 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_74
timestamp 1639504043
transform 1 0 7912 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _0679_
timestamp 1639504043
transform -1 0 9476 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1268_
timestamp 1639504043
transform -1 0 8832 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_clk
timestamp 1639504043
transform 1 0 8280 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A1
timestamp 1639504043
transform 1 0 9568 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_91
timestamp 1639504043
transform 1 0 9476 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1639504043
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0678_
timestamp 1639504043
transform -1 0 10764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0680_
timestamp 1639504043
transform 1 0 10580 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0681_
timestamp 1639504043
transform -1 0 10580 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1418_
timestamp 1639504043
transform 1 0 8924 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1639504043
transform 1 0 10764 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_117
timestamp 1639504043
transform 1 0 11868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1639504043
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1382_
timestamp 1639504043
transform 1 0 12420 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1417_
timestamp 1639504043
transform 1 0 11500 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1639504043
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1639504043
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_130
timestamp 1639504043
transform 1 0 13064 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_142
timestamp 1639504043
transform 1 0 14168 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1639504043
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B1
timestamp 1639504043
transform -1 0 15364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_150
timestamp 1639504043
transform 1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_155
timestamp 1639504043
transform 1 0 15364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _0791_
timestamp 1639504043
transform 1 0 16100 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1411_
timestamp 1639504043
transform 1 0 14536 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__S
timestamp 1639504043
transform 1 0 17940 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1639504043
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_185
timestamp 1639504043
transform 1 0 18124 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1639504043
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1639504043
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1127_
timestamp 1639504043
transform -1 0 17940 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1130_
timestamp 1639504043
transform -1 0 18676 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1378_
timestamp 1639504043
transform 1 0 16652 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1210_
timestamp 1639504043
transform -1 0 20056 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1118_
timestamp 1639504043
transform 1 0 18676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1639504043
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1639504043
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__S
timestamp 1639504043
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A
timestamp 1639504043
transform 1 0 18676 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1253_
timestamp 1639504043
transform 1 0 19872 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1119_
timestamp 1639504043
transform -1 0 19872 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1062_
timestamp 1639504043
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__S
timestamp 1639504043
transform 1 0 19412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1243_
timestamp 1639504043
transform 1 0 20976 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1107_
timestamp 1639504043
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1106_
timestamp 1639504043
transform 1 0 20516 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1639504043
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__S
timestamp 1639504043
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1238_
timestamp 1639504043
transform -1 0 22632 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1639504043
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_227
timestamp 1639504043
transform 1 0 21988 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1639504043
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1639504043
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__S
timestamp 1639504043
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1266_
timestamp 1639504043
transform 1 0 22632 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_238
timestamp 1639504043
transform 1 0 23000 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_234
timestamp 1639504043
transform 1 0 22632 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_231
timestamp 1639504043
transform 1 0 22356 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__S
timestamp 1639504043
transform 1 0 22448 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__S
timestamp 1639504043
transform 1 0 23092 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1247_
timestamp 1639504043
transform 1 0 23460 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_247
timestamp 1639504043
transform 1 0 23828 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_243
timestamp 1639504043
transform 1 0 23460 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__S
timestamp 1639504043
transform 1 0 23276 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__S
timestamp 1639504043
transform 1 0 23920 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_250
timestamp 1639504043
transform 1 0 24104 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1197_
timestamp 1639504043
transform -1 0 25208 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1080_
timestamp 1639504043
transform 1 0 24196 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1639504043
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__S
timestamp 1639504043
transform 1 0 24472 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1639504043
transform -1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1639504043
transform -1 0 26128 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1639504043
transform -1 0 26128 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_268
timestamp 1639504043
transform 1 0 25760 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_267
timestamp 1639504043
transform 1 0 25668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1639504043
transform 1 0 25484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_256
timestamp 1639504043
transform 1 0 24656 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1639504043
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1639504043
transform 1 0 1932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1639504043
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1422_
timestamp 1639504043
transform 1 0 2024 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1639504043
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1639504043
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1639504043
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0669_
timestamp 1639504043
transform 1 0 4324 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_clk
timestamp 1639504043
transform -1 0 4324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_44
timestamp 1639504043
transform 1 0 5152 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_49
timestamp 1639504043
transform 1 0 5612 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0657_
timestamp 1639504043
transform -1 0 5612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1424_
timestamp 1639504043
transform 1 0 5704 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_28_67
timestamp 1639504043
transform 1 0 7268 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1639504043
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1639504043
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1639504043
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0782_
timestamp 1639504043
transform -1 0 11316 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1416_
timestamp 1639504043
transform 1 0 8924 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_28_111
timestamp 1639504043
transform 1 0 11316 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1415_
timestamp 1639504043
transform 1 0 11500 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1639504043
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp 1639504043
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1639504043
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0698_
timestamp 1639504043
transform 1 0 14352 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0781_
timestamp 1639504043
transform 1 0 13064 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1412_
timestamp 1639504043
transform 1 0 15180 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_2  _1126_
timestamp 1639504043
transform 1 0 17572 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1183_
timestamp 1639504043
transform 1 0 18032 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1208_
timestamp 1639504043
transform 1 0 16744 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_206
timestamp 1639504043
transform 1 0 20056 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1639504043
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1125_
timestamp 1639504043
transform -1 0 19136 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1211_
timestamp 1639504043
transform 1 0 19228 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_218
timestamp 1639504043
transform 1 0 21160 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_230
timestamp 1639504043
transform 1 0 22264 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_242
timestamp 1639504043
transform 1 0 23368 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1639504043
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1639504043
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_265
timestamp 1639504043
transform 1 0 25484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1639504043
transform -1 0 26128 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1639504043
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1639504043
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1639504043
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1639504043
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0672_
timestamp 1639504043
transform -1 0 3680 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_28
timestamp 1639504043
transform 1 0 3680 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0665_
timestamp 1639504043
transform 1 0 4600 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0666_
timestamp 1639504043
transform -1 0 4324 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0668_
timestamp 1639504043
transform 1 0 3772 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0670_
timestamp 1639504043
transform -1 0 4600 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1639504043
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0664_
timestamp 1639504043
transform 1 0 5428 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1425_
timestamp 1639504043
transform 1 0 6348 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_29_74
timestamp 1639504043
transform 1 0 7912 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_82
timestamp 1639504043
transform 1 0 8648 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 8096 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A1
timestamp 1639504043
transform 1 0 9568 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_90
timestamp 1639504043
transform 1 0 9384 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1639504043
transform 1 0 9752 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A2
timestamp 1639504043
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_106
timestamp 1639504043
transform 1 0 10856 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_122
timestamp 1639504043
transform 1 0 12328 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1639504043
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0685_
timestamp 1639504043
transform 1 0 11500 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_130
timestamp 1639504043
transform 1 0 13064 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1384_
timestamp 1639504043
transform 1 0 13340 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1639504043
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _0786_
timestamp 1639504043
transform 1 0 14904 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_clk
timestamp 1639504043
transform -1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__S
timestamp 1639504043
transform 1 0 16928 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__S
timestamp 1639504043
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1639504043
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_171
timestamp 1639504043
transform 1 0 16836 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1639504043
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1124_
timestamp 1639504043
transform 1 0 18216 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1639504043
transform -1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1184_
timestamp 1639504043
transform 1 0 17388 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__S
timestamp 1639504043
transform 1 0 19136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_198
timestamp 1639504043
transform 1 0 19320 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_clk
timestamp 1639504043
transform 1 0 18768 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__S
timestamp 1639504043
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_210
timestamp 1639504043
transform 1 0 20424 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_217
timestamp 1639504043
transform 1 0 21068 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_221
timestamp 1639504043
transform 1 0 21436 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1639504043
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0951_
timestamp 1639504043
transform 1 0 20792 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0952_
timestamp 1639504043
transform 1 0 21160 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1239_
timestamp 1639504043
transform 1 0 21804 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__S
timestamp 1639504043
transform 1 0 23276 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_234
timestamp 1639504043
transform 1 0 22632 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_240
timestamp 1639504043
transform 1 0 23184 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_243
timestamp 1639504043
transform 1 0 23460 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1320_
timestamp 1639504043
transform 1 0 24012 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_29_266
timestamp 1639504043
transform 1 0 25576 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1639504043
transform -1 0 26128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1639504043
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1639504043
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1639504043
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1639504043
transform -1 0 4232 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1639504043
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp 1639504043
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_34
timestamp 1639504043
transform 1 0 4232 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1639504043
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0658_
timestamp 1639504043
transform 1 0 5336 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1426_
timestamp 1639504043
transform 1 0 5612 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1639504043
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1305_
timestamp 1639504043
transform 1 0 7176 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_30_102
timestamp 1639504043
transform 1 0 10488 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1639504043
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1383_
timestamp 1639504043
transform -1 0 10488 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_30_114
timestamp 1639504043
transform 1 0 11592 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0667_
timestamp 1639504043
transform -1 0 11592 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0684_
timestamp 1639504043
transform 1 0 11040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1414_
timestamp 1639504043
transform 1 0 11776 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1639504043
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1639504043
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1639504043
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1639504043
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1381_
timestamp 1639504043
transform 1 0 14260 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_A
timestamp 1639504043
transform 1 0 16100 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_160
timestamp 1639504043
transform 1 0 15824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clk
timestamp 1639504043
transform -1 0 16652 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__S
timestamp 1639504043
transform 1 0 17112 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_169
timestamp 1639504043
transform 1 0 16652 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_173
timestamp 1639504043
transform 1 0 17020 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_185
timestamp 1639504043
transform 1 0 18124 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1207_
timestamp 1639504043
transform 1 0 17296 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1639504043
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 1639504043
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_205
timestamp 1639504043
transform 1 0 19964 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1639504043
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _0950_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 20056 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1321_
timestamp 1639504043
transform 1 0 20792 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_30_231
timestamp 1639504043
transform 1 0 22356 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _0953_
timestamp 1639504043
transform 1 0 22724 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1242_
timestamp 1639504043
transform 1 0 23460 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__S
timestamp 1639504043
transform -1 0 25668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_267
timestamp 1639504043
transform 1 0 25668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1639504043
transform -1 0 26128 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1639504043
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0956_
timestamp 1639504043
transform -1 0 25484 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1198_
timestamp 1639504043
transform 1 0 24380 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1639504043
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1639504043
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1356_
timestamp 1639504043
transform 1 0 2116 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1639504043
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0842_
timestamp 1639504043
transform -1 0 4692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0850_
timestamp 1639504043
transform 1 0 3680 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1639504043
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1639504043
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1639504043
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0663_
timestamp 1639504043
transform -1 0 7176 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_31_74
timestamp 1639504043
transform 1 0 7912 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_80
timestamp 1639504043
transform 1 0 8464 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1639504043
transform -1 0 7912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0987_
timestamp 1639504043
transform 1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0988_
timestamp 1639504043
transform 1 0 7176 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A1
timestamp 1639504043
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_101
timestamp 1639504043
transform 1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1306_
timestamp 1639504043
transform 1 0 8832 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A1
timestamp 1639504043
transform 1 0 12328 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_124
timestamp 1639504043
transform 1 0 12512 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1639504043
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0683_
timestamp 1639504043
transform -1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0686_
timestamp 1639504043
transform 1 0 11500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0720_
timestamp 1639504043
transform -1 0 11408 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_143
timestamp 1639504043
transform 1 0 14260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1413_
timestamp 1639504043
transform 1 0 12696 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__S
timestamp 1639504043
transform 1 0 14904 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_149
timestamp 1639504043
transform 1 0 14812 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_152
timestamp 1639504043
transform 1 0 15088 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1639504043
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _0940_
timestamp 1639504043
transform 1 0 15364 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1639504043
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1639504043
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1639504043
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1639504043
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1117_
timestamp 1639504043
transform -1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_193
timestamp 1639504043
transform 1 0 18860 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1639504043
transform 1 0 19412 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_203
timestamp 1639504043
transform 1 0 19780 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0942_
timestamp 1639504043
transform -1 0 19780 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0948_
timestamp 1639504043
transform 1 0 19872 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1639504043
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1639504043
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0949_
timestamp 1639504043
transform -1 0 21712 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1098_
timestamp 1639504043
transform 1 0 21896 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1245_
timestamp 1639504043
transform 1 0 20608 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_248
timestamp 1639504043
transform 1 0 23920 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__and3b_2  _0955_
timestamp 1639504043
transform 1 0 23184 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1104_
timestamp 1639504043
transform -1 0 23184 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1319_
timestamp 1639504043
transform 1 0 24104 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_31_267
timestamp 1639504043
transform 1 0 25668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1639504043
transform -1 0 26128 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1639504043
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1639504043
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1357_
timestamp 1639504043
transform 1 0 1472 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1639504043
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1639504043
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0847_
timestamp 1639504043
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _0848_
timestamp 1639504043
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0849_
timestamp 1639504043
transform 1 0 4508 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B1
timestamp 1639504043
transform 1 0 6256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_43
timestamp 1639504043
transform 1 0 5060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_55
timestamp 1639504043
transform 1 0 6164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_58
timestamp 1639504043
transform 1 0 6440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_62
timestamp 1639504043
transform 1 0 6808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1639504043
transform 1 0 7176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1639504043
transform 1 0 7360 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1639504043
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0662_
timestamp 1639504043
transform -1 0 7176 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1639504043
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_97
timestamp 1639504043
transform 1 0 10028 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1639504043
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A
timestamp 1639504043
transform 1 0 10948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_105
timestamp 1639504043
transform 1 0 10764 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1639504043
transform 1 0 11132 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0660_
timestamp 1639504043
transform 1 0 11408 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0682_
timestamp 1639504043
transform -1 0 11960 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0687_
timestamp 1639504043
transform 1 0 11960 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_130
timestamp 1639504043
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1639504043
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1639504043
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1639504043
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0661_
timestamp 1639504043
transform -1 0 13064 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0938_
timestamp 1639504043
transform 1 0 14352 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__S
timestamp 1639504043
transform 1 0 16376 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1639504043
transform 1 0 15916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1639504043
transform 1 0 16100 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1209_
timestamp 1639504043
transform 1 0 15088 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__S
timestamp 1639504043
transform 1 0 17848 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_177
timestamp 1639504043
transform 1 0 17388 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_181
timestamp 1639504043
transform 1 0 17756 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _0943_
timestamp 1639504043
transform 1 0 18032 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1185_
timestamp 1639504043
transform 1 0 16560 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1639504043
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_208
timestamp 1639504043
transform 1 0 20240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1639504043
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0944_
timestamp 1639504043
transform 1 0 18768 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0945_
timestamp 1639504043
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0946_
timestamp 1639504043
transform 1 0 19964 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__S
timestamp 1639504043
transform 1 0 20424 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1639504043
transform 1 0 20608 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1322_
timestamp 1639504043
transform 1 0 20792 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__a21bo_2  _1091_
timestamp 1639504043
transform 1 0 23552 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1097_
timestamp 1639504043
transform -1 0 23552 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1105_
timestamp 1639504043
transform 1 0 22356 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_266
timestamp 1639504043
transform 1 0 25576 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1639504043
transform -1 0 26128 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1639504043
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1084_
timestamp 1639504043
transform 1 0 25116 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1085_
timestamp 1639504043
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1639504043
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_15
timestamp 1639504043
transform 1 0 2484 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1639504043
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1639504043
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1639504043
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1358_
timestamp 1639504043
transform 1 0 1656 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_clk
timestamp 1639504043
transform -1 0 4324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _0846_
timestamp 1639504043
transform 1 0 3220 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0845_
timestamp 1639504043
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0837_
timestamp 1639504043
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1639504043
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_21
timestamp 1639504043
transform 1 0 3036 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _0841_
timestamp 1639504043
transform 1 0 4048 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0835_
timestamp 1639504043
transform -1 0 4692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0829_
timestamp 1639504043
transform -1 0 4968 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_40
timestamp 1639504043
transform 1 0 4784 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_35
timestamp 1639504043
transform 1 0 4324 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1362_
timestamp 1639504043
transform -1 0 6440 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1639504043
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0827_
timestamp 1639504043
transform -1 0 5520 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1639504043
transform -1 0 5244 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0830_
timestamp 1639504043
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _0836_
timestamp 1639504043
transform 1 0 6440 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1363_
timestamp 1639504043
transform 1 0 6348 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A
timestamp 1639504043
transform 1 0 7912 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__C
timestamp 1639504043
transform 1 0 8740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_76
timestamp 1639504043
transform 1 0 8096 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_82
timestamp 1639504043
transform 1 0 8648 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_72
timestamp 1639504043
transform 1 0 7728 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1639504043
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _0826_
timestamp 1639504043
transform -1 0 8740 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0832_
timestamp 1639504043
transform -1 0 8096 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0834_
timestamp 1639504043
transform -1 0 7728 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0655_
timestamp 1639504043
transform -1 0 9476 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0654_
timestamp 1639504043
transform -1 0 9752 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1639504043
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1639504043
transform 1 0 9660 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_85
timestamp 1639504043
transform 1 0 8924 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_2  _0984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1639504043
transform 1 0 10580 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _0935_
timestamp 1639504043
transform 1 0 9936 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1639504043
transform 1 0 9844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_94
timestamp 1639504043
transform 1 0 9752 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_102
timestamp 1639504043
transform 1 0 10488 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_98
timestamp 1639504043
transform 1 0 10120 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_112
timestamp 1639504043
transform 1 0 11408 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_124
timestamp 1639504043
transform 1 0 12512 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1639504043
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0983_
timestamp 1639504043
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0985_
timestamp 1639504043
transform 1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1307_
timestamp 1639504043
transform 1 0 11500 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_33_130
timestamp 1639504043
transform 1 0 13064 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1639504043
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_141
timestamp 1639504043
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1639504043
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1326_
timestamp 1639504043
transform 1 0 14168 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1639504043
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_150
timestamp 1639504043
transform 1 0 14904 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_157
timestamp 1639504043
transform 1 0 15548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _0653_
timestamp 1639504043
transform -1 0 15548 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0939_
timestamp 1639504043
transform -1 0 14904 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1129_
timestamp 1639504043
transform 1 0 15732 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_34_169
timestamp 1639504043
transform 1 0 16652 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1639504043
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1123_
timestamp 1639504043
transform 1 0 16836 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1212_
timestamp 1639504043
transform 1 0 18216 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1324_
timestamp 1639504043
transform -1 0 19136 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1325_
timestamp 1639504043
transform 1 0 16652 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__S
timestamp 1639504043
transform 1 0 19596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_201
timestamp 1639504043
transform 1 0 19596 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_197
timestamp 1639504043
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1639504043
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0652_
timestamp 1639504043
transform 1 0 19044 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0947_
timestamp 1639504043
transform 1 0 19320 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1254_
timestamp 1639504043
transform 1 0 19688 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1323_
timestamp 1639504043
transform 1 0 19780 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_33_211
timestamp 1639504043
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1639504043
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_225
timestamp 1639504043
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_220
timestamp 1639504043
transform 1 0 21344 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_226
timestamp 1639504043
transform 1 0 21896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1639504043
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0651_
timestamp 1639504043
transform -1 0 22540 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _1111_
timestamp 1639504043
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_231
timestamp 1639504043
transform 1 0 22356 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_239
timestamp 1639504043
transform 1 0 23092 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_247
timestamp 1639504043
transform 1 0 23828 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_240
timestamp 1639504043
transform 1 0 23184 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1639504043
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__or4_2  _0644_
timestamp 1639504043
transform -1 0 23092 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0645_
timestamp 1639504043
transform -1 0 23184 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1077_
timestamp 1639504043
transform 1 0 23552 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1090_
timestamp 1639504043
transform -1 0 24564 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_33_258
timestamp 1639504043
transform 1 0 24840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_266
timestamp 1639504043
transform 1 0 25576 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_256
timestamp 1639504043
transform 1 0 24656 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_268
timestamp 1639504043
transform 1 0 25760 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1639504043
transform -1 0 26128 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1639504043
transform -1 0 26128 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1639504043
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0954_
timestamp 1639504043
transform -1 0 24840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1639504043
transform -1 0 24656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_15
timestamp 1639504043
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1639504043
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1639504043
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_21
timestamp 1639504043
transform 1 0 3036 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_30
timestamp 1639504043
transform 1 0 3864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0844_
timestamp 1639504043
transform 1 0 3128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1361_
timestamp 1639504043
transform -1 0 5704 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1639504043
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0838_
timestamp 1639504043
transform -1 0 6256 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0840_
timestamp 1639504043
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_A
timestamp 1639504043
transform 1 0 7268 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_72
timestamp 1639504043
transform 1 0 7728 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_76
timestamp 1639504043
transform 1 0 8096 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_80
timestamp 1639504043
transform 1 0 8464 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0833_
timestamp 1639504043
transform -1 0 7728 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0927_
timestamp 1639504043
transform 1 0 8188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clk
timestamp 1639504043
transform 1 0 6900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_104
timestamp 1639504043
transform 1 0 10672 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _0825_
timestamp 1639504043
transform 1 0 8832 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0920_
timestamp 1639504043
transform 1 0 10120 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0922_
timestamp 1639504043
transform 1 0 9476 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0924_
timestamp 1639504043
transform 1 0 10396 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A1
timestamp 1639504043
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__B1
timestamp 1639504043
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_122
timestamp 1639504043
transform 1 0 12328 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1639504043
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1036_
timestamp 1639504043
transform -1 0 12880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_2  _1157_
timestamp 1639504043
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1639504043
transform 1 0 13340 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B
timestamp 1639504043
transform 1 0 13984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1639504043
transform 1 0 12880 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_142
timestamp 1639504043
transform 1 0 14168 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0937_
timestamp 1639504043
transform 1 0 13064 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1030_
timestamp 1639504043
transform 1 0 13524 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__S
timestamp 1639504043
transform 1 0 15916 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_149
timestamp 1639504043
transform 1 0 14812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_163
timestamp 1639504043
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1038_
timestamp 1639504043
transform 1 0 14536 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1043_
timestamp 1639504043
transform 1 0 15088 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1044_
timestamp 1639504043
transform 1 0 15640 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1639504043
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1639504043
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_181
timestamp 1639504043
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1639504043
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1116_
timestamp 1639504043
transform -1 0 18584 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_35_190
timestamp 1639504043
transform 1 0 18584 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_202
timestamp 1639504043
transform 1 0 19688 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_214
timestamp 1639504043
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1639504043
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1639504043
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1060_
timestamp 1639504043
transform 1 0 21804 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_35_230
timestamp 1639504043
transform 1 0 22264 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_236
timestamp 1639504043
transform 1 0 22816 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1068_
timestamp 1639504043
transform -1 0 23368 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1318_
timestamp 1639504043
transform 1 0 23368 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_35_259
timestamp 1639504043
transform 1 0 24932 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_267
timestamp 1639504043
transform 1 0 25668 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1639504043
transform -1 0 26128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1639504043
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1639504043
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1359_
timestamp 1639504043
transform 1 0 1932 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1639504043
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1639504043
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1360_
timestamp 1639504043
transform 1 0 3772 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_36_54
timestamp 1639504043
transform 1 0 6072 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_2  _0839_
timestamp 1639504043
transform 1 0 5336 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__S
timestamp 1639504043
transform 1 0 7728 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_66
timestamp 1639504043
transform 1 0 7176 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_77
timestamp 1639504043
transform 1 0 8188 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1639504043
transform -1 0 8832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1639504043
transform -1 0 8188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__A
timestamp 1639504043
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_102
timestamp 1639504043
transform 1 0 10488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1639504043
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1639504043
transform 1 0 9108 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0831_
timestamp 1639504043
transform 1 0 9936 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0923_
timestamp 1639504043
transform -1 0 9936 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1018_
timestamp 1639504043
transform -1 0 10488 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1427_
timestamp 1639504043
transform 1 0 11224 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__A2
timestamp 1639504043
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__S
timestamp 1639504043
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_136
timestamp 1639504043
transform 1 0 13616 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1639504043
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_2  _1156_
timestamp 1639504043
transform 1 0 12788 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1193_
timestamp 1639504043
transform 1 0 14076 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1037_
timestamp 1639504043
transform -1 0 15456 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1050_
timestamp 1639504043
transform 1 0 16284 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1291_
timestamp 1639504043
transform -1 0 16284 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_A
timestamp 1639504043
transform -1 0 17664 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1639504043
transform 1 0 17664 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1051_
timestamp 1639504043
transform -1 0 17480 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clk
timestamp 1639504043
transform -1 0 17204 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__S
timestamp 1639504043
transform 1 0 20240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1639504043
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1639504043
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_205
timestamp 1639504043
transform 1 0 19964 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1639504043
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_210
timestamp 1639504043
transform 1 0 20424 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_222
timestamp 1639504043
transform 1 0 21528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__and3b_2  _0960_
timestamp 1639504043
transform 1 0 21712 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__S
timestamp 1639504043
transform 1 0 23184 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__and3b_2  _0958_
timestamp 1639504043
transform 1 0 22448 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1248_
timestamp 1639504043
transform 1 0 23368 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1639504043
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_263
timestamp 1639504043
transform 1 0 25300 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1639504043
transform -1 0 26128 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1639504043
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0959_
timestamp 1639504043
transform -1 0 25300 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1069_
timestamp 1639504043
transform -1 0 25024 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1639504043
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1639504043
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1639504043
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_27
timestamp 1639504043
transform 1 0 3588 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_35
timestamp 1639504043
transform 1 0 4324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _0843_
timestamp 1639504043
transform -1 0 4324 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_47
timestamp 1639504043
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1639504043
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_57
timestamp 1639504043
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1639504043
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_76
timestamp 1639504043
transform 1 0 8096 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1639504043
transform -1 0 8464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1016_
timestamp 1639504043
transform 1 0 8464 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1215_
timestamp 1639504043
transform -1 0 7728 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_clk
timestamp 1639504043
transform 1 0 7728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _0925_
timestamp 1639504043
transform 1 0 8924 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1017_
timestamp 1639504043
transform 1 0 10488 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1214_
timestamp 1639504043
transform 1 0 9660 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1639504043
transform 1 0 10948 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__S
timestamp 1639504043
transform 1 0 11132 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1639504043
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1639504043
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_120
timestamp 1639504043
transform 1 0 12144 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1639504043
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0936_
timestamp 1639504043
transform 1 0 11868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__S
timestamp 1639504043
transform 1 0 13524 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_132
timestamp 1639504043
transform 1 0 13248 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1194_
timestamp 1639504043
transform -1 0 14536 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__S
timestamp 1639504043
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_164
timestamp 1639504043
transform 1 0 16192 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1201_
timestamp 1639504043
transform -1 0 15364 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1202_
timestamp 1639504043
transform 1 0 15364 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1639504043
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1217_
timestamp 1639504043
transform -1 0 17480 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1218_
timestamp 1639504043
transform 1 0 17480 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_clk
timestamp 1639504043
transform 1 0 18308 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1639504043
transform 1 0 18676 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0963_
timestamp 1639504043
transform 1 0 19688 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1055_
timestamp 1639504043
transform -1 0 19688 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__S
timestamp 1639504043
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1639504043
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1639504043
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1639504043
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0961_
timestamp 1639504043
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1261_
timestamp 1639504043
transform 1 0 20424 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _1061_
timestamp 1639504043
transform -1 0 23828 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _1078_
timestamp 1639504043
transform -1 0 24472 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1267_
timestamp 1639504043
transform 1 0 22264 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_37_254
timestamp 1639504043
transform 1 0 24472 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_266
timestamp 1639504043
transform 1 0 25576 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1639504043
transform -1 0 26128 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_14
timestamp 1639504043
transform 1 0 2392 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1639504043
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1639504043
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1159_
timestamp 1639504043
transform -1 0 2392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1639504043
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1639504043
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1639504043
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1639504043
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1639504043
transform -1 0 6808 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1639504043
transform 1 0 6440 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_53
timestamp 1639504043
transform 1 0 5980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_57
timestamp 1639504043
transform 1 0 6348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1008_
timestamp 1639504043
transform 1 0 6808 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_77
timestamp 1639504043
transform 1 0 8188 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1639504043
transform 1 0 7912 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0823_
timestamp 1639504043
transform 1 0 8280 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _0933_
timestamp 1639504043
transform 1 0 7084 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_38_100
timestamp 1639504043
transform 1 0 10304 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1639504043
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1639504043
transform -1 0 9844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1015_
timestamp 1639504043
transform 1 0 8924 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1020_
timestamp 1639504043
transform 1 0 9844 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__S
timestamp 1639504043
transform 1 0 12328 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_112
timestamp 1639504043
transform 1 0 11408 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_120
timestamp 1639504043
transform 1 0 12144 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_124
timestamp 1639504043
transform 1 0 12512 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__S
timestamp 1639504043
transform 1 0 14444 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1639504043
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1639504043
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_141
timestamp 1639504043
transform 1 0 14076 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1639504043
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0962_
timestamp 1639504043
transform 1 0 13248 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0967_
timestamp 1639504043
transform -1 0 14444 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__S
timestamp 1639504043
transform 1 0 15180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__S
timestamp 1639504043
transform 1 0 15640 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_151
timestamp 1639504043
transform 1 0 14996 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_155
timestamp 1639504043
transform 1 0 15364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1292_
timestamp 1639504043
transform -1 0 16652 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_clk
timestamp 1639504043
transform -1 0 14996 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__S
timestamp 1639504043
transform 1 0 17296 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_169
timestamp 1639504043
transform 1 0 16652 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_175
timestamp 1639504043
transform 1 0 17204 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_178
timestamp 1639504043
transform 1 0 17480 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_184
timestamp 1639504043
transform 1 0 18032 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0966_
timestamp 1639504043
transform 1 0 18124 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__S
timestamp 1639504043
transform 1 0 20056 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1639504043
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0964_
timestamp 1639504043
transform 1 0 20240 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0965_
timestamp 1639504043
transform -1 0 19136 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1188_
timestamp 1639504043
transform 1 0 19228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1316_
timestamp 1639504043
transform 1 0 20516 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1317_
timestamp 1639504043
transform 1 0 22080 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1639504043
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1639504043
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1639504043
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_265
timestamp 1639504043
transform 1 0 25484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1639504043
transform -1 0 26128 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1639504043
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1639504043
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1639504043
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_14
timestamp 1639504043
transform 1 0 2392 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_3
timestamp 1639504043
transform 1 0 1380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1639504043
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1639504043
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1160_
timestamp 1639504043
transform -1 0 2392 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1639504043
transform 1 0 4784 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1639504043
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_39
timestamp 1639504043
transform 1 0 4692 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1639504043
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_29
timestamp 1639504043
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_37
timestamp 1639504043
transform 1 0 4508 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1639504043
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1327_
timestamp 1639504043
transform 1 0 4784 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A3
timestamp 1639504043
transform -1 0 6256 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A
timestamp 1639504043
transform 1 0 4968 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_57
timestamp 1639504043
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1639504043
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _0930_
timestamp 1639504043
transform 1 0 5612 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0934_
timestamp 1639504043
transform -1 0 5612 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1007_
timestamp 1639504043
transform 1 0 6440 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1329_
timestamp 1639504043
transform 1 0 6348 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A2
timestamp 1639504043
transform 1 0 6900 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1639504043
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _0643_
timestamp 1639504043
transform 1 0 8740 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_2  _0929_
timestamp 1639504043
transform 1 0 7084 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _1012_
timestamp 1639504043
transform 1 0 7912 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1216_
timestamp 1639504043
transform 1 0 7912 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__S
timestamp 1639504043
transform 1 0 10488 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_104
timestamp 1639504043
transform 1 0 10672 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1639504043
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _0818_
timestamp 1639504043
transform 1 0 9384 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1639504043
transform 1 0 10488 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0926_
timestamp 1639504043
transform -1 0 10488 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1330_
timestamp 1639504043
transform -1 0 10488 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _1022_
timestamp 1639504043
transform 1 0 10764 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1021_
timestamp 1639504043
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0979_
timestamp 1639504043
transform -1 0 12052 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0816_
timestamp 1639504043
transform 1 0 11040 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1639504043
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1639504043
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_107
timestamp 1639504043
transform 1 0 10948 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1639504043
transform 1 0 10764 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1025_
timestamp 1639504043
transform -1 0 12236 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0977_
timestamp 1639504043
transform 1 0 12144 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0972_
timestamp 1639504043
transform -1 0 12512 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_119
timestamp 1639504043
transform 1 0 12052 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_116
timestamp 1639504043
transform 1 0 11776 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1190_
timestamp 1639504043
transform -1 0 13340 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_40_130
timestamp 1639504043
transform 1 0 13064 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__S
timestamp 1639504043
transform 1 0 12880 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__and3b_2  _0973_
timestamp 1639504043
transform 1 0 14168 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1639504043
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_141
timestamp 1639504043
transform 1 0 14076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1639504043
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_136
timestamp 1639504043
transform 1 0 13616 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__S
timestamp 1639504043
transform 1 0 13708 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_145
timestamp 1639504043
transform 1 0 14444 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_133
timestamp 1639504043
transform 1 0 13340 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__S
timestamp 1639504043
transform 1 0 15640 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_157
timestamp 1639504043
transform 1 0 15548 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_150
timestamp 1639504043
transform 1 0 14904 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__and3b_2  _0968_
timestamp 1639504043
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _0970_
timestamp 1639504043
transform 1 0 15088 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1293_
timestamp 1639504043
transform 1 0 15824 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__S
timestamp 1639504043
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_183
timestamp 1639504043
transform 1 0 17940 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_169
timestamp 1639504043
transform 1 0 16652 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_177
timestamp 1639504043
transform 1 0 17388 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1639504043
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1639504043
transform 1 0 16836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1049_
timestamp 1639504043
transform 1 0 18124 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1219_
timestamp 1639504043
transform 1 0 17112 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1314_
timestamp 1639504043
transform 1 0 17480 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1639504043
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_203
timestamp 1639504043
transform 1 0 19780 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1639504043
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0650_
timestamp 1639504043
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1315_
timestamp 1639504043
transform 1 0 18860 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1639504043
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1639504043
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1639504043
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1639504043
transform 1 0 20884 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1639504043
transform 1 0 21988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1639504043
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1048_
timestamp 1639504043
transform 1 0 20424 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1639504043
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1639504043
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1639504043
transform 1 0 23092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_261
timestamp 1639504043
transform 1 0 25116 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1639504043
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1639504043
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_265
timestamp 1639504043
transform 1 0 25484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1639504043
transform -1 0 26128 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1639504043
transform -1 0 26128 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1639504043
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1639504043
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1639504043
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1639504043
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1639504043
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1639504043
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1639504043
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1639504043
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_57
timestamp 1639504043
transform 1 0 6348 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1639504043
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _0931_
timestamp 1639504043
transform -1 0 6900 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0821_
timestamp 1639504043
transform -1 0 7360 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _0932_
timestamp 1639504043
transform 1 0 7360 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1213_
timestamp 1639504043
transform 1 0 8188 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__C1
timestamp 1639504043
transform 1 0 9292 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__S
timestamp 1639504043
transform 1 0 10212 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__S
timestamp 1639504043
transform -1 0 9660 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_93
timestamp 1639504043
transform 1 0 9660 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _0981_
timestamp 1639504043
transform -1 0 11408 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1011_
timestamp 1639504043
transform -1 0 9292 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1026_
timestamp 1639504043
transform 1 0 10396 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__S
timestamp 1639504043
transform 1 0 12328 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1639504043
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1191_
timestamp 1639504043
transform 1 0 12512 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1192_
timestamp 1639504043
transform 1 0 11500 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0976_
timestamp 1639504043
transform 1 0 13616 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1023_
timestamp 1639504043
transform -1 0 13616 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1195_
timestamp 1639504043
transform -1 0 14720 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0971_
timestamp 1639504043
transform 1 0 15548 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1042_
timestamp 1639504043
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1203_
timestamp 1639504043
transform 1 0 14720 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_41_177
timestamp 1639504043
transform 1 0 17388 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1639504043
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1035_
timestamp 1639504043
transform -1 0 17388 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_189
timestamp 1639504043
transform 1 0 18492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_201
timestamp 1639504043
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_213
timestamp 1639504043
transform 1 0 20700 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1639504043
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1639504043
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1639504043
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1639504043
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1639504043
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_261
timestamp 1639504043
transform 1 0 25116 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1639504043
transform -1 0 26128 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1639504043
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1639504043
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1639504043
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1639504043
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1639504043
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1639504043
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1639504043
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_53
timestamp 1639504043
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1014_
timestamp 1639504043
transform 1 0 6716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A1
timestamp 1639504043
transform 1 0 8556 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1639504043
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1009_
timestamp 1639504043
transform 1 0 7452 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1010_
timestamp 1639504043
transform 1 0 8096 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1013_
timestamp 1639504043
transform -1 0 7452 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A
timestamp 1639504043
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_87
timestamp 1639504043
transform 1 0 9108 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_95
timestamp 1639504043
transform 1 0 9844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1639504043
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1639504043
transform -1 0 10396 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1308_
timestamp 1639504043
transform 1 0 10396 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1189_
timestamp 1639504043
transform 1 0 11960 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_42_130
timestamp 1639504043
transform 1 0 13064 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1639504043
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1639504043
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _0975_
timestamp 1639504043
transform -1 0 14812 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0978_
timestamp 1639504043
transform 1 0 12788 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1027_
timestamp 1639504043
transform 1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__S
timestamp 1639504043
transform 1 0 14812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0974_
timestamp 1639504043
transform 1 0 14996 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1312_
timestamp 1639504043
transform 1 0 15272 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1313_
timestamp 1639504043
transform -1 0 18400 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_42_188
timestamp 1639504043
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1639504043
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1639504043
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1639504043
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1639504043
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1639504043
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1639504043
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1639504043
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_253
timestamp 1639504043
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_257
timestamp 1639504043
transform 1 0 24748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_261
timestamp 1639504043
transform 1 0 25116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1639504043
transform -1 0 26128 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1639504043
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1161_
timestamp 1639504043
transform 1 0 24840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1639504043
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1639504043
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1639504043
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1639504043
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1639504043
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1639504043
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1639504043
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1639504043
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1639504043
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 1639504043
transform -1 0 7636 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1328_
timestamp 1639504043
transform 1 0 7636 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_43_100
timestamp 1639504043
transform 1 0 10304 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_88
timestamp 1639504043
transform 1 0 9200 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1639504043
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0980_
timestamp 1639504043
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0982_
timestamp 1639504043
transform -1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1309_
timestamp 1639504043
transform 1 0 11500 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1310_
timestamp 1639504043
transform 1 0 13064 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1639504043
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1311_
timestamp 1639504043
transform 1 0 14628 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_43_175
timestamp 1639504043
transform 1 0 17204 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_187
timestamp 1639504043
transform 1 0 18308 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1639504043
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0649_
timestamp 1639504043
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_199
timestamp 1639504043
transform 1 0 19412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_211
timestamp 1639504043
transform 1 0 20516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1639504043
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_228
timestamp 1639504043
transform 1 0 22080 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1639504043
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1163_
timestamp 1639504043
transform -1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_236
timestamp 1639504043
transform 1 0 22816 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_240
timestamp 1639504043
transform 1 0 23184 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1165_
timestamp 1639504043
transform 1 0 22908 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_252
timestamp 1639504043
transform 1 0 24288 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_264
timestamp 1639504043
transform 1 0 25392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_268
timestamp 1639504043
transform 1 0 25760 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1639504043
transform -1 0 26128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1166_
timestamp 1639504043
transform 1 0 24840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1167_
timestamp 1639504043
transform 1 0 25116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1639504043
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1639504043
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1639504043
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1639504043
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1639504043
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1639504043
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1639504043
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1639504043
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1639504043
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1639504043
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1639504043
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1639504043
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1639504043
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1639504043
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_109
timestamp 1639504043
transform 1 0 11132 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_115
timestamp 1639504043
transform 1 0 11684 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0646_
timestamp 1639504043
transform 1 0 12512 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1024_
timestamp 1639504043
transform -1 0 12512 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_129
timestamp 1639504043
transform 1 0 12972 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1639504043
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1639504043
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0647_
timestamp 1639504043
transform 1 0 14076 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_44_159
timestamp 1639504043
transform 1 0 15732 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0648_
timestamp 1639504043
transform 1 0 15272 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1029_
timestamp 1639504043
transform 1 0 14536 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1034_
timestamp 1639504043
transform 1 0 16284 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_44_170
timestamp 1639504043
transform 1 0 16744 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_182
timestamp 1639504043
transform 1 0 17848 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1639504043
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1639504043
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1639504043
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1639504043
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1639504043
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1639504043
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1639504043
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1639504043
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1639504043
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 1639504043
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1639504043
transform -1 0 26128 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1639504043
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1639504043
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1639504043
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1639504043
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_27
timestamp 1639504043
transform 1 0 3588 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_29
timestamp 1639504043
transform 1 0 3772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_41
timestamp 1639504043
transform 1 0 4876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1639504043
transform 1 0 3680 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1639504043
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1639504043
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1639504043
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1639504043
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_81
timestamp 1639504043
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_85
timestamp 1639504043
transform 1 0 8924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_97
timestamp 1639504043
transform 1 0 10028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1639504043
transform 1 0 8832 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1639504043
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1639504043
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1639504043
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1639504043
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_137
timestamp 1639504043
transform 1 0 13708 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_141
timestamp 1639504043
transform 1 0 14076 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1639504043
transform 1 0 13984 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_153
timestamp 1639504043
transform 1 0 15180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1639504043
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1639504043
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1639504043
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1639504043
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_193
timestamp 1639504043
transform 1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_197
timestamp 1639504043
transform 1 0 19228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1639504043
transform 1 0 19136 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_209
timestamp 1639504043
transform 1 0 20332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1639504043
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1639504043
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1639504043
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1639504043
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_249
timestamp 1639504043
transform 1 0 24012 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1639504043
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_265
timestamp 1639504043
transform 1 0 25484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1639504043
transform -1 0 26128 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1639504043
transform 1 0 24288 0 -1 27200
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 688 800 808 6 clk
port 0 nsew signal input
rlabel metal2 s 570 28642 626 29442 6 data_req_i
port 1 nsew signal input
rlabel metal2 s 570 0 626 800 6 reset
port 2 nsew signal input
rlabel metal3 s 26498 688 27298 808 6 rxd_uart
port 3 nsew signal input
rlabel metal2 s 1674 28642 1730 29442 6 slave_data_addr_i[0]
port 4 nsew signal input
rlabel metal2 s 4066 28642 4122 29442 6 slave_data_addr_i[1]
port 5 nsew signal input
rlabel metal3 s 26498 8304 27298 8424 6 slave_data_addr_i[2]
port 6 nsew signal input
rlabel metal2 s 8850 28642 8906 29442 6 slave_data_addr_i[3]
port 7 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 slave_data_addr_i[4]
port 8 nsew signal input
rlabel metal3 s 26498 11432 27298 11552 6 slave_data_addr_i[5]
port 9 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 slave_data_addr_i[6]
port 10 nsew signal input
rlabel metal3 s 26498 12928 27298 13048 6 slave_data_addr_i[7]
port 11 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 slave_data_addr_i[8]
port 12 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 slave_data_addr_i[9]
port 13 nsew signal input
rlabel metal3 s 26498 5312 27298 5432 6 slave_data_be_i[0]
port 14 nsew signal input
rlabel metal3 s 26498 6808 27298 6928 6 slave_data_be_i[1]
port 15 nsew signal input
rlabel metal2 s 5262 28642 5318 29442 6 slave_data_be_i[2]
port 16 nsew signal input
rlabel metal2 s 10046 28642 10102 29442 6 slave_data_be_i[3]
port 17 nsew signal input
rlabel metal3 s 26498 2184 27298 2304 6 slave_data_gnt_o
port 18 nsew signal tristate
rlabel metal2 s 2870 28642 2926 29442 6 slave_data_rdata_o[0]
port 19 nsew signal tristate
rlabel metal2 s 12438 0 12494 800 6 slave_data_rdata_o[10]
port 20 nsew signal tristate
rlabel metal2 s 13634 0 13690 800 6 slave_data_rdata_o[11]
port 21 nsew signal tristate
rlabel metal3 s 26498 16056 27298 16176 6 slave_data_rdata_o[12]
port 22 nsew signal tristate
rlabel metal2 s 15934 0 15990 800 6 slave_data_rdata_o[13]
port 23 nsew signal tristate
rlabel metal3 s 26498 17688 27298 17808 6 slave_data_rdata_o[14]
port 24 nsew signal tristate
rlabel metal2 s 17130 0 17186 800 6 slave_data_rdata_o[15]
port 25 nsew signal tristate
rlabel metal2 s 18326 0 18382 800 6 slave_data_rdata_o[16]
port 26 nsew signal tristate
rlabel metal2 s 17130 28642 17186 29442 6 slave_data_rdata_o[17]
port 27 nsew signal tristate
rlabel metal2 s 19522 0 19578 800 6 slave_data_rdata_o[18]
port 28 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 slave_data_rdata_o[19]
port 29 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 slave_data_rdata_o[1]
port 30 nsew signal tristate
rlabel metal2 s 18326 28642 18382 29442 6 slave_data_rdata_o[20]
port 31 nsew signal tristate
rlabel metal2 s 21914 0 21970 800 6 slave_data_rdata_o[21]
port 32 nsew signal tristate
rlabel metal2 s 23110 0 23166 800 6 slave_data_rdata_o[22]
port 33 nsew signal tristate
rlabel metal3 s 0 22992 800 23112 6 slave_data_rdata_o[23]
port 34 nsew signal tristate
rlabel metal3 s 0 24352 800 24472 6 slave_data_rdata_o[24]
port 35 nsew signal tristate
rlabel metal3 s 26498 25304 27298 25424 6 slave_data_rdata_o[25]
port 36 nsew signal tristate
rlabel metal2 s 24306 0 24362 800 6 slave_data_rdata_o[26]
port 37 nsew signal tristate
rlabel metal2 s 21914 28642 21970 29442 6 slave_data_rdata_o[27]
port 38 nsew signal tristate
rlabel metal2 s 25502 0 25558 800 6 slave_data_rdata_o[28]
port 39 nsew signal tristate
rlabel metal2 s 23110 28642 23166 29442 6 slave_data_rdata_o[29]
port 40 nsew signal tristate
rlabel metal2 s 6458 28642 6514 29442 6 slave_data_rdata_o[2]
port 41 nsew signal tristate
rlabel metal2 s 25502 28642 25558 29442 6 slave_data_rdata_o[30]
port 42 nsew signal tristate
rlabel metal3 s 26498 28432 27298 28552 6 slave_data_rdata_o[31]
port 43 nsew signal tristate
rlabel metal2 s 2870 0 2926 800 6 slave_data_rdata_o[3]
port 44 nsew signal tristate
rlabel metal2 s 11242 28642 11298 29442 6 slave_data_rdata_o[4]
port 45 nsew signal tristate
rlabel metal2 s 12438 28642 12494 29442 6 slave_data_rdata_o[5]
port 46 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 slave_data_rdata_o[6]
port 47 nsew signal tristate
rlabel metal2 s 7654 0 7710 800 6 slave_data_rdata_o[7]
port 48 nsew signal tristate
rlabel metal2 s 8850 0 8906 800 6 slave_data_rdata_o[8]
port 49 nsew signal tristate
rlabel metal3 s 0 13200 800 13320 6 slave_data_rdata_o[9]
port 50 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 slave_data_rvalid_o
port 51 nsew signal tristate
rlabel metal2 s 1674 0 1730 800 6 slave_data_wdata_i[0]
port 52 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 slave_data_wdata_i[10]
port 53 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 slave_data_wdata_i[11]
port 54 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 slave_data_wdata_i[12]
port 55 nsew signal input
rlabel metal2 s 14738 28642 14794 29442 6 slave_data_wdata_i[13]
port 56 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 slave_data_wdata_i[14]
port 57 nsew signal input
rlabel metal2 s 15934 28642 15990 29442 6 slave_data_wdata_i[15]
port 58 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 slave_data_wdata_i[16]
port 59 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 slave_data_wdata_i[17]
port 60 nsew signal input
rlabel metal3 s 26498 19184 27298 19304 6 slave_data_wdata_i[18]
port 61 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 slave_data_wdata_i[19]
port 62 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 slave_data_wdata_i[1]
port 63 nsew signal input
rlabel metal2 s 19522 28642 19578 29442 6 slave_data_wdata_i[20]
port 64 nsew signal input
rlabel metal2 s 20718 28642 20774 29442 6 slave_data_wdata_i[21]
port 65 nsew signal input
rlabel metal3 s 26498 20680 27298 20800 6 slave_data_wdata_i[22]
port 66 nsew signal input
rlabel metal3 s 26498 22312 27298 22432 6 slave_data_wdata_i[23]
port 67 nsew signal input
rlabel metal3 s 26498 23808 27298 23928 6 slave_data_wdata_i[24]
port 68 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 slave_data_wdata_i[25]
port 69 nsew signal input
rlabel metal3 s 26498 26936 27298 27056 6 slave_data_wdata_i[26]
port 70 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 slave_data_wdata_i[27]
port 71 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 slave_data_wdata_i[28]
port 72 nsew signal input
rlabel metal2 s 24306 28642 24362 29442 6 slave_data_wdata_i[29]
port 73 nsew signal input
rlabel metal2 s 7654 28642 7710 29442 6 slave_data_wdata_i[2]
port 74 nsew signal input
rlabel metal2 s 26698 28642 26754 29442 6 slave_data_wdata_i[30]
port 75 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 slave_data_wdata_i[31]
port 76 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 slave_data_wdata_i[3]
port 77 nsew signal input
rlabel metal3 s 26498 9936 27298 10056 6 slave_data_wdata_i[4]
port 78 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 slave_data_wdata_i[5]
port 79 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 slave_data_wdata_i[6]
port 80 nsew signal input
rlabel metal2 s 13634 28642 13690 29442 6 slave_data_wdata_i[7]
port 81 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 slave_data_wdata_i[8]
port 82 nsew signal input
rlabel metal3 s 26498 14560 27298 14680 6 slave_data_wdata_i[9]
port 83 nsew signal input
rlabel metal3 s 26498 3680 27298 3800 6 slave_data_we_i
port 84 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 txd_uart
port 85 nsew signal tristate
rlabel metal4 s 5115 2128 5435 27248 6 vccd1
port 86 nsew power input
rlabel metal4 s 13456 2128 13776 27248 6 vccd1
port 86 nsew power input
rlabel metal4 s 21797 2128 22117 27248 6 vccd1
port 86 nsew power input
rlabel metal4 s 9285 2128 9605 27248 6 vssd1
port 87 nsew ground input
rlabel metal4 s 17626 2128 17946 27248 6 vssd1
port 87 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 27298 29442
<< end >>
