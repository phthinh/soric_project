VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ibex_top
  CLASS BLOCK ;
  FOREIGN ibex_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 1400.000 BY 1400.000 ;
  PIN alert_major_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END alert_major_o
  PIN alert_minor_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END alert_minor_o
  PIN boot_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END boot_addr_i[0]
  PIN boot_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 1396.000 429.090 1400.000 ;
    END
  END boot_addr_i[10]
  PIN boot_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END boot_addr_i[11]
  PIN boot_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END boot_addr_i[12]
  PIN boot_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END boot_addr_i[13]
  PIN boot_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 1396.000 605.730 1400.000 ;
    END
  END boot_addr_i[14]
  PIN boot_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 881.320 1400.000 881.920 ;
    END
  END boot_addr_i[15]
  PIN boot_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.200 4.000 637.800 ;
    END
  END boot_addr_i[16]
  PIN boot_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END boot_addr_i[17]
  PIN boot_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 1396.000 734.990 1400.000 ;
    END
  END boot_addr_i[18]
  PIN boot_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 943.200 1400.000 943.800 ;
    END
  END boot_addr_i[19]
  PIN boot_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 1396.000 123.190 1400.000 ;
    END
  END boot_addr_i[1]
  PIN boot_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 1396.000 770.410 1400.000 ;
    END
  END boot_addr_i[20]
  PIN boot_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 0.000 849.990 4.000 ;
    END
  END boot_addr_i[21]
  PIN boot_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 823.520 4.000 824.120 ;
    END
  END boot_addr_i[22]
  PIN boot_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 1396.000 864.250 1400.000 ;
    END
  END boot_addr_i[23]
  PIN boot_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 917.360 4.000 917.960 ;
    END
  END boot_addr_i[24]
  PIN boot_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.760 4.000 938.360 ;
    END
  END boot_addr_i[25]
  PIN boot_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1060.160 1400.000 1060.760 ;
    END
  END boot_addr_i[26]
  PIN boot_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 1396.000 1028.930 1400.000 ;
    END
  END boot_addr_i[27]
  PIN boot_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.920 4.000 1031.520 ;
    END
  END boot_addr_i[28]
  PIN boot_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1072.400 4.000 1073.000 ;
    END
  END boot_addr_i[29]
  PIN boot_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END boot_addr_i[2]
  PIN boot_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 0.000 1083.210 4.000 ;
    END
  END boot_addr_i[30]
  PIN boot_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.510 0.000 1116.790 4.000 ;
    END
  END boot_addr_i[31]
  PIN boot_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END boot_addr_i[3]
  PIN boot_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 1396.000 252.910 1400.000 ;
    END
  END boot_addr_i[4]
  PIN boot_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END boot_addr_i[5]
  PIN boot_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 696.360 1400.000 696.960 ;
    END
  END boot_addr_i[6]
  PIN boot_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END boot_addr_i[7]
  PIN boot_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END boot_addr_i[8]
  PIN boot_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END boot_addr_i[9]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END clk_i
  PIN core_sleep_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END core_sleep_o
  PIN crash_dump_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END crash_dump_o[0]
  PIN crash_dump_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1342.360 4.000 1342.960 ;
    END
  END crash_dump_o[100]
  PIN crash_dump_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1362.080 1400.000 1362.680 ;
    END
  END crash_dump_o[101]
  PIN crash_dump_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1368.880 1400.000 1369.480 ;
    END
  END crash_dump_o[102]
  PIN crash_dump_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1352.560 4.000 1353.160 ;
    END
  END crash_dump_o[103]
  PIN crash_dump_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.030 0.000 1283.310 4.000 ;
    END
  END crash_dump_o[104]
  PIN crash_dump_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.510 1396.000 1346.790 1400.000 ;
    END
  END crash_dump_o[105]
  PIN crash_dump_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.010 1396.000 1358.290 1400.000 ;
    END
  END crash_dump_o[106]
  PIN crash_dump_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1362.760 4.000 1363.360 ;
    END
  END crash_dump_o[107]
  PIN crash_dump_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.070 0.000 1294.350 4.000 ;
    END
  END crash_dump_o[108]
  PIN crash_dump_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.110 0.000 1305.390 4.000 ;
    END
  END crash_dump_o[109]
  PIN crash_dump_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 785.440 1400.000 786.040 ;
    END
  END crash_dump_o[10]
  PIN crash_dump_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 0.000 1316.430 4.000 ;
    END
  END crash_dump_o[110]
  PIN crash_dump_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.970 1396.000 1370.250 1400.000 ;
    END
  END crash_dump_o[111]
  PIN crash_dump_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.190 0.000 1327.470 4.000 ;
    END
  END crash_dump_o[112]
  PIN crash_dump_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.690 0.000 1338.970 4.000 ;
    END
  END crash_dump_o[113]
  PIN crash_dump_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 1396.000 1381.750 1400.000 ;
    END
  END crash_dump_o[114]
  PIN crash_dump_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 0.000 1350.010 4.000 ;
    END
  END crash_dump_o[115]
  PIN crash_dump_o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 4.000 1374.240 ;
    END
  END crash_dump_o[116]
  PIN crash_dump_o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1375.680 1400.000 1376.280 ;
    END
  END crash_dump_o[117]
  PIN crash_dump_o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END crash_dump_o[118]
  PIN crash_dump_o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1382.480 1400.000 1383.080 ;
    END
  END crash_dump_o[119]
  PIN crash_dump_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 812.640 1400.000 813.240 ;
    END
  END crash_dump_o[11]
  PIN crash_dump_o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 0.000 1361.050 4.000 ;
    END
  END crash_dump_o[120]
  PIN crash_dump_o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.430 1396.000 1393.710 1400.000 ;
    END
  END crash_dump_o[121]
  PIN crash_dump_o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 0.000 1372.090 4.000 ;
    END
  END crash_dump_o[122]
  PIN crash_dump_o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.850 0.000 1383.130 4.000 ;
    END
  END crash_dump_o[123]
  PIN crash_dump_o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.890 0.000 1394.170 4.000 ;
    END
  END crash_dump_o[124]
  PIN crash_dump_o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.040 4.000 1394.640 ;
    END
  END crash_dump_o[125]
  PIN crash_dump_o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1389.280 1400.000 1389.880 ;
    END
  END crash_dump_o[126]
  PIN crash_dump_o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1396.080 1400.000 1396.680 ;
    END
  END crash_dump_o[127]
  PIN crash_dump_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END crash_dump_o[12]
  PIN crash_dump_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END crash_dump_o[13]
  PIN crash_dump_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END crash_dump_o[14]
  PIN crash_dump_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 888.800 1400.000 889.400 ;
    END
  END crash_dump_o[15]
  PIN crash_dump_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 0.000 672.430 4.000 ;
    END
  END crash_dump_o[16]
  PIN crash_dump_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 4.000 ;
    END
  END crash_dump_o[17]
  PIN crash_dump_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 0.000 761.210 4.000 ;
    END
  END crash_dump_o[18]
  PIN crash_dump_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 740.560 4.000 741.160 ;
    END
  END crash_dump_o[19]
  PIN crash_dump_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 1396.000 135.150 1400.000 ;
    END
  END crash_dump_o[1]
  PIN crash_dump_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END crash_dump_o[20]
  PIN crash_dump_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 998.280 1400.000 998.880 ;
    END
  END crash_dump_o[21]
  PIN crash_dump_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 1396.000 840.790 1400.000 ;
    END
  END crash_dump_o[22]
  PIN crash_dump_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 1396.000 876.210 1400.000 ;
    END
  END crash_dump_o[23]
  PIN crash_dump_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 1396.000 935.090 1400.000 ;
    END
  END crash_dump_o[24]
  PIN crash_dump_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 1396.000 970.050 1400.000 ;
    END
  END crash_dump_o[25]
  PIN crash_dump_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END crash_dump_o[26]
  PIN crash_dump_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1010.520 4.000 1011.120 ;
    END
  END crash_dump_o[27]
  PIN crash_dump_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.230 0.000 1016.510 4.000 ;
    END
  END crash_dump_o[28]
  PIN crash_dump_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1135.640 1400.000 1136.240 ;
    END
  END crash_dump_o[29]
  PIN crash_dump_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END crash_dump_o[2]
  PIN crash_dump_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1162.840 1400.000 1163.440 ;
    END
  END crash_dump_o[30]
  PIN crash_dump_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1134.960 4.000 1135.560 ;
    END
  END crash_dump_o[31]
  PIN crash_dump_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1217.920 1400.000 1218.520 ;
    END
  END crash_dump_o[32]
  PIN crash_dump_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1224.720 1400.000 1225.320 ;
    END
  END crash_dump_o[33]
  PIN crash_dump_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1231.520 1400.000 1232.120 ;
    END
  END crash_dump_o[34]
  PIN crash_dump_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END crash_dump_o[35]
  PIN crash_dump_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 1396.000 1146.690 1400.000 ;
    END
  END crash_dump_o[36]
  PIN crash_dump_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1238.320 1400.000 1238.920 ;
    END
  END crash_dump_o[37]
  PIN crash_dump_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1186.640 4.000 1187.240 ;
    END
  END crash_dump_o[38]
  PIN crash_dump_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.550 0.000 1127.830 4.000 ;
    END
  END crash_dump_o[39]
  PIN crash_dump_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 600.480 1400.000 601.080 ;
    END
  END crash_dump_o[3]
  PIN crash_dump_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1245.120 1400.000 1245.720 ;
    END
  END crash_dump_o[40]
  PIN crash_dump_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1251.920 1400.000 1252.520 ;
    END
  END crash_dump_o[41]
  PIN crash_dump_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1259.400 1400.000 1260.000 ;
    END
  END crash_dump_o[42]
  PIN crash_dump_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1196.840 4.000 1197.440 ;
    END
  END crash_dump_o[43]
  PIN crash_dump_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1266.200 1400.000 1266.800 ;
    END
  END crash_dump_o[44]
  PIN crash_dump_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.720 4.000 1208.320 ;
    END
  END crash_dump_o[45]
  PIN crash_dump_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1273.000 1400.000 1273.600 ;
    END
  END crash_dump_o[46]
  PIN crash_dump_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.920 4.000 1218.520 ;
    END
  END crash_dump_o[47]
  PIN crash_dump_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.370 1396.000 1158.650 1400.000 ;
    END
  END crash_dump_o[48]
  PIN crash_dump_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1279.800 1400.000 1280.400 ;
    END
  END crash_dump_o[49]
  PIN crash_dump_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END crash_dump_o[4]
  PIN crash_dump_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.590 0.000 1138.870 4.000 ;
    END
  END crash_dump_o[50]
  PIN crash_dump_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 1396.000 1170.150 1400.000 ;
    END
  END crash_dump_o[51]
  PIN crash_dump_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1228.120 4.000 1228.720 ;
    END
  END crash_dump_o[52]
  PIN crash_dump_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1286.600 1400.000 1287.200 ;
    END
  END crash_dump_o[53]
  PIN crash_dump_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 1396.000 1182.110 1400.000 ;
    END
  END crash_dump_o[54]
  PIN crash_dump_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END crash_dump_o[55]
  PIN crash_dump_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1238.320 4.000 1238.920 ;
    END
  END crash_dump_o[56]
  PIN crash_dump_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1249.200 4.000 1249.800 ;
    END
  END crash_dump_o[57]
  PIN crash_dump_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.330 1396.000 1193.610 1400.000 ;
    END
  END crash_dump_o[58]
  PIN crash_dump_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.290 1396.000 1205.570 1400.000 ;
    END
  END crash_dump_o[59]
  PIN crash_dump_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 682.760 1400.000 683.360 ;
    END
  END crash_dump_o[5]
  PIN crash_dump_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.670 0.000 1160.950 4.000 ;
    END
  END crash_dump_o[60]
  PIN crash_dump_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1293.400 1400.000 1294.000 ;
    END
  END crash_dump_o[61]
  PIN crash_dump_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1300.200 1400.000 1300.800 ;
    END
  END crash_dump_o[62]
  PIN crash_dump_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1307.000 1400.000 1307.600 ;
    END
  END crash_dump_o[63]
  PIN crash_dump_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1313.800 1400.000 1314.400 ;
    END
  END crash_dump_o[64]
  PIN crash_dump_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1259.400 4.000 1260.000 ;
    END
  END crash_dump_o[65]
  PIN crash_dump_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1320.600 1400.000 1321.200 ;
    END
  END crash_dump_o[66]
  PIN crash_dump_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.790 1396.000 1217.070 1400.000 ;
    END
  END crash_dump_o[67]
  PIN crash_dump_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1269.600 4.000 1270.200 ;
    END
  END crash_dump_o[68]
  PIN crash_dump_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.800 4.000 1280.400 ;
    END
  END crash_dump_o[69]
  PIN crash_dump_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 1396.000 287.870 1400.000 ;
    END
  END crash_dump_o[6]
  PIN crash_dump_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.710 0.000 1171.990 4.000 ;
    END
  END crash_dump_o[70]
  PIN crash_dump_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.750 1396.000 1229.030 1400.000 ;
    END
  END crash_dump_o[71]
  PIN crash_dump_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.750 0.000 1183.030 4.000 ;
    END
  END crash_dump_o[72]
  PIN crash_dump_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 4.000 ;
    END
  END crash_dump_o[73]
  PIN crash_dump_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.710 1396.000 1240.990 1400.000 ;
    END
  END crash_dump_o[74]
  PIN crash_dump_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.290 0.000 1205.570 4.000 ;
    END
  END crash_dump_o[75]
  PIN crash_dump_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.210 1396.000 1252.490 1400.000 ;
    END
  END crash_dump_o[76]
  PIN crash_dump_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 1396.000 1264.450 1400.000 ;
    END
  END crash_dump_o[77]
  PIN crash_dump_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.670 1396.000 1275.950 1400.000 ;
    END
  END crash_dump_o[78]
  PIN crash_dump_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.630 1396.000 1287.910 1400.000 ;
    END
  END crash_dump_o[79]
  PIN crash_dump_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END crash_dump_o[7]
  PIN crash_dump_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.330 0.000 1216.610 4.000 ;
    END
  END crash_dump_o[80]
  PIN crash_dump_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 0.000 1227.650 4.000 ;
    END
  END crash_dump_o[81]
  PIN crash_dump_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.130 1396.000 1299.410 1400.000 ;
    END
  END crash_dump_o[82]
  PIN crash_dump_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.410 0.000 1238.690 4.000 ;
    END
  END crash_dump_o[83]
  PIN crash_dump_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1327.400 1400.000 1328.000 ;
    END
  END crash_dump_o[84]
  PIN crash_dump_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1290.680 4.000 1291.280 ;
    END
  END crash_dump_o[85]
  PIN crash_dump_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 0.000 1249.730 4.000 ;
    END
  END crash_dump_o[86]
  PIN crash_dump_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1334.880 1400.000 1335.480 ;
    END
  END crash_dump_o[87]
  PIN crash_dump_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1341.680 1400.000 1342.280 ;
    END
  END crash_dump_o[88]
  PIN crash_dump_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.090 1396.000 1311.370 1400.000 ;
    END
  END crash_dump_o[89]
  PIN crash_dump_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 744.640 1400.000 745.240 ;
    END
  END crash_dump_o[8]
  PIN crash_dump_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.050 1396.000 1323.330 1400.000 ;
    END
  END crash_dump_o[90]
  PIN crash_dump_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.950 0.000 1261.230 4.000 ;
    END
  END crash_dump_o[91]
  PIN crash_dump_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.550 1396.000 1334.830 1400.000 ;
    END
  END crash_dump_o[92]
  PIN crash_dump_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.880 4.000 1301.480 ;
    END
  END crash_dump_o[93]
  PIN crash_dump_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1348.480 1400.000 1349.080 ;
    END
  END crash_dump_o[94]
  PIN crash_dump_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1311.080 4.000 1311.680 ;
    END
  END crash_dump_o[95]
  PIN crash_dump_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 0.000 1272.270 4.000 ;
    END
  END crash_dump_o[96]
  PIN crash_dump_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1321.280 4.000 1321.880 ;
    END
  END crash_dump_o[97]
  PIN crash_dump_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1355.280 1400.000 1355.880 ;
    END
  END crash_dump_o[98]
  PIN crash_dump_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.160 4.000 1332.760 ;
    END
  END crash_dump_o[99]
  PIN crash_dump_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 1396.000 393.670 1400.000 ;
    END
  END crash_dump_o[9]
  PIN data_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END data_addr_o[0]
  PIN data_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 1396.000 441.050 1400.000 ;
    END
  END data_addr_o[10]
  PIN data_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 1396.000 476.010 1400.000 ;
    END
  END data_addr_o[11]
  PIN data_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 1396.000 546.850 1400.000 ;
    END
  END data_addr_o[12]
  PIN data_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 854.120 1400.000 854.720 ;
    END
  END data_addr_o[13]
  PIN data_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 1396.000 617.230 1400.000 ;
    END
  END data_addr_o[14]
  PIN data_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 895.600 1400.000 896.200 ;
    END
  END data_addr_o[15]
  PIN data_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 1396.000 676.110 1400.000 ;
    END
  END data_addr_o[16]
  PIN data_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END data_addr_o[17]
  PIN data_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 1396.000 746.950 1400.000 ;
    END
  END data_addr_o[18]
  PIN data_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 950.000 1400.000 950.600 ;
    END
  END data_addr_o[19]
  PIN data_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END data_addr_o[1]
  PIN data_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 1396.000 781.910 1400.000 ;
    END
  END data_addr_o[20]
  PIN data_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1005.080 1400.000 1005.680 ;
    END
  END data_addr_o[21]
  PIN data_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1025.480 1400.000 1026.080 ;
    END
  END data_addr_o[22]
  PIN data_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 1396.000 887.710 1400.000 ;
    END
  END data_addr_o[23]
  PIN data_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1046.560 1400.000 1047.160 ;
    END
  END data_addr_o[24]
  PIN data_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.730 1396.000 982.010 1400.000 ;
    END
  END data_addr_o[25]
  PIN data_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 0.000 983.390 4.000 ;
    END
  END data_addr_o[26]
  PIN data_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.610 1396.000 1040.890 1400.000 ;
    END
  END data_addr_o[27]
  PIN data_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 0.000 1027.550 4.000 ;
    END
  END data_addr_o[28]
  PIN data_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1142.440 1400.000 1143.040 ;
    END
  END data_addr_o[29]
  PIN data_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 572.600 1400.000 573.200 ;
    END
  END data_addr_o[2]
  PIN data_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1103.680 4.000 1104.280 ;
    END
  END data_addr_o[30]
  PIN data_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.950 1396.000 1123.230 1400.000 ;
    END
  END data_addr_o[31]
  PIN data_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END data_addr_o[3]
  PIN data_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 654.880 1400.000 655.480 ;
    END
  END data_addr_o[4]
  PIN data_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END data_addr_o[5]
  PIN data_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 703.160 1400.000 703.760 ;
    END
  END data_addr_o[6]
  PIN data_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END data_addr_o[7]
  PIN data_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.320 4.000 388.920 ;
    END
  END data_addr_o[8]
  PIN data_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END data_addr_o[9]
  PIN data_be_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END data_be_o[0]
  PIN data_be_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 565.800 1400.000 566.400 ;
    END
  END data_be_o[1]
  PIN data_be_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 1396.000 205.530 1400.000 ;
    END
  END data_be_o[2]
  PIN data_be_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 1396.000 228.990 1400.000 ;
    END
  END data_be_o[3]
  PIN data_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 1396.000 5.890 1400.000 ;
    END
  END data_err_i
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 1396.000 17.390 1400.000 ;
    END
  END data_gnt_i
  PIN data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END data_rdata_i[0]
  PIN data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END data_rdata_i[10]
  PIN data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 1396.000 487.970 1400.000 ;
    END
  END data_rdata_i[11]
  PIN data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 820.120 1400.000 820.720 ;
    END
  END data_rdata_i[12]
  PIN data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 860.920 1400.000 861.520 ;
    END
  END data_rdata_i[13]
  PIN data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 867.720 1400.000 868.320 ;
    END
  END data_rdata_i[14]
  PIN data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 902.400 1400.000 903.000 ;
    END
  END data_rdata_i[15]
  PIN data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END data_rdata_i[16]
  PIN data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END data_rdata_i[17]
  PIN data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 1396.000 758.450 1400.000 ;
    END
  END data_rdata_i[18]
  PIN data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 956.800 1400.000 957.400 ;
    END
  END data_rdata_i[19]
  PIN data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END data_rdata_i[1]
  PIN data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END data_rdata_i[20]
  PIN data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 1396.000 817.330 1400.000 ;
    END
  END data_rdata_i[21]
  PIN data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 834.400 4.000 835.000 ;
    END
  END data_rdata_i[22]
  PIN data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END data_rdata_i[23]
  PIN data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 0.000 905.650 4.000 ;
    END
  END data_rdata_i[24]
  PIN data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.530 0.000 949.810 4.000 ;
    END
  END data_rdata_i[25]
  PIN data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1066.960 1400.000 1067.560 ;
    END
  END data_rdata_i[26]
  PIN data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.720 4.000 1021.320 ;
    END
  END data_rdata_i[27]
  PIN data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.030 1396.000 1076.310 1400.000 ;
    END
  END data_rdata_i[28]
  PIN data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1149.240 1400.000 1149.840 ;
    END
  END data_rdata_i[29]
  PIN data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END data_rdata_i[2]
  PIN data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1169.640 1400.000 1170.240 ;
    END
  END data_rdata_i[30]
  PIN data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 1396.000 1134.730 1400.000 ;
    END
  END data_rdata_i[31]
  PIN data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 607.280 1400.000 607.880 ;
    END
  END data_rdata_i[3]
  PIN data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 661.680 1400.000 662.280 ;
    END
  END data_rdata_i[4]
  PIN data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END data_rdata_i[5]
  PIN data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 709.960 1400.000 710.560 ;
    END
  END data_rdata_i[6]
  PIN data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 1396.000 323.290 1400.000 ;
    END
  END data_rdata_i[7]
  PIN data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 1396.000 358.710 1400.000 ;
    END
  END data_rdata_i[8]
  PIN data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END data_rdata_i[9]
  PIN data_rdata_intg_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END data_rdata_intg_i[0]
  PIN data_rdata_intg_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END data_rdata_intg_i[1]
  PIN data_rdata_intg_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 1396.000 217.490 1400.000 ;
    END
  END data_rdata_intg_i[2]
  PIN data_rdata_intg_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 614.080 1400.000 614.680 ;
    END
  END data_rdata_intg_i[3]
  PIN data_rdata_intg_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 669.160 1400.000 669.760 ;
    END
  END data_rdata_intg_i[4]
  PIN data_rdata_intg_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END data_rdata_intg_i[5]
  PIN data_rdata_intg_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1396.000 299.830 1400.000 ;
    END
  END data_rdata_intg_i[6]
  PIN data_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 517.520 1400.000 518.120 ;
    END
  END data_req_o
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 1396.000 29.350 1400.000 ;
    END
  END data_rvalid_i
  PIN data_wdata_intg_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END data_wdata_intg_o[0]
  PIN data_wdata_intg_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 1396.000 146.650 1400.000 ;
    END
  END data_wdata_intg_o[1]
  PIN data_wdata_intg_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END data_wdata_intg_o[2]
  PIN data_wdata_intg_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 620.880 1400.000 621.480 ;
    END
  END data_wdata_intg_o[3]
  PIN data_wdata_intg_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END data_wdata_intg_o[4]
  PIN data_wdata_intg_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END data_wdata_intg_o[5]
  PIN data_wdata_intg_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 1396.000 311.330 1400.000 ;
    END
  END data_wdata_intg_o[6]
  PIN data_wdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 538.600 1400.000 539.200 ;
    END
  END data_wdata_o[0]
  PIN data_wdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 1396.000 452.550 1400.000 ;
    END
  END data_wdata_o[10]
  PIN data_wdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 1396.000 499.930 1400.000 ;
    END
  END data_wdata_o[11]
  PIN data_wdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 826.920 1400.000 827.520 ;
    END
  END data_wdata_o[12]
  PIN data_wdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END data_wdata_o[13]
  PIN data_wdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 1396.000 629.190 1400.000 ;
    END
  END data_wdata_o[14]
  PIN data_wdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 1396.000 664.610 1400.000 ;
    END
  END data_wdata_o[15]
  PIN data_wdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 1396.000 688.070 1400.000 ;
    END
  END data_wdata_o[16]
  PIN data_wdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 1396.000 699.570 1400.000 ;
    END
  END data_wdata_o[17]
  PIN data_wdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END data_wdata_o[18]
  PIN data_wdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END data_wdata_o[19]
  PIN data_wdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END data_wdata_o[1]
  PIN data_wdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 984.680 1400.000 985.280 ;
    END
  END data_wdata_o[20]
  PIN data_wdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END data_wdata_o[21]
  PIN data_wdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 844.600 4.000 845.200 ;
    END
  END data_wdata_o[22]
  PIN data_wdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 1396.000 899.670 1400.000 ;
    END
  END data_wdata_o[23]
  PIN data_wdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 1396.000 946.590 1400.000 ;
    END
  END data_wdata_o[24]
  PIN data_wdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.960 4.000 948.560 ;
    END
  END data_wdata_o[25]
  PIN data_wdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END data_wdata_o[26]
  PIN data_wdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1094.160 1400.000 1094.760 ;
    END
  END data_wdata_o[27]
  PIN data_wdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.800 4.000 1042.400 ;
    END
  END data_wdata_o[28]
  PIN data_wdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END data_wdata_o[29]
  PIN data_wdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END data_wdata_o[2]
  PIN data_wdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1176.440 1400.000 1177.040 ;
    END
  END data_wdata_o[30]
  PIN data_wdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1190.720 1400.000 1191.320 ;
    END
  END data_wdata_o[31]
  PIN data_wdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END data_wdata_o[3]
  PIN data_wdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END data_wdata_o[4]
  PIN data_wdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END data_wdata_o[5]
  PIN data_wdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 716.760 1400.000 717.360 ;
    END
  END data_wdata_o[6]
  PIN data_wdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END data_wdata_o[7]
  PIN data_wdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 751.440 1400.000 752.040 ;
    END
  END data_wdata_o[8]
  PIN data_wdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 771.840 1400.000 772.440 ;
    END
  END data_wdata_o[9]
  PIN data_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 1396.000 40.850 1400.000 ;
    END
  END data_we_o
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END debug_req_i
  PIN eFPGA_delay_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 1396.000 99.730 1400.000 ;
    END
  END eFPGA_delay_o[0]
  PIN eFPGA_delay_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 1396.000 158.610 1400.000 ;
    END
  END eFPGA_delay_o[1]
  PIN eFPGA_delay_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END eFPGA_delay_o[2]
  PIN eFPGA_delay_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 627.680 1400.000 628.280 ;
    END
  END eFPGA_delay_o[3]
  PIN eFPGA_en_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 1396.000 52.810 1400.000 ;
    END
  END eFPGA_en_o
  PIN eFPGA_fpga_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END eFPGA_fpga_done_i
  PIN eFPGA_operand_a_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END eFPGA_operand_a_o[0]
  PIN eFPGA_operand_a_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 792.240 1400.000 792.840 ;
    END
  END eFPGA_operand_a_o[10]
  PIN eFPGA_operand_a_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.960 4.000 523.560 ;
    END
  END eFPGA_operand_a_o[11]
  PIN eFPGA_operand_a_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 1396.000 558.350 1400.000 ;
    END
  END eFPGA_operand_a_o[12]
  PIN eFPGA_operand_a_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END eFPGA_operand_a_o[13]
  PIN eFPGA_operand_a_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 1396.000 640.690 1400.000 ;
    END
  END eFPGA_operand_a_o[14]
  PIN eFPGA_operand_a_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END eFPGA_operand_a_o[15]
  PIN eFPGA_operand_a_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END eFPGA_operand_a_o[16]
  PIN eFPGA_operand_a_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 1396.000 711.530 1400.000 ;
    END
  END eFPGA_operand_a_o[17]
  PIN eFPGA_operand_a_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 4.000 ;
    END
  END eFPGA_operand_a_o[18]
  PIN eFPGA_operand_a_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 964.280 1400.000 964.880 ;
    END
  END eFPGA_operand_a_o[19]
  PIN eFPGA_operand_a_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END eFPGA_operand_a_o[1]
  PIN eFPGA_operand_a_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 1396.000 793.870 1400.000 ;
    END
  END eFPGA_operand_a_o[20]
  PIN eFPGA_operand_a_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1011.880 1400.000 1012.480 ;
    END
  END eFPGA_operand_a_o[21]
  PIN eFPGA_operand_a_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.800 4.000 855.400 ;
    END
  END eFPGA_operand_a_o[22]
  PIN eFPGA_operand_a_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 1396.000 911.630 1400.000 ;
    END
  END eFPGA_operand_a_o[23]
  PIN eFPGA_operand_a_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 0.000 916.690 4.000 ;
    END
  END eFPGA_operand_a_o[24]
  PIN eFPGA_operand_a_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END eFPGA_operand_a_o[25]
  PIN eFPGA_operand_a_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1073.760 1400.000 1074.360 ;
    END
  END eFPGA_operand_a_o[26]
  PIN eFPGA_operand_a_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.110 1396.000 1052.390 1400.000 ;
    END
  END eFPGA_operand_a_o[27]
  PIN eFPGA_operand_a_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1122.040 1400.000 1122.640 ;
    END
  END eFPGA_operand_a_o[28]
  PIN eFPGA_operand_a_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.490 1396.000 1099.770 1400.000 ;
    END
  END eFPGA_operand_a_o[29]
  PIN eFPGA_operand_a_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END eFPGA_operand_a_o[2]
  PIN eFPGA_operand_a_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 1396.000 1111.270 1400.000 ;
    END
  END eFPGA_operand_a_o[30]
  PIN eFPGA_operand_a_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.160 4.000 1145.760 ;
    END
  END eFPGA_operand_a_o[31]
  PIN eFPGA_operand_a_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 634.480 1400.000 635.080 ;
    END
  END eFPGA_operand_a_o[3]
  PIN eFPGA_operand_a_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END eFPGA_operand_a_o[4]
  PIN eFPGA_operand_a_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END eFPGA_operand_a_o[5]
  PIN eFPGA_operand_a_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END eFPGA_operand_a_o[6]
  PIN eFPGA_operand_a_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END eFPGA_operand_a_o[7]
  PIN eFPGA_operand_a_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END eFPGA_operand_a_o[8]
  PIN eFPGA_operand_a_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END eFPGA_operand_a_o[9]
  PIN eFPGA_operand_b_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 545.400 1400.000 546.000 ;
    END
  END eFPGA_operand_b_o[0]
  PIN eFPGA_operand_b_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 799.040 1400.000 799.640 ;
    END
  END eFPGA_operand_b_o[10]
  PIN eFPGA_operand_b_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 1396.000 511.430 1400.000 ;
    END
  END eFPGA_operand_b_o[11]
  PIN eFPGA_operand_b_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 833.720 1400.000 834.320 ;
    END
  END eFPGA_operand_b_o[12]
  PIN eFPGA_operand_b_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END eFPGA_operand_b_o[13]
  PIN eFPGA_operand_b_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 874.520 1400.000 875.120 ;
    END
  END eFPGA_operand_b_o[14]
  PIN eFPGA_operand_b_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END eFPGA_operand_b_o[15]
  PIN eFPGA_operand_b_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END eFPGA_operand_b_o[16]
  PIN eFPGA_operand_b_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 922.800 1400.000 923.400 ;
    END
  END eFPGA_operand_b_o[17]
  PIN eFPGA_operand_b_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END eFPGA_operand_b_o[18]
  PIN eFPGA_operand_b_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 971.080 1400.000 971.680 ;
    END
  END eFPGA_operand_b_o[19]
  PIN eFPGA_operand_b_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 1396.000 170.570 1400.000 ;
    END
  END eFPGA_operand_b_o[1]
  PIN eFPGA_operand_b_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 991.480 1400.000 992.080 ;
    END
  END eFPGA_operand_b_o[20]
  PIN eFPGA_operand_b_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.120 4.000 803.720 ;
    END
  END eFPGA_operand_b_o[21]
  PIN eFPGA_operand_b_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END eFPGA_operand_b_o[22]
  PIN eFPGA_operand_b_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.080 4.000 886.680 ;
    END
  END eFPGA_operand_b_o[23]
  PIN eFPGA_operand_b_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END eFPGA_operand_b_o[24]
  PIN eFPGA_operand_b_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 1396.000 993.970 1400.000 ;
    END
  END eFPGA_operand_b_o[25]
  PIN eFPGA_operand_b_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END eFPGA_operand_b_o[26]
  PIN eFPGA_operand_b_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1100.960 1400.000 1101.560 ;
    END
  END eFPGA_operand_b_o[27]
  PIN eFPGA_operand_b_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1052.000 4.000 1052.600 ;
    END
  END eFPGA_operand_b_o[28]
  PIN eFPGA_operand_b_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1156.040 1400.000 1156.640 ;
    END
  END eFPGA_operand_b_o[29]
  PIN eFPGA_operand_b_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 579.400 1400.000 580.000 ;
    END
  END eFPGA_operand_b_o[2]
  PIN eFPGA_operand_b_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 4.000 ;
    END
  END eFPGA_operand_b_o[30]
  PIN eFPGA_operand_b_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1155.360 4.000 1155.960 ;
    END
  END eFPGA_operand_b_o[31]
  PIN eFPGA_operand_b_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END eFPGA_operand_b_o[3]
  PIN eFPGA_operand_b_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END eFPGA_operand_b_o[4]
  PIN eFPGA_operand_b_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END eFPGA_operand_b_o[5]
  PIN eFPGA_operand_b_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END eFPGA_operand_b_o[6]
  PIN eFPGA_operand_b_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END eFPGA_operand_b_o[7]
  PIN eFPGA_operand_b_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END eFPGA_operand_b_o[8]
  PIN eFPGA_operand_b_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END eFPGA_operand_b_o[9]
  PIN eFPGA_operator_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END eFPGA_operator_o[0]
  PIN eFPGA_operator_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END eFPGA_operator_o[1]
  PIN eFPGA_result_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END eFPGA_result_a_i[0]
  PIN eFPGA_result_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 1396.000 464.510 1400.000 ;
    END
  END eFPGA_result_a_i[10]
  PIN eFPGA_result_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END eFPGA_result_a_i[11]
  PIN eFPGA_result_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END eFPGA_result_a_i[12]
  PIN eFPGA_result_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 4.000 606.520 ;
    END
  END eFPGA_result_a_i[13]
  PIN eFPGA_result_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END eFPGA_result_a_i[14]
  PIN eFPGA_result_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END eFPGA_result_a_i[15]
  PIN eFPGA_result_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END eFPGA_result_a_i[16]
  PIN eFPGA_result_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 929.600 1400.000 930.200 ;
    END
  END eFPGA_result_a_i[17]
  PIN eFPGA_result_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END eFPGA_result_a_i[18]
  PIN eFPGA_result_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END eFPGA_result_a_i[19]
  PIN eFPGA_result_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END eFPGA_result_a_i[1]
  PIN eFPGA_result_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END eFPGA_result_a_i[20]
  PIN eFPGA_result_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 1396.000 829.290 1400.000 ;
    END
  END eFPGA_result_a_i[21]
  PIN eFPGA_result_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 1396.000 852.750 1400.000 ;
    END
  END eFPGA_result_a_i[22]
  PIN eFPGA_result_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 0.000 894.610 4.000 ;
    END
  END eFPGA_result_a_i[23]
  PIN eFPGA_result_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 927.560 4.000 928.160 ;
    END
  END eFPGA_result_a_i[24]
  PIN eFPGA_result_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.570 0.000 960.850 4.000 ;
    END
  END eFPGA_result_a_i[25]
  PIN eFPGA_result_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1080.560 1400.000 1081.160 ;
    END
  END eFPGA_result_a_i[26]
  PIN eFPGA_result_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 4.000 ;
    END
  END eFPGA_result_a_i[27]
  PIN eFPGA_result_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 1396.000 1087.810 1400.000 ;
    END
  END eFPGA_result_a_i[28]
  PIN eFPGA_result_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.850 0.000 1061.130 4.000 ;
    END
  END eFPGA_result_a_i[29]
  PIN eFPGA_result_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 586.200 1400.000 586.800 ;
    END
  END eFPGA_result_a_i[2]
  PIN eFPGA_result_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1113.880 4.000 1114.480 ;
    END
  END eFPGA_result_a_i[30]
  PIN eFPGA_result_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1197.520 1400.000 1198.120 ;
    END
  END eFPGA_result_a_i[31]
  PIN eFPGA_result_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 1396.000 240.950 1400.000 ;
    END
  END eFPGA_result_a_i[3]
  PIN eFPGA_result_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END eFPGA_result_a_i[4]
  PIN eFPGA_result_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 689.560 1400.000 690.160 ;
    END
  END eFPGA_result_a_i[5]
  PIN eFPGA_result_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 723.560 1400.000 724.160 ;
    END
  END eFPGA_result_a_i[6]
  PIN eFPGA_result_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 1396.000 335.250 1400.000 ;
    END
  END eFPGA_result_a_i[7]
  PIN eFPGA_result_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 758.240 1400.000 758.840 ;
    END
  END eFPGA_result_a_i[8]
  PIN eFPGA_result_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END eFPGA_result_a_i[9]
  PIN eFPGA_result_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 552.200 1400.000 552.800 ;
    END
  END eFPGA_result_b_i[0]
  PIN eFPGA_result_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.680 4.000 492.280 ;
    END
  END eFPGA_result_b_i[10]
  PIN eFPGA_result_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 1396.000 523.390 1400.000 ;
    END
  END eFPGA_result_b_i[11]
  PIN eFPGA_result_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 840.520 1400.000 841.120 ;
    END
  END eFPGA_result_b_i[12]
  PIN eFPGA_result_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END eFPGA_result_b_i[13]
  PIN eFPGA_result_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END eFPGA_result_b_i[14]
  PIN eFPGA_result_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 909.200 1400.000 909.800 ;
    END
  END eFPGA_result_b_i[15]
  PIN eFPGA_result_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END eFPGA_result_b_i[16]
  PIN eFPGA_result_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END eFPGA_result_b_i[17]
  PIN eFPGA_result_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 936.400 1400.000 937.000 ;
    END
  END eFPGA_result_b_i[18]
  PIN eFPGA_result_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 977.880 1400.000 978.480 ;
    END
  END eFPGA_result_b_i[19]
  PIN eFPGA_result_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 1396.000 182.070 1400.000 ;
    END
  END eFPGA_result_b_i[1]
  PIN eFPGA_result_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END eFPGA_result_b_i[20]
  PIN eFPGA_result_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1018.680 1400.000 1019.280 ;
    END
  END eFPGA_result_b_i[21]
  PIN eFPGA_result_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 0.000 883.110 4.000 ;
    END
  END eFPGA_result_b_i[22]
  PIN eFPGA_result_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.850 1396.000 923.130 1400.000 ;
    END
  END eFPGA_result_b_i[23]
  PIN eFPGA_result_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 0.000 938.770 4.000 ;
    END
  END eFPGA_result_b_i[24]
  PIN eFPGA_result_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 1396.000 1005.470 1400.000 ;
    END
  END eFPGA_result_b_i[25]
  PIN eFPGA_result_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1087.360 1400.000 1087.960 ;
    END
  END eFPGA_result_b_i[26]
  PIN eFPGA_result_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.070 1396.000 1064.350 1400.000 ;
    END
  END eFPGA_result_b_i[27]
  PIN eFPGA_result_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.770 0.000 1039.050 4.000 ;
    END
  END eFPGA_result_b_i[28]
  PIN eFPGA_result_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1083.280 4.000 1083.880 ;
    END
  END eFPGA_result_b_i[29]
  PIN eFPGA_result_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END eFPGA_result_b_i[2]
  PIN eFPGA_result_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.010 0.000 1105.290 4.000 ;
    END
  END eFPGA_result_b_i[30]
  PIN eFPGA_result_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1204.320 1400.000 1204.920 ;
    END
  END eFPGA_result_b_i[31]
  PIN eFPGA_result_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 641.280 1400.000 641.880 ;
    END
  END eFPGA_result_b_i[3]
  PIN eFPGA_result_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END eFPGA_result_b_i[4]
  PIN eFPGA_result_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 1396.000 264.410 1400.000 ;
    END
  END eFPGA_result_b_i[5]
  PIN eFPGA_result_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END eFPGA_result_b_i[6]
  PIN eFPGA_result_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END eFPGA_result_b_i[7]
  PIN eFPGA_result_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 1396.000 370.210 1400.000 ;
    END
  END eFPGA_result_b_i[8]
  PIN eFPGA_result_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 1396.000 405.630 1400.000 ;
    END
  END eFPGA_result_b_i[9]
  PIN eFPGA_result_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 1396.000 111.690 1400.000 ;
    END
  END eFPGA_result_c_i[0]
  PIN eFPGA_result_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 805.840 1400.000 806.440 ;
    END
  END eFPGA_result_c_i[10]
  PIN eFPGA_result_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 1396.000 534.890 1400.000 ;
    END
  END eFPGA_result_c_i[11]
  PIN eFPGA_result_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 847.320 1400.000 847.920 ;
    END
  END eFPGA_result_c_i[12]
  PIN eFPGA_result_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 1396.000 570.310 1400.000 ;
    END
  END eFPGA_result_c_i[13]
  PIN eFPGA_result_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END eFPGA_result_c_i[14]
  PIN eFPGA_result_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 916.000 1400.000 916.600 ;
    END
  END eFPGA_result_c_i[15]
  PIN eFPGA_result_c_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END eFPGA_result_c_i[16]
  PIN eFPGA_result_c_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END eFPGA_result_c_i[17]
  PIN eFPGA_result_c_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END eFPGA_result_c_i[18]
  PIN eFPGA_result_c_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END eFPGA_result_c_i[19]
  PIN eFPGA_result_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END eFPGA_result_c_i[1]
  PIN eFPGA_result_c_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END eFPGA_result_c_i[20]
  PIN eFPGA_result_c_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END eFPGA_result_c_i[21]
  PIN eFPGA_result_c_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1032.280 1400.000 1032.880 ;
    END
  END eFPGA_result_c_i[22]
  PIN eFPGA_result_c_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.280 4.000 896.880 ;
    END
  END eFPGA_result_c_i[23]
  PIN eFPGA_result_c_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.270 1396.000 958.550 1400.000 ;
    END
  END eFPGA_result_c_i[24]
  PIN eFPGA_result_c_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 1396.000 1017.430 1400.000 ;
    END
  END eFPGA_result_c_i[25]
  PIN eFPGA_result_c_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1000.320 4.000 1000.920 ;
    END
  END eFPGA_result_c_i[26]
  PIN eFPGA_result_c_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1107.760 1400.000 1108.360 ;
    END
  END eFPGA_result_c_i[27]
  PIN eFPGA_result_c_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1128.840 1400.000 1129.440 ;
    END
  END eFPGA_result_c_i[28]
  PIN eFPGA_result_c_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 0.000 1072.170 4.000 ;
    END
  END eFPGA_result_c_i[29]
  PIN eFPGA_result_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END eFPGA_result_c_i[2]
  PIN eFPGA_result_c_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1183.920 1400.000 1184.520 ;
    END
  END eFPGA_result_c_i[30]
  PIN eFPGA_result_c_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1211.120 1400.000 1211.720 ;
    END
  END eFPGA_result_c_i[31]
  PIN eFPGA_result_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 648.080 1400.000 648.680 ;
    END
  END eFPGA_result_c_i[3]
  PIN eFPGA_result_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 675.960 1400.000 676.560 ;
    END
  END eFPGA_result_c_i[4]
  PIN eFPGA_result_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 1396.000 276.370 1400.000 ;
    END
  END eFPGA_result_c_i[5]
  PIN eFPGA_result_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END eFPGA_result_c_i[6]
  PIN eFPGA_result_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 730.360 1400.000 730.960 ;
    END
  END eFPGA_result_c_i[7]
  PIN eFPGA_result_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 1396.000 382.170 1400.000 ;
    END
  END eFPGA_result_c_i[8]
  PIN eFPGA_result_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 1396.000 417.590 1400.000 ;
    END
  END eFPGA_result_c_i[9]
  PIN eFPGA_write_strobe_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END eFPGA_write_strobe_o
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 525.000 1400.000 525.600 ;
    END
  END fetch_enable_i
  PIN hart_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 559.000 1400.000 559.600 ;
    END
  END hart_id_i[0]
  PIN hart_id_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 4.000 503.160 ;
    END
  END hart_id_i[10]
  PIN hart_id_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END hart_id_i[11]
  PIN hart_id_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END hart_id_i[12]
  PIN hart_id_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 1396.000 582.270 1400.000 ;
    END
  END hart_id_i[13]
  PIN hart_id_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 1396.000 652.650 1400.000 ;
    END
  END hart_id_i[14]
  PIN hart_id_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END hart_id_i[15]
  PIN hart_id_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END hart_id_i[16]
  PIN hart_id_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 1396.000 723.030 1400.000 ;
    END
  END hart_id_i[17]
  PIN hart_id_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END hart_id_i[18]
  PIN hart_id_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 0.000 816.870 4.000 ;
    END
  END hart_id_i[19]
  PIN hart_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END hart_id_i[1]
  PIN hart_id_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 1396.000 805.370 1400.000 ;
    END
  END hart_id_i[20]
  PIN hart_id_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END hart_id_i[21]
  PIN hart_id_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1039.760 1400.000 1040.360 ;
    END
  END hart_id_i[22]
  PIN hart_id_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 906.480 4.000 907.080 ;
    END
  END hart_id_i[23]
  PIN hart_id_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1053.360 1400.000 1053.960 ;
    END
  END hart_id_i[24]
  PIN hart_id_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 4.000 ;
    END
  END hart_id_i[25]
  PIN hart_id_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 0.000 994.430 4.000 ;
    END
  END hart_id_i[26]
  PIN hart_id_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1115.240 1400.000 1115.840 ;
    END
  END hart_id_i[27]
  PIN hart_id_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.200 4.000 1062.800 ;
    END
  END hart_id_i[28]
  PIN hart_id_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1093.480 4.000 1094.080 ;
    END
  END hart_id_i[29]
  PIN hart_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 593.680 1400.000 594.280 ;
    END
  END hart_id_i[2]
  PIN hart_id_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.760 4.000 1125.360 ;
    END
  END hart_id_i[30]
  PIN hart_id_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END hart_id_i[31]
  PIN hart_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END hart_id_i[3]
  PIN hart_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END hart_id_i[4]
  PIN hart_id_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END hart_id_i[5]
  PIN hart_id_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 4.000 ;
    END
  END hart_id_i[6]
  PIN hart_id_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 1396.000 346.750 1400.000 ;
    END
  END hart_id_i[7]
  PIN hart_id_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.600 4.000 420.200 ;
    END
  END hart_id_i[8]
  PIN hart_id_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END hart_id_i[9]
  PIN instr_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 30.640 1400.000 31.240 ;
    END
  END instr_addr_o[0]
  PIN instr_addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 215.600 1400.000 216.200 ;
    END
  END instr_addr_o[10]
  PIN instr_addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 229.880 1400.000 230.480 ;
    END
  END instr_addr_o[11]
  PIN instr_addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 243.480 1400.000 244.080 ;
    END
  END instr_addr_o[12]
  PIN instr_addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 257.080 1400.000 257.680 ;
    END
  END instr_addr_o[13]
  PIN instr_addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 270.680 1400.000 271.280 ;
    END
  END instr_addr_o[14]
  PIN instr_addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 284.280 1400.000 284.880 ;
    END
  END instr_addr_o[15]
  PIN instr_addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 298.560 1400.000 299.160 ;
    END
  END instr_addr_o[16]
  PIN instr_addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 312.160 1400.000 312.760 ;
    END
  END instr_addr_o[17]
  PIN instr_addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 325.760 1400.000 326.360 ;
    END
  END instr_addr_o[18]
  PIN instr_addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 339.360 1400.000 339.960 ;
    END
  END instr_addr_o[19]
  PIN instr_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 51.040 1400.000 51.640 ;
    END
  END instr_addr_o[1]
  PIN instr_addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 352.960 1400.000 353.560 ;
    END
  END instr_addr_o[20]
  PIN instr_addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 366.560 1400.000 367.160 ;
    END
  END instr_addr_o[21]
  PIN instr_addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 380.840 1400.000 381.440 ;
    END
  END instr_addr_o[22]
  PIN instr_addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 394.440 1400.000 395.040 ;
    END
  END instr_addr_o[23]
  PIN instr_addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 408.040 1400.000 408.640 ;
    END
  END instr_addr_o[24]
  PIN instr_addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 421.640 1400.000 422.240 ;
    END
  END instr_addr_o[25]
  PIN instr_addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 435.240 1400.000 435.840 ;
    END
  END instr_addr_o[26]
  PIN instr_addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 449.520 1400.000 450.120 ;
    END
  END instr_addr_o[27]
  PIN instr_addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 463.120 1400.000 463.720 ;
    END
  END instr_addr_o[28]
  PIN instr_addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 476.720 1400.000 477.320 ;
    END
  END instr_addr_o[29]
  PIN instr_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 71.440 1400.000 72.040 ;
    END
  END instr_addr_o[2]
  PIN instr_addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 490.320 1400.000 490.920 ;
    END
  END instr_addr_o[30]
  PIN instr_addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 503.920 1400.000 504.520 ;
    END
  END instr_addr_o[31]
  PIN instr_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 92.520 1400.000 93.120 ;
    END
  END instr_addr_o[3]
  PIN instr_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 112.920 1400.000 113.520 ;
    END
  END instr_addr_o[4]
  PIN instr_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 133.320 1400.000 133.920 ;
    END
  END instr_addr_o[5]
  PIN instr_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 154.400 1400.000 155.000 ;
    END
  END instr_addr_o[6]
  PIN instr_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 174.800 1400.000 175.400 ;
    END
  END instr_addr_o[7]
  PIN instr_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 188.400 1400.000 189.000 ;
    END
  END instr_addr_o[8]
  PIN instr_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 202.000 1400.000 202.600 ;
    END
  END instr_addr_o[9]
  PIN instr_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 3.440 1400.000 4.040 ;
    END
  END instr_err_i
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 10.240 1400.000 10.840 ;
    END
  END instr_gnt_i
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 37.440 1400.000 38.040 ;
    END
  END instr_rdata_i[0]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 222.400 1400.000 223.000 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 236.680 1400.000 237.280 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 250.280 1400.000 250.880 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 263.880 1400.000 264.480 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 277.480 1400.000 278.080 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 291.080 1400.000 291.680 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 305.360 1400.000 305.960 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 318.960 1400.000 319.560 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 332.560 1400.000 333.160 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 346.160 1400.000 346.760 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 57.840 1400.000 58.440 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 359.760 1400.000 360.360 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 374.040 1400.000 374.640 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 387.640 1400.000 388.240 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 401.240 1400.000 401.840 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 414.840 1400.000 415.440 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 428.440 1400.000 429.040 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 442.040 1400.000 442.640 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 456.320 1400.000 456.920 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 469.920 1400.000 470.520 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 483.520 1400.000 484.120 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 78.920 1400.000 79.520 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 497.120 1400.000 497.720 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 510.720 1400.000 511.320 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 99.320 1400.000 99.920 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 119.720 1400.000 120.320 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 140.120 1400.000 140.720 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 161.200 1400.000 161.800 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 181.600 1400.000 182.200 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 195.200 1400.000 195.800 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 208.800 1400.000 209.400 ;
    END
  END instr_rdata_i[9]
  PIN instr_rdata_intg_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 44.240 1400.000 44.840 ;
    END
  END instr_rdata_intg_i[0]
  PIN instr_rdata_intg_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 64.640 1400.000 65.240 ;
    END
  END instr_rdata_intg_i[1]
  PIN instr_rdata_intg_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 85.720 1400.000 86.320 ;
    END
  END instr_rdata_intg_i[2]
  PIN instr_rdata_intg_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 106.120 1400.000 106.720 ;
    END
  END instr_rdata_intg_i[3]
  PIN instr_rdata_intg_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 126.520 1400.000 127.120 ;
    END
  END instr_rdata_intg_i[4]
  PIN instr_rdata_intg_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 146.920 1400.000 147.520 ;
    END
  END instr_rdata_intg_i[5]
  PIN instr_rdata_intg_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 168.000 1400.000 168.600 ;
    END
  END instr_rdata_intg_i[6]
  PIN instr_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 17.040 1400.000 17.640 ;
    END
  END instr_req_o
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 23.840 1400.000 24.440 ;
    END
  END instr_rvalid_i
  PIN irq_external_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END irq_external_i
  PIN irq_fast_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END irq_fast_i[0]
  PIN irq_fast_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END irq_fast_i[10]
  PIN irq_fast_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END irq_fast_i[11]
  PIN irq_fast_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END irq_fast_i[12]
  PIN irq_fast_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 1396.000 593.770 1400.000 ;
    END
  END irq_fast_i[13]
  PIN irq_fast_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END irq_fast_i[14]
  PIN irq_fast_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 1396.000 194.030 1400.000 ;
    END
  END irq_fast_i[1]
  PIN irq_fast_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END irq_fast_i[2]
  PIN irq_fast_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END irq_fast_i[3]
  PIN irq_fast_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END irq_fast_i[4]
  PIN irq_fast_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END irq_fast_i[5]
  PIN irq_fast_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END irq_fast_i[6]
  PIN irq_fast_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 737.160 1400.000 737.760 ;
    END
  END irq_fast_i[7]
  PIN irq_fast_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 765.040 1400.000 765.640 ;
    END
  END irq_fast_i[8]
  PIN irq_fast_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 778.640 1400.000 779.240 ;
    END
  END irq_fast_i[9]
  PIN irq_nm_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END irq_nm_i
  PIN irq_software_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1396.000 531.800 1400.000 532.400 ;
    END
  END irq_software_i
  PIN irq_timer_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 1396.000 64.310 1400.000 ;
    END
  END irq_timer_i
  PIN ram_cfg_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 1396.000 76.270 1400.000 ;
    END
  END ram_cfg_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 1396.000 88.230 1400.000 ;
    END
  END rst_ni
  PIN scan_rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END scan_rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END test_en_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 10.640 1222.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.040 10.640 1272.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1321.040 10.640 1322.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.040 10.640 1372.640 1387.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.040 10.640 147.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 10.640 247.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.040 10.640 297.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.040 10.640 347.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 10.640 397.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.040 10.640 447.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.040 10.640 497.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 10.640 547.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.040 10.640 597.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.040 10.640 647.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 10.640 697.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.040 10.640 747.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.040 10.640 797.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 10.640 847.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 896.040 10.640 897.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.040 10.640 947.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.040 10.640 997.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1046.040 10.640 1047.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.040 10.640 1097.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.040 10.640 1147.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1196.040 10.640 1197.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.040 10.640 1247.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1296.040 10.640 1297.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1346.040 10.640 1347.640 1387.440 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 3.825 1396.415 1389.495 ;
      LAYER met1 ;
        RECT 5.520 3.780 1396.475 1389.540 ;
      LAYER met2 ;
        RECT 6.170 1395.720 16.830 1396.565 ;
        RECT 17.670 1395.720 28.790 1396.565 ;
        RECT 29.630 1395.720 40.290 1396.565 ;
        RECT 41.130 1395.720 52.250 1396.565 ;
        RECT 53.090 1395.720 63.750 1396.565 ;
        RECT 64.590 1395.720 75.710 1396.565 ;
        RECT 76.550 1395.720 87.670 1396.565 ;
        RECT 88.510 1395.720 99.170 1396.565 ;
        RECT 100.010 1395.720 111.130 1396.565 ;
        RECT 111.970 1395.720 122.630 1396.565 ;
        RECT 123.470 1395.720 134.590 1396.565 ;
        RECT 135.430 1395.720 146.090 1396.565 ;
        RECT 146.930 1395.720 158.050 1396.565 ;
        RECT 158.890 1395.720 170.010 1396.565 ;
        RECT 170.850 1395.720 181.510 1396.565 ;
        RECT 182.350 1395.720 193.470 1396.565 ;
        RECT 194.310 1395.720 204.970 1396.565 ;
        RECT 205.810 1395.720 216.930 1396.565 ;
        RECT 217.770 1395.720 228.430 1396.565 ;
        RECT 229.270 1395.720 240.390 1396.565 ;
        RECT 241.230 1395.720 252.350 1396.565 ;
        RECT 253.190 1395.720 263.850 1396.565 ;
        RECT 264.690 1395.720 275.810 1396.565 ;
        RECT 276.650 1395.720 287.310 1396.565 ;
        RECT 288.150 1395.720 299.270 1396.565 ;
        RECT 300.110 1395.720 310.770 1396.565 ;
        RECT 311.610 1395.720 322.730 1396.565 ;
        RECT 323.570 1395.720 334.690 1396.565 ;
        RECT 335.530 1395.720 346.190 1396.565 ;
        RECT 347.030 1395.720 358.150 1396.565 ;
        RECT 358.990 1395.720 369.650 1396.565 ;
        RECT 370.490 1395.720 381.610 1396.565 ;
        RECT 382.450 1395.720 393.110 1396.565 ;
        RECT 393.950 1395.720 405.070 1396.565 ;
        RECT 405.910 1395.720 417.030 1396.565 ;
        RECT 417.870 1395.720 428.530 1396.565 ;
        RECT 429.370 1395.720 440.490 1396.565 ;
        RECT 441.330 1395.720 451.990 1396.565 ;
        RECT 452.830 1395.720 463.950 1396.565 ;
        RECT 464.790 1395.720 475.450 1396.565 ;
        RECT 476.290 1395.720 487.410 1396.565 ;
        RECT 488.250 1395.720 499.370 1396.565 ;
        RECT 500.210 1395.720 510.870 1396.565 ;
        RECT 511.710 1395.720 522.830 1396.565 ;
        RECT 523.670 1395.720 534.330 1396.565 ;
        RECT 535.170 1395.720 546.290 1396.565 ;
        RECT 547.130 1395.720 557.790 1396.565 ;
        RECT 558.630 1395.720 569.750 1396.565 ;
        RECT 570.590 1395.720 581.710 1396.565 ;
        RECT 582.550 1395.720 593.210 1396.565 ;
        RECT 594.050 1395.720 605.170 1396.565 ;
        RECT 606.010 1395.720 616.670 1396.565 ;
        RECT 617.510 1395.720 628.630 1396.565 ;
        RECT 629.470 1395.720 640.130 1396.565 ;
        RECT 640.970 1395.720 652.090 1396.565 ;
        RECT 652.930 1395.720 664.050 1396.565 ;
        RECT 664.890 1395.720 675.550 1396.565 ;
        RECT 676.390 1395.720 687.510 1396.565 ;
        RECT 688.350 1395.720 699.010 1396.565 ;
        RECT 699.850 1395.720 710.970 1396.565 ;
        RECT 711.810 1395.720 722.470 1396.565 ;
        RECT 723.310 1395.720 734.430 1396.565 ;
        RECT 735.270 1395.720 746.390 1396.565 ;
        RECT 747.230 1395.720 757.890 1396.565 ;
        RECT 758.730 1395.720 769.850 1396.565 ;
        RECT 770.690 1395.720 781.350 1396.565 ;
        RECT 782.190 1395.720 793.310 1396.565 ;
        RECT 794.150 1395.720 804.810 1396.565 ;
        RECT 805.650 1395.720 816.770 1396.565 ;
        RECT 817.610 1395.720 828.730 1396.565 ;
        RECT 829.570 1395.720 840.230 1396.565 ;
        RECT 841.070 1395.720 852.190 1396.565 ;
        RECT 853.030 1395.720 863.690 1396.565 ;
        RECT 864.530 1395.720 875.650 1396.565 ;
        RECT 876.490 1395.720 887.150 1396.565 ;
        RECT 887.990 1395.720 899.110 1396.565 ;
        RECT 899.950 1395.720 911.070 1396.565 ;
        RECT 911.910 1395.720 922.570 1396.565 ;
        RECT 923.410 1395.720 934.530 1396.565 ;
        RECT 935.370 1395.720 946.030 1396.565 ;
        RECT 946.870 1395.720 957.990 1396.565 ;
        RECT 958.830 1395.720 969.490 1396.565 ;
        RECT 970.330 1395.720 981.450 1396.565 ;
        RECT 982.290 1395.720 993.410 1396.565 ;
        RECT 994.250 1395.720 1004.910 1396.565 ;
        RECT 1005.750 1395.720 1016.870 1396.565 ;
        RECT 1017.710 1395.720 1028.370 1396.565 ;
        RECT 1029.210 1395.720 1040.330 1396.565 ;
        RECT 1041.170 1395.720 1051.830 1396.565 ;
        RECT 1052.670 1395.720 1063.790 1396.565 ;
        RECT 1064.630 1395.720 1075.750 1396.565 ;
        RECT 1076.590 1395.720 1087.250 1396.565 ;
        RECT 1088.090 1395.720 1099.210 1396.565 ;
        RECT 1100.050 1395.720 1110.710 1396.565 ;
        RECT 1111.550 1395.720 1122.670 1396.565 ;
        RECT 1123.510 1395.720 1134.170 1396.565 ;
        RECT 1135.010 1395.720 1146.130 1396.565 ;
        RECT 1146.970 1395.720 1158.090 1396.565 ;
        RECT 1158.930 1395.720 1169.590 1396.565 ;
        RECT 1170.430 1395.720 1181.550 1396.565 ;
        RECT 1182.390 1395.720 1193.050 1396.565 ;
        RECT 1193.890 1395.720 1205.010 1396.565 ;
        RECT 1205.850 1395.720 1216.510 1396.565 ;
        RECT 1217.350 1395.720 1228.470 1396.565 ;
        RECT 1229.310 1395.720 1240.430 1396.565 ;
        RECT 1241.270 1395.720 1251.930 1396.565 ;
        RECT 1252.770 1395.720 1263.890 1396.565 ;
        RECT 1264.730 1395.720 1275.390 1396.565 ;
        RECT 1276.230 1395.720 1287.350 1396.565 ;
        RECT 1288.190 1395.720 1298.850 1396.565 ;
        RECT 1299.690 1395.720 1310.810 1396.565 ;
        RECT 1311.650 1395.720 1322.770 1396.565 ;
        RECT 1323.610 1395.720 1334.270 1396.565 ;
        RECT 1335.110 1395.720 1346.230 1396.565 ;
        RECT 1347.070 1395.720 1357.730 1396.565 ;
        RECT 1358.570 1395.720 1369.690 1396.565 ;
        RECT 1370.530 1395.720 1381.190 1396.565 ;
        RECT 1382.030 1395.720 1393.150 1396.565 ;
        RECT 1393.990 1395.720 1395.090 1396.565 ;
        RECT 5.620 4.280 1395.090 1395.720 ;
        RECT 6.170 3.555 16.370 4.280 ;
        RECT 17.210 3.555 27.410 4.280 ;
        RECT 28.250 3.555 38.450 4.280 ;
        RECT 39.290 3.555 49.490 4.280 ;
        RECT 50.330 3.555 60.530 4.280 ;
        RECT 61.370 3.555 71.570 4.280 ;
        RECT 72.410 3.555 83.070 4.280 ;
        RECT 83.910 3.555 94.110 4.280 ;
        RECT 94.950 3.555 105.150 4.280 ;
        RECT 105.990 3.555 116.190 4.280 ;
        RECT 117.030 3.555 127.230 4.280 ;
        RECT 128.070 3.555 138.270 4.280 ;
        RECT 139.110 3.555 149.310 4.280 ;
        RECT 150.150 3.555 160.810 4.280 ;
        RECT 161.650 3.555 171.850 4.280 ;
        RECT 172.690 3.555 182.890 4.280 ;
        RECT 183.730 3.555 193.930 4.280 ;
        RECT 194.770 3.555 204.970 4.280 ;
        RECT 205.810 3.555 216.010 4.280 ;
        RECT 216.850 3.555 227.510 4.280 ;
        RECT 228.350 3.555 238.550 4.280 ;
        RECT 239.390 3.555 249.590 4.280 ;
        RECT 250.430 3.555 260.630 4.280 ;
        RECT 261.470 3.555 271.670 4.280 ;
        RECT 272.510 3.555 282.710 4.280 ;
        RECT 283.550 3.555 293.750 4.280 ;
        RECT 294.590 3.555 305.250 4.280 ;
        RECT 306.090 3.555 316.290 4.280 ;
        RECT 317.130 3.555 327.330 4.280 ;
        RECT 328.170 3.555 338.370 4.280 ;
        RECT 339.210 3.555 349.410 4.280 ;
        RECT 350.250 3.555 360.450 4.280 ;
        RECT 361.290 3.555 371.490 4.280 ;
        RECT 372.330 3.555 382.990 4.280 ;
        RECT 383.830 3.555 394.030 4.280 ;
        RECT 394.870 3.555 405.070 4.280 ;
        RECT 405.910 3.555 416.110 4.280 ;
        RECT 416.950 3.555 427.150 4.280 ;
        RECT 427.990 3.555 438.190 4.280 ;
        RECT 439.030 3.555 449.690 4.280 ;
        RECT 450.530 3.555 460.730 4.280 ;
        RECT 461.570 3.555 471.770 4.280 ;
        RECT 472.610 3.555 482.810 4.280 ;
        RECT 483.650 3.555 493.850 4.280 ;
        RECT 494.690 3.555 504.890 4.280 ;
        RECT 505.730 3.555 515.930 4.280 ;
        RECT 516.770 3.555 527.430 4.280 ;
        RECT 528.270 3.555 538.470 4.280 ;
        RECT 539.310 3.555 549.510 4.280 ;
        RECT 550.350 3.555 560.550 4.280 ;
        RECT 561.390 3.555 571.590 4.280 ;
        RECT 572.430 3.555 582.630 4.280 ;
        RECT 583.470 3.555 593.670 4.280 ;
        RECT 594.510 3.555 605.170 4.280 ;
        RECT 606.010 3.555 616.210 4.280 ;
        RECT 617.050 3.555 627.250 4.280 ;
        RECT 628.090 3.555 638.290 4.280 ;
        RECT 639.130 3.555 649.330 4.280 ;
        RECT 650.170 3.555 660.370 4.280 ;
        RECT 661.210 3.555 671.870 4.280 ;
        RECT 672.710 3.555 682.910 4.280 ;
        RECT 683.750 3.555 693.950 4.280 ;
        RECT 694.790 3.555 704.990 4.280 ;
        RECT 705.830 3.555 716.030 4.280 ;
        RECT 716.870 3.555 727.070 4.280 ;
        RECT 727.910 3.555 738.110 4.280 ;
        RECT 738.950 3.555 749.610 4.280 ;
        RECT 750.450 3.555 760.650 4.280 ;
        RECT 761.490 3.555 771.690 4.280 ;
        RECT 772.530 3.555 782.730 4.280 ;
        RECT 783.570 3.555 793.770 4.280 ;
        RECT 794.610 3.555 804.810 4.280 ;
        RECT 805.650 3.555 816.310 4.280 ;
        RECT 817.150 3.555 827.350 4.280 ;
        RECT 828.190 3.555 838.390 4.280 ;
        RECT 839.230 3.555 849.430 4.280 ;
        RECT 850.270 3.555 860.470 4.280 ;
        RECT 861.310 3.555 871.510 4.280 ;
        RECT 872.350 3.555 882.550 4.280 ;
        RECT 883.390 3.555 894.050 4.280 ;
        RECT 894.890 3.555 905.090 4.280 ;
        RECT 905.930 3.555 916.130 4.280 ;
        RECT 916.970 3.555 927.170 4.280 ;
        RECT 928.010 3.555 938.210 4.280 ;
        RECT 939.050 3.555 949.250 4.280 ;
        RECT 950.090 3.555 960.290 4.280 ;
        RECT 961.130 3.555 971.790 4.280 ;
        RECT 972.630 3.555 982.830 4.280 ;
        RECT 983.670 3.555 993.870 4.280 ;
        RECT 994.710 3.555 1004.910 4.280 ;
        RECT 1005.750 3.555 1015.950 4.280 ;
        RECT 1016.790 3.555 1026.990 4.280 ;
        RECT 1027.830 3.555 1038.490 4.280 ;
        RECT 1039.330 3.555 1049.530 4.280 ;
        RECT 1050.370 3.555 1060.570 4.280 ;
        RECT 1061.410 3.555 1071.610 4.280 ;
        RECT 1072.450 3.555 1082.650 4.280 ;
        RECT 1083.490 3.555 1093.690 4.280 ;
        RECT 1094.530 3.555 1104.730 4.280 ;
        RECT 1105.570 3.555 1116.230 4.280 ;
        RECT 1117.070 3.555 1127.270 4.280 ;
        RECT 1128.110 3.555 1138.310 4.280 ;
        RECT 1139.150 3.555 1149.350 4.280 ;
        RECT 1150.190 3.555 1160.390 4.280 ;
        RECT 1161.230 3.555 1171.430 4.280 ;
        RECT 1172.270 3.555 1182.470 4.280 ;
        RECT 1183.310 3.555 1193.970 4.280 ;
        RECT 1194.810 3.555 1205.010 4.280 ;
        RECT 1205.850 3.555 1216.050 4.280 ;
        RECT 1216.890 3.555 1227.090 4.280 ;
        RECT 1227.930 3.555 1238.130 4.280 ;
        RECT 1238.970 3.555 1249.170 4.280 ;
        RECT 1250.010 3.555 1260.670 4.280 ;
        RECT 1261.510 3.555 1271.710 4.280 ;
        RECT 1272.550 3.555 1282.750 4.280 ;
        RECT 1283.590 3.555 1293.790 4.280 ;
        RECT 1294.630 3.555 1304.830 4.280 ;
        RECT 1305.670 3.555 1315.870 4.280 ;
        RECT 1316.710 3.555 1326.910 4.280 ;
        RECT 1327.750 3.555 1338.410 4.280 ;
        RECT 1339.250 3.555 1349.450 4.280 ;
        RECT 1350.290 3.555 1360.490 4.280 ;
        RECT 1361.330 3.555 1371.530 4.280 ;
        RECT 1372.370 3.555 1382.570 4.280 ;
        RECT 1383.410 3.555 1393.610 4.280 ;
        RECT 1394.450 3.555 1395.090 4.280 ;
      LAYER met3 ;
        RECT 4.000 1395.680 1395.600 1396.545 ;
        RECT 4.000 1395.040 1396.000 1395.680 ;
        RECT 4.400 1393.640 1396.000 1395.040 ;
        RECT 4.000 1390.280 1396.000 1393.640 ;
        RECT 4.000 1388.880 1395.600 1390.280 ;
        RECT 4.000 1384.840 1396.000 1388.880 ;
        RECT 4.400 1383.480 1396.000 1384.840 ;
        RECT 4.400 1383.440 1395.600 1383.480 ;
        RECT 4.000 1382.080 1395.600 1383.440 ;
        RECT 4.000 1376.680 1396.000 1382.080 ;
        RECT 4.000 1375.280 1395.600 1376.680 ;
        RECT 4.000 1374.640 1396.000 1375.280 ;
        RECT 4.400 1373.240 1396.000 1374.640 ;
        RECT 4.000 1369.880 1396.000 1373.240 ;
        RECT 4.000 1368.480 1395.600 1369.880 ;
        RECT 4.000 1363.760 1396.000 1368.480 ;
        RECT 4.400 1363.080 1396.000 1363.760 ;
        RECT 4.400 1362.360 1395.600 1363.080 ;
        RECT 4.000 1361.680 1395.600 1362.360 ;
        RECT 4.000 1356.280 1396.000 1361.680 ;
        RECT 4.000 1354.880 1395.600 1356.280 ;
        RECT 4.000 1353.560 1396.000 1354.880 ;
        RECT 4.400 1352.160 1396.000 1353.560 ;
        RECT 4.000 1349.480 1396.000 1352.160 ;
        RECT 4.000 1348.080 1395.600 1349.480 ;
        RECT 4.000 1343.360 1396.000 1348.080 ;
        RECT 4.400 1342.680 1396.000 1343.360 ;
        RECT 4.400 1341.960 1395.600 1342.680 ;
        RECT 4.000 1341.280 1395.600 1341.960 ;
        RECT 4.000 1335.880 1396.000 1341.280 ;
        RECT 4.000 1334.480 1395.600 1335.880 ;
        RECT 4.000 1333.160 1396.000 1334.480 ;
        RECT 4.400 1331.760 1396.000 1333.160 ;
        RECT 4.000 1328.400 1396.000 1331.760 ;
        RECT 4.000 1327.000 1395.600 1328.400 ;
        RECT 4.000 1322.280 1396.000 1327.000 ;
        RECT 4.400 1321.600 1396.000 1322.280 ;
        RECT 4.400 1320.880 1395.600 1321.600 ;
        RECT 4.000 1320.200 1395.600 1320.880 ;
        RECT 4.000 1314.800 1396.000 1320.200 ;
        RECT 4.000 1313.400 1395.600 1314.800 ;
        RECT 4.000 1312.080 1396.000 1313.400 ;
        RECT 4.400 1310.680 1396.000 1312.080 ;
        RECT 4.000 1308.000 1396.000 1310.680 ;
        RECT 4.000 1306.600 1395.600 1308.000 ;
        RECT 4.000 1301.880 1396.000 1306.600 ;
        RECT 4.400 1301.200 1396.000 1301.880 ;
        RECT 4.400 1300.480 1395.600 1301.200 ;
        RECT 4.000 1299.800 1395.600 1300.480 ;
        RECT 4.000 1294.400 1396.000 1299.800 ;
        RECT 4.000 1293.000 1395.600 1294.400 ;
        RECT 4.000 1291.680 1396.000 1293.000 ;
        RECT 4.400 1290.280 1396.000 1291.680 ;
        RECT 4.000 1287.600 1396.000 1290.280 ;
        RECT 4.000 1286.200 1395.600 1287.600 ;
        RECT 4.000 1280.800 1396.000 1286.200 ;
        RECT 4.400 1279.400 1395.600 1280.800 ;
        RECT 4.000 1274.000 1396.000 1279.400 ;
        RECT 4.000 1272.600 1395.600 1274.000 ;
        RECT 4.000 1270.600 1396.000 1272.600 ;
        RECT 4.400 1269.200 1396.000 1270.600 ;
        RECT 4.000 1267.200 1396.000 1269.200 ;
        RECT 4.000 1265.800 1395.600 1267.200 ;
        RECT 4.000 1260.400 1396.000 1265.800 ;
        RECT 4.400 1259.000 1395.600 1260.400 ;
        RECT 4.000 1252.920 1396.000 1259.000 ;
        RECT 4.000 1251.520 1395.600 1252.920 ;
        RECT 4.000 1250.200 1396.000 1251.520 ;
        RECT 4.400 1248.800 1396.000 1250.200 ;
        RECT 4.000 1246.120 1396.000 1248.800 ;
        RECT 4.000 1244.720 1395.600 1246.120 ;
        RECT 4.000 1239.320 1396.000 1244.720 ;
        RECT 4.400 1237.920 1395.600 1239.320 ;
        RECT 4.000 1232.520 1396.000 1237.920 ;
        RECT 4.000 1231.120 1395.600 1232.520 ;
        RECT 4.000 1229.120 1396.000 1231.120 ;
        RECT 4.400 1227.720 1396.000 1229.120 ;
        RECT 4.000 1225.720 1396.000 1227.720 ;
        RECT 4.000 1224.320 1395.600 1225.720 ;
        RECT 4.000 1218.920 1396.000 1224.320 ;
        RECT 4.400 1217.520 1395.600 1218.920 ;
        RECT 4.000 1212.120 1396.000 1217.520 ;
        RECT 4.000 1210.720 1395.600 1212.120 ;
        RECT 4.000 1208.720 1396.000 1210.720 ;
        RECT 4.400 1207.320 1396.000 1208.720 ;
        RECT 4.000 1205.320 1396.000 1207.320 ;
        RECT 4.000 1203.920 1395.600 1205.320 ;
        RECT 4.000 1198.520 1396.000 1203.920 ;
        RECT 4.000 1197.840 1395.600 1198.520 ;
        RECT 4.400 1197.120 1395.600 1197.840 ;
        RECT 4.400 1196.440 1396.000 1197.120 ;
        RECT 4.000 1191.720 1396.000 1196.440 ;
        RECT 4.000 1190.320 1395.600 1191.720 ;
        RECT 4.000 1187.640 1396.000 1190.320 ;
        RECT 4.400 1186.240 1396.000 1187.640 ;
        RECT 4.000 1184.920 1396.000 1186.240 ;
        RECT 4.000 1183.520 1395.600 1184.920 ;
        RECT 4.000 1177.440 1396.000 1183.520 ;
        RECT 4.400 1176.040 1395.600 1177.440 ;
        RECT 4.000 1170.640 1396.000 1176.040 ;
        RECT 4.000 1169.240 1395.600 1170.640 ;
        RECT 4.000 1167.240 1396.000 1169.240 ;
        RECT 4.400 1165.840 1396.000 1167.240 ;
        RECT 4.000 1163.840 1396.000 1165.840 ;
        RECT 4.000 1162.440 1395.600 1163.840 ;
        RECT 4.000 1157.040 1396.000 1162.440 ;
        RECT 4.000 1156.360 1395.600 1157.040 ;
        RECT 4.400 1155.640 1395.600 1156.360 ;
        RECT 4.400 1154.960 1396.000 1155.640 ;
        RECT 4.000 1150.240 1396.000 1154.960 ;
        RECT 4.000 1148.840 1395.600 1150.240 ;
        RECT 4.000 1146.160 1396.000 1148.840 ;
        RECT 4.400 1144.760 1396.000 1146.160 ;
        RECT 4.000 1143.440 1396.000 1144.760 ;
        RECT 4.000 1142.040 1395.600 1143.440 ;
        RECT 4.000 1136.640 1396.000 1142.040 ;
        RECT 4.000 1135.960 1395.600 1136.640 ;
        RECT 4.400 1135.240 1395.600 1135.960 ;
        RECT 4.400 1134.560 1396.000 1135.240 ;
        RECT 4.000 1129.840 1396.000 1134.560 ;
        RECT 4.000 1128.440 1395.600 1129.840 ;
        RECT 4.000 1125.760 1396.000 1128.440 ;
        RECT 4.400 1124.360 1396.000 1125.760 ;
        RECT 4.000 1123.040 1396.000 1124.360 ;
        RECT 4.000 1121.640 1395.600 1123.040 ;
        RECT 4.000 1116.240 1396.000 1121.640 ;
        RECT 4.000 1114.880 1395.600 1116.240 ;
        RECT 4.400 1114.840 1395.600 1114.880 ;
        RECT 4.400 1113.480 1396.000 1114.840 ;
        RECT 4.000 1108.760 1396.000 1113.480 ;
        RECT 4.000 1107.360 1395.600 1108.760 ;
        RECT 4.000 1104.680 1396.000 1107.360 ;
        RECT 4.400 1103.280 1396.000 1104.680 ;
        RECT 4.000 1101.960 1396.000 1103.280 ;
        RECT 4.000 1100.560 1395.600 1101.960 ;
        RECT 4.000 1095.160 1396.000 1100.560 ;
        RECT 4.000 1094.480 1395.600 1095.160 ;
        RECT 4.400 1093.760 1395.600 1094.480 ;
        RECT 4.400 1093.080 1396.000 1093.760 ;
        RECT 4.000 1088.360 1396.000 1093.080 ;
        RECT 4.000 1086.960 1395.600 1088.360 ;
        RECT 4.000 1084.280 1396.000 1086.960 ;
        RECT 4.400 1082.880 1396.000 1084.280 ;
        RECT 4.000 1081.560 1396.000 1082.880 ;
        RECT 4.000 1080.160 1395.600 1081.560 ;
        RECT 4.000 1074.760 1396.000 1080.160 ;
        RECT 4.000 1073.400 1395.600 1074.760 ;
        RECT 4.400 1073.360 1395.600 1073.400 ;
        RECT 4.400 1072.000 1396.000 1073.360 ;
        RECT 4.000 1067.960 1396.000 1072.000 ;
        RECT 4.000 1066.560 1395.600 1067.960 ;
        RECT 4.000 1063.200 1396.000 1066.560 ;
        RECT 4.400 1061.800 1396.000 1063.200 ;
        RECT 4.000 1061.160 1396.000 1061.800 ;
        RECT 4.000 1059.760 1395.600 1061.160 ;
        RECT 4.000 1054.360 1396.000 1059.760 ;
        RECT 4.000 1053.000 1395.600 1054.360 ;
        RECT 4.400 1052.960 1395.600 1053.000 ;
        RECT 4.400 1051.600 1396.000 1052.960 ;
        RECT 4.000 1047.560 1396.000 1051.600 ;
        RECT 4.000 1046.160 1395.600 1047.560 ;
        RECT 4.000 1042.800 1396.000 1046.160 ;
        RECT 4.400 1041.400 1396.000 1042.800 ;
        RECT 4.000 1040.760 1396.000 1041.400 ;
        RECT 4.000 1039.360 1395.600 1040.760 ;
        RECT 4.000 1033.280 1396.000 1039.360 ;
        RECT 4.000 1031.920 1395.600 1033.280 ;
        RECT 4.400 1031.880 1395.600 1031.920 ;
        RECT 4.400 1030.520 1396.000 1031.880 ;
        RECT 4.000 1026.480 1396.000 1030.520 ;
        RECT 4.000 1025.080 1395.600 1026.480 ;
        RECT 4.000 1021.720 1396.000 1025.080 ;
        RECT 4.400 1020.320 1396.000 1021.720 ;
        RECT 4.000 1019.680 1396.000 1020.320 ;
        RECT 4.000 1018.280 1395.600 1019.680 ;
        RECT 4.000 1012.880 1396.000 1018.280 ;
        RECT 4.000 1011.520 1395.600 1012.880 ;
        RECT 4.400 1011.480 1395.600 1011.520 ;
        RECT 4.400 1010.120 1396.000 1011.480 ;
        RECT 4.000 1006.080 1396.000 1010.120 ;
        RECT 4.000 1004.680 1395.600 1006.080 ;
        RECT 4.000 1001.320 1396.000 1004.680 ;
        RECT 4.400 999.920 1396.000 1001.320 ;
        RECT 4.000 999.280 1396.000 999.920 ;
        RECT 4.000 997.880 1395.600 999.280 ;
        RECT 4.000 992.480 1396.000 997.880 ;
        RECT 4.000 991.080 1395.600 992.480 ;
        RECT 4.000 990.440 1396.000 991.080 ;
        RECT 4.400 989.040 1396.000 990.440 ;
        RECT 4.000 985.680 1396.000 989.040 ;
        RECT 4.000 984.280 1395.600 985.680 ;
        RECT 4.000 980.240 1396.000 984.280 ;
        RECT 4.400 978.880 1396.000 980.240 ;
        RECT 4.400 978.840 1395.600 978.880 ;
        RECT 4.000 977.480 1395.600 978.840 ;
        RECT 4.000 972.080 1396.000 977.480 ;
        RECT 4.000 970.680 1395.600 972.080 ;
        RECT 4.000 970.040 1396.000 970.680 ;
        RECT 4.400 968.640 1396.000 970.040 ;
        RECT 4.000 965.280 1396.000 968.640 ;
        RECT 4.000 963.880 1395.600 965.280 ;
        RECT 4.000 959.840 1396.000 963.880 ;
        RECT 4.400 958.440 1396.000 959.840 ;
        RECT 4.000 957.800 1396.000 958.440 ;
        RECT 4.000 956.400 1395.600 957.800 ;
        RECT 4.000 951.000 1396.000 956.400 ;
        RECT 4.000 949.600 1395.600 951.000 ;
        RECT 4.000 948.960 1396.000 949.600 ;
        RECT 4.400 947.560 1396.000 948.960 ;
        RECT 4.000 944.200 1396.000 947.560 ;
        RECT 4.000 942.800 1395.600 944.200 ;
        RECT 4.000 938.760 1396.000 942.800 ;
        RECT 4.400 937.400 1396.000 938.760 ;
        RECT 4.400 937.360 1395.600 937.400 ;
        RECT 4.000 936.000 1395.600 937.360 ;
        RECT 4.000 930.600 1396.000 936.000 ;
        RECT 4.000 929.200 1395.600 930.600 ;
        RECT 4.000 928.560 1396.000 929.200 ;
        RECT 4.400 927.160 1396.000 928.560 ;
        RECT 4.000 923.800 1396.000 927.160 ;
        RECT 4.000 922.400 1395.600 923.800 ;
        RECT 4.000 918.360 1396.000 922.400 ;
        RECT 4.400 917.000 1396.000 918.360 ;
        RECT 4.400 916.960 1395.600 917.000 ;
        RECT 4.000 915.600 1395.600 916.960 ;
        RECT 4.000 910.200 1396.000 915.600 ;
        RECT 4.000 908.800 1395.600 910.200 ;
        RECT 4.000 907.480 1396.000 908.800 ;
        RECT 4.400 906.080 1396.000 907.480 ;
        RECT 4.000 903.400 1396.000 906.080 ;
        RECT 4.000 902.000 1395.600 903.400 ;
        RECT 4.000 897.280 1396.000 902.000 ;
        RECT 4.400 896.600 1396.000 897.280 ;
        RECT 4.400 895.880 1395.600 896.600 ;
        RECT 4.000 895.200 1395.600 895.880 ;
        RECT 4.000 889.800 1396.000 895.200 ;
        RECT 4.000 888.400 1395.600 889.800 ;
        RECT 4.000 887.080 1396.000 888.400 ;
        RECT 4.400 885.680 1396.000 887.080 ;
        RECT 4.000 882.320 1396.000 885.680 ;
        RECT 4.000 880.920 1395.600 882.320 ;
        RECT 4.000 876.880 1396.000 880.920 ;
        RECT 4.400 875.520 1396.000 876.880 ;
        RECT 4.400 875.480 1395.600 875.520 ;
        RECT 4.000 874.120 1395.600 875.480 ;
        RECT 4.000 868.720 1396.000 874.120 ;
        RECT 4.000 867.320 1395.600 868.720 ;
        RECT 4.000 866.000 1396.000 867.320 ;
        RECT 4.400 864.600 1396.000 866.000 ;
        RECT 4.000 861.920 1396.000 864.600 ;
        RECT 4.000 860.520 1395.600 861.920 ;
        RECT 4.000 855.800 1396.000 860.520 ;
        RECT 4.400 855.120 1396.000 855.800 ;
        RECT 4.400 854.400 1395.600 855.120 ;
        RECT 4.000 853.720 1395.600 854.400 ;
        RECT 4.000 848.320 1396.000 853.720 ;
        RECT 4.000 846.920 1395.600 848.320 ;
        RECT 4.000 845.600 1396.000 846.920 ;
        RECT 4.400 844.200 1396.000 845.600 ;
        RECT 4.000 841.520 1396.000 844.200 ;
        RECT 4.000 840.120 1395.600 841.520 ;
        RECT 4.000 835.400 1396.000 840.120 ;
        RECT 4.400 834.720 1396.000 835.400 ;
        RECT 4.400 834.000 1395.600 834.720 ;
        RECT 4.000 833.320 1395.600 834.000 ;
        RECT 4.000 827.920 1396.000 833.320 ;
        RECT 4.000 826.520 1395.600 827.920 ;
        RECT 4.000 824.520 1396.000 826.520 ;
        RECT 4.400 823.120 1396.000 824.520 ;
        RECT 4.000 821.120 1396.000 823.120 ;
        RECT 4.000 819.720 1395.600 821.120 ;
        RECT 4.000 814.320 1396.000 819.720 ;
        RECT 4.400 813.640 1396.000 814.320 ;
        RECT 4.400 812.920 1395.600 813.640 ;
        RECT 4.000 812.240 1395.600 812.920 ;
        RECT 4.000 806.840 1396.000 812.240 ;
        RECT 4.000 805.440 1395.600 806.840 ;
        RECT 4.000 804.120 1396.000 805.440 ;
        RECT 4.400 802.720 1396.000 804.120 ;
        RECT 4.000 800.040 1396.000 802.720 ;
        RECT 4.000 798.640 1395.600 800.040 ;
        RECT 4.000 793.920 1396.000 798.640 ;
        RECT 4.400 793.240 1396.000 793.920 ;
        RECT 4.400 792.520 1395.600 793.240 ;
        RECT 4.000 791.840 1395.600 792.520 ;
        RECT 4.000 786.440 1396.000 791.840 ;
        RECT 4.000 785.040 1395.600 786.440 ;
        RECT 4.000 783.040 1396.000 785.040 ;
        RECT 4.400 781.640 1396.000 783.040 ;
        RECT 4.000 779.640 1396.000 781.640 ;
        RECT 4.000 778.240 1395.600 779.640 ;
        RECT 4.000 772.840 1396.000 778.240 ;
        RECT 4.400 771.440 1395.600 772.840 ;
        RECT 4.000 766.040 1396.000 771.440 ;
        RECT 4.000 764.640 1395.600 766.040 ;
        RECT 4.000 762.640 1396.000 764.640 ;
        RECT 4.400 761.240 1396.000 762.640 ;
        RECT 4.000 759.240 1396.000 761.240 ;
        RECT 4.000 757.840 1395.600 759.240 ;
        RECT 4.000 752.440 1396.000 757.840 ;
        RECT 4.400 751.040 1395.600 752.440 ;
        RECT 4.000 745.640 1396.000 751.040 ;
        RECT 4.000 744.240 1395.600 745.640 ;
        RECT 4.000 741.560 1396.000 744.240 ;
        RECT 4.400 740.160 1396.000 741.560 ;
        RECT 4.000 738.160 1396.000 740.160 ;
        RECT 4.000 736.760 1395.600 738.160 ;
        RECT 4.000 731.360 1396.000 736.760 ;
        RECT 4.400 729.960 1395.600 731.360 ;
        RECT 4.000 724.560 1396.000 729.960 ;
        RECT 4.000 723.160 1395.600 724.560 ;
        RECT 4.000 721.160 1396.000 723.160 ;
        RECT 4.400 719.760 1396.000 721.160 ;
        RECT 4.000 717.760 1396.000 719.760 ;
        RECT 4.000 716.360 1395.600 717.760 ;
        RECT 4.000 710.960 1396.000 716.360 ;
        RECT 4.400 709.560 1395.600 710.960 ;
        RECT 4.000 704.160 1396.000 709.560 ;
        RECT 4.000 702.760 1395.600 704.160 ;
        RECT 4.000 700.080 1396.000 702.760 ;
        RECT 4.400 698.680 1396.000 700.080 ;
        RECT 4.000 697.360 1396.000 698.680 ;
        RECT 4.000 695.960 1395.600 697.360 ;
        RECT 4.000 690.560 1396.000 695.960 ;
        RECT 4.000 689.880 1395.600 690.560 ;
        RECT 4.400 689.160 1395.600 689.880 ;
        RECT 4.400 688.480 1396.000 689.160 ;
        RECT 4.000 683.760 1396.000 688.480 ;
        RECT 4.000 682.360 1395.600 683.760 ;
        RECT 4.000 679.680 1396.000 682.360 ;
        RECT 4.400 678.280 1396.000 679.680 ;
        RECT 4.000 676.960 1396.000 678.280 ;
        RECT 4.000 675.560 1395.600 676.960 ;
        RECT 4.000 670.160 1396.000 675.560 ;
        RECT 4.000 669.480 1395.600 670.160 ;
        RECT 4.400 668.760 1395.600 669.480 ;
        RECT 4.400 668.080 1396.000 668.760 ;
        RECT 4.000 662.680 1396.000 668.080 ;
        RECT 4.000 661.280 1395.600 662.680 ;
        RECT 4.000 658.600 1396.000 661.280 ;
        RECT 4.400 657.200 1396.000 658.600 ;
        RECT 4.000 655.880 1396.000 657.200 ;
        RECT 4.000 654.480 1395.600 655.880 ;
        RECT 4.000 649.080 1396.000 654.480 ;
        RECT 4.000 648.400 1395.600 649.080 ;
        RECT 4.400 647.680 1395.600 648.400 ;
        RECT 4.400 647.000 1396.000 647.680 ;
        RECT 4.000 642.280 1396.000 647.000 ;
        RECT 4.000 640.880 1395.600 642.280 ;
        RECT 4.000 638.200 1396.000 640.880 ;
        RECT 4.400 636.800 1396.000 638.200 ;
        RECT 4.000 635.480 1396.000 636.800 ;
        RECT 4.000 634.080 1395.600 635.480 ;
        RECT 4.000 628.680 1396.000 634.080 ;
        RECT 4.000 628.000 1395.600 628.680 ;
        RECT 4.400 627.280 1395.600 628.000 ;
        RECT 4.400 626.600 1396.000 627.280 ;
        RECT 4.000 621.880 1396.000 626.600 ;
        RECT 4.000 620.480 1395.600 621.880 ;
        RECT 4.000 617.120 1396.000 620.480 ;
        RECT 4.400 615.720 1396.000 617.120 ;
        RECT 4.000 615.080 1396.000 615.720 ;
        RECT 4.000 613.680 1395.600 615.080 ;
        RECT 4.000 608.280 1396.000 613.680 ;
        RECT 4.000 606.920 1395.600 608.280 ;
        RECT 4.400 606.880 1395.600 606.920 ;
        RECT 4.400 605.520 1396.000 606.880 ;
        RECT 4.000 601.480 1396.000 605.520 ;
        RECT 4.000 600.080 1395.600 601.480 ;
        RECT 4.000 596.720 1396.000 600.080 ;
        RECT 4.400 595.320 1396.000 596.720 ;
        RECT 4.000 594.680 1396.000 595.320 ;
        RECT 4.000 593.280 1395.600 594.680 ;
        RECT 4.000 587.200 1396.000 593.280 ;
        RECT 4.000 586.520 1395.600 587.200 ;
        RECT 4.400 585.800 1395.600 586.520 ;
        RECT 4.400 585.120 1396.000 585.800 ;
        RECT 4.000 580.400 1396.000 585.120 ;
        RECT 4.000 579.000 1395.600 580.400 ;
        RECT 4.000 575.640 1396.000 579.000 ;
        RECT 4.400 574.240 1396.000 575.640 ;
        RECT 4.000 573.600 1396.000 574.240 ;
        RECT 4.000 572.200 1395.600 573.600 ;
        RECT 4.000 566.800 1396.000 572.200 ;
        RECT 4.000 565.440 1395.600 566.800 ;
        RECT 4.400 565.400 1395.600 565.440 ;
        RECT 4.400 564.040 1396.000 565.400 ;
        RECT 4.000 560.000 1396.000 564.040 ;
        RECT 4.000 558.600 1395.600 560.000 ;
        RECT 4.000 555.240 1396.000 558.600 ;
        RECT 4.400 553.840 1396.000 555.240 ;
        RECT 4.000 553.200 1396.000 553.840 ;
        RECT 4.000 551.800 1395.600 553.200 ;
        RECT 4.000 546.400 1396.000 551.800 ;
        RECT 4.000 545.040 1395.600 546.400 ;
        RECT 4.400 545.000 1395.600 545.040 ;
        RECT 4.400 543.640 1396.000 545.000 ;
        RECT 4.000 539.600 1396.000 543.640 ;
        RECT 4.000 538.200 1395.600 539.600 ;
        RECT 4.000 534.160 1396.000 538.200 ;
        RECT 4.400 532.800 1396.000 534.160 ;
        RECT 4.400 532.760 1395.600 532.800 ;
        RECT 4.000 531.400 1395.600 532.760 ;
        RECT 4.000 526.000 1396.000 531.400 ;
        RECT 4.000 524.600 1395.600 526.000 ;
        RECT 4.000 523.960 1396.000 524.600 ;
        RECT 4.400 522.560 1396.000 523.960 ;
        RECT 4.000 518.520 1396.000 522.560 ;
        RECT 4.000 517.120 1395.600 518.520 ;
        RECT 4.000 513.760 1396.000 517.120 ;
        RECT 4.400 512.360 1396.000 513.760 ;
        RECT 4.000 511.720 1396.000 512.360 ;
        RECT 4.000 510.320 1395.600 511.720 ;
        RECT 4.000 504.920 1396.000 510.320 ;
        RECT 4.000 503.560 1395.600 504.920 ;
        RECT 4.400 503.520 1395.600 503.560 ;
        RECT 4.400 502.160 1396.000 503.520 ;
        RECT 4.000 498.120 1396.000 502.160 ;
        RECT 4.000 496.720 1395.600 498.120 ;
        RECT 4.000 492.680 1396.000 496.720 ;
        RECT 4.400 491.320 1396.000 492.680 ;
        RECT 4.400 491.280 1395.600 491.320 ;
        RECT 4.000 489.920 1395.600 491.280 ;
        RECT 4.000 484.520 1396.000 489.920 ;
        RECT 4.000 483.120 1395.600 484.520 ;
        RECT 4.000 482.480 1396.000 483.120 ;
        RECT 4.400 481.080 1396.000 482.480 ;
        RECT 4.000 477.720 1396.000 481.080 ;
        RECT 4.000 476.320 1395.600 477.720 ;
        RECT 4.000 472.280 1396.000 476.320 ;
        RECT 4.400 470.920 1396.000 472.280 ;
        RECT 4.400 470.880 1395.600 470.920 ;
        RECT 4.000 469.520 1395.600 470.880 ;
        RECT 4.000 464.120 1396.000 469.520 ;
        RECT 4.000 462.720 1395.600 464.120 ;
        RECT 4.000 462.080 1396.000 462.720 ;
        RECT 4.400 460.680 1396.000 462.080 ;
        RECT 4.000 457.320 1396.000 460.680 ;
        RECT 4.000 455.920 1395.600 457.320 ;
        RECT 4.000 451.200 1396.000 455.920 ;
        RECT 4.400 450.520 1396.000 451.200 ;
        RECT 4.400 449.800 1395.600 450.520 ;
        RECT 4.000 449.120 1395.600 449.800 ;
        RECT 4.000 443.040 1396.000 449.120 ;
        RECT 4.000 441.640 1395.600 443.040 ;
        RECT 4.000 441.000 1396.000 441.640 ;
        RECT 4.400 439.600 1396.000 441.000 ;
        RECT 4.000 436.240 1396.000 439.600 ;
        RECT 4.000 434.840 1395.600 436.240 ;
        RECT 4.000 430.800 1396.000 434.840 ;
        RECT 4.400 429.440 1396.000 430.800 ;
        RECT 4.400 429.400 1395.600 429.440 ;
        RECT 4.000 428.040 1395.600 429.400 ;
        RECT 4.000 422.640 1396.000 428.040 ;
        RECT 4.000 421.240 1395.600 422.640 ;
        RECT 4.000 420.600 1396.000 421.240 ;
        RECT 4.400 419.200 1396.000 420.600 ;
        RECT 4.000 415.840 1396.000 419.200 ;
        RECT 4.000 414.440 1395.600 415.840 ;
        RECT 4.000 409.720 1396.000 414.440 ;
        RECT 4.400 409.040 1396.000 409.720 ;
        RECT 4.400 408.320 1395.600 409.040 ;
        RECT 4.000 407.640 1395.600 408.320 ;
        RECT 4.000 402.240 1396.000 407.640 ;
        RECT 4.000 400.840 1395.600 402.240 ;
        RECT 4.000 399.520 1396.000 400.840 ;
        RECT 4.400 398.120 1396.000 399.520 ;
        RECT 4.000 395.440 1396.000 398.120 ;
        RECT 4.000 394.040 1395.600 395.440 ;
        RECT 4.000 389.320 1396.000 394.040 ;
        RECT 4.400 388.640 1396.000 389.320 ;
        RECT 4.400 387.920 1395.600 388.640 ;
        RECT 4.000 387.240 1395.600 387.920 ;
        RECT 4.000 381.840 1396.000 387.240 ;
        RECT 4.000 380.440 1395.600 381.840 ;
        RECT 4.000 379.120 1396.000 380.440 ;
        RECT 4.400 377.720 1396.000 379.120 ;
        RECT 4.000 375.040 1396.000 377.720 ;
        RECT 4.000 373.640 1395.600 375.040 ;
        RECT 4.000 368.240 1396.000 373.640 ;
        RECT 4.400 367.560 1396.000 368.240 ;
        RECT 4.400 366.840 1395.600 367.560 ;
        RECT 4.000 366.160 1395.600 366.840 ;
        RECT 4.000 360.760 1396.000 366.160 ;
        RECT 4.000 359.360 1395.600 360.760 ;
        RECT 4.000 358.040 1396.000 359.360 ;
        RECT 4.400 356.640 1396.000 358.040 ;
        RECT 4.000 353.960 1396.000 356.640 ;
        RECT 4.000 352.560 1395.600 353.960 ;
        RECT 4.000 347.840 1396.000 352.560 ;
        RECT 4.400 347.160 1396.000 347.840 ;
        RECT 4.400 346.440 1395.600 347.160 ;
        RECT 4.000 345.760 1395.600 346.440 ;
        RECT 4.000 340.360 1396.000 345.760 ;
        RECT 4.000 338.960 1395.600 340.360 ;
        RECT 4.000 337.640 1396.000 338.960 ;
        RECT 4.400 336.240 1396.000 337.640 ;
        RECT 4.000 333.560 1396.000 336.240 ;
        RECT 4.000 332.160 1395.600 333.560 ;
        RECT 4.000 326.760 1396.000 332.160 ;
        RECT 4.400 325.360 1395.600 326.760 ;
        RECT 4.000 319.960 1396.000 325.360 ;
        RECT 4.000 318.560 1395.600 319.960 ;
        RECT 4.000 316.560 1396.000 318.560 ;
        RECT 4.400 315.160 1396.000 316.560 ;
        RECT 4.000 313.160 1396.000 315.160 ;
        RECT 4.000 311.760 1395.600 313.160 ;
        RECT 4.000 306.360 1396.000 311.760 ;
        RECT 4.400 304.960 1395.600 306.360 ;
        RECT 4.000 299.560 1396.000 304.960 ;
        RECT 4.000 298.160 1395.600 299.560 ;
        RECT 4.000 296.160 1396.000 298.160 ;
        RECT 4.400 294.760 1396.000 296.160 ;
        RECT 4.000 292.080 1396.000 294.760 ;
        RECT 4.000 290.680 1395.600 292.080 ;
        RECT 4.000 285.280 1396.000 290.680 ;
        RECT 4.400 283.880 1395.600 285.280 ;
        RECT 4.000 278.480 1396.000 283.880 ;
        RECT 4.000 277.080 1395.600 278.480 ;
        RECT 4.000 275.080 1396.000 277.080 ;
        RECT 4.400 273.680 1396.000 275.080 ;
        RECT 4.000 271.680 1396.000 273.680 ;
        RECT 4.000 270.280 1395.600 271.680 ;
        RECT 4.000 264.880 1396.000 270.280 ;
        RECT 4.400 263.480 1395.600 264.880 ;
        RECT 4.000 258.080 1396.000 263.480 ;
        RECT 4.000 256.680 1395.600 258.080 ;
        RECT 4.000 254.680 1396.000 256.680 ;
        RECT 4.400 253.280 1396.000 254.680 ;
        RECT 4.000 251.280 1396.000 253.280 ;
        RECT 4.000 249.880 1395.600 251.280 ;
        RECT 4.000 244.480 1396.000 249.880 ;
        RECT 4.000 243.800 1395.600 244.480 ;
        RECT 4.400 243.080 1395.600 243.800 ;
        RECT 4.400 242.400 1396.000 243.080 ;
        RECT 4.000 237.680 1396.000 242.400 ;
        RECT 4.000 236.280 1395.600 237.680 ;
        RECT 4.000 233.600 1396.000 236.280 ;
        RECT 4.400 232.200 1396.000 233.600 ;
        RECT 4.000 230.880 1396.000 232.200 ;
        RECT 4.000 229.480 1395.600 230.880 ;
        RECT 4.000 223.400 1396.000 229.480 ;
        RECT 4.400 222.000 1395.600 223.400 ;
        RECT 4.000 216.600 1396.000 222.000 ;
        RECT 4.000 215.200 1395.600 216.600 ;
        RECT 4.000 213.200 1396.000 215.200 ;
        RECT 4.400 211.800 1396.000 213.200 ;
        RECT 4.000 209.800 1396.000 211.800 ;
        RECT 4.000 208.400 1395.600 209.800 ;
        RECT 4.000 203.000 1396.000 208.400 ;
        RECT 4.000 202.320 1395.600 203.000 ;
        RECT 4.400 201.600 1395.600 202.320 ;
        RECT 4.400 200.920 1396.000 201.600 ;
        RECT 4.000 196.200 1396.000 200.920 ;
        RECT 4.000 194.800 1395.600 196.200 ;
        RECT 4.000 192.120 1396.000 194.800 ;
        RECT 4.400 190.720 1396.000 192.120 ;
        RECT 4.000 189.400 1396.000 190.720 ;
        RECT 4.000 188.000 1395.600 189.400 ;
        RECT 4.000 182.600 1396.000 188.000 ;
        RECT 4.000 181.920 1395.600 182.600 ;
        RECT 4.400 181.200 1395.600 181.920 ;
        RECT 4.400 180.520 1396.000 181.200 ;
        RECT 4.000 175.800 1396.000 180.520 ;
        RECT 4.000 174.400 1395.600 175.800 ;
        RECT 4.000 171.720 1396.000 174.400 ;
        RECT 4.400 170.320 1396.000 171.720 ;
        RECT 4.000 169.000 1396.000 170.320 ;
        RECT 4.000 167.600 1395.600 169.000 ;
        RECT 4.000 162.200 1396.000 167.600 ;
        RECT 4.000 160.840 1395.600 162.200 ;
        RECT 4.400 160.800 1395.600 160.840 ;
        RECT 4.400 159.440 1396.000 160.800 ;
        RECT 4.000 155.400 1396.000 159.440 ;
        RECT 4.000 154.000 1395.600 155.400 ;
        RECT 4.000 150.640 1396.000 154.000 ;
        RECT 4.400 149.240 1396.000 150.640 ;
        RECT 4.000 147.920 1396.000 149.240 ;
        RECT 4.000 146.520 1395.600 147.920 ;
        RECT 4.000 141.120 1396.000 146.520 ;
        RECT 4.000 140.440 1395.600 141.120 ;
        RECT 4.400 139.720 1395.600 140.440 ;
        RECT 4.400 139.040 1396.000 139.720 ;
        RECT 4.000 134.320 1396.000 139.040 ;
        RECT 4.000 132.920 1395.600 134.320 ;
        RECT 4.000 130.240 1396.000 132.920 ;
        RECT 4.400 128.840 1396.000 130.240 ;
        RECT 4.000 127.520 1396.000 128.840 ;
        RECT 4.000 126.120 1395.600 127.520 ;
        RECT 4.000 120.720 1396.000 126.120 ;
        RECT 4.000 119.360 1395.600 120.720 ;
        RECT 4.400 119.320 1395.600 119.360 ;
        RECT 4.400 117.960 1396.000 119.320 ;
        RECT 4.000 113.920 1396.000 117.960 ;
        RECT 4.000 112.520 1395.600 113.920 ;
        RECT 4.000 109.160 1396.000 112.520 ;
        RECT 4.400 107.760 1396.000 109.160 ;
        RECT 4.000 107.120 1396.000 107.760 ;
        RECT 4.000 105.720 1395.600 107.120 ;
        RECT 4.000 100.320 1396.000 105.720 ;
        RECT 4.000 98.960 1395.600 100.320 ;
        RECT 4.400 98.920 1395.600 98.960 ;
        RECT 4.400 97.560 1396.000 98.920 ;
        RECT 4.000 93.520 1396.000 97.560 ;
        RECT 4.000 92.120 1395.600 93.520 ;
        RECT 4.000 88.760 1396.000 92.120 ;
        RECT 4.400 87.360 1396.000 88.760 ;
        RECT 4.000 86.720 1396.000 87.360 ;
        RECT 4.000 85.320 1395.600 86.720 ;
        RECT 4.000 79.920 1396.000 85.320 ;
        RECT 4.000 78.520 1395.600 79.920 ;
        RECT 4.000 77.880 1396.000 78.520 ;
        RECT 4.400 76.480 1396.000 77.880 ;
        RECT 4.000 72.440 1396.000 76.480 ;
        RECT 4.000 71.040 1395.600 72.440 ;
        RECT 4.000 67.680 1396.000 71.040 ;
        RECT 4.400 66.280 1396.000 67.680 ;
        RECT 4.000 65.640 1396.000 66.280 ;
        RECT 4.000 64.240 1395.600 65.640 ;
        RECT 4.000 58.840 1396.000 64.240 ;
        RECT 4.000 57.480 1395.600 58.840 ;
        RECT 4.400 57.440 1395.600 57.480 ;
        RECT 4.400 56.080 1396.000 57.440 ;
        RECT 4.000 52.040 1396.000 56.080 ;
        RECT 4.000 50.640 1395.600 52.040 ;
        RECT 4.000 47.280 1396.000 50.640 ;
        RECT 4.400 45.880 1396.000 47.280 ;
        RECT 4.000 45.240 1396.000 45.880 ;
        RECT 4.000 43.840 1395.600 45.240 ;
        RECT 4.000 38.440 1396.000 43.840 ;
        RECT 4.000 37.040 1395.600 38.440 ;
        RECT 4.000 36.400 1396.000 37.040 ;
        RECT 4.400 35.000 1396.000 36.400 ;
        RECT 4.000 31.640 1396.000 35.000 ;
        RECT 4.000 30.240 1395.600 31.640 ;
        RECT 4.000 26.200 1396.000 30.240 ;
        RECT 4.400 24.840 1396.000 26.200 ;
        RECT 4.400 24.800 1395.600 24.840 ;
        RECT 4.000 23.440 1395.600 24.800 ;
        RECT 4.000 18.040 1396.000 23.440 ;
        RECT 4.000 16.640 1395.600 18.040 ;
        RECT 4.000 16.000 1396.000 16.640 ;
        RECT 4.400 14.600 1396.000 16.000 ;
        RECT 4.000 11.240 1396.000 14.600 ;
        RECT 4.000 9.840 1395.600 11.240 ;
        RECT 4.000 5.800 1396.000 9.840 ;
        RECT 4.400 4.440 1396.000 5.800 ;
        RECT 4.400 4.400 1395.600 4.440 ;
        RECT 4.000 3.575 1395.600 4.400 ;
      LAYER met4 ;
        RECT 439.135 10.240 445.640 1380.225 ;
        RECT 448.040 10.240 470.640 1380.225 ;
        RECT 473.040 10.240 495.640 1380.225 ;
        RECT 498.040 10.240 520.640 1380.225 ;
        RECT 523.040 10.240 545.640 1380.225 ;
        RECT 548.040 10.240 570.640 1380.225 ;
        RECT 573.040 10.240 595.640 1380.225 ;
        RECT 598.040 10.240 620.640 1380.225 ;
        RECT 623.040 10.240 645.640 1380.225 ;
        RECT 648.040 10.240 670.640 1380.225 ;
        RECT 673.040 10.240 695.640 1380.225 ;
        RECT 698.040 10.240 720.640 1380.225 ;
        RECT 723.040 10.240 745.640 1380.225 ;
        RECT 748.040 10.240 770.640 1380.225 ;
        RECT 773.040 10.240 795.640 1380.225 ;
        RECT 798.040 10.240 820.640 1380.225 ;
        RECT 823.040 10.240 845.640 1380.225 ;
        RECT 848.040 10.240 870.640 1380.225 ;
        RECT 873.040 10.240 895.640 1380.225 ;
        RECT 898.040 10.240 920.640 1380.225 ;
        RECT 923.040 10.240 945.640 1380.225 ;
        RECT 948.040 10.240 970.640 1380.225 ;
        RECT 973.040 10.240 995.640 1380.225 ;
        RECT 998.040 10.240 1020.640 1380.225 ;
        RECT 1023.040 10.240 1045.640 1380.225 ;
        RECT 1048.040 10.240 1070.640 1380.225 ;
        RECT 1073.040 10.240 1095.640 1380.225 ;
        RECT 1098.040 10.240 1120.640 1380.225 ;
        RECT 1123.040 10.240 1145.640 1380.225 ;
        RECT 1148.040 10.240 1170.640 1380.225 ;
        RECT 1173.040 10.240 1195.640 1380.225 ;
        RECT 1198.040 10.240 1220.640 1380.225 ;
        RECT 1223.040 10.240 1245.640 1380.225 ;
        RECT 1248.040 10.240 1270.640 1380.225 ;
        RECT 1273.040 10.240 1295.640 1380.225 ;
        RECT 1298.040 10.240 1320.640 1380.225 ;
        RECT 1323.040 10.240 1323.585 1380.225 ;
        RECT 439.135 7.655 1323.585 10.240 ;
  END
END ibex_top
END LIBRARY

