magic
tech sky130A
magscale 1 2
timestamp 1640734220
<< locali >>
rect 26341 25891 26375 28713
rect 3801 23511 3835 23749
rect 26341 20043 26375 24497
rect 19073 18819 19107 18921
rect 9781 18071 9815 18241
rect 6193 17527 6227 17833
rect 15025 16099 15059 16201
rect 26341 15215 26375 15861
rect 3617 13311 3651 13413
rect 17233 12835 17267 12937
rect 21925 12631 21959 12733
rect 10609 11543 10643 11713
rect 12357 10455 12391 10761
rect 21649 10659 21683 10761
rect 15945 10455 15979 10625
rect 17233 9027 17267 9129
rect 12633 8347 12667 8517
rect 8493 5559 8527 5661
rect 18705 5151 18739 5253
<< viali >>
rect 26341 28713 26375 28747
rect 9781 26945 9815 26979
rect 14105 26945 14139 26979
rect 9965 26741 9999 26775
rect 14289 26741 14323 26775
rect 13645 26537 13679 26571
rect 6837 26469 6871 26503
rect 9505 26469 9539 26503
rect 11069 26469 11103 26503
rect 13553 26469 13587 26503
rect 10149 26401 10183 26435
rect 10885 26401 10919 26435
rect 14657 26401 14691 26435
rect 7021 26333 7055 26367
rect 7297 26333 7331 26367
rect 9413 26333 9447 26367
rect 10575 26333 10609 26367
rect 10977 26333 11011 26367
rect 14347 26333 14381 26367
rect 14749 26333 14783 26367
rect 15209 26333 15243 26367
rect 9321 26265 9355 26299
rect 9965 26265 9999 26299
rect 10333 26265 10367 26299
rect 13185 26265 13219 26299
rect 14105 26265 14139 26299
rect 14841 26265 14875 26299
rect 15025 26265 15059 26299
rect 7205 26197 7239 26231
rect 9873 26197 9907 26231
rect 2237 25993 2271 26027
rect 7757 25993 7791 26027
rect 9689 25993 9723 26027
rect 11253 25993 11287 26027
rect 10118 25925 10152 25959
rect 11529 25925 11563 25959
rect 11713 25925 11747 25959
rect 11897 25925 11931 25959
rect 14648 25925 14682 25959
rect 2053 25857 2087 25891
rect 4353 25857 4387 25891
rect 6633 25857 6667 25891
rect 8033 25857 8067 25891
rect 8309 25857 8343 25891
rect 8565 25857 8599 25891
rect 12817 25857 12851 25891
rect 13084 25857 13118 25891
rect 14381 25857 14415 25891
rect 16937 25857 16971 25891
rect 23949 25857 23983 25891
rect 24961 25857 24995 25891
rect 25237 25857 25271 25891
rect 26341 25857 26375 25891
rect 6377 25789 6411 25823
rect 9873 25789 9907 25823
rect 12173 25789 12207 25823
rect 16681 25789 16715 25823
rect 25513 25789 25547 25823
rect 8217 25721 8251 25755
rect 12541 25721 12575 25755
rect 12633 25653 12667 25687
rect 14197 25653 14231 25687
rect 15761 25653 15795 25687
rect 18061 25653 18095 25687
rect 7205 25449 7239 25483
rect 8309 25449 8343 25483
rect 9413 25449 9447 25483
rect 10701 25449 10735 25483
rect 11345 25449 11379 25483
rect 13093 25449 13127 25483
rect 13185 25449 13219 25483
rect 14105 25449 14139 25483
rect 16681 25449 16715 25483
rect 5641 25381 5675 25415
rect 8493 25381 8527 25415
rect 9229 25381 9263 25415
rect 5825 25313 5859 25347
rect 7849 25313 7883 25347
rect 8769 25313 8803 25347
rect 8953 25313 8987 25347
rect 10241 25313 10275 25347
rect 13829 25313 13863 25347
rect 14749 25313 14783 25347
rect 14933 25313 14967 25347
rect 15025 25313 15059 25347
rect 19349 25313 19383 25347
rect 5457 25245 5491 25279
rect 5641 25245 5675 25279
rect 7481 25245 7515 25279
rect 7665 25245 7699 25279
rect 7757 25245 7791 25279
rect 7941 25245 7975 25279
rect 8125 25245 8159 25279
rect 10609 25245 10643 25279
rect 11345 25245 11379 25279
rect 11437 25245 11471 25279
rect 12909 25245 12943 25279
rect 13645 25245 13679 25279
rect 15392 25245 15426 25279
rect 16221 25245 16255 25279
rect 16497 25245 16531 25279
rect 17015 25245 17049 25279
rect 17325 25245 17359 25279
rect 17417 25245 17451 25279
rect 17694 25245 17728 25279
rect 18061 25245 18095 25279
rect 18153 25245 18187 25279
rect 6092 25177 6126 25211
rect 10057 25177 10091 25211
rect 14473 25177 14507 25211
rect 15669 25177 15703 25211
rect 16773 25177 16807 25211
rect 19616 25177 19650 25211
rect 9597 25109 9631 25143
rect 9965 25109 9999 25143
rect 10425 25109 10459 25143
rect 11713 25109 11747 25143
rect 13553 25109 13587 25143
rect 14565 25109 14599 25143
rect 15485 25109 15519 25143
rect 16405 25109 16439 25143
rect 17601 25109 17635 25143
rect 20729 25109 20763 25143
rect 6469 24905 6503 24939
rect 7941 24905 7975 24939
rect 8953 24905 8987 24939
rect 11253 24905 11287 24939
rect 15485 24905 15519 24939
rect 16037 24905 16071 24939
rect 18061 24905 18095 24939
rect 19717 24905 19751 24939
rect 7205 24837 7239 24871
rect 9321 24837 9355 24871
rect 10140 24837 10174 24871
rect 12449 24837 12483 24871
rect 18613 24837 18647 24871
rect 20729 24837 20763 24871
rect 6193 24769 6227 24803
rect 6653 24769 6687 24803
rect 6745 24769 6779 24803
rect 6837 24769 6871 24803
rect 6929 24769 6963 24803
rect 7113 24769 7147 24803
rect 7297 24769 7331 24803
rect 7573 24769 7607 24803
rect 7849 24769 7883 24803
rect 8861 24769 8895 24803
rect 11529 24769 11563 24803
rect 11771 24769 11805 24803
rect 12081 24769 12115 24803
rect 12173 24769 12207 24803
rect 12265 24769 12299 24803
rect 13829 24769 13863 24803
rect 14013 24769 14047 24803
rect 14197 24769 14231 24803
rect 14473 24769 14507 24803
rect 14749 24769 14783 24803
rect 15117 24769 15151 24803
rect 15209 24769 15243 24803
rect 16681 24769 16715 24803
rect 16937 24769 16971 24803
rect 18245 24769 18279 24803
rect 18429 24769 18463 24803
rect 19533 24769 19567 24803
rect 20051 24769 20085 24803
rect 20361 24769 20395 24803
rect 20545 24769 20579 24803
rect 20913 24769 20947 24803
rect 7389 24701 7423 24735
rect 9413 24701 9447 24735
rect 9505 24701 9539 24735
rect 9873 24701 9907 24735
rect 14565 24701 14599 24735
rect 16497 24701 16531 24735
rect 18889 24701 18923 24735
rect 20453 24701 20487 24735
rect 12633 24633 12667 24667
rect 14933 24633 14967 24667
rect 16221 24633 16255 24667
rect 19257 24633 19291 24667
rect 19349 24633 19383 24667
rect 5825 24565 5859 24599
rect 6101 24565 6135 24599
rect 8125 24565 8159 24599
rect 14381 24565 14415 24599
rect 14749 24565 14783 24599
rect 15209 24565 15243 24599
rect 19901 24565 19935 24599
rect 26341 24497 26375 24531
rect 7481 24361 7515 24395
rect 9689 24361 9723 24395
rect 11529 24361 11563 24395
rect 13645 24361 13679 24395
rect 16957 24361 16991 24395
rect 18337 24361 18371 24395
rect 6837 24293 6871 24327
rect 7757 24293 7791 24327
rect 9505 24293 9539 24327
rect 12633 24293 12667 24327
rect 17785 24293 17819 24327
rect 18889 24293 18923 24327
rect 21005 24293 21039 24327
rect 6653 24225 6687 24259
rect 10149 24225 10183 24259
rect 12357 24225 12391 24259
rect 15485 24225 15519 24259
rect 16313 24225 16347 24259
rect 16405 24225 16439 24259
rect 17417 24225 17451 24259
rect 17509 24225 17543 24259
rect 19625 24225 19659 24259
rect 21189 24225 21223 24259
rect 21281 24225 21315 24259
rect 23305 24225 23339 24259
rect 3801 24157 3835 24191
rect 5825 24157 5859 24191
rect 6009 24157 6043 24191
rect 6101 24157 6135 24191
rect 6469 24157 6503 24191
rect 6929 24157 6963 24191
rect 7297 24157 7331 24191
rect 7481 24157 7515 24191
rect 7573 24157 7607 24191
rect 9873 24157 9907 24191
rect 11898 24157 11932 24191
rect 12265 24157 12299 24191
rect 13737 24157 13771 24191
rect 14105 24157 14139 24191
rect 14197 24157 14231 24191
rect 14564 24157 14598 24191
rect 15026 24157 15060 24191
rect 15393 24157 15427 24191
rect 17325 24157 17359 24191
rect 17969 24157 18003 24191
rect 18153 24157 18187 24191
rect 19349 24157 19383 24191
rect 21648 24157 21682 24191
rect 22903 24157 22937 24191
rect 23213 24157 23247 24191
rect 4068 24089 4102 24123
rect 9229 24089 9263 24123
rect 10394 24089 10428 24123
rect 13001 24089 13035 24123
rect 13921 24089 13955 24123
rect 14841 24089 14875 24123
rect 18521 24089 18555 24123
rect 19870 24089 19904 24123
rect 22661 24089 22695 24123
rect 5181 24021 5215 24055
rect 5641 24021 5675 24055
rect 7113 24021 7147 24055
rect 10057 24021 10091 24055
rect 11805 24021 11839 24055
rect 12541 24021 12575 24055
rect 14657 24021 14691 24055
rect 16497 24021 16531 24055
rect 16865 24021 16899 24055
rect 18981 24021 19015 24055
rect 19533 24021 19567 24055
rect 21741 24021 21775 24055
rect 1593 23817 1627 23851
rect 4353 23817 4387 23851
rect 6469 23817 6503 23851
rect 9781 23817 9815 23851
rect 10425 23817 10459 23851
rect 12357 23817 12391 23851
rect 13829 23817 13863 23851
rect 15393 23817 15427 23851
rect 16773 23817 16807 23851
rect 17417 23817 17451 23851
rect 18429 23817 18463 23851
rect 19717 23817 19751 23851
rect 20085 23817 20119 23851
rect 20545 23817 20579 23851
rect 22017 23817 22051 23851
rect 23489 23817 23523 23851
rect 2728 23749 2762 23783
rect 3801 23749 3835 23783
rect 3985 23749 4019 23783
rect 10793 23749 10827 23783
rect 17233 23749 17267 23783
rect 20913 23749 20947 23783
rect 21097 23749 21131 23783
rect 21281 23749 21315 23783
rect 22354 23749 22388 23783
rect 23857 23749 23891 23783
rect 24041 23749 24075 23783
rect 2973 23613 3007 23647
rect 4169 23681 4203 23715
rect 4445 23681 4479 23715
rect 4721 23681 4755 23715
rect 4988 23681 5022 23715
rect 6837 23681 6871 23715
rect 6929 23681 6963 23715
rect 7205 23681 7239 23715
rect 7481 23681 7515 23715
rect 8125 23681 8159 23715
rect 8309 23681 8343 23715
rect 10333 23681 10367 23715
rect 11897 23681 11931 23715
rect 12173 23681 12207 23715
rect 12449 23681 12483 23715
rect 12705 23681 12739 23715
rect 14013 23681 14047 23715
rect 14269 23681 14303 23715
rect 18337 23681 18371 23715
rect 18797 23681 18831 23715
rect 19625 23681 19659 23715
rect 20453 23681 20487 23715
rect 21833 23681 21867 23715
rect 23673 23681 23707 23715
rect 6653 23613 6687 23647
rect 7297 23613 7331 23647
rect 9321 23613 9355 23647
rect 10609 23613 10643 23647
rect 19901 23613 19935 23647
rect 20637 23613 20671 23647
rect 22109 23613 22143 23647
rect 6101 23545 6135 23579
rect 7665 23545 7699 23579
rect 9689 23545 9723 23579
rect 9965 23545 9999 23579
rect 12081 23545 12115 23579
rect 16865 23545 16899 23579
rect 18613 23545 18647 23579
rect 19257 23545 19291 23579
rect 3801 23477 3835 23511
rect 7481 23477 7515 23511
rect 7941 23477 7975 23511
rect 8125 23477 8159 23511
rect 19165 23477 19199 23511
rect 7389 23273 7423 23307
rect 8125 23273 8159 23307
rect 9781 23273 9815 23307
rect 12633 23273 12667 23307
rect 13921 23273 13955 23307
rect 15025 23273 15059 23307
rect 21925 23273 21959 23307
rect 4169 23205 4203 23239
rect 8401 23205 8435 23239
rect 19993 23205 20027 23239
rect 21833 23205 21867 23239
rect 22109 23205 22143 23239
rect 4261 23137 4295 23171
rect 4629 23137 4663 23171
rect 5273 23137 5307 23171
rect 6009 23137 6043 23171
rect 8217 23137 8251 23171
rect 13277 23137 13311 23171
rect 13553 23137 13587 23171
rect 14749 23137 14783 23171
rect 21465 23137 21499 23171
rect 22569 23137 22603 23171
rect 22661 23137 22695 23171
rect 23673 23137 23707 23171
rect 25145 23137 25179 23171
rect 4077 23069 4111 23103
rect 4721 23069 4755 23103
rect 5641 23069 5675 23103
rect 5733 23069 5767 23103
rect 7665 23069 7699 23103
rect 7849 23069 7883 23103
rect 7941 23069 7975 23103
rect 8309 23069 8343 23103
rect 9965 23069 9999 23103
rect 13737 23069 13771 23103
rect 14473 23069 14507 23103
rect 19809 23069 19843 23103
rect 20177 23069 20211 23103
rect 21373 23069 21407 23103
rect 23271 23069 23305 23103
rect 23581 23069 23615 23103
rect 4445 23001 4479 23035
rect 5917 23001 5951 23035
rect 6254 23001 6288 23035
rect 9045 23001 9079 23035
rect 9229 23001 9263 23035
rect 13093 23001 13127 23035
rect 16405 23001 16439 23035
rect 16589 23001 16623 23035
rect 23029 23001 23063 23035
rect 4721 22933 4755 22967
rect 13001 22933 13035 22967
rect 14105 22933 14139 22967
rect 14565 22933 14599 22967
rect 16681 22933 16715 22967
rect 22477 22933 22511 22967
rect 5549 22729 5583 22763
rect 9229 22729 9263 22763
rect 9321 22729 9355 22763
rect 10149 22729 10183 22763
rect 13829 22729 13863 22763
rect 22293 22729 22327 22763
rect 22661 22729 22695 22763
rect 24133 22729 24167 22763
rect 5641 22661 5675 22695
rect 7021 22661 7055 22695
rect 8033 22661 8067 22695
rect 9045 22661 9079 22695
rect 9597 22661 9631 22695
rect 13369 22661 13403 22695
rect 14105 22661 14139 22695
rect 14289 22661 14323 22695
rect 17141 22661 17175 22695
rect 17509 22661 17543 22695
rect 17693 22661 17727 22695
rect 21833 22661 21867 22695
rect 22998 22661 23032 22695
rect 3341 22593 3375 22627
rect 3608 22593 3642 22627
rect 6837 22593 6871 22627
rect 7481 22593 7515 22627
rect 7573 22593 7607 22627
rect 8309 22593 8343 22627
rect 8677 22593 8711 22627
rect 8769 22593 8803 22627
rect 9413 22593 9447 22627
rect 9873 22593 9907 22627
rect 10057 22593 10091 22627
rect 10333 22593 10367 22627
rect 16957 22593 16991 22627
rect 17233 22593 17267 22627
rect 18521 22593 18555 22627
rect 22477 22593 22511 22627
rect 22753 22593 22787 22627
rect 8401 22525 8435 22559
rect 16221 22525 16255 22559
rect 7205 22457 7239 22491
rect 8309 22457 8343 22491
rect 9781 22457 9815 22491
rect 13737 22457 13771 22491
rect 15945 22457 15979 22491
rect 17325 22457 17359 22491
rect 22201 22457 22235 22491
rect 4721 22389 4755 22423
rect 6101 22389 6135 22423
rect 7297 22389 7331 22423
rect 7757 22389 7791 22423
rect 8861 22389 8895 22423
rect 15761 22389 15795 22423
rect 16773 22389 16807 22423
rect 18337 22389 18371 22423
rect 4353 22185 4387 22219
rect 11253 22185 11287 22219
rect 17141 22185 17175 22219
rect 22293 22185 22327 22219
rect 23489 22185 23523 22219
rect 6929 22049 6963 22083
rect 8769 22049 8803 22083
rect 9505 22049 9539 22083
rect 12357 22049 12391 22083
rect 15761 22049 15795 22083
rect 22201 22049 22235 22083
rect 22845 22049 22879 22083
rect 1961 21981 1995 22015
rect 3801 21981 3835 22015
rect 4174 21981 4208 22015
rect 8953 21981 8987 22015
rect 9045 21981 9079 22015
rect 9229 21981 9263 22015
rect 11069 21981 11103 22015
rect 11713 21981 11747 22015
rect 11805 21981 11839 22015
rect 11989 21981 12023 22015
rect 12541 21981 12575 22015
rect 12633 21981 12667 22015
rect 15485 21981 15519 22015
rect 17325 21981 17359 22015
rect 17601 21981 17635 22015
rect 19257 21981 19291 22015
rect 22753 21981 22787 22015
rect 23581 21981 23615 22015
rect 23765 21981 23799 22015
rect 2228 21913 2262 21947
rect 3985 21913 4019 21947
rect 4077 21913 4111 21947
rect 7113 21913 7147 21947
rect 8502 21913 8536 21947
rect 9772 21913 9806 21947
rect 12265 21913 12299 21947
rect 16006 21913 16040 21947
rect 17868 21913 17902 21947
rect 19502 21913 19536 21947
rect 3341 21845 3375 21879
rect 7389 21845 7423 21879
rect 9413 21845 9447 21879
rect 10885 21845 10919 21879
rect 12725 21845 12759 21879
rect 15669 21845 15703 21879
rect 17509 21845 17543 21879
rect 18981 21845 19015 21879
rect 20637 21845 20671 21879
rect 22661 21845 22695 21879
rect 2697 21641 2731 21675
rect 3709 21641 3743 21675
rect 8585 21641 8619 21675
rect 9505 21641 9539 21675
rect 10425 21641 10459 21675
rect 11621 21641 11655 21675
rect 16681 21641 16715 21675
rect 17141 21641 17175 21675
rect 17969 21641 18003 21675
rect 18613 21641 18647 21675
rect 20821 21641 20855 21675
rect 4077 21573 4111 21607
rect 9781 21573 9815 21607
rect 12734 21573 12768 21607
rect 17509 21573 17543 21607
rect 2881 21505 2915 21539
rect 2973 21505 3007 21539
rect 3249 21505 3283 21539
rect 3525 21505 3559 21539
rect 8769 21505 8803 21539
rect 8861 21505 8895 21539
rect 9045 21505 9079 21539
rect 9689 21505 9723 21539
rect 10241 21505 10275 21539
rect 13001 21505 13035 21539
rect 15292 21505 15326 21539
rect 17049 21505 17083 21539
rect 18521 21505 18555 21539
rect 19441 21505 19475 21539
rect 19718 21505 19752 21539
rect 20264 21505 20298 21539
rect 20671 21505 20705 21539
rect 21465 21505 21499 21539
rect 21649 21505 21683 21539
rect 22018 21505 22052 21539
rect 22385 21505 22419 21539
rect 22569 21505 22603 21539
rect 23087 21505 23121 21539
rect 23489 21505 23523 21539
rect 4169 21437 4203 21471
rect 4261 21437 4295 21471
rect 9965 21437 9999 21471
rect 15025 21437 15059 21471
rect 17325 21437 17359 21471
rect 18705 21437 18739 21471
rect 19349 21437 19383 21471
rect 20085 21437 20119 21471
rect 20177 21437 20211 21471
rect 20380 21437 20414 21471
rect 21281 21437 21315 21471
rect 22477 21437 22511 21471
rect 23397 21437 23431 21471
rect 4721 21369 4755 21403
rect 4905 21369 4939 21403
rect 9229 21369 9263 21403
rect 10057 21369 10091 21403
rect 17877 21369 17911 21403
rect 18153 21369 18187 21403
rect 19073 21369 19107 21403
rect 21833 21369 21867 21403
rect 3157 21301 3191 21335
rect 3341 21301 3375 21335
rect 7389 21301 7423 21335
rect 8953 21301 8987 21335
rect 16405 21301 16439 21335
rect 19349 21301 19383 21335
rect 19625 21301 19659 21335
rect 22753 21301 22787 21335
rect 22937 21301 22971 21335
rect 3801 21097 3835 21131
rect 4997 21097 5031 21131
rect 9873 21097 9907 21131
rect 10057 21097 10091 21131
rect 17509 21097 17543 21131
rect 17969 21097 18003 21131
rect 19257 21097 19291 21131
rect 20545 21097 20579 21131
rect 23949 21097 23983 21131
rect 18613 21029 18647 21063
rect 18705 21029 18739 21063
rect 19073 21029 19107 21063
rect 20453 21029 20487 21063
rect 1501 20961 1535 20995
rect 3341 20961 3375 20995
rect 4445 20961 4479 20995
rect 7941 20961 7975 20995
rect 8309 20961 8343 20995
rect 8677 20961 8711 20995
rect 11989 20961 12023 20995
rect 18245 20961 18279 20995
rect 19717 20961 19751 20995
rect 19809 20961 19843 20995
rect 3433 20893 3467 20927
rect 4629 20893 4663 20927
rect 6377 20893 6411 20927
rect 8033 20893 8067 20927
rect 8585 20893 8619 20927
rect 9965 20893 9999 20927
rect 11621 20893 11655 20927
rect 11804 20893 11838 20927
rect 11897 20893 11931 20927
rect 12173 20893 12207 20927
rect 12449 20893 12483 20927
rect 14473 20893 14507 20927
rect 18889 20893 18923 20927
rect 22201 20893 22235 20927
rect 22477 20893 22511 20927
rect 22569 20893 22603 20927
rect 22836 20893 22870 20927
rect 1768 20825 1802 20859
rect 4169 20825 4203 20859
rect 4261 20825 4295 20859
rect 6110 20825 6144 20859
rect 7674 20825 7708 20859
rect 12357 20825 12391 20859
rect 12716 20825 12750 20859
rect 14740 20825 14774 20859
rect 20085 20825 20119 20859
rect 21956 20825 21990 20859
rect 2881 20757 2915 20791
rect 4813 20757 4847 20791
rect 6561 20757 6595 20791
rect 9689 20757 9723 20791
rect 13829 20757 13863 20791
rect 15853 20757 15887 20791
rect 19625 20757 19659 20791
rect 20821 20757 20855 20791
rect 22293 20757 22327 20791
rect 2513 20553 2547 20587
rect 3157 20553 3191 20587
rect 4169 20553 4203 20587
rect 4353 20553 4387 20587
rect 4721 20553 4755 20587
rect 7389 20553 7423 20587
rect 9137 20553 9171 20587
rect 9597 20553 9631 20587
rect 10609 20553 10643 20587
rect 13645 20553 13679 20587
rect 14473 20553 14507 20587
rect 15301 20553 15335 20587
rect 16129 20553 16163 20587
rect 19073 20553 19107 20587
rect 20729 20553 20763 20587
rect 20913 20553 20947 20587
rect 21373 20553 21407 20587
rect 22569 20553 22603 20587
rect 6193 20485 6227 20519
rect 7297 20485 7331 20519
rect 19717 20485 19751 20519
rect 19901 20485 19935 20519
rect 23213 20485 23247 20519
rect 23397 20485 23431 20519
rect 23581 20485 23615 20519
rect 2697 20417 2731 20451
rect 2789 20417 2823 20451
rect 3065 20417 3099 20451
rect 3525 20417 3559 20451
rect 3985 20417 4019 20451
rect 4813 20417 4847 20451
rect 5182 20417 5216 20451
rect 5365 20417 5399 20451
rect 5457 20417 5491 20451
rect 5640 20417 5674 20451
rect 6009 20417 6043 20451
rect 6561 20417 6595 20451
rect 6837 20417 6871 20451
rect 6930 20417 6964 20451
rect 7113 20417 7147 20451
rect 8585 20417 8619 20451
rect 9045 20417 9079 20451
rect 10057 20417 10091 20451
rect 10149 20417 10183 20451
rect 12265 20417 12299 20451
rect 12532 20417 12566 20451
rect 13829 20417 13863 20451
rect 13994 20417 14028 20451
rect 14105 20417 14139 20451
rect 14381 20417 14415 20451
rect 14657 20417 14691 20451
rect 14840 20417 14874 20451
rect 15209 20417 15243 20451
rect 15485 20417 15519 20451
rect 15650 20417 15684 20451
rect 15853 20417 15887 20451
rect 16037 20417 16071 20451
rect 20085 20417 20119 20451
rect 21281 20417 21315 20451
rect 22477 20417 22511 20451
rect 3617 20349 3651 20383
rect 3801 20349 3835 20383
rect 4537 20349 4571 20383
rect 4997 20349 5031 20383
rect 5089 20349 5123 20383
rect 5733 20349 5767 20383
rect 5825 20349 5859 20383
rect 6745 20349 6779 20383
rect 8493 20349 8527 20383
rect 9229 20349 9263 20383
rect 9781 20349 9815 20383
rect 14197 20349 14231 20383
rect 14933 20349 14967 20383
rect 15025 20349 15059 20383
rect 15761 20349 15795 20383
rect 21465 20349 21499 20383
rect 21925 20349 21959 20383
rect 22753 20349 22787 20383
rect 2973 20281 3007 20315
rect 8217 20281 8251 20315
rect 8677 20281 8711 20315
rect 9873 20281 9907 20315
rect 6469 20213 6503 20247
rect 8585 20213 8619 20247
rect 10333 20213 10367 20247
rect 22109 20213 22143 20247
rect 5457 20009 5491 20043
rect 9413 20009 9447 20043
rect 9689 20009 9723 20043
rect 10701 20009 10735 20043
rect 13185 20009 13219 20043
rect 22385 20009 22419 20043
rect 25329 20009 25363 20043
rect 26341 20009 26375 20043
rect 3157 19941 3191 19975
rect 7757 19941 7791 19975
rect 8953 19941 8987 19975
rect 22109 19941 22143 19975
rect 3801 19873 3835 19907
rect 3893 19873 3927 19907
rect 6837 19873 6871 19907
rect 7941 19873 7975 19907
rect 10057 19873 10091 19907
rect 14933 19873 14967 19907
rect 15025 19873 15059 19907
rect 15485 19873 15519 19907
rect 17601 19873 17635 19907
rect 21741 19873 21775 19907
rect 22937 19873 22971 19907
rect 1777 19805 1811 19839
rect 3525 19805 3559 19839
rect 4077 19805 4111 19839
rect 4169 19805 4203 19839
rect 6570 19805 6604 19839
rect 7573 19805 7607 19839
rect 8125 19805 8159 19839
rect 8309 19805 8343 19839
rect 8401 19805 8435 19839
rect 9137 19805 9171 19839
rect 9781 19805 9815 19839
rect 10333 19805 10367 19839
rect 11805 19805 11839 19839
rect 14657 19805 14691 19839
rect 14822 19805 14856 19839
rect 15209 19805 15243 19839
rect 25145 19805 25179 19839
rect 2044 19737 2078 19771
rect 9321 19737 9355 19771
rect 12072 19737 12106 19771
rect 15393 19737 15427 19771
rect 15730 19737 15764 19771
rect 17509 19737 17543 19771
rect 18337 19737 18371 19771
rect 3341 19669 3375 19703
rect 4353 19669 4387 19703
rect 7481 19669 7515 19703
rect 8585 19669 8619 19703
rect 10241 19669 10275 19703
rect 16865 19669 16899 19703
rect 17049 19669 17083 19703
rect 17417 19669 17451 19703
rect 18061 19669 18095 19703
rect 18429 19669 18463 19703
rect 22201 19669 22235 19703
rect 22753 19669 22787 19703
rect 22845 19669 22879 19703
rect 25053 19669 25087 19703
rect 4353 19465 4387 19499
rect 4537 19465 4571 19499
rect 6101 19465 6135 19499
rect 7481 19465 7515 19499
rect 10517 19465 10551 19499
rect 12173 19465 12207 19499
rect 12633 19465 12667 19499
rect 15577 19465 15611 19499
rect 17509 19465 17543 19499
rect 20361 19465 20395 19499
rect 22293 19465 22327 19499
rect 22569 19465 22603 19499
rect 3893 19397 3927 19431
rect 8493 19397 8527 19431
rect 9045 19397 9079 19431
rect 9382 19397 9416 19431
rect 19226 19397 19260 19431
rect 23029 19397 23063 19431
rect 2973 19329 3007 19363
rect 3065 19329 3099 19363
rect 3985 19329 4019 19363
rect 4988 19329 5022 19363
rect 6377 19329 6411 19363
rect 6561 19329 6595 19363
rect 6745 19329 6779 19363
rect 6930 19329 6964 19363
rect 7113 19329 7147 19363
rect 7389 19353 7423 19387
rect 7665 19329 7699 19363
rect 8309 19329 8343 19363
rect 8677 19329 8711 19363
rect 8861 19329 8895 19363
rect 10701 19329 10735 19363
rect 11529 19329 11563 19363
rect 11712 19329 11746 19363
rect 11805 19329 11839 19363
rect 12081 19329 12115 19363
rect 12357 19329 12391 19363
rect 12817 19329 12851 19363
rect 13369 19329 13403 19363
rect 14013 19329 14047 19363
rect 14196 19329 14230 19363
rect 14565 19329 14599 19363
rect 16865 19329 16899 19363
rect 18622 19329 18656 19363
rect 22937 19329 22971 19363
rect 3341 19261 3375 19295
rect 3525 19261 3559 19295
rect 3801 19261 3835 19295
rect 4721 19261 4755 19295
rect 6837 19261 6871 19295
rect 8125 19261 8159 19295
rect 9137 19261 9171 19295
rect 11897 19261 11931 19295
rect 14289 19261 14323 19295
rect 14381 19261 14415 19295
rect 18889 19261 18923 19295
rect 18981 19261 19015 19295
rect 22385 19261 22419 19295
rect 23121 19261 23155 19295
rect 3249 19193 3283 19227
rect 7205 19193 7239 19227
rect 13553 19193 13587 19227
rect 2789 19125 2823 19159
rect 7941 19125 7975 19159
rect 10793 19125 10827 19159
rect 12541 19125 12575 19159
rect 14657 19125 14691 19159
rect 3525 18921 3559 18955
rect 6193 18921 6227 18955
rect 7665 18921 7699 18955
rect 9137 18921 9171 18955
rect 10241 18921 10275 18955
rect 11713 18921 11747 18955
rect 15669 18921 15703 18955
rect 15945 18921 15979 18955
rect 17233 18921 17267 18955
rect 18061 18921 18095 18955
rect 19073 18921 19107 18955
rect 20637 18921 20671 18955
rect 21281 18921 21315 18955
rect 8033 18853 8067 18887
rect 21097 18853 21131 18887
rect 6929 18785 6963 18819
rect 8769 18785 8803 18819
rect 9873 18785 9907 18819
rect 10701 18785 10735 18819
rect 10793 18785 10827 18819
rect 11161 18785 11195 18819
rect 12725 18785 12759 18819
rect 12817 18785 12851 18819
rect 16589 18785 16623 18819
rect 17693 18785 17727 18819
rect 17785 18785 17819 18819
rect 18613 18785 18647 18819
rect 19073 18785 19107 18819
rect 2145 18717 2179 18751
rect 6377 18717 6411 18751
rect 6653 18717 6687 18751
rect 6745 18717 6779 18751
rect 7481 18717 7515 18751
rect 7849 18717 7883 18751
rect 8401 18717 8435 18751
rect 8585 18717 8619 18751
rect 8953 18717 8987 18751
rect 9229 18717 9263 18751
rect 9413 18717 9447 18751
rect 9505 18717 9539 18751
rect 9631 18711 9665 18745
rect 10425 18717 10459 18751
rect 10517 18717 10551 18751
rect 11253 18717 11287 18751
rect 12541 18717 12575 18751
rect 12910 18717 12944 18751
rect 13093 18717 13127 18751
rect 15577 18717 15611 18751
rect 15853 18717 15887 18751
rect 16129 18717 16163 18751
rect 16865 18717 16899 18751
rect 17417 18717 17451 18751
rect 17600 18717 17634 18751
rect 17969 18717 18003 18751
rect 18245 18717 18279 18751
rect 18410 18711 18444 18745
rect 18521 18717 18555 18751
rect 18797 18717 18831 18751
rect 19257 18717 19291 18751
rect 22661 18717 22695 18751
rect 24225 18717 24259 18751
rect 2412 18649 2446 18683
rect 8309 18649 8343 18683
rect 15310 18649 15344 18683
rect 19513 18649 19547 18683
rect 20913 18649 20947 18683
rect 22394 18649 22428 18683
rect 23958 18649 23992 18683
rect 7389 18581 7423 18615
rect 9965 18581 9999 18615
rect 11345 18581 11379 18615
rect 12449 18581 12483 18615
rect 14197 18581 14231 18615
rect 16313 18581 16347 18615
rect 16773 18581 16807 18615
rect 18889 18581 18923 18615
rect 22845 18581 22879 18615
rect 3249 18377 3283 18411
rect 3525 18377 3559 18411
rect 8677 18377 8711 18411
rect 9597 18377 9631 18411
rect 12081 18377 12115 18411
rect 13553 18377 13587 18411
rect 15577 18377 15611 18411
rect 19809 18377 19843 18411
rect 21189 18377 21223 18411
rect 2136 18309 2170 18343
rect 4997 18309 5031 18343
rect 5181 18309 5215 18343
rect 9229 18309 9263 18343
rect 12440 18309 12474 18343
rect 23121 18309 23155 18343
rect 1869 18241 1903 18275
rect 3709 18241 3743 18275
rect 3801 18241 3835 18275
rect 4077 18241 4111 18275
rect 6561 18241 6595 18275
rect 7021 18241 7055 18275
rect 8861 18241 8895 18275
rect 9689 18241 9723 18275
rect 9781 18241 9815 18275
rect 9965 18241 9999 18275
rect 10241 18241 10275 18275
rect 10333 18241 10367 18275
rect 11713 18241 11747 18275
rect 11897 18241 11931 18275
rect 14453 18241 14487 18275
rect 17509 18241 17543 18275
rect 17674 18244 17708 18278
rect 17792 18241 17826 18275
rect 18061 18241 18095 18275
rect 18337 18241 18371 18275
rect 18797 18241 18831 18275
rect 20177 18241 20211 18275
rect 20269 18241 20303 18275
rect 21373 18241 21407 18275
rect 21465 18241 21499 18275
rect 21557 18241 21591 18275
rect 22017 18241 22051 18275
rect 22385 18241 22419 18275
rect 22568 18241 22602 18275
rect 22661 18241 22695 18275
rect 22937 18241 22971 18275
rect 9413 18105 9447 18139
rect 12173 18173 12207 18207
rect 14197 18173 14231 18207
rect 17877 18173 17911 18207
rect 19717 18173 19751 18207
rect 20453 18173 20487 18207
rect 22753 18173 22787 18207
rect 10149 18105 10183 18139
rect 18245 18105 18279 18139
rect 18521 18105 18555 18139
rect 18613 18105 18647 18139
rect 21833 18105 21867 18139
rect 23213 18105 23247 18139
rect 3985 18037 4019 18071
rect 6745 18037 6779 18071
rect 6837 18037 6871 18071
rect 7665 18037 7699 18071
rect 9045 18037 9079 18071
rect 9781 18037 9815 18071
rect 10425 18037 10459 18071
rect 4629 17833 4663 17867
rect 4813 17833 4847 17867
rect 6193 17833 6227 17867
rect 9965 17833 9999 17867
rect 10333 17833 10367 17867
rect 15485 17833 15519 17867
rect 20177 17833 20211 17867
rect 22017 17833 22051 17867
rect 3801 17765 3835 17799
rect 3341 17697 3375 17731
rect 4445 17697 4479 17731
rect 3065 17629 3099 17663
rect 3157 17629 3191 17663
rect 3433 17629 3467 17663
rect 4261 17561 4295 17595
rect 13001 17765 13035 17799
rect 17693 17765 17727 17799
rect 21281 17765 21315 17799
rect 8217 17697 8251 17731
rect 9873 17697 9907 17731
rect 11621 17697 11655 17731
rect 13553 17697 13587 17731
rect 14105 17697 14139 17731
rect 20085 17697 20119 17731
rect 20729 17697 20763 17731
rect 21649 17697 21683 17731
rect 21741 17697 21775 17731
rect 24409 17697 24443 17731
rect 9321 17629 9355 17663
rect 9781 17629 9815 17663
rect 10609 17629 10643 17663
rect 13185 17629 13219 17663
rect 13333 17626 13367 17660
rect 13461 17629 13495 17663
rect 13737 17629 13771 17663
rect 17049 17629 17083 17663
rect 17233 17629 17267 17663
rect 19073 17629 19107 17663
rect 21097 17629 21131 17663
rect 21373 17629 21407 17663
rect 21521 17623 21555 17657
rect 21925 17629 21959 17663
rect 22201 17629 22235 17663
rect 22477 17629 22511 17663
rect 22625 17626 22659 17660
rect 22753 17629 22787 17663
rect 22845 17629 22879 17663
rect 23029 17629 23063 17663
rect 7950 17561 7984 17595
rect 9137 17561 9171 17595
rect 9505 17561 9539 17595
rect 11866 17561 11900 17595
rect 13921 17561 13955 17595
rect 14350 17561 14384 17595
rect 18806 17561 18840 17595
rect 23213 17561 23247 17595
rect 24654 17561 24688 17595
rect 2881 17493 2915 17527
rect 4169 17493 4203 17527
rect 6193 17493 6227 17527
rect 6285 17493 6319 17527
rect 6837 17493 6871 17527
rect 9597 17493 9631 17527
rect 10149 17493 10183 17527
rect 10793 17493 10827 17527
rect 20545 17493 20579 17527
rect 20637 17493 20671 17527
rect 22385 17493 22419 17527
rect 25789 17493 25823 17527
rect 3801 17289 3835 17323
rect 5549 17289 5583 17323
rect 11253 17289 11287 17323
rect 17325 17289 17359 17323
rect 18337 17289 18371 17323
rect 20545 17289 20579 17323
rect 21189 17289 21223 17323
rect 21833 17289 21867 17323
rect 22661 17289 22695 17323
rect 2136 17221 2170 17255
rect 4261 17221 4295 17255
rect 7582 17221 7616 17255
rect 7941 17221 7975 17255
rect 14197 17221 14231 17255
rect 17509 17221 17543 17255
rect 22201 17221 22235 17255
rect 23121 17221 23155 17255
rect 1869 17153 1903 17187
rect 4169 17153 4203 17187
rect 4629 17153 4663 17187
rect 4905 17153 4939 17187
rect 4997 17153 5031 17187
rect 5641 17153 5675 17187
rect 5825 17153 5859 17187
rect 6010 17153 6044 17187
rect 6193 17153 6227 17187
rect 7849 17153 7883 17187
rect 8125 17153 8159 17187
rect 8511 17153 8545 17187
rect 8677 17153 8711 17187
rect 8861 17153 8895 17187
rect 9026 17153 9060 17187
rect 9229 17153 9263 17187
rect 9413 17153 9447 17187
rect 9689 17153 9723 17187
rect 9872 17153 9906 17187
rect 10241 17153 10275 17187
rect 11069 17153 11103 17187
rect 13461 17153 13495 17187
rect 13609 17156 13643 17190
rect 13737 17153 13771 17187
rect 14013 17153 14047 17187
rect 17693 17179 17727 17213
rect 17876 17153 17910 17187
rect 18061 17153 18095 17187
rect 18245 17153 18279 17187
rect 18705 17153 18739 17187
rect 20729 17153 20763 17187
rect 23029 17153 23063 17187
rect 4353 17085 4387 17119
rect 4721 17085 4755 17119
rect 5917 17085 5951 17119
rect 8309 17085 8343 17119
rect 8401 17085 8435 17119
rect 9137 17085 9171 17119
rect 9965 17085 9999 17119
rect 10057 17085 10091 17119
rect 13829 17085 13863 17119
rect 17969 17085 18003 17119
rect 22293 17085 22327 17119
rect 22477 17085 22511 17119
rect 23213 17085 23247 17119
rect 6469 17017 6503 17051
rect 9597 17017 9631 17051
rect 18521 17017 18555 17051
rect 21649 17017 21683 17051
rect 3249 16949 3283 16983
rect 5181 16949 5215 16983
rect 10333 16949 10367 16983
rect 13001 16949 13035 16983
rect 13277 16949 13311 16983
rect 3525 16745 3559 16779
rect 6193 16745 6227 16779
rect 8401 16745 8435 16779
rect 8769 16745 8803 16779
rect 9045 16745 9079 16779
rect 12633 16745 12667 16779
rect 13553 16745 13587 16779
rect 20913 16745 20947 16779
rect 22477 16745 22511 16779
rect 4629 16677 4663 16711
rect 15761 16677 15795 16711
rect 16589 16677 16623 16711
rect 2145 16609 2179 16643
rect 4261 16609 4295 16643
rect 4445 16609 4479 16643
rect 4813 16609 4847 16643
rect 7849 16609 7883 16643
rect 9413 16609 9447 16643
rect 13277 16609 13311 16643
rect 16129 16609 16163 16643
rect 16957 16609 16991 16643
rect 17785 16609 17819 16643
rect 17877 16609 17911 16643
rect 18245 16609 18279 16643
rect 18981 16609 19015 16643
rect 19257 16609 19291 16643
rect 21097 16609 21131 16643
rect 23121 16609 23155 16643
rect 23213 16609 23247 16643
rect 4169 16541 4203 16575
rect 8217 16541 8251 16575
rect 9321 16541 9355 16575
rect 10977 16541 11011 16575
rect 15577 16541 15611 16575
rect 15853 16541 15887 16575
rect 16018 16541 16052 16575
rect 16221 16541 16255 16575
rect 16405 16541 16439 16575
rect 16681 16541 16715 16575
rect 16864 16541 16898 16575
rect 17049 16541 17083 16575
rect 17233 16541 17267 16575
rect 17509 16541 17543 16575
rect 17692 16541 17726 16575
rect 18061 16541 18095 16575
rect 19513 16541 19547 16575
rect 22845 16541 22879 16575
rect 23028 16541 23062 16575
rect 23397 16541 23431 16575
rect 2412 16473 2446 16507
rect 5080 16473 5114 16507
rect 7582 16473 7616 16507
rect 9658 16473 9692 16507
rect 23581 16473 23615 16507
rect 3801 16405 3835 16439
rect 6469 16405 6503 16439
rect 9137 16405 9171 16439
rect 10793 16405 10827 16439
rect 11069 16405 11103 16439
rect 12725 16405 12759 16439
rect 13093 16405 13127 16439
rect 13185 16405 13219 16439
rect 15485 16405 15519 16439
rect 17325 16405 17359 16439
rect 18337 16405 18371 16439
rect 18705 16405 18739 16439
rect 18797 16405 18831 16439
rect 20637 16405 20671 16439
rect 21281 16405 21315 16439
rect 21373 16405 21407 16439
rect 21741 16405 21775 16439
rect 3249 16201 3283 16235
rect 3893 16201 3927 16235
rect 4261 16201 4295 16235
rect 6469 16201 6503 16235
rect 7297 16201 7331 16235
rect 11529 16201 11563 16235
rect 12449 16201 12483 16235
rect 13093 16201 13127 16235
rect 13553 16201 13587 16235
rect 14381 16201 14415 16235
rect 15025 16201 15059 16235
rect 16313 16201 16347 16235
rect 18061 16201 18095 16235
rect 18429 16201 18463 16235
rect 18889 16201 18923 16235
rect 19533 16201 19567 16235
rect 21005 16201 21039 16235
rect 3801 16133 3835 16167
rect 10048 16133 10082 16167
rect 16926 16133 16960 16167
rect 20821 16133 20855 16167
rect 24308 16133 24342 16167
rect 1869 16065 1903 16099
rect 2136 16065 2170 16099
rect 4353 16065 4387 16099
rect 6561 16065 6595 16099
rect 6837 16065 6871 16099
rect 6930 16065 6964 16099
rect 7113 16065 7147 16099
rect 7389 16065 7423 16099
rect 7665 16065 7699 16099
rect 7775 16065 7809 16099
rect 7941 16065 7975 16099
rect 8309 16065 8343 16099
rect 8953 16065 8987 16099
rect 9136 16065 9170 16099
rect 9321 16065 9355 16099
rect 9505 16065 9539 16099
rect 9781 16065 9815 16099
rect 11713 16065 11747 16099
rect 12633 16065 12667 16099
rect 13001 16065 13035 16099
rect 13921 16065 13955 16099
rect 14565 16065 14599 16099
rect 15025 16065 15059 16099
rect 15301 16065 15335 16099
rect 15466 16065 15500 16099
rect 15577 16065 15611 16099
rect 15853 16065 15887 16099
rect 16129 16065 16163 16099
rect 16681 16065 16715 16099
rect 18797 16065 18831 16099
rect 19717 16065 19751 16099
rect 19901 16065 19935 16099
rect 19993 16065 20027 16099
rect 20177 16065 20211 16099
rect 20453 16065 20487 16099
rect 21373 16065 21407 16099
rect 22376 16065 22410 16099
rect 24041 16065 24075 16099
rect 3709 15997 3743 16031
rect 6745 15997 6779 16031
rect 7573 15997 7607 16031
rect 9229 15997 9263 16031
rect 9689 15997 9723 16031
rect 12357 15997 12391 16031
rect 12817 15997 12851 16031
rect 14013 15997 14047 16031
rect 14105 15997 14139 16031
rect 15669 15997 15703 16031
rect 18981 15997 19015 16031
rect 20361 15997 20395 16031
rect 21281 15997 21315 16031
rect 22109 15997 22143 16031
rect 13461 15929 13495 15963
rect 20453 15929 20487 15963
rect 8033 15861 8067 15895
rect 11161 15861 11195 15895
rect 15209 15861 15243 15895
rect 15945 15861 15979 15895
rect 18245 15861 18279 15895
rect 21281 15861 21315 15895
rect 23489 15861 23523 15895
rect 25421 15861 25455 15895
rect 26341 15861 26375 15895
rect 2881 15657 2915 15691
rect 3341 15657 3375 15691
rect 7757 15657 7791 15691
rect 11345 15657 11379 15691
rect 13461 15657 13495 15691
rect 14749 15657 14783 15691
rect 16957 15657 16991 15691
rect 18521 15657 18555 15691
rect 20453 15657 20487 15691
rect 22017 15657 22051 15691
rect 22845 15657 22879 15691
rect 7665 15589 7699 15623
rect 12357 15589 12391 15623
rect 22293 15589 22327 15623
rect 22753 15589 22787 15623
rect 3433 15521 3467 15555
rect 7113 15521 7147 15555
rect 9965 15521 9999 15555
rect 12817 15521 12851 15555
rect 14841 15521 14875 15555
rect 20637 15521 20671 15555
rect 21189 15521 21223 15555
rect 23397 15521 23431 15555
rect 3065 15453 3099 15487
rect 3157 15453 3191 15487
rect 10221 15453 10255 15487
rect 12633 15453 12667 15487
rect 13737 15453 13771 15487
rect 14565 15453 14599 15487
rect 15577 15453 15611 15487
rect 17141 15453 17175 15487
rect 17397 15453 17431 15487
rect 18889 15453 18923 15487
rect 19257 15453 19291 15487
rect 20545 15453 20579 15487
rect 21005 15453 21039 15487
rect 21373 15453 21407 15487
rect 21556 15453 21590 15487
rect 21649 15453 21683 15487
rect 21741 15453 21775 15487
rect 21925 15453 21959 15487
rect 7297 15385 7331 15419
rect 15844 15385 15878 15419
rect 18705 15385 18739 15419
rect 19073 15385 19107 15419
rect 7205 15317 7239 15351
rect 9873 15317 9907 15351
rect 12449 15317 12483 15351
rect 13001 15317 13035 15351
rect 13093 15317 13127 15351
rect 13553 15317 13587 15351
rect 19441 15317 19475 15351
rect 21005 15317 21039 15351
rect 23213 15317 23247 15351
rect 23305 15317 23339 15351
rect 26341 15181 26375 15215
rect 7297 15113 7331 15147
rect 7665 15113 7699 15147
rect 12725 15113 12759 15147
rect 18153 15113 18187 15147
rect 18981 15113 19015 15147
rect 23305 15113 23339 15147
rect 23673 15113 23707 15147
rect 8125 15045 8159 15079
rect 21649 15045 21683 15079
rect 22170 15045 22204 15079
rect 4261 14977 4295 15011
rect 4630 14977 4664 15011
rect 4813 14977 4847 15011
rect 5089 14977 5123 15011
rect 6653 14977 6687 15011
rect 7039 14977 7073 15011
rect 7205 14977 7239 15011
rect 9689 14977 9723 15011
rect 9854 14977 9888 15011
rect 10057 14977 10091 15011
rect 10241 14977 10275 15011
rect 10701 14977 10735 15011
rect 12173 14977 12207 15011
rect 12632 14977 12666 15011
rect 12909 14977 12943 15011
rect 15117 14977 15151 15011
rect 16773 14977 16807 15011
rect 17049 14977 17083 15011
rect 18303 14977 18337 15011
rect 18613 14977 18647 15011
rect 18797 14977 18831 15011
rect 20913 14977 20947 15011
rect 21078 14977 21112 15011
rect 21189 14977 21223 15011
rect 21465 14977 21499 15011
rect 21925 14977 21959 15011
rect 23489 14977 23523 15011
rect 4445 14909 4479 14943
rect 4537 14909 4571 14943
rect 6469 14909 6503 14943
rect 6837 14909 6871 14943
rect 6929 14909 6963 14943
rect 7757 14909 7791 14943
rect 7941 14909 7975 14943
rect 9965 14909 9999 14943
rect 12265 14909 12299 14943
rect 14657 14909 14691 14943
rect 15209 14909 15243 14943
rect 15301 14909 15335 14943
rect 18705 14909 18739 14943
rect 21281 14909 21315 14943
rect 16957 14841 16991 14875
rect 4169 14773 4203 14807
rect 4905 14773 4939 14807
rect 9505 14773 9539 14807
rect 10333 14773 10367 14807
rect 10517 14773 10551 14807
rect 12081 14773 12115 14807
rect 14749 14773 14783 14807
rect 17233 14773 17267 14807
rect 20729 14773 20763 14807
rect 5181 14569 5215 14603
rect 7389 14569 7423 14603
rect 12265 14569 12299 14603
rect 12909 14569 12943 14603
rect 13093 14569 13127 14603
rect 14841 14569 14875 14603
rect 5457 14501 5491 14535
rect 13921 14501 13955 14535
rect 20637 14501 20671 14535
rect 13277 14433 13311 14467
rect 14197 14433 14231 14467
rect 14381 14433 14415 14467
rect 3801 14365 3835 14399
rect 4068 14365 4102 14399
rect 6570 14365 6604 14399
rect 6837 14365 6871 14399
rect 8769 14365 8803 14399
rect 10425 14365 10459 14399
rect 10681 14365 10715 14399
rect 12173 14365 12207 14399
rect 12449 14365 12483 14399
rect 12817 14365 12851 14399
rect 13369 14365 13403 14399
rect 13679 14365 13713 14399
rect 14473 14365 14507 14399
rect 20453 14365 20487 14399
rect 22201 14365 22235 14399
rect 22569 14365 22603 14399
rect 22753 14365 22787 14399
rect 23397 14365 23431 14399
rect 23489 14365 23523 14399
rect 8502 14297 8536 14331
rect 12633 14297 12667 14331
rect 22293 14297 22327 14331
rect 22845 14297 22879 14331
rect 23029 14297 23063 14331
rect 23213 14297 23247 14331
rect 11805 14229 11839 14263
rect 11989 14229 12023 14263
rect 19993 14229 20027 14263
rect 2881 14025 2915 14059
rect 4813 14025 4847 14059
rect 8401 14025 8435 14059
rect 9505 14025 9539 14059
rect 13185 14025 13219 14059
rect 16129 14025 16163 14059
rect 17233 14025 17267 14059
rect 19073 14025 19107 14059
rect 19625 14025 19659 14059
rect 19993 14025 20027 14059
rect 20821 14025 20855 14059
rect 22293 14025 22327 14059
rect 8309 13957 8343 13991
rect 8769 13957 8803 13991
rect 13461 13957 13495 13991
rect 14657 13957 14691 13991
rect 14841 13957 14875 13991
rect 17785 13957 17819 13991
rect 18889 13957 18923 13991
rect 23121 13957 23155 13991
rect 1768 13889 1802 13923
rect 3433 13889 3467 13923
rect 3700 13889 3734 13923
rect 6929 13889 6963 13923
rect 7113 13889 7147 13923
rect 7205 13889 7239 13923
rect 7333 13892 7367 13926
rect 7481 13889 7515 13923
rect 7573 13889 7607 13923
rect 7756 13889 7790 13923
rect 7941 13889 7975 13923
rect 8125 13889 8159 13923
rect 9413 13889 9447 13923
rect 11713 13889 11747 13923
rect 12725 13889 12759 13923
rect 13369 13889 13403 13923
rect 13645 13889 13679 13923
rect 13829 13889 13863 13923
rect 14163 13889 14197 13923
rect 14473 13889 14507 13923
rect 14565 13889 14599 13923
rect 20453 13889 20487 13923
rect 21833 13889 21867 13923
rect 22017 13889 22051 13923
rect 22109 13889 22143 13923
rect 23029 13889 23063 13923
rect 1501 13821 1535 13855
rect 6745 13821 6779 13855
rect 7849 13821 7883 13855
rect 8861 13821 8895 13855
rect 8953 13821 8987 13855
rect 13921 13821 13955 13855
rect 15025 13821 15059 13855
rect 19441 13821 19475 13855
rect 19533 13821 19567 13855
rect 20177 13821 20211 13855
rect 20361 13821 20395 13855
rect 22569 13821 22603 13855
rect 23213 13821 23247 13855
rect 17049 13753 17083 13787
rect 9229 13685 9263 13719
rect 11529 13685 11563 13719
rect 12909 13685 12943 13719
rect 21557 13685 21591 13719
rect 21833 13685 21867 13719
rect 22661 13685 22695 13719
rect 5181 13481 5215 13515
rect 10793 13481 10827 13515
rect 13553 13481 13587 13515
rect 14197 13481 14231 13515
rect 14565 13481 14599 13515
rect 16313 13481 16347 13515
rect 17969 13481 18003 13515
rect 19349 13481 19383 13515
rect 20177 13481 20211 13515
rect 21005 13481 21039 13515
rect 23397 13481 23431 13515
rect 2881 13413 2915 13447
rect 3617 13413 3651 13447
rect 9321 13413 9355 13447
rect 14289 13413 14323 13447
rect 18889 13413 18923 13447
rect 3801 13345 3835 13379
rect 7941 13345 7975 13379
rect 8493 13345 8527 13379
rect 9413 13345 9447 13379
rect 11989 13345 12023 13379
rect 12081 13345 12115 13379
rect 12541 13345 12575 13379
rect 15117 13345 15151 13379
rect 15669 13345 15703 13379
rect 15761 13345 15795 13379
rect 16865 13345 16899 13379
rect 17417 13345 17451 13379
rect 17509 13345 17543 13379
rect 18429 13345 18463 13379
rect 18521 13345 18555 13379
rect 19901 13345 19935 13379
rect 20729 13345 20763 13379
rect 1501 13277 1535 13311
rect 3341 13277 3375 13311
rect 3525 13277 3559 13311
rect 3617 13277 3651 13311
rect 8217 13277 8251 13311
rect 8401 13277 8435 13311
rect 8586 13277 8620 13311
rect 8769 13277 8803 13311
rect 9137 13277 9171 13311
rect 11713 13277 11747 13311
rect 11896 13277 11930 13311
rect 12265 13277 12299 13311
rect 13369 13277 13403 13311
rect 14473 13277 14507 13311
rect 15393 13277 15427 13311
rect 15541 13277 15575 13311
rect 15945 13277 15979 13311
rect 17141 13277 17175 13311
rect 17324 13277 17358 13311
rect 17693 13277 17727 13311
rect 19073 13277 19107 13311
rect 20545 13277 20579 13311
rect 21189 13277 21223 13311
rect 21372 13277 21406 13311
rect 21462 13277 21496 13311
rect 21557 13277 21591 13311
rect 21741 13277 21775 13311
rect 22017 13277 22051 13311
rect 23581 13277 23615 13311
rect 23765 13277 23799 13311
rect 1768 13209 1802 13243
rect 4046 13209 4080 13243
rect 7674 13209 7708 13243
rect 9680 13209 9714 13243
rect 12449 13209 12483 13243
rect 16773 13209 16807 13243
rect 17877 13209 17911 13243
rect 19717 13209 19751 13243
rect 21925 13209 21959 13243
rect 22262 13209 22296 13243
rect 3157 13141 3191 13175
rect 6561 13141 6595 13175
rect 8125 13141 8159 13175
rect 9045 13141 9079 13175
rect 11437 13141 11471 13175
rect 14933 13141 14967 13175
rect 15025 13141 15059 13175
rect 16037 13141 16071 13175
rect 16681 13141 16715 13175
rect 18337 13141 18371 13175
rect 19809 13141 19843 13175
rect 20637 13141 20671 13175
rect 23673 13141 23707 13175
rect 2145 12937 2179 12971
rect 3433 12937 3467 12971
rect 6469 12937 6503 12971
rect 7941 12937 7975 12971
rect 8769 12937 8803 12971
rect 9597 12937 9631 12971
rect 15117 12937 15151 12971
rect 17233 12937 17267 12971
rect 17693 12937 17727 12971
rect 18061 12937 18095 12971
rect 19533 12937 19567 12971
rect 22937 12937 22971 12971
rect 4445 12869 4479 12903
rect 7604 12869 7638 12903
rect 8309 12869 8343 12903
rect 13430 12869 13464 12903
rect 16230 12869 16264 12903
rect 24010 12869 24044 12903
rect 2329 12801 2363 12835
rect 2421 12801 2455 12835
rect 2789 12801 2823 12835
rect 2972 12801 3006 12835
rect 3341 12801 3375 12835
rect 3614 12801 3648 12835
rect 3800 12801 3834 12835
rect 3893 12801 3927 12835
rect 4169 12801 4203 12835
rect 4629 12801 4663 12835
rect 4998 12801 5032 12835
rect 5181 12801 5215 12835
rect 5457 12801 5491 12835
rect 5825 12801 5859 12835
rect 7849 12801 7883 12835
rect 8953 12801 8987 12835
rect 9136 12801 9170 12835
rect 9505 12801 9539 12835
rect 9781 12801 9815 12835
rect 9964 12801 9998 12835
rect 10057 12801 10091 12835
rect 10333 12801 10367 12835
rect 10609 12801 10643 12835
rect 10792 12801 10826 12835
rect 10885 12801 10919 12835
rect 11161 12801 11195 12835
rect 11621 12801 11655 12835
rect 11877 12801 11911 12835
rect 13185 12801 13219 12835
rect 16497 12801 16531 12835
rect 16681 12801 16715 12835
rect 17233 12801 17267 12835
rect 18153 12801 18187 12835
rect 18409 12801 18443 12835
rect 19959 12801 19993 12835
rect 20453 12801 20487 12835
rect 20637 12801 20671 12835
rect 20821 12801 20855 12835
rect 21281 12801 21315 12835
rect 21649 12801 21683 12835
rect 22201 12801 22235 12835
rect 22293 12801 22327 12835
rect 22476 12801 22510 12835
rect 22569 12801 22603 12835
rect 22845 12801 22879 12835
rect 23142 12801 23176 12835
rect 23489 12801 23523 12835
rect 23673 12801 23707 12835
rect 23765 12801 23799 12835
rect 2697 12733 2731 12767
rect 3065 12733 3099 12767
rect 3157 12733 3191 12767
rect 3985 12733 4019 12767
rect 4813 12733 4847 12767
rect 4905 12733 4939 12767
rect 8401 12733 8435 12767
rect 8585 12733 8619 12767
rect 9229 12733 9263 12767
rect 9321 12733 9355 12767
rect 10149 12733 10183 12767
rect 10977 12733 11011 12767
rect 16773 12733 16807 12767
rect 17417 12733 17451 12767
rect 17601 12733 17635 12767
rect 20269 12733 20303 12767
rect 20361 12733 20395 12767
rect 21465 12733 21499 12767
rect 21925 12733 21959 12767
rect 22661 12733 22695 12767
rect 5273 12665 5307 12699
rect 5641 12665 5675 12699
rect 10517 12665 10551 12699
rect 14565 12665 14599 12699
rect 19717 12665 19751 12699
rect 21557 12665 21591 12699
rect 23213 12665 23247 12699
rect 2605 12597 2639 12631
rect 4261 12597 4295 12631
rect 11253 12597 11287 12631
rect 13001 12597 13035 12631
rect 16681 12597 16715 12631
rect 17049 12597 17083 12631
rect 21925 12597 21959 12631
rect 22017 12597 22051 12631
rect 25145 12597 25179 12631
rect 2329 12393 2363 12427
rect 2789 12393 2823 12427
rect 3341 12393 3375 12427
rect 5273 12393 5307 12427
rect 5457 12393 5491 12427
rect 6561 12393 6595 12427
rect 7941 12393 7975 12427
rect 8217 12393 8251 12427
rect 8493 12393 8527 12427
rect 8677 12393 8711 12427
rect 9505 12393 9539 12427
rect 14933 12393 14967 12427
rect 16957 12393 16991 12427
rect 18613 12393 18647 12427
rect 21281 12393 21315 12427
rect 21649 12393 21683 12427
rect 22385 12393 22419 12427
rect 6193 12325 6227 12359
rect 21925 12325 21959 12359
rect 22477 12325 22511 12359
rect 2973 12257 3007 12291
rect 10149 12257 10183 12291
rect 10425 12257 10459 12291
rect 11253 12257 11287 12291
rect 14841 12257 14875 12291
rect 15485 12257 15519 12291
rect 16405 12257 16439 12291
rect 20545 12257 20579 12291
rect 21005 12257 21039 12291
rect 22937 12257 22971 12291
rect 23029 12257 23063 12291
rect 2513 12189 2547 12223
rect 2605 12189 2639 12223
rect 2881 12189 2915 12223
rect 3157 12189 3191 12223
rect 3893 12189 3927 12223
rect 4160 12189 4194 12223
rect 5641 12189 5675 12223
rect 6377 12189 6411 12223
rect 8401 12189 8435 12223
rect 8953 12189 8987 12223
rect 9413 12189 9447 12223
rect 9873 12189 9907 12223
rect 10885 12189 10919 12223
rect 11050 12189 11084 12223
rect 11161 12189 11195 12223
rect 11437 12189 11471 12223
rect 11713 12189 11747 12223
rect 15301 12189 15335 12223
rect 15393 12189 15427 12223
rect 15945 12189 15979 12223
rect 16037 12189 16071 12223
rect 16497 12189 16531 12223
rect 17141 12189 17175 12223
rect 17325 12189 17359 12223
rect 17601 12189 17635 12223
rect 17693 12189 17727 12223
rect 18060 12189 18094 12223
rect 19533 12189 19567 12223
rect 19993 12189 20027 12223
rect 20177 12189 20211 12223
rect 20637 12189 20671 12223
rect 20821 12189 20855 12223
rect 21281 12189 21315 12223
rect 21465 12189 21499 12223
rect 22017 12189 22051 12223
rect 22845 12189 22879 12223
rect 5917 12121 5951 12155
rect 6101 12121 6135 12155
rect 7849 12121 7883 12155
rect 11621 12121 11655 12155
rect 11958 12121 11992 12155
rect 17049 12121 17083 12155
rect 18337 12121 18371 12155
rect 18521 12121 18555 12155
rect 9137 12053 9171 12087
rect 9229 12053 9263 12087
rect 9965 12053 9999 12087
rect 10701 12053 10735 12087
rect 13093 12053 13127 12087
rect 15853 12053 15887 12087
rect 16589 12053 16623 12087
rect 18153 12053 18187 12087
rect 19349 12053 19383 12087
rect 20453 12053 20487 12087
rect 2881 11849 2915 11883
rect 5181 11849 5215 11883
rect 7205 11849 7239 11883
rect 9413 11849 9447 11883
rect 10425 11849 10459 11883
rect 13369 11849 13403 11883
rect 16405 11849 16439 11883
rect 17693 11849 17727 11883
rect 20453 11849 20487 11883
rect 22937 11849 22971 11883
rect 10057 11781 10091 11815
rect 10241 11781 10275 11815
rect 13553 11781 13587 11815
rect 1768 11713 1802 11747
rect 3801 11713 3835 11747
rect 4068 11713 4102 11747
rect 5365 11713 5399 11747
rect 5457 11713 5491 11747
rect 5825 11713 5859 11747
rect 6837 11713 6871 11747
rect 6929 11713 6963 11747
rect 9505 11713 9539 11747
rect 10609 11713 10643 11747
rect 10885 11713 10919 11747
rect 11989 11713 12023 11747
rect 12256 11713 12290 11747
rect 13737 11713 13771 11747
rect 14933 11713 14967 11747
rect 15117 11713 15151 11747
rect 15485 11713 15519 11747
rect 15945 11713 15979 11747
rect 16313 11713 16347 11747
rect 16865 11713 16899 11747
rect 17233 11713 17267 11747
rect 17601 11713 17635 11747
rect 18061 11713 18095 11747
rect 20361 11713 20395 11747
rect 20637 11713 20671 11747
rect 23029 11713 23063 11747
rect 1501 11645 1535 11679
rect 7113 11645 7147 11679
rect 9689 11645 9723 11679
rect 15853 11645 15887 11679
rect 17417 11645 17451 11679
rect 15393 11577 15427 11611
rect 16957 11577 16991 11611
rect 17877 11577 17911 11611
rect 5641 11509 5675 11543
rect 9045 11509 9079 11543
rect 9873 11509 9907 11543
rect 10241 11509 10275 11543
rect 10609 11509 10643 11543
rect 10701 11509 10735 11543
rect 16221 11509 16255 11543
rect 20269 11509 20303 11543
rect 2421 11305 2455 11339
rect 4537 11305 4571 11339
rect 7481 11305 7515 11339
rect 15301 11305 15335 11339
rect 21465 11305 21499 11339
rect 15025 11237 15059 11271
rect 15945 11237 15979 11271
rect 17325 11237 17359 11271
rect 21005 11237 21039 11271
rect 2881 11169 2915 11203
rect 2973 11169 3007 11203
rect 4169 11169 4203 11203
rect 5641 11169 5675 11203
rect 9229 11169 9263 11203
rect 10149 11169 10183 11203
rect 10793 11169 10827 11203
rect 15669 11169 15703 11203
rect 20729 11169 20763 11203
rect 23029 11169 23063 11203
rect 23305 11169 23339 11203
rect 2605 11101 2639 11135
rect 2697 11101 2731 11135
rect 3893 11101 3927 11135
rect 4076 11101 4110 11135
rect 4261 11101 4295 11135
rect 4445 11101 4479 11135
rect 5273 11101 5307 11135
rect 5456 11101 5490 11135
rect 5549 11101 5583 11135
rect 5825 11101 5859 11135
rect 6101 11101 6135 11135
rect 7849 11101 7883 11135
rect 9505 11101 9539 11135
rect 15393 11101 15427 11135
rect 15577 11101 15611 11135
rect 16037 11101 16071 11135
rect 16681 11101 16715 11135
rect 16773 11101 16807 11135
rect 16957 11101 16991 11135
rect 17233 11101 17267 11135
rect 19717 11101 19751 11135
rect 19901 11101 19935 11135
rect 20269 11101 20303 11135
rect 20453 11101 20487 11135
rect 21373 11101 21407 11135
rect 22845 11101 22879 11135
rect 6346 11033 6380 11067
rect 10241 11033 10275 11067
rect 10333 11033 10367 11067
rect 17141 11033 17175 11067
rect 20085 11033 20119 11067
rect 22293 11033 22327 11067
rect 22937 11033 22971 11067
rect 5917 10965 5951 10999
rect 7665 10965 7699 10999
rect 9413 10965 9447 10999
rect 9873 10965 9907 10999
rect 10701 10965 10735 10999
rect 20545 10965 20579 10999
rect 21649 10965 21683 10999
rect 22477 10965 22511 10999
rect 2881 10761 2915 10795
rect 7757 10761 7791 10795
rect 9321 10761 9355 10795
rect 12265 10761 12299 10795
rect 12357 10761 12391 10795
rect 13829 10761 13863 10795
rect 17141 10761 17175 10795
rect 19349 10761 19383 10795
rect 20545 10761 20579 10795
rect 21649 10761 21683 10795
rect 22201 10761 22235 10795
rect 6193 10693 6227 10727
rect 3065 10625 3099 10659
rect 4629 10625 4663 10659
rect 4812 10625 4846 10659
rect 4905 10625 4939 10659
rect 4997 10625 5031 10659
rect 5181 10625 5215 10659
rect 5457 10625 5491 10659
rect 5605 10625 5639 10659
rect 5825 10625 5859 10659
rect 6009 10625 6043 10659
rect 6377 10625 6411 10659
rect 6633 10625 6667 10659
rect 7941 10625 7975 10659
rect 8197 10625 8231 10659
rect 9505 10625 9539 10659
rect 9688 10625 9722 10659
rect 10057 10625 10091 10659
rect 10333 10625 10367 10659
rect 10516 10625 10550 10659
rect 10609 10625 10643 10659
rect 10885 10625 10919 10659
rect 12081 10625 12115 10659
rect 3249 10557 3283 10591
rect 5733 10557 5767 10591
rect 9781 10557 9815 10591
rect 9873 10557 9907 10591
rect 10701 10557 10735 10591
rect 12716 10625 12750 10659
rect 15301 10625 15335 10659
rect 15577 10625 15611 10659
rect 15945 10625 15979 10659
rect 16497 10625 16531 10659
rect 17049 10625 17083 10659
rect 17509 10625 17543 10659
rect 17693 10625 17727 10659
rect 18061 10625 18095 10659
rect 18797 10625 18831 10659
rect 19441 10625 19475 10659
rect 20637 10625 20671 10659
rect 21189 10625 21223 10659
rect 21373 10625 21407 10659
rect 21649 10625 21683 10659
rect 23029 10625 23063 10659
rect 23121 10625 23155 10659
rect 23489 10625 23523 10659
rect 23581 10625 23615 10659
rect 23765 10625 23799 10659
rect 12449 10557 12483 10591
rect 15577 10489 15611 10523
rect 17233 10557 17267 10591
rect 19165 10557 19199 10591
rect 20361 10557 20395 10591
rect 21557 10557 21591 10591
rect 22293 10557 22327 10591
rect 22385 10557 22419 10591
rect 23305 10557 23339 10591
rect 18613 10489 18647 10523
rect 21005 10489 21039 10523
rect 23949 10489 23983 10523
rect 5273 10421 5307 10455
rect 10149 10421 10183 10455
rect 10977 10421 11011 10455
rect 12357 10421 12391 10455
rect 15209 10421 15243 10455
rect 15761 10421 15795 10455
rect 15945 10421 15979 10455
rect 16129 10421 16163 10455
rect 16313 10421 16347 10455
rect 16681 10421 16715 10455
rect 17877 10421 17911 10455
rect 18981 10421 19015 10455
rect 19809 10421 19843 10455
rect 19993 10421 20027 10455
rect 20085 10421 20119 10455
rect 21833 10421 21867 10455
rect 22661 10421 22695 10455
rect 2881 10217 2915 10251
rect 7205 10217 7239 10251
rect 12265 10217 12299 10251
rect 12633 10217 12667 10251
rect 17049 10217 17083 10251
rect 19349 10217 19383 10251
rect 3985 10149 4019 10183
rect 9045 10149 9079 10183
rect 21557 10149 21591 10183
rect 1501 10081 1535 10115
rect 3525 10081 3559 10115
rect 8493 10081 8527 10115
rect 14657 10081 14691 10115
rect 15485 10081 15519 10115
rect 15669 10081 15703 10115
rect 16313 10081 16347 10115
rect 17509 10081 17543 10115
rect 17693 10081 17727 10115
rect 18429 10081 18463 10115
rect 18981 10081 19015 10115
rect 19993 10081 20027 10115
rect 20177 10081 20211 10115
rect 21189 10081 21223 10115
rect 21281 10081 21315 10115
rect 22017 10081 22051 10115
rect 22201 10081 22235 10115
rect 23305 10081 23339 10115
rect 23581 10081 23615 10115
rect 3341 10013 3375 10047
rect 3801 10013 3835 10047
rect 5733 10013 5767 10047
rect 5825 10013 5859 10047
rect 8217 10013 8251 10047
rect 8401 10013 8435 10047
rect 8586 10013 8620 10047
rect 8769 10013 8803 10047
rect 10158 10013 10192 10047
rect 10425 10013 10459 10047
rect 10885 10013 10919 10047
rect 11141 10013 11175 10047
rect 12449 10013 12483 10047
rect 13553 10013 13587 10047
rect 13645 10013 13679 10047
rect 14289 10013 14323 10047
rect 16497 10013 16531 10047
rect 17417 10013 17451 10047
rect 18889 10013 18923 10047
rect 19533 10013 19567 10047
rect 19625 10013 19659 10047
rect 20269 10013 20303 10047
rect 21741 10013 21775 10047
rect 22293 10013 22327 10047
rect 23121 10013 23155 10047
rect 23765 10013 23799 10047
rect 23949 10013 23983 10047
rect 24593 10013 24627 10047
rect 1768 9945 1802 9979
rect 6092 9945 6126 9979
rect 14105 9945 14139 9979
rect 14933 9945 14967 9979
rect 15761 9945 15795 9979
rect 16589 9945 16623 9979
rect 18245 9945 18279 9979
rect 21097 9945 21131 9979
rect 23213 9945 23247 9979
rect 3157 9877 3191 9911
rect 5549 9877 5583 9911
rect 8125 9877 8159 9911
rect 13277 9877 13311 9911
rect 13829 9877 13863 9911
rect 14473 9877 14507 9911
rect 14841 9877 14875 9911
rect 15301 9877 15335 9911
rect 16129 9877 16163 9911
rect 16957 9877 16991 9911
rect 17877 9877 17911 9911
rect 18337 9877 18371 9911
rect 18705 9877 18739 9911
rect 20637 9877 20671 9911
rect 20729 9877 20763 9911
rect 22661 9877 22695 9911
rect 22753 9877 22787 9911
rect 24133 9877 24167 9911
rect 24409 9877 24443 9911
rect 2513 9673 2547 9707
rect 11345 9673 11379 9707
rect 15209 9673 15243 9707
rect 16681 9673 16715 9707
rect 17325 9673 17359 9707
rect 18521 9673 18555 9707
rect 18981 9673 19015 9707
rect 19441 9673 19475 9707
rect 20821 9673 20855 9707
rect 22293 9673 22327 9707
rect 23029 9673 23063 9707
rect 23121 9673 23155 9707
rect 14381 9605 14415 9639
rect 15117 9605 15151 9639
rect 16037 9605 16071 9639
rect 18061 9605 18095 9639
rect 19993 9605 20027 9639
rect 20913 9605 20947 9639
rect 22201 9605 22235 9639
rect 2697 9537 2731 9571
rect 2789 9537 2823 9571
rect 3065 9537 3099 9571
rect 3341 9537 3375 9571
rect 3617 9537 3651 9571
rect 4261 9537 4295 9571
rect 4445 9537 4479 9571
rect 9882 9537 9916 9571
rect 10149 9537 10183 9571
rect 10609 9537 10643 9571
rect 10793 9537 10827 9571
rect 11161 9537 11195 9571
rect 11529 9537 11563 9571
rect 11796 9537 11830 9571
rect 13369 9537 13403 9571
rect 13737 9537 13771 9571
rect 15669 9537 15703 9571
rect 15853 9537 15887 9571
rect 17233 9537 17267 9571
rect 19073 9537 19107 9571
rect 23673 9537 23707 9571
rect 2973 9469 3007 9503
rect 3433 9469 3467 9503
rect 13185 9469 13219 9503
rect 14105 9469 14139 9503
rect 14289 9469 14323 9503
rect 15025 9469 15059 9503
rect 17417 9469 17451 9503
rect 18153 9469 18187 9503
rect 18245 9469 18279 9503
rect 18797 9469 18831 9503
rect 20085 9469 20119 9503
rect 20177 9469 20211 9503
rect 21005 9469 21039 9503
rect 21373 9469 21407 9503
rect 21557 9469 21591 9503
rect 22385 9469 22419 9503
rect 23213 9469 23247 9503
rect 23489 9469 23523 9503
rect 4077 9401 4111 9435
rect 10793 9401 10827 9435
rect 12909 9401 12943 9435
rect 13921 9401 13955 9435
rect 17693 9401 17727 9435
rect 3157 9333 3191 9367
rect 3801 9333 3835 9367
rect 8769 9333 8803 9367
rect 10425 9333 10459 9367
rect 13553 9333 13587 9367
rect 14749 9333 14783 9367
rect 15577 9333 15611 9367
rect 16405 9333 16439 9367
rect 16865 9333 16899 9367
rect 19625 9333 19659 9367
rect 20453 9333 20487 9367
rect 21833 9333 21867 9367
rect 22661 9333 22695 9367
rect 23857 9333 23891 9367
rect 2605 9129 2639 9163
rect 3249 9129 3283 9163
rect 3893 9129 3927 9163
rect 6009 9129 6043 9163
rect 7849 9129 7883 9163
rect 12081 9129 12115 9163
rect 17233 9129 17267 9163
rect 17325 9129 17359 9163
rect 18889 9129 18923 9163
rect 20637 9129 20671 9163
rect 23305 9129 23339 9163
rect 4537 9061 4571 9095
rect 12357 9061 12391 9095
rect 12725 9061 12759 9095
rect 3341 8993 3375 9027
rect 3801 8993 3835 9027
rect 11805 8993 11839 9027
rect 14657 8993 14691 9027
rect 15209 8993 15243 9027
rect 17233 8993 17267 9027
rect 17601 8993 17635 9027
rect 18337 8993 18371 9027
rect 19717 8993 19751 9027
rect 19901 8993 19935 9027
rect 20085 8993 20119 9027
rect 23029 8993 23063 9027
rect 2421 8925 2455 8959
rect 2973 8925 3007 8959
rect 3065 8925 3099 8959
rect 3617 8925 3651 8959
rect 4077 8925 4111 8959
rect 4169 8925 4203 8959
rect 4721 8925 4755 8959
rect 5181 8925 5215 8959
rect 6193 8925 6227 8959
rect 7481 8925 7515 8959
rect 7665 8925 7699 8959
rect 12541 8925 12575 8959
rect 12633 8925 12667 8959
rect 12817 8925 12851 8959
rect 13001 8925 13035 8959
rect 13185 8925 13219 8959
rect 13369 8925 13403 8959
rect 13645 8925 13679 8959
rect 13921 8925 13955 8959
rect 14473 8925 14507 8959
rect 14565 8925 14599 8959
rect 14933 8925 14967 8959
rect 17785 8925 17819 8959
rect 18521 8925 18555 8959
rect 18705 8925 18739 8959
rect 19073 8925 19107 8959
rect 19625 8925 19659 8959
rect 20269 8925 20303 8959
rect 20453 8925 20487 8959
rect 20821 8925 20855 8959
rect 22845 8925 22879 8959
rect 22937 8925 22971 8959
rect 23489 8925 23523 8959
rect 11437 8857 11471 8891
rect 11897 8857 11931 8891
rect 17877 8857 17911 8891
rect 20913 8857 20947 8891
rect 21097 8857 21131 8891
rect 21649 8857 21683 8891
rect 22293 8857 22327 8891
rect 2789 8789 2823 8823
rect 3525 8789 3559 8823
rect 4353 8789 4387 8823
rect 5365 8789 5399 8823
rect 7389 8789 7423 8823
rect 11713 8789 11747 8823
rect 13553 8789 13587 8823
rect 13737 8789 13771 8823
rect 14105 8789 14139 8823
rect 15117 8789 15151 8823
rect 18245 8789 18279 8823
rect 19257 8789 19291 8823
rect 22477 8789 22511 8823
rect 1593 8585 1627 8619
rect 4445 8585 4479 8619
rect 6009 8585 6043 8619
rect 9321 8585 9355 8619
rect 11805 8585 11839 8619
rect 12449 8585 12483 8619
rect 12817 8585 12851 8619
rect 13093 8585 13127 8619
rect 13737 8585 13771 8619
rect 14289 8585 14323 8619
rect 15669 8585 15703 8619
rect 19073 8585 19107 8619
rect 12633 8517 12667 8551
rect 13829 8517 13863 8551
rect 2706 8449 2740 8483
rect 2973 8449 3007 8483
rect 3065 8449 3099 8483
rect 3332 8449 3366 8483
rect 4629 8449 4663 8483
rect 4885 8449 4919 8483
rect 6745 8449 6779 8483
rect 7113 8449 7147 8483
rect 7380 8449 7414 8483
rect 8861 8449 8895 8483
rect 9045 8449 9079 8483
rect 9229 8449 9263 8483
rect 11897 8449 11931 8483
rect 6561 8381 6595 8415
rect 11345 8381 11379 8415
rect 11713 8381 11747 8415
rect 13277 8449 13311 8483
rect 14473 8449 14507 8483
rect 12909 8381 12943 8415
rect 13553 8381 13587 8415
rect 8493 8313 8527 8347
rect 8861 8313 8895 8347
rect 12633 8313 12667 8347
rect 14841 8313 14875 8347
rect 6929 8245 6963 8279
rect 12265 8245 12299 8279
rect 14197 8245 14231 8279
rect 14657 8245 14691 8279
rect 16129 8245 16163 8279
rect 22109 8245 22143 8279
rect 4537 8041 4571 8075
rect 5365 8041 5399 8075
rect 6469 8041 6503 8075
rect 8125 8041 8159 8075
rect 8585 8041 8619 8075
rect 9229 8041 9263 8075
rect 9781 8041 9815 8075
rect 10241 8041 10275 8075
rect 13277 8041 13311 8075
rect 18153 8041 18187 8075
rect 7389 7973 7423 8007
rect 7665 7973 7699 8007
rect 9045 7973 9079 8007
rect 14105 7973 14139 8007
rect 3525 7905 3559 7939
rect 4813 7905 4847 7939
rect 5181 7905 5215 7939
rect 7021 7905 7055 7939
rect 8217 7905 8251 7939
rect 9321 7905 9355 7939
rect 12265 7905 12299 7939
rect 12449 7905 12483 7939
rect 14565 7905 14599 7939
rect 14657 7905 14691 7939
rect 15577 7905 15611 7939
rect 16773 7905 16807 7939
rect 18889 7905 18923 7939
rect 19717 7905 19751 7939
rect 21281 7905 21315 7939
rect 21557 7905 21591 7939
rect 22753 7905 22787 7939
rect 2881 7837 2915 7871
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 3617 7837 3651 7871
rect 3985 7837 4019 7871
rect 4358 7837 4392 7871
rect 4997 7837 5031 7871
rect 5549 7837 5583 7871
rect 5825 7837 5859 7871
rect 6193 7837 6227 7871
rect 6377 7837 6411 7871
rect 6837 7837 6871 7871
rect 7481 7837 7515 7871
rect 7849 7837 7883 7871
rect 7941 7837 7975 7871
rect 8677 7837 8711 7871
rect 8769 7837 8803 7871
rect 9229 7837 9263 7871
rect 9597 7837 9631 7871
rect 9873 7837 9907 7871
rect 12081 7837 12115 7871
rect 13829 7837 13863 7871
rect 14473 7837 14507 7871
rect 16037 7837 16071 7871
rect 16589 7837 16623 7871
rect 17234 7837 17268 7871
rect 17601 7837 17635 7871
rect 17693 7837 17727 7871
rect 18429 7837 18463 7871
rect 18705 7837 18739 7871
rect 21741 7837 21775 7871
rect 22569 7837 22603 7871
rect 23029 7837 23063 7871
rect 4169 7769 4203 7803
rect 4261 7769 4295 7803
rect 6009 7769 6043 7803
rect 6929 7769 6963 7803
rect 9505 7769 9539 7803
rect 12541 7769 12575 7803
rect 15301 7769 15335 7803
rect 16681 7769 16715 7803
rect 17049 7769 17083 7803
rect 17785 7769 17819 7803
rect 18199 7769 18233 7803
rect 21649 7769 21683 7803
rect 2697 7701 2731 7735
rect 3065 7701 3099 7735
rect 3893 7701 3927 7735
rect 5733 7701 5767 7735
rect 8401 7701 8435 7735
rect 10057 7701 10091 7735
rect 12909 7701 12943 7735
rect 14933 7701 14967 7735
rect 15393 7701 15427 7735
rect 15945 7701 15979 7735
rect 16221 7701 16255 7735
rect 18521 7701 18555 7735
rect 22109 7701 22143 7735
rect 22201 7701 22235 7735
rect 22661 7701 22695 7735
rect 23213 7701 23247 7735
rect 4537 7497 4571 7531
rect 9321 7497 9355 7531
rect 11529 7497 11563 7531
rect 15954 7497 15988 7531
rect 16497 7497 16531 7531
rect 18245 7497 18279 7531
rect 18613 7497 18647 7531
rect 19450 7497 19484 7531
rect 20177 7497 20211 7531
rect 4997 7429 5031 7463
rect 6009 7429 6043 7463
rect 6377 7429 6411 7463
rect 7297 7429 7331 7463
rect 7757 7429 7791 7463
rect 7941 7429 7975 7463
rect 8309 7429 8343 7463
rect 8493 7429 8527 7463
rect 9045 7429 9079 7463
rect 16926 7429 16960 7463
rect 21382 7429 21416 7463
rect 22210 7429 22244 7463
rect 23204 7429 23238 7463
rect 3157 7361 3191 7395
rect 3413 7361 3447 7395
rect 4813 7361 4847 7395
rect 6561 7361 6595 7395
rect 6745 7361 6779 7395
rect 7015 7361 7049 7395
rect 7481 7361 7515 7395
rect 8769 7361 8803 7395
rect 9137 7361 9171 7395
rect 9413 7361 9447 7395
rect 9689 7361 9723 7395
rect 10241 7361 10275 7395
rect 10425 7361 10459 7395
rect 10701 7361 10735 7395
rect 10885 7361 10919 7395
rect 11161 7361 11195 7395
rect 11713 7361 11747 7395
rect 11989 7361 12023 7395
rect 12081 7361 12115 7395
rect 13737 7361 13771 7395
rect 14013 7361 14047 7395
rect 14280 7361 14314 7395
rect 15577 7361 15611 7395
rect 16221 7361 16255 7395
rect 16313 7361 16347 7395
rect 19073 7361 19107 7395
rect 20269 7361 20303 7395
rect 21005 7361 21039 7395
rect 21649 7361 21683 7395
rect 21833 7361 21867 7395
rect 22477 7361 22511 7395
rect 22569 7361 22603 7395
rect 22937 7361 22971 7395
rect 6837 7293 6871 7327
rect 7389 7293 7423 7327
rect 8585 7293 8619 7327
rect 9505 7293 9539 7327
rect 10517 7293 10551 7327
rect 16681 7293 16715 7327
rect 18705 7293 18739 7327
rect 18889 7293 18923 7327
rect 20361 7293 20395 7327
rect 8125 7225 8159 7259
rect 9873 7225 9907 7259
rect 19809 7225 19843 7259
rect 7757 7157 7791 7191
rect 10057 7157 10091 7191
rect 11069 7157 11103 7191
rect 11345 7157 11379 7191
rect 11805 7157 11839 7191
rect 12265 7157 12299 7191
rect 13921 7157 13955 7191
rect 15393 7157 15427 7191
rect 15945 7157 15979 7191
rect 18061 7157 18095 7191
rect 19441 7157 19475 7191
rect 19625 7157 19659 7191
rect 21373 7157 21407 7191
rect 22201 7157 22235 7191
rect 22753 7157 22787 7191
rect 24317 7157 24351 7191
rect 6745 6953 6779 6987
rect 8125 6953 8159 6987
rect 10333 6953 10367 6987
rect 12449 6953 12483 6987
rect 14197 6953 14231 6987
rect 14381 6953 14415 6987
rect 15577 6953 15611 6987
rect 17141 6953 17175 6987
rect 19441 6953 19475 6987
rect 23305 6953 23339 6987
rect 9137 6885 9171 6919
rect 16773 6885 16807 6919
rect 12173 6817 12207 6851
rect 14933 6817 14967 6851
rect 6561 6749 6595 6783
rect 7297 6749 7331 6783
rect 8217 6749 8251 6783
rect 8493 6749 8527 6783
rect 8953 6749 8987 6783
rect 10609 6749 10643 6783
rect 11906 6749 11940 6783
rect 12265 6749 12299 6783
rect 12541 6749 12575 6783
rect 12817 6749 12851 6783
rect 12909 6749 12943 6783
rect 15117 6749 15151 6783
rect 15301 6749 15335 6783
rect 15669 6749 15703 6783
rect 15853 6749 15887 6783
rect 17049 6749 17083 6783
rect 17141 6749 17175 6783
rect 18705 6749 18739 6783
rect 19257 6749 19291 6783
rect 19533 6749 19567 6783
rect 23121 6749 23155 6783
rect 23455 6749 23489 6783
rect 23765 6749 23799 6783
rect 23857 6749 23891 6783
rect 9965 6681 9999 6715
rect 10379 6681 10413 6715
rect 14372 6681 14406 6715
rect 14749 6681 14783 6715
rect 15393 6681 15427 6715
rect 18438 6681 18472 6715
rect 18889 6681 18923 6715
rect 19073 6681 19107 6715
rect 19778 6681 19812 6715
rect 22854 6681 22888 6715
rect 7113 6613 7147 6647
rect 8401 6613 8435 6647
rect 10793 6613 10827 6647
rect 12725 6613 12759 6647
rect 17325 6613 17359 6647
rect 20913 6613 20947 6647
rect 21741 6613 21775 6647
rect 6009 6409 6043 6443
rect 7021 6409 7055 6443
rect 7481 6409 7515 6443
rect 10977 6409 11011 6443
rect 11897 6409 11931 6443
rect 11989 6409 12023 6443
rect 14749 6409 14783 6443
rect 19441 6409 19475 6443
rect 20729 6409 20763 6443
rect 6561 6341 6595 6375
rect 8217 6341 8251 6375
rect 14841 6341 14875 6375
rect 18521 6341 18555 6375
rect 23489 6341 23523 6375
rect 23857 6341 23891 6375
rect 6745 6273 6779 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 7389 6273 7423 6307
rect 7757 6273 7791 6307
rect 10609 6273 10643 6307
rect 10793 6273 10827 6307
rect 11161 6273 11195 6307
rect 18336 6273 18370 6307
rect 18613 6273 18647 6307
rect 18797 6273 18831 6307
rect 18981 6273 19015 6307
rect 19257 6273 19291 6307
rect 19993 6273 20027 6307
rect 20879 6273 20913 6307
rect 21281 6273 21315 6307
rect 22386 6273 22420 6307
rect 22753 6273 22787 6307
rect 22845 6273 22879 6307
rect 23397 6273 23431 6307
rect 23673 6273 23707 6307
rect 6377 6205 6411 6239
rect 12173 6205 12207 6239
rect 17877 6205 17911 6239
rect 17969 6205 18003 6239
rect 21189 6205 21223 6239
rect 22201 6205 22235 6239
rect 23305 6205 23339 6239
rect 6193 6137 6227 6171
rect 11529 6137 11563 6171
rect 23029 6137 23063 6171
rect 7849 6069 7883 6103
rect 8125 6069 8159 6103
rect 11345 6069 11379 6103
rect 20177 6069 20211 6103
rect 23397 6069 23431 6103
rect 5181 5865 5215 5899
rect 5549 5865 5583 5899
rect 10149 5865 10183 5899
rect 21649 5865 21683 5899
rect 5641 5797 5675 5831
rect 7389 5797 7423 5831
rect 8401 5797 8435 5831
rect 9965 5797 9999 5831
rect 6837 5729 6871 5763
rect 6929 5729 6963 5763
rect 7113 5729 7147 5763
rect 8033 5729 8067 5763
rect 10885 5729 10919 5763
rect 21465 5729 21499 5763
rect 5365 5661 5399 5695
rect 5825 5661 5859 5695
rect 6101 5661 6135 5695
rect 6285 5661 6319 5695
rect 7021 5661 7055 5695
rect 7293 5671 7327 5705
rect 8217 5661 8251 5695
rect 8493 5661 8527 5695
rect 8769 5661 8803 5695
rect 8953 5661 8987 5695
rect 9137 5661 9171 5695
rect 9321 5661 9355 5695
rect 9781 5661 9815 5695
rect 10609 5661 10643 5695
rect 18613 5661 18647 5695
rect 21649 5661 21683 5695
rect 6009 5593 6043 5627
rect 6469 5593 6503 5627
rect 21373 5593 21407 5627
rect 6653 5525 6687 5559
rect 7757 5525 7791 5559
rect 7849 5525 7883 5559
rect 8493 5525 8527 5559
rect 8677 5525 8711 5559
rect 10241 5525 10275 5559
rect 10701 5525 10735 5559
rect 11437 5525 11471 5559
rect 13093 5525 13127 5559
rect 13829 5525 13863 5559
rect 18797 5525 18831 5559
rect 21833 5525 21867 5559
rect 4813 5321 4847 5355
rect 6193 5321 6227 5355
rect 6561 5321 6595 5355
rect 8769 5321 8803 5355
rect 11621 5321 11655 5355
rect 13553 5321 13587 5355
rect 14381 5321 14415 5355
rect 15393 5321 15427 5355
rect 17969 5321 18003 5355
rect 18889 5321 18923 5355
rect 19441 5321 19475 5355
rect 21005 5321 21039 5355
rect 22753 5321 22787 5355
rect 8309 5253 8343 5287
rect 10434 5253 10468 5287
rect 18705 5253 18739 5287
rect 21833 5253 21867 5287
rect 22201 5253 22235 5287
rect 24317 5253 24351 5287
rect 3433 5185 3467 5219
rect 3700 5185 3734 5219
rect 5181 5185 5215 5219
rect 5273 5185 5307 5219
rect 5825 5185 5859 5219
rect 6377 5185 6411 5219
rect 7021 5185 7055 5219
rect 7389 5185 7423 5219
rect 7481 5185 7515 5219
rect 7629 5185 7663 5219
rect 7754 5185 7788 5219
rect 8033 5185 8067 5219
rect 8585 5185 8619 5219
rect 9137 5185 9171 5219
rect 9413 5185 9447 5219
rect 10057 5185 10091 5219
rect 10793 5185 10827 5219
rect 11253 5185 11287 5219
rect 11805 5185 11839 5219
rect 12817 5185 12851 5219
rect 12909 5185 12943 5219
rect 13645 5185 13679 5219
rect 15485 5185 15519 5219
rect 16681 5185 16715 5219
rect 16866 5185 16900 5219
rect 17509 5185 17543 5219
rect 18613 5185 18647 5219
rect 20143 5185 20177 5219
rect 21373 5185 21407 5219
rect 22845 5185 22879 5219
rect 23213 5185 23247 5219
rect 23455 5185 23489 5219
rect 23949 5185 23983 5219
rect 24133 5185 24167 5219
rect 5641 5117 5675 5151
rect 5733 5117 5767 5151
rect 6929 5117 6963 5151
rect 7113 5117 7147 5151
rect 7205 5117 7239 5151
rect 7849 5117 7883 5151
rect 8401 5117 8435 5151
rect 13829 5117 13863 5151
rect 14473 5117 14507 5151
rect 14657 5117 14691 5151
rect 14933 5117 14967 5151
rect 15669 5117 15703 5151
rect 17233 5117 17267 5151
rect 17325 5117 17359 5151
rect 18061 5117 18095 5151
rect 18245 5117 18279 5151
rect 18705 5117 18739 5151
rect 19533 5117 19567 5151
rect 19625 5117 19659 5151
rect 20453 5117 20487 5151
rect 20545 5117 20579 5151
rect 21281 5117 21315 5151
rect 22937 5117 22971 5151
rect 23765 5117 23799 5151
rect 23857 5117 23891 5151
rect 5089 5049 5123 5083
rect 8953 5049 8987 5083
rect 10609 5049 10643 5083
rect 10977 5049 11011 5083
rect 13185 5049 13219 5083
rect 19901 5049 19935 5083
rect 6745 4981 6779 5015
rect 8125 4981 8159 5015
rect 8309 4981 8343 5015
rect 9229 4981 9263 5015
rect 10425 4981 10459 5015
rect 11069 4981 11103 5015
rect 12633 4981 12667 5015
rect 13093 4981 13127 5015
rect 14013 4981 14047 5015
rect 15025 4981 15059 5015
rect 16221 4981 16255 5015
rect 17601 4981 17635 5015
rect 18429 4981 18463 5015
rect 19073 4981 19107 5015
rect 21373 4981 21407 5015
rect 22385 4981 22419 5015
rect 3617 4777 3651 4811
rect 5273 4777 5307 4811
rect 6745 4777 6779 4811
rect 7573 4777 7607 4811
rect 8677 4777 8711 4811
rect 10241 4777 10275 4811
rect 12081 4777 12115 4811
rect 13553 4777 13587 4811
rect 14657 4777 14691 4811
rect 15577 4777 15611 4811
rect 17509 4777 17543 4811
rect 18797 4777 18831 4811
rect 20545 4777 20579 4811
rect 21281 4777 21315 4811
rect 21741 4777 21775 4811
rect 24133 4777 24167 4811
rect 5549 4709 5583 4743
rect 8217 4709 8251 4743
rect 9045 4709 9079 4743
rect 9965 4709 9999 4743
rect 10149 4709 10183 4743
rect 16221 4709 16255 4743
rect 19441 4709 19475 4743
rect 6009 4641 6043 4675
rect 7021 4641 7055 4675
rect 10793 4641 10827 4675
rect 11713 4641 11747 4675
rect 12725 4641 12759 4675
rect 15025 4641 15059 4675
rect 16405 4641 16439 4675
rect 20177 4641 20211 4675
rect 21649 4641 21683 4675
rect 22477 4641 22511 4675
rect 22753 4641 22787 4675
rect 3433 4573 3467 4607
rect 3893 4573 3927 4607
rect 4160 4573 4194 4607
rect 5733 4573 5767 4607
rect 5917 4573 5951 4607
rect 6193 4573 6227 4607
rect 6561 4573 6595 4607
rect 6929 4573 6963 4607
rect 7113 4573 7147 4607
rect 7205 4573 7239 4607
rect 7389 4573 7423 4607
rect 7481 4573 7515 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 8309 4573 8343 4607
rect 8585 4573 8619 4607
rect 10609 4573 10643 4607
rect 11311 4573 11345 4607
rect 11621 4573 11655 4607
rect 12541 4573 12575 4607
rect 13001 4573 13035 4607
rect 13277 4573 13311 4607
rect 13921 4573 13955 4607
rect 14289 4573 14323 4607
rect 14933 4573 14967 4607
rect 15117 4573 15151 4607
rect 15427 4573 15461 4607
rect 15853 4573 15887 4607
rect 16681 4573 16715 4607
rect 17141 4573 17175 4607
rect 17785 4573 17819 4607
rect 17877 4573 17911 4607
rect 19073 4573 19107 4607
rect 20729 4573 20763 4607
rect 20913 4573 20947 4607
rect 21005 4573 21039 4607
rect 21465 4573 21499 4607
rect 21741 4573 21775 4607
rect 22293 4573 22327 4607
rect 24593 4573 24627 4607
rect 10701 4505 10735 4539
rect 11069 4505 11103 4539
rect 13544 4505 13578 4539
rect 14666 4505 14700 4539
rect 16037 4505 16071 4539
rect 18429 4505 18463 4539
rect 18806 4505 18840 4539
rect 19993 4505 20027 4539
rect 23020 4505 23054 4539
rect 6193 4437 6227 4471
rect 8401 4437 8435 4471
rect 12173 4437 12207 4471
rect 12633 4437 12667 4471
rect 13185 4437 13219 4471
rect 16589 4437 16623 4471
rect 17049 4437 17083 4471
rect 17518 4437 17552 4471
rect 18061 4437 18095 4471
rect 19625 4437 19659 4471
rect 20085 4437 20119 4471
rect 21925 4437 21959 4471
rect 22385 4437 22419 4471
rect 24409 4437 24443 4471
rect 6837 4233 6871 4267
rect 7205 4233 7239 4267
rect 7757 4233 7791 4267
rect 9698 4233 9732 4267
rect 10425 4233 10459 4267
rect 11980 4233 12014 4267
rect 12826 4233 12860 4267
rect 13737 4233 13771 4267
rect 16948 4233 16982 4267
rect 20002 4233 20036 4267
rect 21382 4233 21416 4267
rect 22302 4233 22336 4267
rect 3525 4165 3559 4199
rect 9321 4165 9355 4199
rect 11345 4165 11379 4199
rect 12357 4165 12391 4199
rect 12449 4165 12483 4199
rect 17325 4165 17359 4199
rect 18306 4165 18340 4199
rect 19625 4165 19659 4199
rect 21005 4165 21039 4199
rect 21925 4165 21959 4199
rect 22661 4165 22695 4199
rect 23765 4165 23799 4199
rect 3157 4097 3191 4131
rect 3341 4097 3375 4131
rect 3709 4097 3743 4131
rect 5825 4097 5859 4131
rect 6101 4097 6135 4131
rect 7573 4097 7607 4131
rect 7849 4097 7883 4131
rect 10977 4097 11011 4131
rect 11161 4097 11195 4131
rect 13587 4097 13621 4131
rect 13921 4097 13955 4131
rect 14177 4097 14211 4131
rect 15485 4097 15519 4131
rect 16095 4097 16129 4131
rect 16405 4097 16439 4131
rect 17417 4097 17451 4131
rect 20545 4097 20579 4131
rect 20913 4097 20947 4131
rect 22903 4097 22937 4131
rect 23397 4097 23431 4131
rect 23581 4097 23615 4131
rect 6193 4029 6227 4063
rect 6561 4029 6595 4063
rect 6745 4029 6779 4063
rect 10517 4029 10551 4063
rect 10701 4029 10735 4063
rect 13185 4029 13219 4063
rect 13277 4029 13311 4063
rect 16497 4029 16531 4063
rect 17509 4029 17543 4063
rect 18061 4029 18095 4063
rect 20729 4029 20763 4063
rect 23213 4029 23247 4063
rect 23305 4029 23339 4063
rect 7389 3961 7423 3995
rect 10057 3961 10091 3995
rect 17785 3961 17819 3995
rect 19441 3961 19475 3995
rect 20545 3961 20579 3995
rect 22477 3961 22511 3995
rect 2973 3893 3007 3927
rect 7941 3893 7975 3927
rect 8861 3893 8895 3927
rect 9689 3893 9723 3927
rect 9873 3893 9907 3927
rect 11805 3893 11839 3927
rect 11989 3893 12023 3927
rect 12817 3893 12851 3927
rect 13001 3893 13035 3927
rect 15301 3893 15335 3927
rect 15669 3893 15703 3927
rect 15945 3893 15979 3927
rect 16773 3893 16807 3927
rect 16957 3893 16991 3927
rect 17417 3893 17451 3927
rect 19993 3893 20027 3927
rect 20177 3893 20211 3927
rect 21373 3893 21407 3927
rect 21557 3893 21591 3927
rect 22293 3893 22327 3927
rect 6285 3689 6319 3723
rect 6837 3689 6871 3723
rect 8401 3689 8435 3723
rect 8769 3689 8803 3723
rect 11253 3689 11287 3723
rect 11989 3689 12023 3723
rect 14841 3689 14875 3723
rect 15209 3689 15243 3723
rect 17049 3689 17083 3723
rect 21005 3689 21039 3723
rect 21189 3689 21223 3723
rect 21741 3689 21775 3723
rect 23581 3689 23615 3723
rect 14105 3621 14139 3655
rect 16773 3621 16807 3655
rect 8217 3553 8251 3587
rect 9873 3553 9907 3587
rect 11437 3553 11471 3587
rect 15393 3553 15427 3587
rect 18429 3553 18463 3587
rect 19349 3553 19383 3587
rect 21281 3553 21315 3587
rect 7961 3485 7995 3519
rect 8585 3485 8619 3519
rect 8769 3485 8803 3519
rect 9137 3485 9171 3519
rect 9229 3485 9263 3519
rect 9597 3485 9631 3519
rect 11529 3485 11563 3519
rect 11896 3485 11930 3519
rect 12173 3485 12207 3519
rect 13921 3485 13955 3519
rect 14347 3485 14381 3519
rect 14657 3485 14691 3519
rect 14749 3485 14783 3519
rect 14841 3485 14875 3519
rect 15025 3485 15059 3519
rect 15660 3485 15694 3519
rect 18889 3485 18923 3519
rect 21373 3485 21407 3519
rect 21925 3485 21959 3519
rect 22201 3485 22235 3519
rect 24041 3485 24075 3519
rect 25145 3485 25179 3519
rect 10140 3417 10174 3451
rect 12440 3417 12474 3451
rect 18162 3417 18196 3451
rect 19616 3417 19650 3451
rect 21465 3417 21499 3451
rect 21649 3417 21683 3451
rect 22446 3417 22480 3451
rect 9045 3349 9079 3383
rect 9781 3349 9815 3383
rect 13553 3349 13587 3383
rect 13737 3349 13771 3383
rect 19073 3349 19107 3383
rect 20729 3349 20763 3383
rect 22109 3349 22143 3383
rect 7757 3145 7791 3179
rect 8861 3145 8895 3179
rect 9229 3145 9263 3179
rect 10977 3145 11011 3179
rect 12449 3145 12483 3179
rect 14473 3145 14507 3179
rect 16865 3145 16899 3179
rect 19533 3145 19567 3179
rect 21189 3145 21223 3179
rect 21465 3145 21499 3179
rect 6622 3077 6656 3111
rect 9137 3077 9171 3111
rect 11529 3077 11563 3111
rect 14841 3077 14875 3111
rect 15025 3077 15059 3111
rect 20054 3077 20088 3111
rect 6377 3009 6411 3043
rect 8769 3009 8803 3043
rect 9413 3009 9447 3043
rect 9680 3009 9714 3043
rect 11161 3009 11195 3043
rect 11713 3009 11747 3043
rect 12633 3009 12667 3043
rect 13093 3009 13127 3043
rect 13360 3009 13394 3043
rect 14657 3009 14691 3043
rect 16681 3009 16715 3043
rect 19349 3009 19383 3043
rect 19809 3009 19843 3043
rect 21373 3009 21407 3043
rect 8677 2941 8711 2975
rect 11897 2941 11931 2975
rect 8401 2873 8435 2907
rect 10793 2873 10827 2907
rect 21833 2805 21867 2839
rect 22753 2805 22787 2839
rect 9873 2601 9907 2635
rect 13461 2601 13495 2635
rect 20453 2533 20487 2567
rect 10057 2397 10091 2431
rect 13185 2397 13219 2431
rect 13369 2397 13403 2431
rect 20177 2397 20211 2431
rect 20545 2397 20579 2431
rect 20729 2397 20763 2431
<< metal1 >>
rect 26326 28744 26332 28756
rect 26287 28716 26332 28744
rect 26326 28704 26332 28716
rect 26384 28704 26390 28756
rect 1104 27226 26220 27248
rect 1104 27174 9322 27226
rect 9374 27174 9386 27226
rect 9438 27174 9450 27226
rect 9502 27174 9514 27226
rect 9566 27174 9578 27226
rect 9630 27174 17694 27226
rect 17746 27174 17758 27226
rect 17810 27174 17822 27226
rect 17874 27174 17886 27226
rect 17938 27174 17950 27226
rect 18002 27174 26220 27226
rect 1104 27152 26220 27174
rect 9766 26976 9772 26988
rect 9727 26948 9772 26976
rect 9766 26936 9772 26948
rect 9824 26936 9830 26988
rect 14090 26976 14096 26988
rect 14051 26948 14096 26976
rect 14090 26936 14096 26948
rect 14148 26936 14154 26988
rect 9950 26772 9956 26784
rect 9911 26744 9956 26772
rect 9950 26732 9956 26744
rect 10008 26732 10014 26784
rect 14277 26775 14335 26781
rect 14277 26741 14289 26775
rect 14323 26772 14335 26775
rect 14642 26772 14648 26784
rect 14323 26744 14648 26772
rect 14323 26741 14335 26744
rect 14277 26735 14335 26741
rect 14642 26732 14648 26744
rect 14700 26732 14706 26784
rect 1104 26682 26220 26704
rect 1104 26630 5136 26682
rect 5188 26630 5200 26682
rect 5252 26630 5264 26682
rect 5316 26630 5328 26682
rect 5380 26630 5392 26682
rect 5444 26630 13508 26682
rect 13560 26630 13572 26682
rect 13624 26630 13636 26682
rect 13688 26630 13700 26682
rect 13752 26630 13764 26682
rect 13816 26630 21880 26682
rect 21932 26630 21944 26682
rect 21996 26630 22008 26682
rect 22060 26630 22072 26682
rect 22124 26630 22136 26682
rect 22188 26630 26220 26682
rect 1104 26608 26220 26630
rect 13633 26571 13691 26577
rect 13633 26537 13645 26571
rect 13679 26568 13691 26571
rect 14090 26568 14096 26580
rect 13679 26540 14096 26568
rect 13679 26537 13691 26540
rect 13633 26531 13691 26537
rect 14090 26528 14096 26540
rect 14148 26528 14154 26580
rect 6825 26503 6883 26509
rect 6825 26469 6837 26503
rect 6871 26500 6883 26503
rect 7006 26500 7012 26512
rect 6871 26472 7012 26500
rect 6871 26469 6883 26472
rect 6825 26463 6883 26469
rect 7006 26460 7012 26472
rect 7064 26460 7070 26512
rect 9214 26460 9220 26512
rect 9272 26500 9278 26512
rect 9493 26503 9551 26509
rect 9493 26500 9505 26503
rect 9272 26472 9505 26500
rect 9272 26460 9278 26472
rect 9493 26469 9505 26472
rect 9539 26469 9551 26503
rect 10686 26500 10692 26512
rect 9493 26463 9551 26469
rect 10152 26472 10692 26500
rect 10152 26441 10180 26472
rect 10686 26460 10692 26472
rect 10744 26500 10750 26512
rect 11057 26503 11115 26509
rect 11057 26500 11069 26503
rect 10744 26472 11069 26500
rect 10744 26460 10750 26472
rect 11057 26469 11069 26472
rect 11103 26469 11115 26503
rect 11057 26463 11115 26469
rect 13541 26503 13599 26509
rect 13541 26469 13553 26503
rect 13587 26500 13599 26503
rect 13906 26500 13912 26512
rect 13587 26472 13912 26500
rect 13587 26469 13599 26472
rect 13541 26463 13599 26469
rect 13906 26460 13912 26472
rect 13964 26460 13970 26512
rect 14734 26500 14740 26512
rect 14660 26472 14740 26500
rect 10137 26435 10195 26441
rect 10137 26401 10149 26435
rect 10183 26401 10195 26435
rect 10137 26395 10195 26401
rect 10873 26435 10931 26441
rect 10873 26401 10885 26435
rect 10919 26432 10931 26435
rect 11238 26432 11244 26444
rect 10919 26404 11244 26432
rect 10919 26401 10931 26404
rect 10873 26395 10931 26401
rect 11238 26392 11244 26404
rect 11296 26392 11302 26444
rect 14660 26441 14688 26472
rect 14734 26460 14740 26472
rect 14792 26460 14798 26512
rect 14645 26435 14703 26441
rect 14645 26401 14657 26435
rect 14691 26401 14703 26435
rect 14645 26395 14703 26401
rect 7009 26367 7067 26373
rect 7009 26333 7021 26367
rect 7055 26364 7067 26367
rect 7098 26364 7104 26376
rect 7055 26336 7104 26364
rect 7055 26333 7067 26336
rect 7009 26327 7067 26333
rect 7098 26324 7104 26336
rect 7156 26324 7162 26376
rect 7282 26364 7288 26376
rect 7243 26336 7288 26364
rect 7282 26324 7288 26336
rect 7340 26324 7346 26376
rect 9401 26367 9459 26373
rect 9401 26333 9413 26367
rect 9447 26364 9459 26367
rect 9674 26364 9680 26376
rect 9447 26336 9680 26364
rect 9447 26333 9459 26336
rect 9401 26327 9459 26333
rect 9674 26324 9680 26336
rect 9732 26324 9738 26376
rect 10563 26367 10621 26373
rect 10563 26333 10575 26367
rect 10609 26364 10621 26367
rect 10962 26364 10968 26376
rect 10609 26336 10824 26364
rect 10923 26336 10968 26364
rect 10609 26333 10621 26336
rect 10563 26327 10621 26333
rect 9122 26256 9128 26308
rect 9180 26296 9186 26308
rect 9309 26299 9367 26305
rect 9309 26296 9321 26299
rect 9180 26268 9321 26296
rect 9180 26256 9186 26268
rect 9309 26265 9321 26268
rect 9355 26265 9367 26299
rect 9309 26259 9367 26265
rect 9953 26299 10011 26305
rect 9953 26265 9965 26299
rect 9999 26296 10011 26299
rect 10321 26299 10379 26305
rect 10321 26296 10333 26299
rect 9999 26268 10333 26296
rect 9999 26265 10011 26268
rect 9953 26259 10011 26265
rect 10321 26265 10333 26268
rect 10367 26265 10379 26299
rect 10796 26296 10824 26336
rect 10962 26324 10968 26336
rect 11020 26324 11026 26376
rect 14335 26367 14393 26373
rect 14335 26333 14347 26367
rect 14381 26364 14393 26367
rect 14737 26367 14795 26373
rect 14381 26336 14596 26364
rect 14381 26333 14393 26336
rect 14335 26327 14393 26333
rect 11882 26296 11888 26308
rect 10796 26268 11888 26296
rect 10321 26259 10379 26265
rect 11882 26256 11888 26268
rect 11940 26256 11946 26308
rect 12434 26256 12440 26308
rect 12492 26296 12498 26308
rect 13173 26299 13231 26305
rect 13173 26296 13185 26299
rect 12492 26268 13185 26296
rect 12492 26256 12498 26268
rect 13173 26265 13185 26268
rect 13219 26265 13231 26299
rect 14090 26296 14096 26308
rect 14051 26268 14096 26296
rect 13173 26259 13231 26265
rect 14090 26256 14096 26268
rect 14148 26256 14154 26308
rect 14568 26296 14596 26336
rect 14737 26333 14749 26367
rect 14783 26364 14795 26367
rect 15102 26364 15108 26376
rect 14783 26336 15108 26364
rect 14783 26333 14795 26336
rect 14737 26327 14795 26333
rect 15102 26324 15108 26336
rect 15160 26364 15166 26376
rect 15197 26367 15255 26373
rect 15197 26364 15209 26367
rect 15160 26336 15209 26364
rect 15160 26324 15166 26336
rect 15197 26333 15209 26336
rect 15243 26333 15255 26367
rect 15197 26327 15255 26333
rect 14829 26299 14887 26305
rect 14829 26296 14841 26299
rect 14568 26268 14841 26296
rect 14829 26265 14841 26268
rect 14875 26296 14887 26299
rect 14918 26296 14924 26308
rect 14875 26268 14924 26296
rect 14875 26265 14887 26268
rect 14829 26259 14887 26265
rect 14918 26256 14924 26268
rect 14976 26256 14982 26308
rect 15013 26299 15071 26305
rect 15013 26265 15025 26299
rect 15059 26265 15071 26299
rect 15013 26259 15071 26265
rect 7190 26228 7196 26240
rect 7151 26200 7196 26228
rect 7190 26188 7196 26200
rect 7248 26188 7254 26240
rect 9858 26228 9864 26240
rect 9819 26200 9864 26228
rect 9858 26188 9864 26200
rect 9916 26188 9922 26240
rect 14734 26188 14740 26240
rect 14792 26228 14798 26240
rect 15028 26228 15056 26259
rect 14792 26200 15056 26228
rect 14792 26188 14798 26200
rect 1104 26138 26220 26160
rect 1104 26086 9322 26138
rect 9374 26086 9386 26138
rect 9438 26086 9450 26138
rect 9502 26086 9514 26138
rect 9566 26086 9578 26138
rect 9630 26086 17694 26138
rect 17746 26086 17758 26138
rect 17810 26086 17822 26138
rect 17874 26086 17886 26138
rect 17938 26086 17950 26138
rect 18002 26086 26220 26138
rect 1104 26064 26220 26086
rect 1394 25984 1400 26036
rect 1452 26024 1458 26036
rect 2225 26027 2283 26033
rect 2225 26024 2237 26027
rect 1452 25996 2237 26024
rect 1452 25984 1458 25996
rect 2225 25993 2237 25996
rect 2271 25993 2283 26027
rect 2225 25987 2283 25993
rect 7098 25984 7104 26036
rect 7156 26024 7162 26036
rect 7745 26027 7803 26033
rect 7745 26024 7757 26027
rect 7156 25996 7757 26024
rect 7156 25984 7162 25996
rect 7745 25993 7757 25996
rect 7791 26024 7803 26027
rect 7834 26024 7840 26036
rect 7791 25996 7840 26024
rect 7791 25993 7803 25996
rect 7745 25987 7803 25993
rect 7834 25984 7840 25996
rect 7892 25984 7898 26036
rect 9674 26024 9680 26036
rect 9587 25996 9680 26024
rect 9674 25984 9680 25996
rect 9732 26024 9738 26036
rect 11238 26024 11244 26036
rect 9732 25996 11008 26024
rect 11199 25996 11244 26024
rect 9732 25984 9738 25996
rect 10980 25968 11008 25996
rect 11238 25984 11244 25996
rect 11296 26024 11302 26036
rect 11296 25996 11744 26024
rect 11296 25984 11302 25996
rect 8312 25928 9628 25956
rect 474 25848 480 25900
rect 532 25888 538 25900
rect 1578 25888 1584 25900
rect 532 25860 1584 25888
rect 532 25848 538 25860
rect 1578 25848 1584 25860
rect 1636 25888 1642 25900
rect 2041 25891 2099 25897
rect 2041 25888 2053 25891
rect 1636 25860 2053 25888
rect 1636 25848 1642 25860
rect 2041 25857 2053 25860
rect 2087 25857 2099 25891
rect 2041 25851 2099 25857
rect 3326 25848 3332 25900
rect 3384 25888 3390 25900
rect 4246 25888 4252 25900
rect 3384 25860 4252 25888
rect 3384 25848 3390 25860
rect 4246 25848 4252 25860
rect 4304 25888 4310 25900
rect 4341 25891 4399 25897
rect 4341 25888 4353 25891
rect 4304 25860 4353 25888
rect 4304 25848 4310 25860
rect 4341 25857 4353 25860
rect 4387 25857 4399 25891
rect 4341 25851 4399 25857
rect 5626 25848 5632 25900
rect 5684 25888 5690 25900
rect 6621 25891 6679 25897
rect 6621 25888 6633 25891
rect 5684 25860 6633 25888
rect 5684 25848 5690 25860
rect 6621 25857 6633 25860
rect 6667 25857 6679 25891
rect 8018 25888 8024 25900
rect 7979 25860 8024 25888
rect 6621 25851 6679 25857
rect 8018 25848 8024 25860
rect 8076 25848 8082 25900
rect 8312 25897 8340 25928
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25857 8355 25891
rect 8553 25891 8611 25897
rect 8553 25888 8565 25891
rect 8297 25851 8355 25857
rect 8404 25860 8565 25888
rect 5810 25780 5816 25832
rect 5868 25820 5874 25832
rect 6365 25823 6423 25829
rect 6365 25820 6377 25823
rect 5868 25792 6377 25820
rect 5868 25780 5874 25792
rect 6365 25789 6377 25792
rect 6411 25789 6423 25823
rect 8404 25820 8432 25860
rect 8553 25857 8565 25860
rect 8599 25857 8611 25891
rect 8553 25851 8611 25857
rect 9600 25832 9628 25928
rect 9950 25916 9956 25968
rect 10008 25956 10014 25968
rect 10106 25959 10164 25965
rect 10106 25956 10118 25959
rect 10008 25928 10118 25956
rect 10008 25916 10014 25928
rect 10106 25925 10118 25928
rect 10152 25925 10164 25959
rect 10106 25919 10164 25925
rect 10962 25916 10968 25968
rect 11020 25956 11026 25968
rect 11716 25965 11744 25996
rect 15010 25984 15016 26036
rect 15068 26024 15074 26036
rect 21266 26024 21272 26036
rect 15068 25996 21272 26024
rect 15068 25984 15074 25996
rect 21266 25984 21272 25996
rect 21324 25984 21330 26036
rect 11517 25959 11575 25965
rect 11517 25956 11529 25959
rect 11020 25928 11529 25956
rect 11020 25916 11026 25928
rect 11517 25925 11529 25928
rect 11563 25925 11575 25959
rect 11517 25919 11575 25925
rect 11701 25959 11759 25965
rect 11701 25925 11713 25959
rect 11747 25925 11759 25959
rect 11882 25956 11888 25968
rect 11843 25928 11888 25956
rect 11701 25919 11759 25925
rect 11882 25916 11888 25928
rect 11940 25916 11946 25968
rect 13998 25956 14004 25968
rect 12820 25928 14004 25956
rect 12820 25897 12848 25928
rect 13998 25916 14004 25928
rect 14056 25956 14062 25968
rect 14642 25965 14648 25968
rect 14636 25956 14648 25965
rect 14056 25928 14412 25956
rect 14603 25928 14648 25956
rect 14056 25916 14062 25928
rect 13078 25897 13084 25900
rect 12805 25891 12863 25897
rect 12805 25857 12817 25891
rect 12851 25857 12863 25891
rect 12805 25851 12863 25857
rect 13072 25851 13084 25897
rect 13136 25888 13142 25900
rect 14384 25897 14412 25928
rect 14636 25919 14648 25928
rect 14642 25916 14648 25919
rect 14700 25916 14706 25968
rect 16114 25916 16120 25968
rect 16172 25956 16178 25968
rect 17218 25956 17224 25968
rect 16172 25928 17224 25956
rect 16172 25916 16178 25928
rect 17218 25916 17224 25928
rect 17276 25916 17282 25968
rect 14369 25891 14427 25897
rect 13136 25860 13172 25888
rect 13078 25848 13084 25851
rect 13136 25848 13142 25860
rect 14369 25857 14381 25891
rect 14415 25857 14427 25891
rect 14369 25851 14427 25857
rect 16758 25848 16764 25900
rect 16816 25888 16822 25900
rect 16925 25891 16983 25897
rect 16925 25888 16937 25891
rect 16816 25860 16937 25888
rect 16816 25848 16822 25860
rect 16925 25857 16937 25860
rect 16971 25857 16983 25891
rect 23934 25888 23940 25900
rect 23895 25860 23940 25888
rect 16925 25851 16983 25857
rect 23934 25848 23940 25860
rect 23992 25848 23998 25900
rect 24946 25888 24952 25900
rect 24907 25860 24952 25888
rect 24946 25848 24952 25860
rect 25004 25848 25010 25900
rect 25225 25891 25283 25897
rect 25225 25857 25237 25891
rect 25271 25888 25283 25891
rect 26329 25891 26387 25897
rect 26329 25888 26341 25891
rect 25271 25860 26341 25888
rect 25271 25857 25283 25860
rect 25225 25851 25283 25857
rect 26329 25857 26341 25860
rect 26375 25857 26387 25891
rect 26329 25851 26387 25857
rect 6365 25783 6423 25789
rect 8220 25792 8432 25820
rect 8220 25761 8248 25792
rect 9582 25780 9588 25832
rect 9640 25820 9646 25832
rect 9861 25823 9919 25829
rect 9861 25820 9873 25823
rect 9640 25792 9873 25820
rect 9640 25780 9646 25792
rect 9861 25789 9873 25792
rect 9907 25789 9919 25823
rect 9861 25783 9919 25789
rect 12161 25823 12219 25829
rect 12161 25789 12173 25823
rect 12207 25820 12219 25823
rect 12434 25820 12440 25832
rect 12207 25792 12440 25820
rect 12207 25789 12219 25792
rect 12161 25783 12219 25789
rect 12434 25780 12440 25792
rect 12492 25780 12498 25832
rect 16666 25820 16672 25832
rect 16627 25792 16672 25820
rect 16666 25780 16672 25792
rect 16724 25780 16730 25832
rect 25501 25823 25559 25829
rect 25501 25789 25513 25823
rect 25547 25820 25559 25823
rect 26878 25820 26884 25832
rect 25547 25792 26884 25820
rect 25547 25789 25559 25792
rect 25501 25783 25559 25789
rect 26878 25780 26884 25792
rect 26936 25780 26942 25832
rect 8205 25755 8263 25761
rect 8205 25721 8217 25755
rect 8251 25721 8263 25755
rect 8205 25715 8263 25721
rect 12529 25755 12587 25761
rect 12529 25721 12541 25755
rect 12575 25752 12587 25755
rect 12575 25724 12848 25752
rect 12575 25721 12587 25724
rect 12529 25715 12587 25721
rect 12618 25684 12624 25696
rect 12579 25656 12624 25684
rect 12618 25644 12624 25656
rect 12676 25644 12682 25696
rect 12820 25684 12848 25724
rect 13170 25684 13176 25696
rect 12820 25656 13176 25684
rect 13170 25644 13176 25656
rect 13228 25644 13234 25696
rect 14185 25687 14243 25693
rect 14185 25653 14197 25687
rect 14231 25684 14243 25687
rect 14734 25684 14740 25696
rect 14231 25656 14740 25684
rect 14231 25653 14243 25656
rect 14185 25647 14243 25653
rect 14734 25644 14740 25656
rect 14792 25644 14798 25696
rect 15746 25684 15752 25696
rect 15707 25656 15752 25684
rect 15746 25644 15752 25656
rect 15804 25644 15810 25696
rect 18046 25684 18052 25696
rect 18007 25656 18052 25684
rect 18046 25644 18052 25656
rect 18104 25644 18110 25696
rect 1104 25594 26220 25616
rect 1104 25542 5136 25594
rect 5188 25542 5200 25594
rect 5252 25542 5264 25594
rect 5316 25542 5328 25594
rect 5380 25542 5392 25594
rect 5444 25542 13508 25594
rect 13560 25542 13572 25594
rect 13624 25542 13636 25594
rect 13688 25542 13700 25594
rect 13752 25542 13764 25594
rect 13816 25542 21880 25594
rect 21932 25542 21944 25594
rect 21996 25542 22008 25594
rect 22060 25542 22072 25594
rect 22124 25542 22136 25594
rect 22188 25542 26220 25594
rect 1104 25520 26220 25542
rect 7193 25483 7251 25489
rect 7193 25449 7205 25483
rect 7239 25480 7251 25483
rect 7282 25480 7288 25492
rect 7239 25452 7288 25480
rect 7239 25449 7251 25452
rect 7193 25443 7251 25449
rect 7282 25440 7288 25452
rect 7340 25440 7346 25492
rect 8018 25440 8024 25492
rect 8076 25480 8082 25492
rect 8297 25483 8355 25489
rect 8297 25480 8309 25483
rect 8076 25452 8309 25480
rect 8076 25440 8082 25452
rect 8297 25449 8309 25452
rect 8343 25449 8355 25483
rect 8297 25443 8355 25449
rect 9401 25483 9459 25489
rect 9401 25449 9413 25483
rect 9447 25480 9459 25483
rect 9766 25480 9772 25492
rect 9447 25452 9772 25480
rect 9447 25449 9459 25452
rect 9401 25443 9459 25449
rect 9766 25440 9772 25452
rect 9824 25440 9830 25492
rect 10686 25480 10692 25492
rect 10647 25452 10692 25480
rect 10686 25440 10692 25452
rect 10744 25440 10750 25492
rect 11330 25480 11336 25492
rect 11291 25452 11336 25480
rect 11330 25440 11336 25452
rect 11388 25440 11394 25492
rect 13078 25480 13084 25492
rect 13039 25452 13084 25480
rect 13078 25440 13084 25452
rect 13136 25440 13142 25492
rect 13170 25440 13176 25492
rect 13228 25480 13234 25492
rect 13228 25452 13273 25480
rect 13228 25440 13234 25452
rect 13906 25440 13912 25492
rect 13964 25480 13970 25492
rect 14093 25483 14151 25489
rect 14093 25480 14105 25483
rect 13964 25452 14105 25480
rect 13964 25440 13970 25452
rect 14093 25449 14105 25452
rect 14139 25449 14151 25483
rect 14093 25443 14151 25449
rect 16669 25483 16727 25489
rect 16669 25449 16681 25483
rect 16715 25480 16727 25483
rect 16758 25480 16764 25492
rect 16715 25452 16764 25480
rect 16715 25449 16727 25452
rect 16669 25443 16727 25449
rect 16758 25440 16764 25452
rect 16816 25440 16822 25492
rect 17144 25452 19380 25480
rect 5626 25412 5632 25424
rect 5587 25384 5632 25412
rect 5626 25372 5632 25384
rect 5684 25372 5690 25424
rect 8478 25412 8484 25424
rect 8439 25384 8484 25412
rect 8478 25372 8484 25384
rect 8536 25372 8542 25424
rect 9214 25412 9220 25424
rect 9175 25384 9220 25412
rect 9214 25372 9220 25384
rect 9272 25372 9278 25424
rect 5810 25344 5816 25356
rect 5771 25316 5816 25344
rect 5810 25304 5816 25316
rect 5868 25304 5874 25356
rect 7190 25304 7196 25356
rect 7248 25344 7254 25356
rect 7837 25347 7895 25353
rect 7837 25344 7849 25347
rect 7248 25316 7849 25344
rect 7248 25304 7254 25316
rect 7837 25313 7849 25316
rect 7883 25313 7895 25347
rect 7837 25307 7895 25313
rect 8757 25347 8815 25353
rect 8757 25313 8769 25347
rect 8803 25344 8815 25347
rect 8941 25347 8999 25353
rect 8941 25344 8953 25347
rect 8803 25316 8953 25344
rect 8803 25313 8815 25316
rect 8757 25307 8815 25313
rect 8941 25313 8953 25316
rect 8987 25344 8999 25347
rect 9858 25344 9864 25356
rect 8987 25316 9864 25344
rect 8987 25313 8999 25316
rect 8941 25307 8999 25313
rect 9858 25304 9864 25316
rect 9916 25304 9922 25356
rect 10229 25347 10287 25353
rect 10229 25313 10241 25347
rect 10275 25344 10287 25347
rect 10704 25344 10732 25440
rect 11882 25344 11888 25356
rect 10275 25316 10732 25344
rect 11348 25316 11888 25344
rect 10275 25313 10287 25316
rect 10229 25307 10287 25313
rect 5445 25279 5503 25285
rect 5445 25245 5457 25279
rect 5491 25276 5503 25279
rect 5534 25276 5540 25288
rect 5491 25248 5540 25276
rect 5491 25245 5503 25248
rect 5445 25239 5503 25245
rect 5534 25236 5540 25248
rect 5592 25236 5598 25288
rect 5629 25279 5687 25285
rect 5629 25245 5641 25279
rect 5675 25276 5687 25279
rect 7469 25279 7527 25285
rect 7469 25276 7481 25279
rect 5675 25248 7481 25276
rect 5675 25245 5687 25248
rect 5629 25239 5687 25245
rect 7469 25245 7481 25248
rect 7515 25245 7527 25279
rect 7469 25239 7527 25245
rect 7653 25279 7711 25285
rect 7653 25245 7665 25279
rect 7699 25245 7711 25279
rect 7653 25239 7711 25245
rect 6080 25211 6138 25217
rect 6080 25177 6092 25211
rect 6126 25208 6138 25211
rect 6454 25208 6460 25220
rect 6126 25180 6460 25208
rect 6126 25177 6138 25180
rect 6080 25171 6138 25177
rect 6454 25168 6460 25180
rect 6512 25168 6518 25220
rect 7006 25168 7012 25220
rect 7064 25208 7070 25220
rect 7668 25208 7696 25239
rect 7742 25236 7748 25288
rect 7800 25276 7806 25288
rect 7926 25276 7932 25288
rect 7800 25248 7845 25276
rect 7887 25248 7932 25276
rect 7800 25236 7806 25248
rect 7926 25236 7932 25248
rect 7984 25236 7990 25288
rect 8110 25276 8116 25288
rect 8071 25248 8116 25276
rect 8110 25236 8116 25248
rect 8168 25236 8174 25288
rect 9766 25236 9772 25288
rect 9824 25276 9830 25288
rect 11348 25285 11376 25316
rect 11882 25304 11888 25316
rect 11940 25344 11946 25356
rect 12158 25344 12164 25356
rect 11940 25316 12164 25344
rect 11940 25304 11946 25316
rect 12158 25304 12164 25316
rect 12216 25304 12222 25356
rect 13817 25347 13875 25353
rect 13817 25313 13829 25347
rect 13863 25344 13875 25347
rect 14737 25347 14795 25353
rect 14737 25344 14749 25347
rect 13863 25316 14749 25344
rect 13863 25313 13875 25316
rect 13817 25307 13875 25313
rect 14737 25313 14749 25316
rect 14783 25313 14795 25347
rect 14918 25344 14924 25356
rect 14879 25316 14924 25344
rect 14737 25307 14795 25313
rect 10597 25279 10655 25285
rect 10597 25276 10609 25279
rect 9824 25248 10609 25276
rect 9824 25236 9830 25248
rect 10597 25245 10609 25248
rect 10643 25245 10655 25279
rect 10597 25239 10655 25245
rect 11333 25279 11391 25285
rect 11333 25245 11345 25279
rect 11379 25245 11391 25279
rect 11333 25239 11391 25245
rect 11422 25236 11428 25288
rect 11480 25276 11486 25288
rect 11480 25248 11525 25276
rect 11480 25236 11486 25248
rect 12618 25236 12624 25288
rect 12676 25276 12682 25288
rect 12897 25279 12955 25285
rect 12897 25276 12909 25279
rect 12676 25248 12909 25276
rect 12676 25236 12682 25248
rect 12897 25245 12909 25248
rect 12943 25245 12955 25279
rect 12897 25239 12955 25245
rect 13633 25279 13691 25285
rect 13633 25245 13645 25279
rect 13679 25276 13691 25279
rect 14090 25276 14096 25288
rect 13679 25248 14096 25276
rect 13679 25245 13691 25248
rect 13633 25239 13691 25245
rect 14090 25236 14096 25248
rect 14148 25236 14154 25288
rect 14752 25276 14780 25307
rect 14918 25304 14924 25316
rect 14976 25304 14982 25356
rect 15013 25347 15071 25353
rect 15013 25313 15025 25347
rect 15059 25344 15071 25347
rect 15194 25344 15200 25356
rect 15059 25316 15200 25344
rect 15059 25313 15071 25316
rect 15013 25307 15071 25313
rect 15194 25304 15200 25316
rect 15252 25344 15258 25356
rect 15746 25344 15752 25356
rect 15252 25316 15752 25344
rect 15252 25304 15258 25316
rect 15746 25304 15752 25316
rect 15804 25304 15810 25356
rect 16224 25316 16620 25344
rect 15380 25279 15438 25285
rect 14752 25248 15056 25276
rect 15028 25220 15056 25248
rect 15380 25245 15392 25279
rect 15426 25276 15438 25279
rect 15470 25276 15476 25288
rect 15426 25248 15476 25276
rect 15426 25245 15438 25248
rect 15380 25239 15438 25245
rect 15470 25236 15476 25248
rect 15528 25236 15534 25288
rect 16224 25285 16252 25316
rect 16209 25279 16267 25285
rect 16209 25245 16221 25279
rect 16255 25245 16267 25279
rect 16482 25276 16488 25288
rect 16443 25248 16488 25276
rect 16209 25239 16267 25245
rect 16482 25236 16488 25248
rect 16540 25236 16546 25288
rect 16592 25276 16620 25316
rect 16666 25304 16672 25356
rect 16724 25344 16730 25356
rect 17144 25344 17172 25452
rect 18138 25412 18144 25424
rect 16724 25316 17172 25344
rect 17236 25384 18144 25412
rect 16724 25304 16730 25316
rect 16850 25276 16856 25288
rect 16592 25248 16856 25276
rect 16850 25236 16856 25248
rect 16908 25236 16914 25288
rect 17003 25279 17061 25285
rect 17003 25245 17015 25279
rect 17049 25276 17061 25279
rect 17236 25276 17264 25384
rect 18138 25372 18144 25384
rect 18196 25372 18202 25424
rect 19352 25356 19380 25452
rect 19334 25344 19340 25356
rect 19247 25316 19340 25344
rect 19334 25304 19340 25316
rect 19392 25304 19398 25356
rect 17049 25248 17264 25276
rect 17313 25279 17371 25285
rect 17049 25245 17061 25248
rect 17003 25239 17061 25245
rect 17313 25245 17325 25279
rect 17359 25245 17371 25279
rect 17313 25239 17371 25245
rect 17405 25279 17463 25285
rect 17405 25245 17417 25279
rect 17451 25276 17463 25279
rect 17494 25276 17500 25288
rect 17451 25248 17500 25276
rect 17451 25245 17463 25248
rect 17405 25239 17463 25245
rect 7064 25180 7696 25208
rect 7064 25168 7070 25180
rect 9214 25168 9220 25220
rect 9272 25208 9278 25220
rect 10045 25211 10103 25217
rect 9272 25180 9628 25208
rect 9272 25168 9278 25180
rect 9600 25149 9628 25180
rect 10045 25177 10057 25211
rect 10091 25208 10103 25211
rect 11514 25208 11520 25220
rect 10091 25180 11520 25208
rect 10091 25177 10103 25180
rect 10045 25171 10103 25177
rect 11514 25168 11520 25180
rect 11572 25168 11578 25220
rect 14461 25211 14519 25217
rect 14461 25177 14473 25211
rect 14507 25208 14519 25211
rect 14734 25208 14740 25220
rect 14507 25180 14740 25208
rect 14507 25177 14519 25180
rect 14461 25171 14519 25177
rect 14734 25168 14740 25180
rect 14792 25168 14798 25220
rect 15010 25168 15016 25220
rect 15068 25208 15074 25220
rect 15657 25211 15715 25217
rect 15657 25208 15669 25211
rect 15068 25180 15669 25208
rect 15068 25168 15074 25180
rect 15657 25177 15669 25180
rect 15703 25177 15715 25211
rect 16758 25208 16764 25220
rect 16719 25180 16764 25208
rect 15657 25171 15715 25177
rect 16758 25168 16764 25180
rect 16816 25168 16822 25220
rect 17328 25208 17356 25239
rect 17494 25236 17500 25248
rect 17552 25236 17558 25288
rect 17586 25236 17592 25288
rect 17644 25276 17650 25288
rect 17682 25279 17740 25285
rect 17682 25276 17694 25279
rect 17644 25248 17694 25276
rect 17644 25236 17650 25248
rect 17682 25245 17694 25248
rect 17728 25245 17740 25279
rect 18046 25276 18052 25288
rect 18007 25248 18052 25276
rect 17682 25239 17740 25245
rect 18046 25236 18052 25248
rect 18104 25236 18110 25288
rect 18138 25236 18144 25288
rect 18196 25276 18202 25288
rect 18598 25276 18604 25288
rect 18196 25248 18604 25276
rect 18196 25236 18202 25248
rect 18598 25236 18604 25248
rect 18656 25236 18662 25288
rect 19604 25211 19662 25217
rect 17328 25180 18184 25208
rect 18156 25152 18184 25180
rect 19604 25177 19616 25211
rect 19650 25208 19662 25211
rect 19702 25208 19708 25220
rect 19650 25180 19708 25208
rect 19650 25177 19662 25180
rect 19604 25171 19662 25177
rect 19702 25168 19708 25180
rect 19760 25168 19766 25220
rect 9585 25143 9643 25149
rect 9585 25109 9597 25143
rect 9631 25109 9643 25143
rect 9950 25140 9956 25152
rect 9911 25112 9956 25140
rect 9585 25103 9643 25109
rect 9950 25100 9956 25112
rect 10008 25100 10014 25152
rect 10410 25140 10416 25152
rect 10371 25112 10416 25140
rect 10410 25100 10416 25112
rect 10468 25100 10474 25152
rect 11698 25140 11704 25152
rect 11659 25112 11704 25140
rect 11698 25100 11704 25112
rect 11756 25100 11762 25152
rect 13170 25100 13176 25152
rect 13228 25140 13234 25152
rect 13541 25143 13599 25149
rect 13541 25140 13553 25143
rect 13228 25112 13553 25140
rect 13228 25100 13234 25112
rect 13541 25109 13553 25112
rect 13587 25109 13599 25143
rect 13541 25103 13599 25109
rect 14553 25143 14611 25149
rect 14553 25109 14565 25143
rect 14599 25140 14611 25143
rect 15473 25143 15531 25149
rect 15473 25140 15485 25143
rect 14599 25112 15485 25140
rect 14599 25109 14611 25112
rect 14553 25103 14611 25109
rect 15473 25109 15485 25112
rect 15519 25109 15531 25143
rect 15473 25103 15531 25109
rect 16393 25143 16451 25149
rect 16393 25109 16405 25143
rect 16439 25140 16451 25143
rect 16574 25140 16580 25152
rect 16439 25112 16580 25140
rect 16439 25109 16451 25112
rect 16393 25103 16451 25109
rect 16574 25100 16580 25112
rect 16632 25100 16638 25152
rect 17402 25100 17408 25152
rect 17460 25140 17466 25152
rect 17589 25143 17647 25149
rect 17589 25140 17601 25143
rect 17460 25112 17601 25140
rect 17460 25100 17466 25112
rect 17589 25109 17601 25112
rect 17635 25109 17647 25143
rect 17589 25103 17647 25109
rect 18138 25100 18144 25152
rect 18196 25100 18202 25152
rect 20714 25140 20720 25152
rect 20675 25112 20720 25140
rect 20714 25100 20720 25112
rect 20772 25100 20778 25152
rect 1104 25050 26220 25072
rect 1104 24998 9322 25050
rect 9374 24998 9386 25050
rect 9438 24998 9450 25050
rect 9502 24998 9514 25050
rect 9566 24998 9578 25050
rect 9630 24998 17694 25050
rect 17746 24998 17758 25050
rect 17810 24998 17822 25050
rect 17874 24998 17886 25050
rect 17938 24998 17950 25050
rect 18002 24998 26220 25050
rect 1104 24976 26220 24998
rect 6454 24936 6460 24948
rect 6415 24908 6460 24936
rect 6454 24896 6460 24908
rect 6512 24896 6518 24948
rect 7929 24939 7987 24945
rect 6748 24908 7604 24936
rect 6748 24868 6776 24908
rect 7190 24868 7196 24880
rect 6564 24840 6776 24868
rect 6181 24803 6239 24809
rect 6181 24769 6193 24803
rect 6227 24800 6239 24803
rect 6564 24800 6592 24840
rect 6748 24809 6776 24840
rect 6840 24840 7196 24868
rect 6840 24809 6868 24840
rect 7190 24828 7196 24840
rect 7248 24828 7254 24880
rect 6227 24772 6592 24800
rect 6641 24803 6699 24809
rect 6227 24769 6239 24772
rect 6181 24763 6239 24769
rect 6641 24769 6653 24803
rect 6687 24769 6699 24803
rect 6641 24763 6699 24769
rect 6733 24803 6791 24809
rect 6733 24769 6745 24803
rect 6779 24769 6791 24803
rect 6733 24763 6791 24769
rect 6825 24803 6883 24809
rect 6825 24769 6837 24803
rect 6871 24769 6883 24803
rect 6825 24763 6883 24769
rect 6656 24732 6684 24763
rect 6914 24760 6920 24812
rect 6972 24800 6978 24812
rect 7576 24809 7604 24908
rect 7929 24905 7941 24939
rect 7975 24936 7987 24939
rect 8110 24936 8116 24948
rect 7975 24908 8116 24936
rect 7975 24905 7987 24908
rect 7929 24899 7987 24905
rect 8110 24896 8116 24908
rect 8168 24896 8174 24948
rect 8478 24896 8484 24948
rect 8536 24936 8542 24948
rect 8941 24939 8999 24945
rect 8941 24936 8953 24939
rect 8536 24908 8953 24936
rect 8536 24896 8542 24908
rect 8941 24905 8953 24908
rect 8987 24905 8999 24939
rect 8941 24899 8999 24905
rect 11241 24939 11299 24945
rect 11241 24905 11253 24939
rect 11287 24936 11299 24939
rect 11330 24936 11336 24948
rect 11287 24908 11336 24936
rect 11287 24905 11299 24908
rect 11241 24899 11299 24905
rect 11330 24896 11336 24908
rect 11388 24936 11394 24948
rect 11388 24908 12112 24936
rect 11388 24896 11394 24908
rect 9306 24868 9312 24880
rect 9267 24840 9312 24868
rect 9306 24828 9312 24840
rect 9364 24868 9370 24880
rect 9950 24868 9956 24880
rect 9364 24840 9956 24868
rect 9364 24828 9370 24840
rect 9950 24828 9956 24840
rect 10008 24828 10014 24880
rect 10128 24871 10186 24877
rect 10128 24837 10140 24871
rect 10174 24868 10186 24871
rect 10410 24868 10416 24880
rect 10174 24840 10416 24868
rect 10174 24837 10186 24840
rect 10128 24831 10186 24837
rect 10410 24828 10416 24840
rect 10468 24828 10474 24880
rect 12084 24868 12112 24908
rect 14274 24896 14280 24948
rect 14332 24936 14338 24948
rect 14918 24936 14924 24948
rect 14332 24908 14924 24936
rect 14332 24896 14338 24908
rect 14918 24896 14924 24908
rect 14976 24896 14982 24948
rect 15470 24936 15476 24948
rect 15431 24908 15476 24936
rect 15470 24896 15476 24908
rect 15528 24896 15534 24948
rect 16025 24939 16083 24945
rect 16025 24905 16037 24939
rect 16071 24936 16083 24939
rect 16482 24936 16488 24948
rect 16071 24908 16488 24936
rect 16071 24905 16083 24908
rect 16025 24899 16083 24905
rect 16482 24896 16488 24908
rect 16540 24896 16546 24948
rect 18049 24939 18107 24945
rect 18049 24905 18061 24939
rect 18095 24936 18107 24939
rect 18138 24936 18144 24948
rect 18095 24908 18144 24936
rect 18095 24905 18107 24908
rect 18049 24899 18107 24905
rect 18138 24896 18144 24908
rect 18196 24896 18202 24948
rect 19702 24936 19708 24948
rect 19663 24908 19708 24936
rect 19702 24896 19708 24908
rect 19760 24896 19766 24948
rect 20272 24908 20852 24936
rect 12437 24871 12495 24877
rect 12437 24868 12449 24871
rect 12084 24840 12449 24868
rect 7101 24803 7159 24809
rect 6972 24772 7017 24800
rect 6972 24760 6978 24772
rect 7101 24769 7113 24803
rect 7147 24800 7159 24803
rect 7285 24803 7343 24809
rect 7285 24800 7297 24803
rect 7147 24772 7297 24800
rect 7147 24769 7159 24772
rect 7101 24763 7159 24769
rect 7285 24769 7297 24772
rect 7331 24769 7343 24803
rect 7285 24763 7343 24769
rect 7561 24803 7619 24809
rect 7561 24769 7573 24803
rect 7607 24769 7619 24803
rect 7834 24800 7840 24812
rect 7795 24772 7840 24800
rect 7561 24763 7619 24769
rect 7006 24732 7012 24744
rect 6656 24704 7012 24732
rect 7006 24692 7012 24704
rect 7064 24692 7070 24744
rect 7377 24735 7435 24741
rect 7377 24701 7389 24735
rect 7423 24701 7435 24735
rect 7576 24732 7604 24763
rect 7834 24760 7840 24772
rect 7892 24760 7898 24812
rect 8849 24803 8907 24809
rect 8849 24769 8861 24803
rect 8895 24800 8907 24803
rect 10686 24800 10692 24812
rect 8895 24772 10692 24800
rect 8895 24769 8907 24772
rect 8849 24763 8907 24769
rect 7742 24732 7748 24744
rect 7576 24704 7748 24732
rect 7377 24695 7435 24701
rect 7024 24664 7052 24692
rect 7392 24664 7420 24695
rect 7742 24692 7748 24704
rect 7800 24692 7806 24744
rect 9122 24692 9128 24744
rect 9180 24732 9186 24744
rect 9508 24741 9536 24772
rect 10686 24760 10692 24772
rect 10744 24760 10750 24812
rect 11514 24800 11520 24812
rect 11475 24772 11520 24800
rect 11514 24760 11520 24772
rect 11572 24760 11578 24812
rect 12084 24809 12112 24840
rect 12437 24837 12449 24840
rect 12483 24837 12495 24871
rect 12437 24831 12495 24837
rect 14292 24840 14596 24868
rect 11759 24803 11817 24809
rect 11759 24769 11771 24803
rect 11805 24800 11817 24803
rect 12069 24803 12127 24809
rect 11805 24772 12020 24800
rect 11805 24769 11817 24772
rect 11759 24763 11817 24769
rect 9401 24735 9459 24741
rect 9401 24732 9413 24735
rect 9180 24704 9413 24732
rect 9180 24692 9186 24704
rect 9401 24701 9413 24704
rect 9447 24701 9459 24735
rect 9401 24695 9459 24701
rect 9493 24735 9551 24741
rect 9493 24701 9505 24735
rect 9539 24701 9551 24735
rect 9493 24695 9551 24701
rect 9582 24692 9588 24744
rect 9640 24732 9646 24744
rect 9861 24735 9919 24741
rect 9861 24732 9873 24735
rect 9640 24704 9873 24732
rect 9640 24692 9646 24704
rect 9861 24701 9873 24704
rect 9907 24701 9919 24735
rect 9861 24695 9919 24701
rect 7024 24636 7420 24664
rect 11992 24664 12020 24772
rect 12069 24769 12081 24803
rect 12115 24769 12127 24803
rect 12069 24763 12127 24769
rect 12158 24760 12164 24812
rect 12216 24800 12222 24812
rect 12253 24803 12311 24809
rect 12253 24800 12265 24803
rect 12216 24772 12265 24800
rect 12216 24760 12222 24772
rect 12253 24769 12265 24772
rect 12299 24769 12311 24803
rect 12253 24763 12311 24769
rect 13817 24803 13875 24809
rect 13817 24769 13829 24803
rect 13863 24769 13875 24803
rect 13817 24763 13875 24769
rect 13832 24732 13860 24763
rect 13906 24760 13912 24812
rect 13964 24800 13970 24812
rect 14001 24803 14059 24809
rect 14001 24800 14013 24803
rect 13964 24772 14013 24800
rect 13964 24760 13970 24772
rect 14001 24769 14013 24772
rect 14047 24769 14059 24803
rect 14001 24763 14059 24769
rect 14185 24803 14243 24809
rect 14185 24769 14197 24803
rect 14231 24800 14243 24803
rect 14292 24800 14320 24840
rect 14461 24803 14519 24809
rect 14461 24800 14473 24803
rect 14231 24772 14320 24800
rect 14384 24772 14473 24800
rect 14231 24769 14243 24772
rect 14185 24763 14243 24769
rect 14090 24732 14096 24744
rect 13832 24704 14096 24732
rect 12342 24664 12348 24676
rect 11992 24636 12348 24664
rect 12342 24624 12348 24636
rect 12400 24664 12406 24676
rect 12621 24667 12679 24673
rect 12621 24664 12633 24667
rect 12400 24636 12633 24664
rect 12400 24624 12406 24636
rect 12621 24633 12633 24636
rect 12667 24633 12679 24667
rect 12621 24627 12679 24633
rect 5626 24556 5632 24608
rect 5684 24596 5690 24608
rect 5813 24599 5871 24605
rect 5813 24596 5825 24599
rect 5684 24568 5825 24596
rect 5684 24556 5690 24568
rect 5813 24565 5825 24568
rect 5859 24565 5871 24599
rect 5813 24559 5871 24565
rect 6089 24599 6147 24605
rect 6089 24565 6101 24599
rect 6135 24596 6147 24599
rect 7098 24596 7104 24608
rect 6135 24568 7104 24596
rect 6135 24565 6147 24568
rect 6089 24559 6147 24565
rect 7098 24556 7104 24568
rect 7156 24596 7162 24608
rect 7926 24596 7932 24608
rect 7156 24568 7932 24596
rect 7156 24556 7162 24568
rect 7926 24556 7932 24568
rect 7984 24556 7990 24608
rect 8018 24556 8024 24608
rect 8076 24596 8082 24608
rect 8113 24599 8171 24605
rect 8113 24596 8125 24599
rect 8076 24568 8125 24596
rect 8076 24556 8082 24568
rect 8113 24565 8125 24568
rect 8159 24565 8171 24599
rect 8113 24559 8171 24565
rect 11698 24556 11704 24608
rect 11756 24596 11762 24608
rect 13832 24596 13860 24704
rect 14090 24692 14096 24704
rect 14148 24732 14154 24744
rect 14384 24732 14412 24772
rect 14461 24769 14473 24772
rect 14507 24769 14519 24803
rect 14568 24800 14596 24840
rect 14752 24840 15240 24868
rect 14752 24809 14780 24840
rect 15212 24812 15240 24840
rect 16574 24828 16580 24880
rect 16632 24868 16638 24880
rect 18156 24868 18184 24896
rect 18598 24868 18604 24880
rect 16632 24840 16804 24868
rect 18156 24840 18460 24868
rect 18559 24840 18604 24868
rect 16632 24828 16638 24840
rect 14737 24803 14795 24809
rect 14568 24772 14688 24800
rect 14461 24763 14519 24769
rect 14660 24744 14688 24772
rect 14737 24769 14749 24803
rect 14783 24769 14795 24803
rect 15102 24800 15108 24812
rect 15063 24772 15108 24800
rect 14737 24763 14795 24769
rect 15102 24760 15108 24772
rect 15160 24760 15166 24812
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 16666 24800 16672 24812
rect 15252 24772 15297 24800
rect 16627 24772 16672 24800
rect 15252 24760 15258 24772
rect 16666 24760 16672 24772
rect 16724 24760 16730 24812
rect 16776 24800 16804 24840
rect 16925 24803 16983 24809
rect 16925 24800 16937 24803
rect 16776 24772 16937 24800
rect 16925 24769 16937 24772
rect 16971 24769 16983 24803
rect 16925 24763 16983 24769
rect 17310 24760 17316 24812
rect 17368 24800 17374 24812
rect 17494 24800 17500 24812
rect 17368 24772 17500 24800
rect 17368 24760 17374 24772
rect 17494 24760 17500 24772
rect 17552 24800 17558 24812
rect 18432 24809 18460 24840
rect 18598 24828 18604 24840
rect 18656 24828 18662 24880
rect 18233 24803 18291 24809
rect 18233 24800 18245 24803
rect 17552 24772 18245 24800
rect 17552 24760 17558 24772
rect 18233 24769 18245 24772
rect 18279 24769 18291 24803
rect 18233 24763 18291 24769
rect 18417 24803 18475 24809
rect 18417 24769 18429 24803
rect 18463 24769 18475 24803
rect 19521 24803 19579 24809
rect 19521 24800 19533 24803
rect 18417 24763 18475 24769
rect 19352 24772 19533 24800
rect 14550 24732 14556 24744
rect 14148 24704 14412 24732
rect 14511 24704 14556 24732
rect 14148 24692 14154 24704
rect 14550 24692 14556 24704
rect 14608 24692 14614 24744
rect 14642 24692 14648 24744
rect 14700 24732 14706 24744
rect 15120 24732 15148 24760
rect 14700 24704 15148 24732
rect 16485 24735 16543 24741
rect 14700 24692 14706 24704
rect 16485 24701 16497 24735
rect 16531 24732 16543 24735
rect 16574 24732 16580 24744
rect 16531 24704 16580 24732
rect 16531 24701 16543 24704
rect 16485 24695 16543 24701
rect 16574 24692 16580 24704
rect 16632 24692 16638 24744
rect 18506 24692 18512 24744
rect 18564 24732 18570 24744
rect 18877 24735 18935 24741
rect 18877 24732 18889 24735
rect 18564 24704 18889 24732
rect 18564 24692 18570 24704
rect 18877 24701 18889 24704
rect 18923 24701 18935 24735
rect 18877 24695 18935 24701
rect 14921 24667 14979 24673
rect 14921 24633 14933 24667
rect 14967 24664 14979 24667
rect 16206 24664 16212 24676
rect 14967 24636 16068 24664
rect 16167 24636 16212 24664
rect 14967 24633 14979 24636
rect 14921 24627 14979 24633
rect 14366 24596 14372 24608
rect 11756 24568 13860 24596
rect 14327 24568 14372 24596
rect 11756 24556 11762 24568
rect 14366 24556 14372 24568
rect 14424 24556 14430 24608
rect 14737 24599 14795 24605
rect 14737 24565 14749 24599
rect 14783 24596 14795 24599
rect 14826 24596 14832 24608
rect 14783 24568 14832 24596
rect 14783 24565 14795 24568
rect 14737 24559 14795 24565
rect 14826 24556 14832 24568
rect 14884 24556 14890 24608
rect 14936 24596 14964 24627
rect 15010 24596 15016 24608
rect 14936 24568 15016 24596
rect 15010 24556 15016 24568
rect 15068 24556 15074 24608
rect 15194 24556 15200 24608
rect 15252 24596 15258 24608
rect 16040 24596 16068 24636
rect 16206 24624 16212 24636
rect 16264 24624 16270 24676
rect 19242 24664 19248 24676
rect 19203 24636 19248 24664
rect 19242 24624 19248 24636
rect 19300 24624 19306 24676
rect 19352 24673 19380 24772
rect 19521 24769 19533 24772
rect 19567 24769 19579 24803
rect 19521 24763 19579 24769
rect 20039 24803 20097 24809
rect 20039 24769 20051 24803
rect 20085 24800 20097 24803
rect 20272 24800 20300 24908
rect 20714 24868 20720 24880
rect 20456 24840 20720 24868
rect 20085 24772 20300 24800
rect 20349 24803 20407 24809
rect 20085 24769 20097 24772
rect 20039 24763 20097 24769
rect 20349 24769 20361 24803
rect 20395 24800 20407 24803
rect 20456 24800 20484 24840
rect 20714 24828 20720 24840
rect 20772 24828 20778 24880
rect 20395 24772 20484 24800
rect 20533 24803 20591 24809
rect 20395 24769 20407 24772
rect 20349 24763 20407 24769
rect 20533 24769 20545 24803
rect 20579 24769 20591 24803
rect 20824 24800 20852 24908
rect 20901 24803 20959 24809
rect 20901 24800 20913 24803
rect 20824 24772 20913 24800
rect 20533 24763 20591 24769
rect 20901 24769 20913 24772
rect 20947 24800 20959 24803
rect 21174 24800 21180 24812
rect 20947 24772 21180 24800
rect 20947 24769 20959 24772
rect 20901 24763 20959 24769
rect 20441 24735 20499 24741
rect 20441 24732 20453 24735
rect 20364 24704 20453 24732
rect 19337 24667 19395 24673
rect 19337 24633 19349 24667
rect 19383 24633 19395 24667
rect 20364 24664 20392 24704
rect 20441 24701 20453 24704
rect 20487 24732 20499 24735
rect 20548 24732 20576 24763
rect 21174 24760 21180 24772
rect 21232 24760 21238 24812
rect 20487 24704 20576 24732
rect 20487 24701 20499 24704
rect 20441 24695 20499 24701
rect 19337 24627 19395 24633
rect 19628 24636 20392 24664
rect 17310 24596 17316 24608
rect 15252 24568 15297 24596
rect 16040 24568 17316 24596
rect 15252 24556 15258 24568
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 17586 24556 17592 24608
rect 17644 24596 17650 24608
rect 19628 24596 19656 24636
rect 17644 24568 19656 24596
rect 17644 24556 17650 24568
rect 19702 24556 19708 24608
rect 19760 24596 19766 24608
rect 19889 24599 19947 24605
rect 19889 24596 19901 24599
rect 19760 24568 19901 24596
rect 19760 24556 19766 24568
rect 19889 24565 19901 24568
rect 19935 24565 19947 24599
rect 19889 24559 19947 24565
rect 26326 24528 26332 24540
rect 1104 24506 26220 24528
rect 1104 24454 5136 24506
rect 5188 24454 5200 24506
rect 5252 24454 5264 24506
rect 5316 24454 5328 24506
rect 5380 24454 5392 24506
rect 5444 24454 13508 24506
rect 13560 24454 13572 24506
rect 13624 24454 13636 24506
rect 13688 24454 13700 24506
rect 13752 24454 13764 24506
rect 13816 24454 21880 24506
rect 21932 24454 21944 24506
rect 21996 24454 22008 24506
rect 22060 24454 22072 24506
rect 22124 24454 22136 24506
rect 22188 24454 26220 24506
rect 26287 24500 26332 24528
rect 26326 24488 26332 24500
rect 26384 24488 26390 24540
rect 1104 24432 26220 24454
rect 5534 24352 5540 24404
rect 5592 24392 5598 24404
rect 7466 24392 7472 24404
rect 5592 24364 7328 24392
rect 7379 24364 7472 24392
rect 5592 24352 5598 24364
rect 6825 24327 6883 24333
rect 6825 24293 6837 24327
rect 6871 24324 6883 24327
rect 7006 24324 7012 24336
rect 6871 24296 7012 24324
rect 6871 24293 6883 24296
rect 6825 24287 6883 24293
rect 7006 24284 7012 24296
rect 7064 24284 7070 24336
rect 7300 24324 7328 24364
rect 7466 24352 7472 24364
rect 7524 24392 7530 24404
rect 7834 24392 7840 24404
rect 7524 24364 7840 24392
rect 7524 24352 7530 24364
rect 7834 24352 7840 24364
rect 7892 24352 7898 24404
rect 9214 24352 9220 24404
rect 9272 24392 9278 24404
rect 9677 24395 9735 24401
rect 9272 24364 9536 24392
rect 9272 24352 9278 24364
rect 7745 24327 7803 24333
rect 7745 24324 7757 24327
rect 7300 24296 7757 24324
rect 7745 24293 7757 24296
rect 7791 24324 7803 24327
rect 9306 24324 9312 24336
rect 7791 24296 9312 24324
rect 7791 24293 7803 24296
rect 7745 24287 7803 24293
rect 9306 24284 9312 24296
rect 9364 24284 9370 24336
rect 9508 24333 9536 24364
rect 9677 24361 9689 24395
rect 9723 24392 9735 24395
rect 9766 24392 9772 24404
rect 9723 24364 9772 24392
rect 9723 24361 9735 24364
rect 9677 24355 9735 24361
rect 9766 24352 9772 24364
rect 9824 24352 9830 24404
rect 11422 24352 11428 24404
rect 11480 24392 11486 24404
rect 11517 24395 11575 24401
rect 11517 24392 11529 24395
rect 11480 24364 11529 24392
rect 11480 24352 11486 24364
rect 11517 24361 11529 24364
rect 11563 24361 11575 24395
rect 11517 24355 11575 24361
rect 13633 24395 13691 24401
rect 13633 24361 13645 24395
rect 13679 24392 13691 24395
rect 14550 24392 14556 24404
rect 13679 24364 14556 24392
rect 13679 24361 13691 24364
rect 13633 24355 13691 24361
rect 9493 24327 9551 24333
rect 9493 24293 9505 24327
rect 9539 24293 9551 24327
rect 9493 24287 9551 24293
rect 6641 24259 6699 24265
rect 6641 24225 6653 24259
rect 6687 24256 6699 24259
rect 7098 24256 7104 24268
rect 6687 24228 7104 24256
rect 6687 24225 6699 24228
rect 6641 24219 6699 24225
rect 7098 24216 7104 24228
rect 7156 24216 7162 24268
rect 7190 24216 7196 24268
rect 7248 24256 7254 24268
rect 8018 24256 8024 24268
rect 7248 24228 8024 24256
rect 7248 24216 7254 24228
rect 8018 24216 8024 24228
rect 8076 24216 8082 24268
rect 9214 24216 9220 24268
rect 9272 24256 9278 24268
rect 9582 24256 9588 24268
rect 9272 24228 9588 24256
rect 9272 24216 9278 24228
rect 9582 24216 9588 24228
rect 9640 24256 9646 24268
rect 10137 24259 10195 24265
rect 10137 24256 10149 24259
rect 9640 24228 10149 24256
rect 9640 24216 9646 24228
rect 10137 24225 10149 24228
rect 10183 24225 10195 24259
rect 11532 24256 11560 24355
rect 14550 24352 14556 24364
rect 14608 24352 14614 24404
rect 14826 24352 14832 24404
rect 14884 24392 14890 24404
rect 15194 24392 15200 24404
rect 14884 24364 15200 24392
rect 14884 24352 14890 24364
rect 15194 24352 15200 24364
rect 15252 24352 15258 24404
rect 16206 24352 16212 24404
rect 16264 24392 16270 24404
rect 16945 24395 17003 24401
rect 16945 24392 16957 24395
rect 16264 24364 16957 24392
rect 16264 24352 16270 24364
rect 16945 24361 16957 24364
rect 16991 24361 17003 24395
rect 18325 24395 18383 24401
rect 18325 24392 18337 24395
rect 16945 24355 17003 24361
rect 17512 24364 18337 24392
rect 12618 24324 12624 24336
rect 12579 24296 12624 24324
rect 12618 24284 12624 24296
rect 12676 24284 12682 24336
rect 14366 24284 14372 24336
rect 14424 24324 14430 24336
rect 15102 24324 15108 24336
rect 14424 24296 15108 24324
rect 14424 24284 14430 24296
rect 15102 24284 15108 24296
rect 15160 24324 15166 24336
rect 17512 24324 17540 24364
rect 18325 24361 18337 24364
rect 18371 24392 18383 24395
rect 19426 24392 19432 24404
rect 18371 24364 19432 24392
rect 18371 24361 18383 24364
rect 18325 24355 18383 24361
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 15160 24296 17540 24324
rect 15160 24284 15166 24296
rect 12342 24256 12348 24268
rect 11532 24228 12020 24256
rect 12303 24228 12348 24256
rect 10137 24219 10195 24225
rect 3789 24191 3847 24197
rect 3789 24157 3801 24191
rect 3835 24188 3847 24191
rect 5718 24188 5724 24200
rect 3835 24160 5724 24188
rect 3835 24157 3847 24160
rect 3789 24151 3847 24157
rect 5718 24148 5724 24160
rect 5776 24148 5782 24200
rect 5813 24191 5871 24197
rect 5813 24157 5825 24191
rect 5859 24157 5871 24191
rect 5994 24188 6000 24200
rect 5955 24160 6000 24188
rect 5813 24151 5871 24157
rect 4062 24129 4068 24132
rect 4056 24083 4068 24129
rect 4120 24120 4126 24132
rect 5828 24120 5856 24151
rect 5994 24148 6000 24160
rect 6052 24148 6058 24200
rect 6089 24191 6147 24197
rect 6089 24157 6101 24191
rect 6135 24188 6147 24191
rect 6457 24191 6515 24197
rect 6457 24188 6469 24191
rect 6135 24160 6469 24188
rect 6135 24157 6147 24160
rect 6089 24151 6147 24157
rect 6457 24157 6469 24160
rect 6503 24157 6515 24191
rect 6457 24151 6515 24157
rect 6917 24191 6975 24197
rect 6917 24157 6929 24191
rect 6963 24188 6975 24191
rect 7282 24188 7288 24200
rect 6963 24160 7288 24188
rect 6963 24157 6975 24160
rect 6917 24151 6975 24157
rect 7282 24148 7288 24160
rect 7340 24148 7346 24200
rect 7374 24148 7380 24200
rect 7432 24188 7438 24200
rect 7469 24191 7527 24197
rect 7469 24188 7481 24191
rect 7432 24160 7481 24188
rect 7432 24148 7438 24160
rect 7469 24157 7481 24160
rect 7515 24157 7527 24191
rect 7469 24151 7527 24157
rect 7558 24148 7564 24200
rect 7616 24188 7622 24200
rect 7616 24160 7661 24188
rect 7616 24148 7622 24160
rect 9766 24148 9772 24200
rect 9824 24188 9830 24200
rect 9861 24191 9919 24197
rect 9861 24188 9873 24191
rect 9824 24160 9873 24188
rect 9824 24148 9830 24160
rect 9861 24157 9873 24160
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 11698 24148 11704 24200
rect 11756 24188 11762 24200
rect 11886 24191 11944 24197
rect 11886 24188 11898 24191
rect 11756 24160 11898 24188
rect 11756 24148 11762 24160
rect 11886 24157 11898 24160
rect 11932 24157 11944 24191
rect 11992 24188 12020 24228
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 15470 24256 15476 24268
rect 13740 24228 15240 24256
rect 15431 24228 15476 24256
rect 13740 24197 13768 24228
rect 12253 24191 12311 24197
rect 12253 24188 12265 24191
rect 11992 24160 12265 24188
rect 11886 24151 11944 24157
rect 12253 24157 12265 24160
rect 12299 24157 12311 24191
rect 12253 24151 12311 24157
rect 13725 24191 13783 24197
rect 13725 24157 13737 24191
rect 13771 24157 13783 24191
rect 14090 24188 14096 24200
rect 14051 24160 14096 24188
rect 13725 24151 13783 24157
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 14185 24191 14243 24197
rect 14185 24157 14197 24191
rect 14231 24157 14243 24191
rect 14185 24151 14243 24157
rect 14552 24191 14610 24197
rect 14552 24157 14564 24191
rect 14598 24188 14610 24191
rect 14642 24188 14648 24200
rect 14598 24160 14648 24188
rect 14598 24157 14610 24160
rect 14552 24151 14610 24157
rect 7650 24120 7656 24132
rect 4120 24092 4156 24120
rect 5828 24092 7656 24120
rect 4062 24080 4068 24083
rect 4120 24080 4126 24092
rect 7650 24080 7656 24092
rect 7708 24080 7714 24132
rect 9217 24123 9275 24129
rect 9217 24089 9229 24123
rect 9263 24120 9275 24123
rect 9674 24120 9680 24132
rect 9263 24092 9680 24120
rect 9263 24089 9275 24092
rect 9217 24083 9275 24089
rect 9674 24080 9680 24092
rect 9732 24080 9738 24132
rect 10382 24123 10440 24129
rect 10382 24120 10394 24123
rect 10060 24092 10394 24120
rect 4246 24012 4252 24064
rect 4304 24052 4310 24064
rect 5169 24055 5227 24061
rect 5169 24052 5181 24055
rect 4304 24024 5181 24052
rect 4304 24012 4310 24024
rect 5169 24021 5181 24024
rect 5215 24021 5227 24055
rect 5169 24015 5227 24021
rect 5258 24012 5264 24064
rect 5316 24052 5322 24064
rect 5629 24055 5687 24061
rect 5629 24052 5641 24055
rect 5316 24024 5641 24052
rect 5316 24012 5322 24024
rect 5629 24021 5641 24024
rect 5675 24021 5687 24055
rect 7098 24052 7104 24064
rect 7059 24024 7104 24052
rect 5629 24015 5687 24021
rect 7098 24012 7104 24024
rect 7156 24012 7162 24064
rect 10060 24061 10088 24092
rect 10382 24089 10394 24092
rect 10428 24089 10440 24123
rect 12986 24120 12992 24132
rect 12947 24092 12992 24120
rect 10382 24083 10440 24089
rect 12986 24080 12992 24092
rect 13044 24080 13050 24132
rect 13906 24120 13912 24132
rect 13867 24092 13912 24120
rect 13906 24080 13912 24092
rect 13964 24120 13970 24132
rect 14200 24120 14228 24151
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 15010 24148 15016 24200
rect 15068 24188 15074 24200
rect 15212 24188 15240 24228
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 16316 24265 16344 24296
rect 17512 24268 17540 24296
rect 17586 24284 17592 24336
rect 17644 24324 17650 24336
rect 17773 24327 17831 24333
rect 17773 24324 17785 24327
rect 17644 24296 17785 24324
rect 17644 24284 17650 24296
rect 17773 24293 17785 24296
rect 17819 24293 17831 24327
rect 18874 24324 18880 24336
rect 18835 24296 18880 24324
rect 17773 24287 17831 24293
rect 18874 24284 18880 24296
rect 18932 24284 18938 24336
rect 19334 24284 19340 24336
rect 19392 24324 19398 24336
rect 20993 24327 21051 24333
rect 19392 24296 19656 24324
rect 19392 24284 19398 24296
rect 16301 24259 16359 24265
rect 16301 24225 16313 24259
rect 16347 24225 16359 24259
rect 16301 24219 16359 24225
rect 16393 24259 16451 24265
rect 16393 24225 16405 24259
rect 16439 24256 16451 24259
rect 16758 24256 16764 24268
rect 16439 24228 16764 24256
rect 16439 24225 16451 24228
rect 16393 24219 16451 24225
rect 16758 24216 16764 24228
rect 16816 24216 16822 24268
rect 17402 24256 17408 24268
rect 17363 24228 17408 24256
rect 17402 24216 17408 24228
rect 17460 24216 17466 24268
rect 17494 24216 17500 24268
rect 17552 24256 17558 24268
rect 18690 24256 18696 24268
rect 17552 24228 17645 24256
rect 17880 24228 18696 24256
rect 17552 24216 17558 24228
rect 15378 24188 15384 24200
rect 15068 24160 15113 24188
rect 15212 24160 15384 24188
rect 15068 24148 15074 24160
rect 15378 24148 15384 24160
rect 15436 24148 15442 24200
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24188 17371 24191
rect 17880 24188 17908 24228
rect 18690 24216 18696 24228
rect 18748 24216 18754 24268
rect 19628 24265 19656 24296
rect 20993 24293 21005 24327
rect 21039 24324 21051 24327
rect 21082 24324 21088 24336
rect 21039 24296 21088 24324
rect 21039 24293 21051 24296
rect 20993 24287 21051 24293
rect 21082 24284 21088 24296
rect 21140 24324 21146 24336
rect 21140 24296 21312 24324
rect 21140 24284 21146 24296
rect 19613 24259 19671 24265
rect 19613 24225 19625 24259
rect 19659 24225 19671 24259
rect 21174 24256 21180 24268
rect 21135 24228 21180 24256
rect 19613 24219 19671 24225
rect 17359 24160 17908 24188
rect 17957 24191 18015 24197
rect 17359 24157 17371 24160
rect 17313 24151 17371 24157
rect 17957 24157 17969 24191
rect 18003 24188 18015 24191
rect 18046 24188 18052 24200
rect 18003 24160 18052 24188
rect 18003 24157 18015 24160
rect 17957 24151 18015 24157
rect 18046 24148 18052 24160
rect 18104 24148 18110 24200
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24188 18199 24191
rect 18598 24188 18604 24200
rect 18187 24160 18604 24188
rect 18187 24157 18199 24160
rect 18141 24151 18199 24157
rect 18598 24148 18604 24160
rect 18656 24148 18662 24200
rect 19337 24191 19395 24197
rect 19337 24188 19349 24191
rect 18984 24160 19349 24188
rect 14826 24120 14832 24132
rect 13964 24092 14228 24120
rect 14787 24092 14832 24120
rect 13964 24080 13970 24092
rect 14826 24080 14832 24092
rect 14884 24080 14890 24132
rect 16574 24080 16580 24132
rect 16632 24120 16638 24132
rect 18506 24120 18512 24132
rect 16632 24092 18512 24120
rect 16632 24080 16638 24092
rect 18506 24080 18512 24092
rect 18564 24080 18570 24132
rect 10045 24055 10103 24061
rect 10045 24021 10057 24055
rect 10091 24021 10103 24055
rect 11790 24052 11796 24064
rect 11751 24024 11796 24052
rect 10045 24015 10103 24021
rect 11790 24012 11796 24024
rect 11848 24012 11854 24064
rect 11882 24012 11888 24064
rect 11940 24052 11946 24064
rect 12529 24055 12587 24061
rect 12529 24052 12541 24055
rect 11940 24024 12541 24052
rect 11940 24012 11946 24024
rect 12529 24021 12541 24024
rect 12575 24021 12587 24055
rect 14642 24052 14648 24064
rect 14603 24024 14648 24052
rect 12529 24015 12587 24021
rect 14642 24012 14648 24024
rect 14700 24012 14706 24064
rect 16482 24012 16488 24064
rect 16540 24052 16546 24064
rect 16850 24052 16856 24064
rect 16540 24024 16585 24052
rect 16811 24024 16856 24052
rect 16540 24012 16546 24024
rect 16850 24012 16856 24024
rect 16908 24012 16914 24064
rect 18984 24061 19012 24160
rect 19337 24157 19349 24160
rect 19383 24157 19395 24191
rect 19628 24188 19656 24219
rect 21174 24216 21180 24228
rect 21232 24216 21238 24268
rect 21284 24265 21312 24296
rect 21269 24259 21327 24265
rect 21269 24225 21281 24259
rect 21315 24225 21327 24259
rect 23293 24259 23351 24265
rect 23293 24256 23305 24259
rect 21269 24219 21327 24225
rect 22480 24228 23305 24256
rect 21636 24191 21694 24197
rect 19628 24160 20024 24188
rect 19337 24151 19395 24157
rect 19858 24123 19916 24129
rect 19858 24120 19870 24123
rect 19536 24092 19870 24120
rect 19536 24061 19564 24092
rect 19858 24089 19870 24092
rect 19904 24089 19916 24123
rect 19996 24120 20024 24160
rect 21636 24157 21648 24191
rect 21682 24188 21694 24191
rect 21910 24188 21916 24200
rect 21682 24160 21916 24188
rect 21682 24157 21694 24160
rect 21636 24151 21694 24157
rect 21910 24148 21916 24160
rect 21968 24188 21974 24200
rect 22480 24188 22508 24228
rect 23293 24225 23305 24228
rect 23339 24225 23351 24259
rect 23293 24219 23351 24225
rect 21968 24160 22508 24188
rect 22891 24191 22949 24197
rect 21968 24148 21974 24160
rect 22891 24157 22903 24191
rect 22937 24188 22949 24191
rect 23198 24188 23204 24200
rect 22937 24160 23060 24188
rect 23159 24160 23204 24188
rect 22937 24157 22949 24160
rect 22891 24151 22949 24157
rect 22094 24120 22100 24132
rect 19996 24092 22100 24120
rect 19858 24083 19916 24089
rect 22094 24080 22100 24092
rect 22152 24080 22158 24132
rect 22554 24080 22560 24132
rect 22612 24120 22618 24132
rect 22649 24123 22707 24129
rect 22649 24120 22661 24123
rect 22612 24092 22661 24120
rect 22612 24080 22618 24092
rect 22649 24089 22661 24092
rect 22695 24089 22707 24123
rect 23032 24120 23060 24160
rect 23198 24148 23204 24160
rect 23256 24148 23262 24200
rect 24026 24120 24032 24132
rect 23032 24092 24032 24120
rect 22649 24083 22707 24089
rect 24026 24080 24032 24092
rect 24084 24080 24090 24132
rect 18969 24055 19027 24061
rect 18969 24021 18981 24055
rect 19015 24021 19027 24055
rect 18969 24015 19027 24021
rect 19521 24055 19579 24061
rect 19521 24021 19533 24055
rect 19567 24021 19579 24055
rect 19521 24015 19579 24021
rect 20530 24012 20536 24064
rect 20588 24052 20594 24064
rect 21729 24055 21787 24061
rect 21729 24052 21741 24055
rect 20588 24024 21741 24052
rect 20588 24012 20594 24024
rect 21729 24021 21741 24024
rect 21775 24021 21787 24055
rect 21729 24015 21787 24021
rect 1104 23962 26220 23984
rect 1104 23910 9322 23962
rect 9374 23910 9386 23962
rect 9438 23910 9450 23962
rect 9502 23910 9514 23962
rect 9566 23910 9578 23962
rect 9630 23910 17694 23962
rect 17746 23910 17758 23962
rect 17810 23910 17822 23962
rect 17874 23910 17886 23962
rect 17938 23910 17950 23962
rect 18002 23910 26220 23962
rect 1104 23888 26220 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 4246 23808 4252 23860
rect 4304 23848 4310 23860
rect 4341 23851 4399 23857
rect 4341 23848 4353 23851
rect 4304 23820 4353 23848
rect 4304 23808 4310 23820
rect 4341 23817 4353 23820
rect 4387 23817 4399 23851
rect 4341 23811 4399 23817
rect 4448 23820 5948 23848
rect 2716 23783 2774 23789
rect 2716 23749 2728 23783
rect 2762 23780 2774 23783
rect 3789 23783 3847 23789
rect 3789 23780 3801 23783
rect 2762 23752 3801 23780
rect 2762 23749 2774 23752
rect 2716 23743 2774 23749
rect 3789 23749 3801 23752
rect 3835 23749 3847 23783
rect 3789 23743 3847 23749
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 4062 23780 4068 23792
rect 4019 23752 4068 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 4062 23740 4068 23752
rect 4120 23740 4126 23792
rect 4448 23724 4476 23820
rect 5810 23780 5816 23792
rect 4724 23752 5816 23780
rect 4154 23712 4160 23724
rect 4115 23684 4160 23712
rect 4154 23672 4160 23684
rect 4212 23672 4218 23724
rect 4430 23712 4436 23724
rect 4391 23684 4436 23712
rect 4430 23672 4436 23684
rect 4488 23672 4494 23724
rect 4724 23721 4752 23752
rect 5810 23740 5816 23752
rect 5868 23740 5874 23792
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23681 4767 23715
rect 4709 23675 4767 23681
rect 4976 23715 5034 23721
rect 4976 23681 4988 23715
rect 5022 23712 5034 23715
rect 5258 23712 5264 23724
rect 5022 23684 5264 23712
rect 5022 23681 5034 23684
rect 4976 23675 5034 23681
rect 2961 23647 3019 23653
rect 2961 23613 2973 23647
rect 3007 23644 3019 23647
rect 4724 23644 4752 23675
rect 5258 23672 5264 23684
rect 5316 23672 5322 23724
rect 5920 23712 5948 23820
rect 5994 23808 6000 23860
rect 6052 23848 6058 23860
rect 6457 23851 6515 23857
rect 6457 23848 6469 23851
rect 6052 23820 6469 23848
rect 6052 23808 6058 23820
rect 6457 23817 6469 23820
rect 6503 23817 6515 23851
rect 8110 23848 8116 23860
rect 6457 23811 6515 23817
rect 6932 23820 8116 23848
rect 6822 23712 6828 23724
rect 5920 23684 6828 23712
rect 6822 23672 6828 23684
rect 6880 23672 6886 23724
rect 6932 23721 6960 23820
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 9766 23848 9772 23860
rect 9727 23820 9772 23848
rect 9766 23808 9772 23820
rect 9824 23808 9830 23860
rect 10413 23851 10471 23857
rect 10413 23817 10425 23851
rect 10459 23848 10471 23851
rect 11790 23848 11796 23860
rect 10459 23820 11796 23848
rect 10459 23817 10471 23820
rect 10413 23811 10471 23817
rect 11790 23808 11796 23820
rect 11848 23808 11854 23860
rect 12345 23851 12403 23857
rect 12345 23817 12357 23851
rect 12391 23848 12403 23851
rect 12434 23848 12440 23860
rect 12391 23820 12440 23848
rect 12391 23817 12403 23820
rect 12345 23811 12403 23817
rect 12434 23808 12440 23820
rect 12492 23848 12498 23860
rect 12986 23848 12992 23860
rect 12492 23820 12992 23848
rect 12492 23808 12498 23820
rect 12986 23808 12992 23820
rect 13044 23808 13050 23860
rect 13817 23851 13875 23857
rect 13817 23817 13829 23851
rect 13863 23848 13875 23851
rect 13906 23848 13912 23860
rect 13863 23820 13912 23848
rect 13863 23817 13875 23820
rect 13817 23811 13875 23817
rect 13906 23808 13912 23820
rect 13964 23808 13970 23860
rect 15378 23848 15384 23860
rect 15339 23820 15384 23848
rect 15378 23808 15384 23820
rect 15436 23808 15442 23860
rect 16758 23848 16764 23860
rect 16719 23820 16764 23848
rect 16758 23808 16764 23820
rect 16816 23808 16822 23860
rect 17405 23851 17463 23857
rect 17405 23817 17417 23851
rect 17451 23848 17463 23851
rect 17494 23848 17500 23860
rect 17451 23820 17500 23848
rect 17451 23817 17463 23820
rect 17405 23811 17463 23817
rect 17494 23808 17500 23820
rect 17552 23808 17558 23860
rect 18417 23851 18475 23857
rect 18417 23817 18429 23851
rect 18463 23848 18475 23851
rect 19334 23848 19340 23860
rect 18463 23820 19340 23848
rect 18463 23817 18475 23820
rect 18417 23811 18475 23817
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 19702 23848 19708 23860
rect 19663 23820 19708 23848
rect 19702 23808 19708 23820
rect 19760 23808 19766 23860
rect 20073 23851 20131 23857
rect 20073 23817 20085 23851
rect 20119 23817 20131 23851
rect 20530 23848 20536 23860
rect 20491 23820 20536 23848
rect 20073 23811 20131 23817
rect 7282 23740 7288 23792
rect 7340 23740 7346 23792
rect 10778 23780 10784 23792
rect 10739 23752 10784 23780
rect 10778 23740 10784 23752
rect 10836 23740 10842 23792
rect 12452 23752 14044 23780
rect 6917 23715 6975 23721
rect 6917 23681 6929 23715
rect 6963 23681 6975 23715
rect 7190 23712 7196 23724
rect 7151 23684 7196 23712
rect 6917 23675 6975 23681
rect 7190 23672 7196 23684
rect 7248 23672 7254 23724
rect 7300 23712 7328 23740
rect 7469 23715 7527 23721
rect 7469 23712 7481 23715
rect 7300 23684 7481 23712
rect 7469 23681 7481 23684
rect 7515 23681 7527 23715
rect 7469 23675 7527 23681
rect 8113 23715 8171 23721
rect 8113 23681 8125 23715
rect 8159 23681 8171 23715
rect 8113 23675 8171 23681
rect 8297 23715 8355 23721
rect 8297 23681 8309 23715
rect 8343 23712 8355 23715
rect 8570 23712 8576 23724
rect 8343 23684 8576 23712
rect 8343 23681 8355 23684
rect 8297 23675 8355 23681
rect 3007 23616 4752 23644
rect 6641 23647 6699 23653
rect 3007 23613 3019 23616
rect 2961 23607 3019 23613
rect 6641 23613 6653 23647
rect 6687 23644 6699 23647
rect 7285 23647 7343 23653
rect 7285 23644 7297 23647
rect 6687 23616 7297 23644
rect 6687 23613 6699 23616
rect 6641 23607 6699 23613
rect 7285 23613 7297 23616
rect 7331 23644 7343 23647
rect 7374 23644 7380 23656
rect 7331 23616 7380 23644
rect 7331 23613 7343 23616
rect 7285 23607 7343 23613
rect 6089 23579 6147 23585
rect 6089 23545 6101 23579
rect 6135 23576 6147 23579
rect 6656 23576 6684 23607
rect 7374 23604 7380 23616
rect 7432 23644 7438 23656
rect 8128 23644 8156 23675
rect 8570 23672 8576 23684
rect 8628 23672 8634 23724
rect 10321 23715 10379 23721
rect 10321 23681 10333 23715
rect 10367 23712 10379 23715
rect 10686 23712 10692 23724
rect 10367 23684 10692 23712
rect 10367 23681 10379 23684
rect 10321 23675 10379 23681
rect 10686 23672 10692 23684
rect 10744 23672 10750 23724
rect 7432 23616 8156 23644
rect 9309 23647 9367 23653
rect 7432 23604 7438 23616
rect 9309 23613 9321 23647
rect 9355 23644 9367 23647
rect 9766 23644 9772 23656
rect 9355 23616 9772 23644
rect 9355 23613 9367 23616
rect 9309 23607 9367 23613
rect 9766 23604 9772 23616
rect 9824 23604 9830 23656
rect 10042 23604 10048 23656
rect 10100 23644 10106 23656
rect 10597 23647 10655 23653
rect 10597 23644 10609 23647
rect 10100 23616 10609 23644
rect 10100 23604 10106 23616
rect 10597 23613 10609 23616
rect 10643 23644 10655 23647
rect 10796 23644 10824 23740
rect 11882 23712 11888 23724
rect 11843 23684 11888 23712
rect 11882 23672 11888 23684
rect 11940 23672 11946 23724
rect 12158 23712 12164 23724
rect 12119 23684 12164 23712
rect 12158 23672 12164 23684
rect 12216 23672 12222 23724
rect 12452 23721 12480 23752
rect 14016 23724 14044 23752
rect 16574 23740 16580 23792
rect 16632 23780 16638 23792
rect 17221 23783 17279 23789
rect 17221 23780 17233 23783
rect 16632 23752 17233 23780
rect 16632 23740 16638 23752
rect 17221 23749 17233 23752
rect 17267 23749 17279 23783
rect 17221 23743 17279 23749
rect 18874 23740 18880 23792
rect 18932 23780 18938 23792
rect 20088 23780 20116 23811
rect 20530 23808 20536 23820
rect 20588 23808 20594 23860
rect 21174 23848 21180 23860
rect 20916 23820 21180 23848
rect 20916 23789 20944 23820
rect 21174 23808 21180 23820
rect 21232 23808 21238 23860
rect 22005 23851 22063 23857
rect 22005 23817 22017 23851
rect 22051 23817 22063 23851
rect 22005 23811 22063 23817
rect 18932 23752 20116 23780
rect 20901 23783 20959 23789
rect 18932 23740 18938 23752
rect 20901 23749 20913 23783
rect 20947 23749 20959 23783
rect 21082 23780 21088 23792
rect 21043 23752 21088 23780
rect 20901 23743 20959 23749
rect 21082 23740 21088 23752
rect 21140 23740 21146 23792
rect 21269 23783 21327 23789
rect 21269 23749 21281 23783
rect 21315 23780 21327 23783
rect 21910 23780 21916 23792
rect 21315 23752 21916 23780
rect 21315 23749 21327 23752
rect 21269 23743 21327 23749
rect 21910 23740 21916 23752
rect 21968 23740 21974 23792
rect 22020 23780 22048 23811
rect 23198 23808 23204 23860
rect 23256 23848 23262 23860
rect 23477 23851 23535 23857
rect 23477 23848 23489 23851
rect 23256 23820 23489 23848
rect 23256 23808 23262 23820
rect 23477 23817 23489 23820
rect 23523 23817 23535 23851
rect 23477 23811 23535 23817
rect 22342 23783 22400 23789
rect 22342 23780 22354 23783
rect 22020 23752 22354 23780
rect 22342 23749 22354 23752
rect 22388 23749 22400 23783
rect 23492 23780 23520 23811
rect 23845 23783 23903 23789
rect 23845 23780 23857 23783
rect 23492 23752 23857 23780
rect 22342 23743 22400 23749
rect 23845 23749 23857 23752
rect 23891 23749 23903 23783
rect 24026 23780 24032 23792
rect 23987 23752 24032 23780
rect 23845 23743 23903 23749
rect 24026 23740 24032 23752
rect 24084 23740 24090 23792
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23681 12495 23715
rect 12693 23715 12751 23721
rect 12693 23712 12705 23715
rect 12437 23675 12495 23681
rect 12544 23684 12705 23712
rect 12544 23644 12572 23684
rect 12693 23681 12705 23684
rect 12739 23681 12751 23715
rect 13998 23712 14004 23724
rect 13959 23684 14004 23712
rect 12693 23675 12751 23681
rect 13998 23672 14004 23684
rect 14056 23672 14062 23724
rect 14090 23672 14096 23724
rect 14148 23712 14154 23724
rect 14257 23715 14315 23721
rect 14257 23712 14269 23715
rect 14148 23684 14269 23712
rect 14148 23672 14154 23684
rect 14257 23681 14269 23684
rect 14303 23681 14315 23715
rect 18322 23712 18328 23724
rect 18283 23684 18328 23712
rect 14257 23675 14315 23681
rect 18322 23672 18328 23684
rect 18380 23672 18386 23724
rect 18785 23715 18843 23721
rect 18785 23681 18797 23715
rect 18831 23681 18843 23715
rect 18785 23675 18843 23681
rect 19613 23715 19671 23721
rect 19613 23681 19625 23715
rect 19659 23712 19671 23715
rect 19978 23712 19984 23724
rect 19659 23684 19984 23712
rect 19659 23681 19671 23684
rect 19613 23675 19671 23681
rect 18800 23644 18828 23675
rect 19978 23672 19984 23684
rect 20036 23672 20042 23724
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23712 20499 23715
rect 20806 23712 20812 23724
rect 20487 23684 20812 23712
rect 20487 23681 20499 23684
rect 20441 23675 20499 23681
rect 20806 23672 20812 23684
rect 20864 23672 20870 23724
rect 21726 23672 21732 23724
rect 21784 23712 21790 23724
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 21784 23684 21833 23712
rect 21784 23672 21790 23684
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 21928 23712 21956 23740
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 21928 23684 23673 23712
rect 21821 23675 21879 23681
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 19702 23644 19708 23656
rect 10643 23616 10824 23644
rect 12406 23616 12572 23644
rect 17144 23616 19708 23644
rect 10643 23613 10655 23616
rect 10597 23607 10655 23613
rect 6135 23548 6684 23576
rect 7653 23579 7711 23585
rect 6135 23545 6147 23548
rect 6089 23539 6147 23545
rect 7653 23545 7665 23579
rect 7699 23576 7711 23579
rect 8202 23576 8208 23588
rect 7699 23548 8208 23576
rect 7699 23545 7711 23548
rect 7653 23539 7711 23545
rect 8202 23536 8208 23548
rect 8260 23536 8266 23588
rect 9677 23579 9735 23585
rect 9677 23545 9689 23579
rect 9723 23576 9735 23579
rect 9953 23579 10011 23585
rect 9953 23576 9965 23579
rect 9723 23548 9965 23576
rect 9723 23545 9735 23548
rect 9677 23539 9735 23545
rect 9953 23545 9965 23548
rect 9999 23545 10011 23579
rect 9953 23539 10011 23545
rect 12069 23579 12127 23585
rect 12069 23545 12081 23579
rect 12115 23576 12127 23579
rect 12406 23576 12434 23616
rect 16850 23576 16856 23588
rect 12115 23548 12434 23576
rect 16811 23548 16856 23576
rect 12115 23545 12127 23548
rect 12069 23539 12127 23545
rect 16850 23536 16856 23548
rect 16908 23536 16914 23588
rect 3789 23511 3847 23517
rect 3789 23477 3801 23511
rect 3835 23508 3847 23511
rect 6730 23508 6736 23520
rect 3835 23480 6736 23508
rect 3835 23477 3847 23480
rect 3789 23471 3847 23477
rect 6730 23468 6736 23480
rect 6788 23468 6794 23520
rect 7466 23508 7472 23520
rect 7427 23480 7472 23508
rect 7466 23468 7472 23480
rect 7524 23468 7530 23520
rect 7742 23468 7748 23520
rect 7800 23508 7806 23520
rect 7929 23511 7987 23517
rect 7929 23508 7941 23511
rect 7800 23480 7941 23508
rect 7800 23468 7806 23480
rect 7929 23477 7941 23480
rect 7975 23477 7987 23511
rect 8110 23508 8116 23520
rect 8071 23480 8116 23508
rect 7929 23471 7987 23477
rect 8110 23468 8116 23480
rect 8168 23468 8174 23520
rect 12158 23468 12164 23520
rect 12216 23508 12222 23520
rect 17144 23508 17172 23616
rect 19702 23604 19708 23616
rect 19760 23604 19766 23656
rect 19889 23647 19947 23653
rect 19889 23613 19901 23647
rect 19935 23644 19947 23647
rect 20530 23644 20536 23656
rect 19935 23616 20536 23644
rect 19935 23613 19947 23616
rect 19889 23607 19947 23613
rect 18506 23536 18512 23588
rect 18564 23576 18570 23588
rect 18601 23579 18659 23585
rect 18601 23576 18613 23579
rect 18564 23548 18613 23576
rect 18564 23536 18570 23548
rect 18601 23545 18613 23548
rect 18647 23545 18659 23579
rect 19242 23576 19248 23588
rect 19203 23548 19248 23576
rect 18601 23539 18659 23545
rect 19242 23536 19248 23548
rect 19300 23536 19306 23588
rect 12216 23480 17172 23508
rect 19153 23511 19211 23517
rect 12216 23468 12222 23480
rect 19153 23477 19165 23511
rect 19199 23508 19211 23511
rect 19426 23508 19432 23520
rect 19199 23480 19432 23508
rect 19199 23477 19211 23480
rect 19153 23471 19211 23477
rect 19426 23468 19432 23480
rect 19484 23508 19490 23520
rect 19904 23508 19932 23607
rect 20530 23604 20536 23616
rect 20588 23644 20594 23656
rect 20625 23647 20683 23653
rect 20625 23644 20637 23647
rect 20588 23616 20637 23644
rect 20588 23604 20594 23616
rect 20625 23613 20637 23616
rect 20671 23613 20683 23647
rect 22094 23644 22100 23656
rect 22007 23616 22100 23644
rect 20625 23607 20683 23613
rect 22094 23604 22100 23616
rect 22152 23604 22158 23656
rect 19484 23480 19932 23508
rect 22112 23508 22140 23604
rect 22738 23508 22744 23520
rect 22112 23480 22744 23508
rect 19484 23468 19490 23480
rect 22738 23468 22744 23480
rect 22796 23468 22802 23520
rect 1104 23418 26220 23440
rect 1104 23366 5136 23418
rect 5188 23366 5200 23418
rect 5252 23366 5264 23418
rect 5316 23366 5328 23418
rect 5380 23366 5392 23418
rect 5444 23366 13508 23418
rect 13560 23366 13572 23418
rect 13624 23366 13636 23418
rect 13688 23366 13700 23418
rect 13752 23366 13764 23418
rect 13816 23366 21880 23418
rect 21932 23366 21944 23418
rect 21996 23366 22008 23418
rect 22060 23366 22072 23418
rect 22124 23366 22136 23418
rect 22188 23366 26220 23418
rect 1104 23344 26220 23366
rect 7098 23304 7104 23316
rect 4724 23276 7104 23304
rect 4154 23236 4160 23248
rect 4115 23208 4160 23236
rect 4154 23196 4160 23208
rect 4212 23196 4218 23248
rect 4249 23171 4307 23177
rect 4249 23137 4261 23171
rect 4295 23168 4307 23171
rect 4430 23168 4436 23180
rect 4295 23140 4436 23168
rect 4295 23137 4307 23140
rect 4249 23131 4307 23137
rect 4430 23128 4436 23140
rect 4488 23128 4494 23180
rect 4617 23171 4675 23177
rect 4617 23137 4629 23171
rect 4663 23168 4675 23171
rect 4724 23168 4752 23276
rect 7098 23264 7104 23276
rect 7156 23264 7162 23316
rect 7190 23264 7196 23316
rect 7248 23304 7254 23316
rect 7377 23307 7435 23313
rect 7377 23304 7389 23307
rect 7248 23276 7389 23304
rect 7248 23264 7254 23276
rect 7377 23273 7389 23276
rect 7423 23273 7435 23307
rect 8113 23307 8171 23313
rect 8113 23304 8125 23307
rect 7377 23267 7435 23273
rect 7484 23276 8125 23304
rect 7006 23196 7012 23248
rect 7064 23236 7070 23248
rect 7484 23236 7512 23276
rect 8113 23273 8125 23276
rect 8159 23273 8171 23307
rect 9766 23304 9772 23316
rect 9727 23276 9772 23304
rect 8113 23267 8171 23273
rect 9766 23264 9772 23276
rect 9824 23264 9830 23316
rect 12618 23304 12624 23316
rect 12579 23276 12624 23304
rect 12618 23264 12624 23276
rect 12676 23264 12682 23316
rect 13909 23307 13967 23313
rect 13909 23273 13921 23307
rect 13955 23304 13967 23307
rect 14090 23304 14096 23316
rect 13955 23276 14096 23304
rect 13955 23273 13967 23276
rect 13909 23267 13967 23273
rect 14090 23264 14096 23276
rect 14148 23264 14154 23316
rect 15013 23307 15071 23313
rect 15013 23273 15025 23307
rect 15059 23304 15071 23307
rect 15102 23304 15108 23316
rect 15059 23276 15108 23304
rect 15059 23273 15071 23276
rect 15013 23267 15071 23273
rect 8389 23239 8447 23245
rect 8389 23236 8401 23239
rect 7064 23208 7512 23236
rect 7852 23208 8401 23236
rect 7064 23196 7070 23208
rect 4663 23140 4752 23168
rect 5261 23171 5319 23177
rect 4663 23137 4675 23140
rect 4617 23131 4675 23137
rect 5261 23137 5273 23171
rect 5307 23168 5319 23171
rect 5534 23168 5540 23180
rect 5307 23140 5540 23168
rect 5307 23137 5319 23140
rect 5261 23131 5319 23137
rect 5534 23128 5540 23140
rect 5592 23128 5598 23180
rect 5810 23128 5816 23180
rect 5868 23168 5874 23180
rect 5997 23171 6055 23177
rect 5997 23168 6009 23171
rect 5868 23140 6009 23168
rect 5868 23128 5874 23140
rect 5997 23137 6009 23140
rect 6043 23137 6055 23171
rect 5997 23131 6055 23137
rect 7852 23112 7880 23208
rect 8389 23205 8401 23208
rect 8435 23205 8447 23239
rect 8389 23199 8447 23205
rect 8202 23128 8208 23180
rect 8260 23168 8266 23180
rect 8260 23140 8305 23168
rect 8260 23128 8266 23140
rect 10778 23128 10784 23180
rect 10836 23168 10842 23180
rect 13265 23171 13323 23177
rect 13265 23168 13277 23171
rect 10836 23140 13277 23168
rect 10836 23128 10842 23140
rect 13265 23137 13277 23140
rect 13311 23168 13323 23171
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 13311 23140 13553 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 13541 23137 13553 23140
rect 13587 23168 13599 23171
rect 14737 23171 14795 23177
rect 14737 23168 14749 23171
rect 13587 23140 14749 23168
rect 13587 23137 13599 23140
rect 13541 23131 13599 23137
rect 14737 23137 14749 23140
rect 14783 23168 14795 23171
rect 15028 23168 15056 23267
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 21726 23264 21732 23316
rect 21784 23304 21790 23316
rect 21913 23307 21971 23313
rect 21913 23304 21925 23307
rect 21784 23276 21925 23304
rect 21784 23264 21790 23276
rect 21913 23273 21925 23276
rect 21959 23273 21971 23307
rect 21913 23267 21971 23273
rect 19981 23239 20039 23245
rect 19981 23205 19993 23239
rect 20027 23236 20039 23239
rect 20622 23236 20628 23248
rect 20027 23208 20628 23236
rect 20027 23205 20039 23208
rect 19981 23199 20039 23205
rect 20622 23196 20628 23208
rect 20680 23236 20686 23248
rect 21821 23239 21879 23245
rect 20680 23208 21496 23236
rect 20680 23196 20686 23208
rect 21468 23180 21496 23208
rect 21821 23205 21833 23239
rect 21867 23236 21879 23239
rect 22097 23239 22155 23245
rect 22097 23236 22109 23239
rect 21867 23208 22109 23236
rect 21867 23205 21879 23208
rect 21821 23199 21879 23205
rect 22097 23205 22109 23208
rect 22143 23205 22155 23239
rect 22097 23199 22155 23205
rect 21450 23168 21456 23180
rect 14783 23140 15056 23168
rect 21363 23140 21456 23168
rect 14783 23137 14795 23140
rect 14737 23131 14795 23137
rect 21450 23128 21456 23140
rect 21508 23128 21514 23180
rect 22554 23168 22560 23180
rect 22515 23140 22560 23168
rect 22554 23128 22560 23140
rect 22612 23128 22618 23180
rect 22649 23171 22707 23177
rect 22649 23137 22661 23171
rect 22695 23137 22707 23171
rect 22649 23131 22707 23137
rect 23661 23171 23719 23177
rect 23661 23137 23673 23171
rect 23707 23168 23719 23171
rect 24026 23168 24032 23180
rect 23707 23140 24032 23168
rect 23707 23137 23719 23140
rect 23661 23131 23719 23137
rect 4065 23103 4123 23109
rect 4065 23069 4077 23103
rect 4111 23069 4123 23103
rect 4706 23100 4712 23112
rect 4667 23072 4712 23100
rect 4065 23063 4123 23069
rect 4080 22964 4108 23063
rect 4706 23060 4712 23072
rect 4764 23060 4770 23112
rect 5626 23100 5632 23112
rect 5587 23072 5632 23100
rect 5626 23060 5632 23072
rect 5684 23060 5690 23112
rect 5721 23103 5779 23109
rect 5721 23069 5733 23103
rect 5767 23100 5779 23103
rect 7653 23103 7711 23109
rect 7653 23100 7665 23103
rect 5767 23072 7665 23100
rect 5767 23069 5779 23072
rect 5721 23063 5779 23069
rect 7653 23069 7665 23072
rect 7699 23069 7711 23103
rect 7834 23100 7840 23112
rect 7747 23072 7840 23100
rect 7653 23063 7711 23069
rect 7834 23060 7840 23072
rect 7892 23060 7898 23112
rect 7926 23060 7932 23112
rect 7984 23100 7990 23112
rect 8220 23100 8248 23128
rect 8297 23103 8355 23109
rect 8297 23100 8309 23103
rect 7984 23072 8029 23100
rect 8220 23072 8309 23100
rect 7984 23060 7990 23072
rect 8297 23069 8309 23072
rect 8343 23069 8355 23103
rect 9950 23100 9956 23112
rect 9911 23072 9956 23100
rect 8297 23063 8355 23069
rect 9950 23060 9956 23072
rect 10008 23100 10014 23112
rect 12158 23100 12164 23112
rect 10008 23072 12164 23100
rect 10008 23060 10014 23072
rect 12158 23060 12164 23072
rect 12216 23060 12222 23112
rect 13725 23103 13783 23109
rect 13725 23069 13737 23103
rect 13771 23100 13783 23103
rect 13814 23100 13820 23112
rect 13771 23072 13820 23100
rect 13771 23069 13783 23072
rect 13725 23063 13783 23069
rect 13814 23060 13820 23072
rect 13872 23060 13878 23112
rect 14461 23103 14519 23109
rect 14461 23069 14473 23103
rect 14507 23100 14519 23103
rect 14550 23100 14556 23112
rect 14507 23072 14556 23100
rect 14507 23069 14519 23072
rect 14461 23063 14519 23069
rect 14550 23060 14556 23072
rect 14608 23060 14614 23112
rect 19702 23060 19708 23112
rect 19760 23100 19766 23112
rect 19797 23103 19855 23109
rect 19797 23100 19809 23103
rect 19760 23072 19809 23100
rect 19760 23060 19766 23072
rect 19797 23069 19809 23072
rect 19843 23069 19855 23103
rect 19797 23063 19855 23069
rect 20165 23103 20223 23109
rect 20165 23069 20177 23103
rect 20211 23100 20223 23103
rect 20530 23100 20536 23112
rect 20211 23072 20536 23100
rect 20211 23069 20223 23072
rect 20165 23063 20223 23069
rect 20530 23060 20536 23072
rect 20588 23100 20594 23112
rect 21361 23103 21419 23109
rect 21361 23100 21373 23103
rect 20588 23072 21373 23100
rect 20588 23060 20594 23072
rect 21361 23069 21373 23072
rect 21407 23100 21419 23103
rect 22664 23100 22692 23131
rect 24026 23128 24032 23140
rect 24084 23128 24090 23180
rect 25130 23168 25136 23180
rect 25091 23140 25136 23168
rect 25130 23128 25136 23140
rect 25188 23128 25194 23180
rect 21407 23072 22692 23100
rect 23259 23103 23317 23109
rect 21407 23069 21419 23072
rect 21361 23063 21419 23069
rect 23259 23069 23271 23103
rect 23305 23100 23317 23103
rect 23566 23100 23572 23112
rect 23305 23069 23336 23100
rect 23527 23072 23572 23100
rect 23259 23063 23336 23069
rect 4433 23035 4491 23041
rect 4433 23001 4445 23035
rect 4479 23032 4491 23035
rect 5905 23035 5963 23041
rect 4479 23004 5212 23032
rect 4479 23001 4491 23004
rect 4433 22995 4491 23001
rect 4709 22967 4767 22973
rect 4709 22964 4721 22967
rect 4080 22936 4721 22964
rect 4709 22933 4721 22936
rect 4755 22933 4767 22967
rect 5184 22964 5212 23004
rect 5905 23001 5917 23035
rect 5951 23032 5963 23035
rect 6242 23035 6300 23041
rect 6242 23032 6254 23035
rect 5951 23004 6254 23032
rect 5951 23001 5963 23004
rect 5905 22995 5963 23001
rect 6242 23001 6254 23004
rect 6288 23001 6300 23035
rect 6242 22995 6300 23001
rect 6914 22992 6920 23044
rect 6972 23032 6978 23044
rect 9033 23035 9091 23041
rect 9033 23032 9045 23035
rect 6972 23004 9045 23032
rect 6972 22992 6978 23004
rect 9033 23001 9045 23004
rect 9079 23001 9091 23035
rect 9214 23032 9220 23044
rect 9175 23004 9220 23032
rect 9033 22995 9091 23001
rect 9214 22992 9220 23004
rect 9272 22992 9278 23044
rect 13081 23035 13139 23041
rect 13081 23001 13093 23035
rect 13127 23032 13139 23035
rect 14642 23032 14648 23044
rect 13127 23004 14648 23032
rect 13127 23001 13139 23004
rect 13081 22995 13139 23001
rect 14642 22992 14648 23004
rect 14700 22992 14706 23044
rect 16393 23035 16451 23041
rect 16393 23001 16405 23035
rect 16439 23032 16451 23035
rect 16577 23035 16635 23041
rect 16577 23032 16589 23035
rect 16439 23004 16589 23032
rect 16439 23001 16451 23004
rect 16393 22995 16451 23001
rect 16577 23001 16589 23004
rect 16623 23032 16635 23035
rect 18046 23032 18052 23044
rect 16623 23004 18052 23032
rect 16623 23001 16635 23004
rect 16577 22995 16635 23001
rect 18046 22992 18052 23004
rect 18104 22992 18110 23044
rect 23014 23032 23020 23044
rect 22975 23004 23020 23032
rect 23014 22992 23020 23004
rect 23072 22992 23078 23044
rect 23308 23032 23336 23063
rect 23566 23060 23572 23072
rect 23624 23060 23630 23112
rect 23474 23032 23480 23044
rect 23308 23004 23480 23032
rect 23474 22992 23480 23004
rect 23532 22992 23538 23044
rect 9858 22964 9864 22976
rect 5184 22936 9864 22964
rect 4709 22927 4767 22933
rect 9858 22924 9864 22936
rect 9916 22924 9922 22976
rect 12802 22924 12808 22976
rect 12860 22964 12866 22976
rect 12989 22967 13047 22973
rect 12989 22964 13001 22967
rect 12860 22936 13001 22964
rect 12860 22924 12866 22936
rect 12989 22933 13001 22936
rect 13035 22933 13047 22967
rect 14090 22964 14096 22976
rect 14051 22936 14096 22964
rect 12989 22927 13047 22933
rect 14090 22924 14096 22936
rect 14148 22924 14154 22976
rect 14553 22967 14611 22973
rect 14553 22933 14565 22967
rect 14599 22964 14611 22967
rect 14826 22964 14832 22976
rect 14599 22936 14832 22964
rect 14599 22933 14611 22936
rect 14553 22927 14611 22933
rect 14826 22924 14832 22936
rect 14884 22924 14890 22976
rect 16666 22964 16672 22976
rect 16627 22936 16672 22964
rect 16666 22924 16672 22936
rect 16724 22964 16730 22976
rect 18322 22964 18328 22976
rect 16724 22936 18328 22964
rect 16724 22924 16730 22936
rect 18322 22924 18328 22936
rect 18380 22924 18386 22976
rect 22462 22964 22468 22976
rect 22423 22936 22468 22964
rect 22462 22924 22468 22936
rect 22520 22924 22526 22976
rect 1104 22874 26220 22896
rect 1104 22822 9322 22874
rect 9374 22822 9386 22874
rect 9438 22822 9450 22874
rect 9502 22822 9514 22874
rect 9566 22822 9578 22874
rect 9630 22822 17694 22874
rect 17746 22822 17758 22874
rect 17810 22822 17822 22874
rect 17874 22822 17886 22874
rect 17938 22822 17950 22874
rect 18002 22822 26220 22874
rect 1104 22800 26220 22822
rect 5534 22760 5540 22772
rect 5447 22732 5540 22760
rect 5534 22720 5540 22732
rect 5592 22760 5598 22772
rect 5810 22760 5816 22772
rect 5592 22732 5816 22760
rect 5592 22720 5598 22732
rect 5810 22720 5816 22732
rect 5868 22720 5874 22772
rect 7834 22760 7840 22772
rect 7024 22732 7840 22760
rect 5552 22692 5580 22720
rect 3344 22664 5580 22692
rect 5629 22695 5687 22701
rect 3344 22636 3372 22664
rect 5629 22661 5641 22695
rect 5675 22692 5687 22695
rect 6914 22692 6920 22704
rect 5675 22664 6920 22692
rect 5675 22661 5687 22664
rect 5629 22655 5687 22661
rect 6914 22652 6920 22664
rect 6972 22652 6978 22704
rect 7024 22701 7052 22732
rect 7834 22720 7840 22732
rect 7892 22720 7898 22772
rect 8294 22720 8300 22772
rect 8352 22760 8358 22772
rect 8846 22760 8852 22772
rect 8352 22732 8852 22760
rect 8352 22720 8358 22732
rect 8846 22720 8852 22732
rect 8904 22720 8910 22772
rect 8938 22720 8944 22772
rect 8996 22760 9002 22772
rect 9217 22763 9275 22769
rect 9217 22760 9229 22763
rect 8996 22732 9229 22760
rect 8996 22720 9002 22732
rect 9217 22729 9229 22732
rect 9263 22729 9275 22763
rect 9217 22723 9275 22729
rect 9309 22763 9367 22769
rect 9309 22729 9321 22763
rect 9355 22729 9367 22763
rect 9309 22723 9367 22729
rect 7009 22695 7067 22701
rect 7009 22661 7021 22695
rect 7055 22661 7067 22695
rect 7009 22655 7067 22661
rect 7190 22652 7196 22704
rect 7248 22692 7254 22704
rect 7248 22664 7604 22692
rect 7248 22652 7254 22664
rect 3326 22624 3332 22636
rect 3239 22596 3332 22624
rect 3326 22584 3332 22596
rect 3384 22584 3390 22636
rect 3596 22627 3654 22633
rect 3596 22593 3608 22627
rect 3642 22624 3654 22627
rect 4338 22624 4344 22636
rect 3642 22596 4344 22624
rect 3642 22593 3654 22596
rect 3596 22587 3654 22593
rect 4338 22584 4344 22596
rect 4396 22584 4402 22636
rect 6825 22627 6883 22633
rect 6825 22593 6837 22627
rect 6871 22624 6883 22627
rect 7098 22624 7104 22636
rect 6871 22596 7104 22624
rect 6871 22593 6883 22596
rect 6825 22587 6883 22593
rect 7098 22584 7104 22596
rect 7156 22584 7162 22636
rect 7576 22633 7604 22664
rect 7650 22652 7656 22704
rect 7708 22692 7714 22704
rect 8021 22695 8079 22701
rect 8021 22692 8033 22695
rect 7708 22664 8033 22692
rect 7708 22652 7714 22664
rect 8021 22661 8033 22664
rect 8067 22692 8079 22695
rect 9033 22695 9091 22701
rect 9033 22692 9045 22695
rect 8067 22664 9045 22692
rect 8067 22661 8079 22664
rect 8021 22655 8079 22661
rect 9033 22661 9045 22664
rect 9079 22661 9091 22695
rect 9033 22655 9091 22661
rect 9122 22652 9128 22704
rect 9180 22692 9186 22704
rect 9324 22692 9352 22723
rect 9950 22720 9956 22772
rect 10008 22760 10014 22772
rect 10137 22763 10195 22769
rect 10137 22760 10149 22763
rect 10008 22732 10149 22760
rect 10008 22720 10014 22732
rect 10137 22729 10149 22732
rect 10183 22729 10195 22763
rect 13814 22760 13820 22772
rect 13775 22732 13820 22760
rect 10137 22723 10195 22729
rect 13814 22720 13820 22732
rect 13872 22720 13878 22772
rect 22281 22763 22339 22769
rect 22281 22729 22293 22763
rect 22327 22729 22339 22763
rect 22281 22723 22339 22729
rect 22649 22763 22707 22769
rect 22649 22729 22661 22763
rect 22695 22729 22707 22763
rect 22649 22723 22707 22729
rect 9180 22664 9352 22692
rect 9585 22695 9643 22701
rect 9180 22652 9186 22664
rect 9585 22661 9597 22695
rect 9631 22692 9643 22695
rect 9631 22664 10364 22692
rect 9631 22661 9643 22664
rect 9585 22655 9643 22661
rect 10336 22636 10364 22664
rect 12986 22652 12992 22704
rect 13044 22692 13050 22704
rect 13357 22695 13415 22701
rect 13357 22692 13369 22695
rect 13044 22664 13369 22692
rect 13044 22652 13050 22664
rect 13357 22661 13369 22664
rect 13403 22661 13415 22695
rect 13357 22655 13415 22661
rect 13998 22652 14004 22704
rect 14056 22692 14062 22704
rect 14093 22695 14151 22701
rect 14093 22692 14105 22695
rect 14056 22664 14105 22692
rect 14056 22652 14062 22664
rect 14093 22661 14105 22664
rect 14139 22661 14151 22695
rect 14093 22655 14151 22661
rect 14277 22695 14335 22701
rect 14277 22661 14289 22695
rect 14323 22692 14335 22695
rect 16666 22692 16672 22704
rect 14323 22664 16672 22692
rect 14323 22661 14335 22664
rect 14277 22655 14335 22661
rect 16666 22652 16672 22664
rect 16724 22652 16730 22704
rect 17126 22692 17132 22704
rect 17039 22664 17132 22692
rect 17126 22652 17132 22664
rect 17184 22692 17190 22704
rect 17497 22695 17555 22701
rect 17497 22692 17509 22695
rect 17184 22664 17509 22692
rect 17184 22652 17190 22664
rect 17497 22661 17509 22664
rect 17543 22661 17555 22695
rect 17497 22655 17555 22661
rect 17681 22695 17739 22701
rect 17681 22661 17693 22695
rect 17727 22692 17739 22695
rect 19150 22692 19156 22704
rect 17727 22664 19156 22692
rect 17727 22661 17739 22664
rect 17681 22655 17739 22661
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22593 7527 22627
rect 7469 22587 7527 22593
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 8294 22624 8300 22636
rect 8255 22596 8300 22624
rect 7561 22587 7619 22593
rect 7484 22556 7512 22587
rect 8294 22584 8300 22596
rect 8352 22584 8358 22636
rect 8662 22624 8668 22636
rect 8623 22596 8668 22624
rect 8662 22584 8668 22596
rect 8720 22584 8726 22636
rect 8757 22627 8815 22633
rect 8757 22593 8769 22627
rect 8803 22593 8815 22627
rect 8757 22587 8815 22593
rect 9401 22627 9459 22633
rect 9401 22593 9413 22627
rect 9447 22593 9459 22627
rect 9401 22587 9459 22593
rect 9861 22627 9919 22633
rect 9861 22593 9873 22627
rect 9907 22624 9919 22627
rect 10042 22624 10048 22636
rect 9907 22596 10048 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 8386 22556 8392 22568
rect 7484 22528 7696 22556
rect 8347 22528 8392 22556
rect 7193 22491 7251 22497
rect 7193 22457 7205 22491
rect 7239 22488 7251 22491
rect 7558 22488 7564 22500
rect 7239 22460 7564 22488
rect 7239 22457 7251 22460
rect 7193 22451 7251 22457
rect 7558 22448 7564 22460
rect 7616 22448 7622 22500
rect 7668 22488 7696 22528
rect 8386 22516 8392 22528
rect 8444 22556 8450 22568
rect 8772 22556 8800 22587
rect 8444 22528 8800 22556
rect 8444 22516 8450 22528
rect 8297 22491 8355 22497
rect 8297 22488 8309 22491
rect 7668 22460 8309 22488
rect 8297 22457 8309 22460
rect 8343 22488 8355 22491
rect 8570 22488 8576 22500
rect 8343 22460 8576 22488
rect 8343 22457 8355 22460
rect 8297 22451 8355 22457
rect 8570 22448 8576 22460
rect 8628 22448 8634 22500
rect 8662 22448 8668 22500
rect 8720 22488 8726 22500
rect 9416 22488 9444 22587
rect 10042 22584 10048 22596
rect 10100 22584 10106 22636
rect 10318 22624 10324 22636
rect 10231 22596 10324 22624
rect 10318 22584 10324 22596
rect 10376 22584 10382 22636
rect 11882 22584 11888 22636
rect 11940 22624 11946 22636
rect 16945 22627 17003 22633
rect 16945 22624 16957 22627
rect 11940 22596 16957 22624
rect 11940 22584 11946 22596
rect 16945 22593 16957 22596
rect 16991 22593 17003 22627
rect 16945 22587 17003 22593
rect 17221 22627 17279 22633
rect 17221 22593 17233 22627
rect 17267 22624 17279 22627
rect 17696 22624 17724 22655
rect 19150 22652 19156 22664
rect 19208 22652 19214 22704
rect 21450 22652 21456 22704
rect 21508 22692 21514 22704
rect 21821 22695 21879 22701
rect 21821 22692 21833 22695
rect 21508 22664 21833 22692
rect 21508 22652 21514 22664
rect 21821 22661 21833 22664
rect 21867 22661 21879 22695
rect 21821 22655 21879 22661
rect 18506 22624 18512 22636
rect 17267 22596 17724 22624
rect 18467 22596 18512 22624
rect 17267 22593 17279 22596
rect 17221 22587 17279 22593
rect 18506 22584 18512 22596
rect 18564 22584 18570 22636
rect 22296 22624 22324 22723
rect 22664 22692 22692 22723
rect 23566 22720 23572 22772
rect 23624 22760 23630 22772
rect 24121 22763 24179 22769
rect 24121 22760 24133 22763
rect 23624 22732 24133 22760
rect 23624 22720 23630 22732
rect 24121 22729 24133 22732
rect 24167 22729 24179 22763
rect 24121 22723 24179 22729
rect 22986 22695 23044 22701
rect 22986 22692 22998 22695
rect 22664 22664 22998 22692
rect 22986 22661 22998 22664
rect 23032 22661 23044 22695
rect 22986 22655 23044 22661
rect 22465 22627 22523 22633
rect 22465 22624 22477 22627
rect 22296 22596 22477 22624
rect 22465 22593 22477 22596
rect 22511 22593 22523 22627
rect 22738 22624 22744 22636
rect 22699 22596 22744 22624
rect 22465 22587 22523 22593
rect 22738 22584 22744 22596
rect 22796 22584 22802 22636
rect 10060 22556 10088 22584
rect 10410 22556 10416 22568
rect 10060 22528 10416 22556
rect 10410 22516 10416 22528
rect 10468 22516 10474 22568
rect 15286 22516 15292 22568
rect 15344 22556 15350 22568
rect 16206 22556 16212 22568
rect 15344 22528 16212 22556
rect 15344 22516 15350 22528
rect 16206 22516 16212 22528
rect 16264 22516 16270 22568
rect 9769 22491 9827 22497
rect 9769 22488 9781 22491
rect 8720 22460 9781 22488
rect 8720 22448 8726 22460
rect 9769 22457 9781 22460
rect 9815 22457 9827 22491
rect 9769 22451 9827 22457
rect 13725 22491 13783 22497
rect 13725 22457 13737 22491
rect 13771 22488 13783 22491
rect 14090 22488 14096 22500
rect 13771 22460 14096 22488
rect 13771 22457 13783 22460
rect 13725 22451 13783 22457
rect 14090 22448 14096 22460
rect 14148 22448 14154 22500
rect 15933 22491 15991 22497
rect 15933 22457 15945 22491
rect 15979 22488 15991 22491
rect 16666 22488 16672 22500
rect 15979 22460 16672 22488
rect 15979 22457 15991 22460
rect 15933 22451 15991 22457
rect 16666 22448 16672 22460
rect 16724 22448 16730 22500
rect 17310 22488 17316 22500
rect 17271 22460 17316 22488
rect 17310 22448 17316 22460
rect 17368 22448 17374 22500
rect 22189 22491 22247 22497
rect 22189 22457 22201 22491
rect 22235 22488 22247 22491
rect 22278 22488 22284 22500
rect 22235 22460 22284 22488
rect 22235 22457 22247 22460
rect 22189 22451 22247 22457
rect 22278 22448 22284 22460
rect 22336 22448 22342 22500
rect 4706 22420 4712 22432
rect 4667 22392 4712 22420
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 5626 22380 5632 22432
rect 5684 22420 5690 22432
rect 6086 22420 6092 22432
rect 5684 22392 6092 22420
rect 5684 22380 5690 22392
rect 6086 22380 6092 22392
rect 6144 22380 6150 22432
rect 7006 22380 7012 22432
rect 7064 22420 7070 22432
rect 7285 22423 7343 22429
rect 7285 22420 7297 22423
rect 7064 22392 7297 22420
rect 7064 22380 7070 22392
rect 7285 22389 7297 22392
rect 7331 22389 7343 22423
rect 7285 22383 7343 22389
rect 7745 22423 7803 22429
rect 7745 22389 7757 22423
rect 7791 22420 7803 22423
rect 8110 22420 8116 22432
rect 7791 22392 8116 22420
rect 7791 22389 7803 22392
rect 7745 22383 7803 22389
rect 8110 22380 8116 22392
rect 8168 22380 8174 22432
rect 8849 22423 8907 22429
rect 8849 22389 8861 22423
rect 8895 22420 8907 22423
rect 8938 22420 8944 22432
rect 8895 22392 8944 22420
rect 8895 22389 8907 22392
rect 8849 22383 8907 22389
rect 8938 22380 8944 22392
rect 8996 22380 9002 22432
rect 15470 22380 15476 22432
rect 15528 22420 15534 22432
rect 15749 22423 15807 22429
rect 15749 22420 15761 22423
rect 15528 22392 15761 22420
rect 15528 22380 15534 22392
rect 15749 22389 15761 22392
rect 15795 22389 15807 22423
rect 16758 22420 16764 22432
rect 16719 22392 16764 22420
rect 15749 22383 15807 22389
rect 16758 22380 16764 22392
rect 16816 22380 16822 22432
rect 18322 22420 18328 22432
rect 18283 22392 18328 22420
rect 18322 22380 18328 22392
rect 18380 22380 18386 22432
rect 1104 22330 26220 22352
rect 1104 22278 5136 22330
rect 5188 22278 5200 22330
rect 5252 22278 5264 22330
rect 5316 22278 5328 22330
rect 5380 22278 5392 22330
rect 5444 22278 13508 22330
rect 13560 22278 13572 22330
rect 13624 22278 13636 22330
rect 13688 22278 13700 22330
rect 13752 22278 13764 22330
rect 13816 22278 21880 22330
rect 21932 22278 21944 22330
rect 21996 22278 22008 22330
rect 22060 22278 22072 22330
rect 22124 22278 22136 22330
rect 22188 22278 26220 22330
rect 1104 22256 26220 22278
rect 4338 22216 4344 22228
rect 4299 22188 4344 22216
rect 4338 22176 4344 22188
rect 4396 22176 4402 22228
rect 7098 22176 7104 22228
rect 7156 22216 7162 22228
rect 9766 22216 9772 22228
rect 7156 22188 9772 22216
rect 7156 22176 7162 22188
rect 9766 22176 9772 22188
rect 9824 22176 9830 22228
rect 11241 22219 11299 22225
rect 11241 22185 11253 22219
rect 11287 22185 11299 22219
rect 17126 22216 17132 22228
rect 17087 22188 17132 22216
rect 11241 22179 11299 22185
rect 6086 22108 6092 22160
rect 6144 22148 6150 22160
rect 7742 22148 7748 22160
rect 6144 22120 7748 22148
rect 6144 22108 6150 22120
rect 7742 22108 7748 22120
rect 7800 22108 7806 22160
rect 3970 22040 3976 22092
rect 4028 22040 4034 22092
rect 6914 22080 6920 22092
rect 6875 22052 6920 22080
rect 6914 22040 6920 22052
rect 6972 22040 6978 22092
rect 8757 22083 8815 22089
rect 8757 22049 8769 22083
rect 8803 22080 8815 22083
rect 9306 22080 9312 22092
rect 8803 22052 9312 22080
rect 8803 22049 8815 22052
rect 8757 22043 8815 22049
rect 9306 22040 9312 22052
rect 9364 22080 9370 22092
rect 9493 22083 9551 22089
rect 9493 22080 9505 22083
rect 9364 22052 9505 22080
rect 9364 22040 9370 22052
rect 9493 22049 9505 22052
rect 9539 22049 9551 22083
rect 11256 22080 11284 22179
rect 17126 22176 17132 22188
rect 17184 22176 17190 22228
rect 22278 22216 22284 22228
rect 22239 22188 22284 22216
rect 22278 22176 22284 22188
rect 22336 22176 22342 22228
rect 23474 22216 23480 22228
rect 23435 22188 23480 22216
rect 23474 22176 23480 22188
rect 23532 22176 23538 22228
rect 12342 22080 12348 22092
rect 11256 22052 12112 22080
rect 12303 22052 12348 22080
rect 9493 22043 9551 22049
rect 1486 21972 1492 22024
rect 1544 22012 1550 22024
rect 1949 22015 2007 22021
rect 1949 22012 1961 22015
rect 1544 21984 1961 22012
rect 1544 21972 1550 21984
rect 1949 21981 1961 21984
rect 1995 22012 2007 22015
rect 3326 22012 3332 22024
rect 1995 21984 3332 22012
rect 1995 21981 2007 21984
rect 1949 21975 2007 21981
rect 3326 21972 3332 21984
rect 3384 21972 3390 22024
rect 3418 21972 3424 22024
rect 3476 22012 3482 22024
rect 3789 22015 3847 22021
rect 3789 22012 3801 22015
rect 3476 21984 3801 22012
rect 3476 21972 3482 21984
rect 3789 21981 3801 21984
rect 3835 21981 3847 22015
rect 3988 22012 4016 22040
rect 4162 22015 4220 22021
rect 4162 22012 4174 22015
rect 3988 21984 4174 22012
rect 3789 21975 3847 21981
rect 4162 21981 4174 21984
rect 4208 21981 4220 22015
rect 4162 21975 4220 21981
rect 8846 21972 8852 22024
rect 8904 22012 8910 22024
rect 8941 22015 8999 22021
rect 8941 22012 8953 22015
rect 8904 21984 8953 22012
rect 8904 21972 8910 21984
rect 8941 21981 8953 21984
rect 8987 21981 8999 22015
rect 8941 21975 8999 21981
rect 9033 22015 9091 22021
rect 9033 21981 9045 22015
rect 9079 22012 9091 22015
rect 9122 22012 9128 22024
rect 9079 21984 9128 22012
rect 9079 21981 9091 21984
rect 9033 21975 9091 21981
rect 9122 21972 9128 21984
rect 9180 22012 9186 22024
rect 9217 22015 9275 22021
rect 9217 22012 9229 22015
rect 9180 21984 9229 22012
rect 9180 21972 9186 21984
rect 9217 21981 9229 21984
rect 9263 21981 9275 22015
rect 10042 22012 10048 22024
rect 9217 21975 9275 21981
rect 9646 21984 10048 22012
rect 2216 21947 2274 21953
rect 2216 21913 2228 21947
rect 2262 21944 2274 21947
rect 2682 21944 2688 21956
rect 2262 21916 2688 21944
rect 2262 21913 2274 21916
rect 2216 21907 2274 21913
rect 2682 21904 2688 21916
rect 2740 21904 2746 21956
rect 3694 21904 3700 21956
rect 3752 21944 3758 21956
rect 3973 21947 4031 21953
rect 3973 21944 3985 21947
rect 3752 21916 3985 21944
rect 3752 21904 3758 21916
rect 3973 21913 3985 21916
rect 4019 21913 4031 21947
rect 3973 21907 4031 21913
rect 4065 21947 4123 21953
rect 4065 21913 4077 21947
rect 4111 21944 4123 21947
rect 4706 21944 4712 21956
rect 4111 21916 4712 21944
rect 4111 21913 4123 21916
rect 4065 21907 4123 21913
rect 4706 21904 4712 21916
rect 4764 21904 4770 21956
rect 7101 21947 7159 21953
rect 7101 21913 7113 21947
rect 7147 21944 7159 21947
rect 7650 21944 7656 21956
rect 7147 21916 7656 21944
rect 7147 21913 7159 21916
rect 7101 21907 7159 21913
rect 7650 21904 7656 21916
rect 7708 21904 7714 21956
rect 8294 21904 8300 21956
rect 8352 21944 8358 21956
rect 8490 21947 8548 21953
rect 8490 21944 8502 21947
rect 8352 21916 8502 21944
rect 8352 21904 8358 21916
rect 8490 21913 8502 21916
rect 8536 21913 8548 21947
rect 9646 21944 9674 21984
rect 10042 21972 10048 21984
rect 10100 21972 10106 22024
rect 10318 21972 10324 22024
rect 10376 22012 10382 22024
rect 11057 22015 11115 22021
rect 11057 22012 11069 22015
rect 10376 21984 11069 22012
rect 10376 21972 10382 21984
rect 11057 21981 11069 21984
rect 11103 21981 11115 22015
rect 11057 21975 11115 21981
rect 11146 21972 11152 22024
rect 11204 22012 11210 22024
rect 11701 22015 11759 22021
rect 11701 22012 11713 22015
rect 11204 21984 11713 22012
rect 11204 21972 11210 21984
rect 11701 21981 11713 21984
rect 11747 22012 11759 22015
rect 11793 22015 11851 22021
rect 11793 22012 11805 22015
rect 11747 21984 11805 22012
rect 11747 21981 11759 21984
rect 11701 21975 11759 21981
rect 11793 21981 11805 21984
rect 11839 21981 11851 22015
rect 11793 21975 11851 21981
rect 11882 21972 11888 22024
rect 11940 22012 11946 22024
rect 11977 22015 12035 22021
rect 11977 22012 11989 22015
rect 11940 21984 11989 22012
rect 11940 21972 11946 21984
rect 11977 21981 11989 21984
rect 12023 21981 12035 22015
rect 12084 22012 12112 22052
rect 12342 22040 12348 22052
rect 12400 22080 12406 22092
rect 12434 22080 12440 22092
rect 12400 22052 12440 22080
rect 12400 22040 12406 22052
rect 12434 22040 12440 22052
rect 12492 22040 12498 22092
rect 12544 22052 12756 22080
rect 12544 22021 12572 22052
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 12084 21984 12541 22012
rect 11977 21975 12035 21981
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 12621 22015 12679 22021
rect 12621 21981 12633 22015
rect 12667 21981 12679 22015
rect 12728 22012 12756 22052
rect 13998 22040 14004 22092
rect 14056 22080 14062 22092
rect 15010 22080 15016 22092
rect 14056 22052 15016 22080
rect 14056 22040 14062 22052
rect 15010 22040 15016 22052
rect 15068 22080 15074 22092
rect 15749 22083 15807 22089
rect 15749 22080 15761 22083
rect 15068 22052 15761 22080
rect 15068 22040 15074 22052
rect 15749 22049 15761 22052
rect 15795 22049 15807 22083
rect 15749 22043 15807 22049
rect 22189 22083 22247 22089
rect 22189 22049 22201 22083
rect 22235 22080 22247 22083
rect 22830 22080 22836 22092
rect 22235 22052 22836 22080
rect 22235 22049 22247 22052
rect 22189 22043 22247 22049
rect 22830 22040 22836 22052
rect 22888 22040 22894 22092
rect 15286 22012 15292 22024
rect 12728 21984 15292 22012
rect 12621 21975 12679 21981
rect 8490 21907 8548 21913
rect 9416 21916 9674 21944
rect 9760 21947 9818 21953
rect 3326 21876 3332 21888
rect 3287 21848 3332 21876
rect 3326 21836 3332 21848
rect 3384 21836 3390 21888
rect 7377 21879 7435 21885
rect 7377 21845 7389 21879
rect 7423 21876 7435 21879
rect 8386 21876 8392 21888
rect 7423 21848 8392 21876
rect 7423 21845 7435 21848
rect 7377 21839 7435 21845
rect 8386 21836 8392 21848
rect 8444 21836 8450 21888
rect 9122 21836 9128 21888
rect 9180 21876 9186 21888
rect 9416 21885 9444 21916
rect 9760 21913 9772 21947
rect 9806 21913 9818 21947
rect 12253 21947 12311 21953
rect 9760 21907 9818 21913
rect 10888 21916 12020 21944
rect 9401 21879 9459 21885
rect 9401 21876 9413 21879
rect 9180 21848 9413 21876
rect 9180 21836 9186 21848
rect 9401 21845 9413 21848
rect 9447 21845 9459 21879
rect 9401 21839 9459 21845
rect 9674 21836 9680 21888
rect 9732 21876 9738 21888
rect 9784 21876 9812 21907
rect 10888 21885 10916 21916
rect 11992 21888 12020 21916
rect 12253 21913 12265 21947
rect 12299 21944 12311 21947
rect 12636 21944 12664 21975
rect 15286 21972 15292 21984
rect 15344 21972 15350 22024
rect 15470 22012 15476 22024
rect 15431 21984 15476 22012
rect 15470 21972 15476 21984
rect 15528 21972 15534 22024
rect 17310 22012 17316 22024
rect 17271 21984 17316 22012
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 17589 22015 17647 22021
rect 17589 21981 17601 22015
rect 17635 22012 17647 22015
rect 19242 22012 19248 22024
rect 17635 21984 19248 22012
rect 17635 21981 17647 21984
rect 17589 21975 17647 21981
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 22741 22015 22799 22021
rect 22741 21981 22753 22015
rect 22787 22012 22799 22015
rect 23014 22012 23020 22024
rect 22787 21984 23020 22012
rect 22787 21981 22799 21984
rect 22741 21975 22799 21981
rect 23014 21972 23020 21984
rect 23072 21972 23078 22024
rect 23566 22012 23572 22024
rect 23527 21984 23572 22012
rect 23566 21972 23572 21984
rect 23624 21972 23630 22024
rect 23753 22015 23811 22021
rect 23753 21981 23765 22015
rect 23799 22012 23811 22015
rect 24026 22012 24032 22024
rect 23799 21984 24032 22012
rect 23799 21981 23811 21984
rect 23753 21975 23811 21981
rect 24026 21972 24032 21984
rect 24084 21972 24090 22024
rect 15994 21947 16052 21953
rect 15994 21944 16006 21947
rect 12299 21916 12664 21944
rect 15672 21916 16006 21944
rect 12299 21913 12311 21916
rect 12253 21907 12311 21913
rect 9732 21848 9812 21876
rect 10873 21879 10931 21885
rect 9732 21836 9738 21848
rect 10873 21845 10885 21879
rect 10919 21845 10931 21879
rect 10873 21839 10931 21845
rect 11974 21836 11980 21888
rect 12032 21836 12038 21888
rect 12710 21876 12716 21888
rect 12671 21848 12716 21876
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 15672 21885 15700 21916
rect 15994 21913 16006 21916
rect 16040 21913 16052 21947
rect 15994 21907 16052 21913
rect 17856 21947 17914 21953
rect 17856 21913 17868 21947
rect 17902 21944 17914 21947
rect 18322 21944 18328 21956
rect 17902 21916 18328 21944
rect 17902 21913 17914 21916
rect 17856 21907 17914 21913
rect 18322 21904 18328 21916
rect 18380 21904 18386 21956
rect 19058 21904 19064 21956
rect 19116 21944 19122 21956
rect 19490 21947 19548 21953
rect 19490 21944 19502 21947
rect 19116 21916 19502 21944
rect 19116 21904 19122 21916
rect 19490 21913 19502 21916
rect 19536 21913 19548 21947
rect 19490 21907 19548 21913
rect 15657 21879 15715 21885
rect 15657 21845 15669 21879
rect 15703 21845 15715 21879
rect 17494 21876 17500 21888
rect 17455 21848 17500 21876
rect 15657 21839 15715 21845
rect 17494 21836 17500 21848
rect 17552 21836 17558 21888
rect 18969 21879 19027 21885
rect 18969 21845 18981 21879
rect 19015 21876 19027 21879
rect 19242 21876 19248 21888
rect 19015 21848 19248 21876
rect 19015 21845 19027 21848
rect 18969 21839 19027 21845
rect 19242 21836 19248 21848
rect 19300 21836 19306 21888
rect 19334 21836 19340 21888
rect 19392 21876 19398 21888
rect 20070 21876 20076 21888
rect 19392 21848 20076 21876
rect 19392 21836 19398 21848
rect 20070 21836 20076 21848
rect 20128 21876 20134 21888
rect 20625 21879 20683 21885
rect 20625 21876 20637 21879
rect 20128 21848 20637 21876
rect 20128 21836 20134 21848
rect 20625 21845 20637 21848
rect 20671 21845 20683 21879
rect 22646 21876 22652 21888
rect 22607 21848 22652 21876
rect 20625 21839 20683 21845
rect 22646 21836 22652 21848
rect 22704 21836 22710 21888
rect 1104 21786 26220 21808
rect 1104 21734 9322 21786
rect 9374 21734 9386 21786
rect 9438 21734 9450 21786
rect 9502 21734 9514 21786
rect 9566 21734 9578 21786
rect 9630 21734 17694 21786
rect 17746 21734 17758 21786
rect 17810 21734 17822 21786
rect 17874 21734 17886 21786
rect 17938 21734 17950 21786
rect 18002 21734 26220 21786
rect 1104 21712 26220 21734
rect 2682 21672 2688 21684
rect 2643 21644 2688 21672
rect 2682 21632 2688 21644
rect 2740 21632 2746 21684
rect 3694 21672 3700 21684
rect 3655 21644 3700 21672
rect 3694 21632 3700 21644
rect 3752 21632 3758 21684
rect 7926 21632 7932 21684
rect 7984 21672 7990 21684
rect 8573 21675 8631 21681
rect 8573 21672 8585 21675
rect 7984 21644 8585 21672
rect 7984 21632 7990 21644
rect 8573 21641 8585 21644
rect 8619 21641 8631 21675
rect 8573 21635 8631 21641
rect 9493 21675 9551 21681
rect 9493 21641 9505 21675
rect 9539 21672 9551 21675
rect 9674 21672 9680 21684
rect 9539 21644 9680 21672
rect 9539 21641 9551 21644
rect 9493 21635 9551 21641
rect 3326 21604 3332 21616
rect 3239 21576 3332 21604
rect 2866 21536 2872 21548
rect 2827 21508 2872 21536
rect 2866 21496 2872 21508
rect 2924 21496 2930 21548
rect 2958 21496 2964 21548
rect 3016 21536 3022 21548
rect 3252 21545 3280 21576
rect 3326 21564 3332 21576
rect 3384 21604 3390 21616
rect 4065 21607 4123 21613
rect 4065 21604 4077 21607
rect 3384 21576 4077 21604
rect 3384 21564 3390 21576
rect 4065 21573 4077 21576
rect 4111 21573 4123 21607
rect 8588 21604 8616 21635
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 10413 21675 10471 21681
rect 10413 21672 10425 21675
rect 10100 21644 10425 21672
rect 10100 21632 10106 21644
rect 10413 21641 10425 21644
rect 10459 21672 10471 21675
rect 11146 21672 11152 21684
rect 10459 21644 11152 21672
rect 10459 21641 10471 21644
rect 10413 21635 10471 21641
rect 11146 21632 11152 21644
rect 11204 21632 11210 21684
rect 11609 21675 11667 21681
rect 11609 21641 11621 21675
rect 11655 21672 11667 21675
rect 12342 21672 12348 21684
rect 11655 21644 12348 21672
rect 11655 21641 11667 21644
rect 11609 21635 11667 21641
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 12434 21632 12440 21684
rect 12492 21672 12498 21684
rect 14182 21672 14188 21684
rect 12492 21644 14188 21672
rect 12492 21632 12498 21644
rect 14182 21632 14188 21644
rect 14240 21632 14246 21684
rect 16666 21672 16672 21684
rect 16627 21644 16672 21672
rect 16666 21632 16672 21644
rect 16724 21632 16730 21684
rect 16758 21632 16764 21684
rect 16816 21672 16822 21684
rect 17129 21675 17187 21681
rect 17129 21672 17141 21675
rect 16816 21644 17141 21672
rect 16816 21632 16822 21644
rect 17129 21641 17141 21644
rect 17175 21641 17187 21675
rect 17129 21635 17187 21641
rect 17957 21675 18015 21681
rect 17957 21641 17969 21675
rect 18003 21672 18015 21675
rect 18506 21672 18512 21684
rect 18003 21644 18512 21672
rect 18003 21641 18015 21644
rect 17957 21635 18015 21641
rect 18506 21632 18512 21644
rect 18564 21632 18570 21684
rect 18601 21675 18659 21681
rect 18601 21641 18613 21675
rect 18647 21672 18659 21675
rect 20809 21675 20867 21681
rect 20809 21672 20821 21675
rect 18647 21644 20821 21672
rect 18647 21641 18659 21644
rect 18601 21635 18659 21641
rect 20809 21641 20821 21644
rect 20855 21641 20867 21675
rect 20809 21635 20867 21641
rect 21468 21644 22416 21672
rect 9769 21607 9827 21613
rect 8588 21576 9720 21604
rect 4065 21567 4123 21573
rect 3237 21539 3295 21545
rect 3016 21508 3061 21536
rect 3016 21496 3022 21508
rect 3237 21505 3249 21539
rect 3283 21505 3295 21539
rect 3237 21499 3295 21505
rect 3513 21539 3571 21545
rect 3513 21505 3525 21539
rect 3559 21536 3571 21539
rect 3559 21508 3740 21536
rect 3559 21505 3571 21508
rect 3513 21499 3571 21505
rect 3712 21400 3740 21508
rect 8662 21496 8668 21548
rect 8720 21536 8726 21548
rect 8757 21539 8815 21545
rect 8757 21536 8769 21539
rect 8720 21508 8769 21536
rect 8720 21496 8726 21508
rect 8757 21505 8769 21508
rect 8803 21505 8815 21539
rect 8757 21499 8815 21505
rect 8846 21496 8852 21548
rect 8904 21536 8910 21548
rect 8904 21508 8949 21536
rect 8904 21496 8910 21508
rect 9030 21496 9036 21548
rect 9088 21536 9094 21548
rect 9692 21545 9720 21576
rect 9769 21573 9781 21607
rect 9815 21604 9827 21607
rect 9858 21604 9864 21616
rect 9815 21576 9864 21604
rect 9815 21573 9827 21576
rect 9769 21567 9827 21573
rect 9858 21564 9864 21576
rect 9916 21564 9922 21616
rect 11882 21604 11888 21616
rect 10060 21576 11888 21604
rect 9677 21539 9735 21545
rect 9088 21508 9133 21536
rect 9088 21496 9094 21508
rect 9677 21505 9689 21539
rect 9723 21536 9735 21539
rect 10060 21536 10088 21576
rect 11882 21564 11888 21576
rect 11940 21564 11946 21616
rect 12710 21564 12716 21616
rect 12768 21613 12774 21616
rect 12768 21604 12780 21613
rect 12768 21576 12813 21604
rect 12768 21567 12780 21576
rect 12768 21564 12774 21567
rect 16206 21564 16212 21616
rect 16264 21604 16270 21616
rect 17497 21607 17555 21613
rect 17497 21604 17509 21607
rect 16264 21576 17509 21604
rect 16264 21564 16270 21576
rect 17497 21573 17509 21576
rect 17543 21573 17555 21607
rect 17497 21567 17555 21573
rect 19260 21576 20484 21604
rect 10226 21536 10232 21548
rect 9723 21508 10088 21536
rect 10139 21508 10232 21536
rect 9723 21505 9735 21508
rect 9677 21499 9735 21505
rect 10226 21496 10232 21508
rect 10284 21536 10290 21548
rect 11974 21536 11980 21548
rect 10284 21508 11980 21536
rect 10284 21496 10290 21508
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21536 13047 21539
rect 13998 21536 14004 21548
rect 13035 21508 14004 21536
rect 13035 21505 13047 21508
rect 12989 21499 13047 21505
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 15280 21539 15338 21545
rect 15280 21505 15292 21539
rect 15326 21536 15338 21539
rect 16114 21536 16120 21548
rect 15326 21508 16120 21536
rect 15326 21505 15338 21508
rect 15280 21499 15338 21505
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21536 17095 21539
rect 17126 21536 17132 21548
rect 17083 21508 17132 21536
rect 17083 21505 17095 21508
rect 17037 21499 17095 21505
rect 17126 21496 17132 21508
rect 17184 21496 17190 21548
rect 18322 21496 18328 21548
rect 18380 21536 18386 21548
rect 18509 21539 18567 21545
rect 18509 21536 18521 21539
rect 18380 21508 18521 21536
rect 18380 21496 18386 21508
rect 18509 21505 18521 21508
rect 18555 21505 18567 21539
rect 19150 21536 19156 21548
rect 19063 21508 19156 21536
rect 18509 21499 18567 21505
rect 4154 21468 4160 21480
rect 4115 21440 4160 21468
rect 4154 21428 4160 21440
rect 4212 21428 4218 21480
rect 4249 21471 4307 21477
rect 4249 21437 4261 21471
rect 4295 21468 4307 21471
rect 9953 21471 10011 21477
rect 4295 21440 4476 21468
rect 4295 21437 4307 21440
rect 4249 21431 4307 21437
rect 4448 21412 4476 21440
rect 9953 21437 9965 21471
rect 9999 21437 10011 21471
rect 15010 21468 15016 21480
rect 14971 21440 15016 21468
rect 9953 21431 10011 21437
rect 3160 21372 3740 21400
rect 3160 21344 3188 21372
rect 4430 21360 4436 21412
rect 4488 21400 4494 21412
rect 4709 21403 4767 21409
rect 4709 21400 4721 21403
rect 4488 21372 4721 21400
rect 4488 21360 4494 21372
rect 4709 21369 4721 21372
rect 4755 21400 4767 21403
rect 4893 21403 4951 21409
rect 4893 21400 4905 21403
rect 4755 21372 4905 21400
rect 4755 21369 4767 21372
rect 4709 21363 4767 21369
rect 4893 21369 4905 21372
rect 4939 21400 4951 21403
rect 9122 21400 9128 21412
rect 4939 21372 9128 21400
rect 4939 21369 4951 21372
rect 4893 21363 4951 21369
rect 9122 21360 9128 21372
rect 9180 21360 9186 21412
rect 9217 21403 9275 21409
rect 9217 21369 9229 21403
rect 9263 21400 9275 21403
rect 9968 21400 9996 21431
rect 15010 21428 15016 21440
rect 15068 21428 15074 21480
rect 17313 21471 17371 21477
rect 17313 21437 17325 21471
rect 17359 21468 17371 21471
rect 17494 21468 17500 21480
rect 17359 21440 17500 21468
rect 17359 21437 17371 21440
rect 17313 21431 17371 21437
rect 17494 21428 17500 21440
rect 17552 21468 17558 21480
rect 18693 21471 18751 21477
rect 18693 21468 18705 21471
rect 17552 21440 18705 21468
rect 17552 21428 17558 21440
rect 18693 21437 18705 21440
rect 18739 21468 18751 21471
rect 18874 21468 18880 21480
rect 18739 21440 18880 21468
rect 18739 21437 18751 21440
rect 18693 21431 18751 21437
rect 18874 21428 18880 21440
rect 18932 21428 18938 21480
rect 9263 21372 9996 21400
rect 9263 21369 9275 21372
rect 9217 21363 9275 21369
rect 10042 21360 10048 21412
rect 10100 21400 10106 21412
rect 19076 21409 19104 21508
rect 19150 21496 19156 21508
rect 19208 21536 19214 21548
rect 19260 21536 19288 21576
rect 19426 21536 19432 21548
rect 19208 21508 19288 21536
rect 19387 21508 19432 21536
rect 19208 21496 19214 21508
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 19702 21496 19708 21548
rect 19760 21536 19766 21548
rect 20252 21540 20310 21545
rect 20180 21539 20310 21540
rect 20180 21536 20264 21539
rect 19760 21512 20264 21536
rect 19760 21508 20208 21512
rect 19760 21496 19766 21508
rect 20252 21505 20264 21512
rect 20298 21505 20310 21539
rect 20456 21536 20484 21576
rect 20659 21539 20717 21545
rect 20659 21536 20671 21539
rect 20456 21508 20671 21536
rect 20252 21499 20310 21505
rect 20659 21505 20671 21508
rect 20705 21505 20717 21539
rect 20659 21499 20717 21505
rect 21358 21496 21364 21548
rect 21416 21536 21422 21548
rect 21468 21545 21496 21644
rect 21560 21576 21772 21604
rect 21453 21539 21511 21545
rect 21453 21536 21465 21539
rect 21416 21508 21465 21536
rect 21416 21496 21422 21508
rect 21453 21505 21465 21508
rect 21499 21505 21511 21539
rect 21453 21499 21511 21505
rect 19242 21428 19248 21480
rect 19300 21468 19306 21480
rect 19337 21471 19395 21477
rect 19337 21468 19349 21471
rect 19300 21440 19349 21468
rect 19300 21428 19306 21440
rect 19337 21437 19349 21440
rect 19383 21468 19395 21471
rect 20070 21468 20076 21480
rect 19383 21440 19840 21468
rect 20031 21440 20076 21468
rect 19383 21437 19395 21440
rect 19337 21431 19395 21437
rect 17865 21403 17923 21409
rect 10100 21372 10145 21400
rect 10100 21360 10106 21372
rect 17865 21369 17877 21403
rect 17911 21400 17923 21403
rect 18141 21403 18199 21409
rect 18141 21400 18153 21403
rect 17911 21372 18153 21400
rect 17911 21369 17923 21372
rect 17865 21363 17923 21369
rect 18141 21369 18153 21372
rect 18187 21369 18199 21403
rect 18141 21363 18199 21369
rect 19061 21403 19119 21409
rect 19061 21369 19073 21403
rect 19107 21369 19119 21403
rect 19812 21400 19840 21440
rect 20070 21428 20076 21440
rect 20128 21428 20134 21480
rect 20162 21428 20168 21480
rect 20220 21468 20226 21480
rect 20368 21471 20426 21477
rect 20220 21440 20265 21468
rect 20220 21428 20226 21440
rect 20368 21437 20380 21471
rect 20414 21468 20426 21471
rect 21266 21468 21272 21480
rect 20414 21440 20484 21468
rect 21179 21440 21272 21468
rect 20414 21437 20426 21440
rect 20368 21431 20426 21437
rect 20456 21400 20484 21440
rect 21266 21428 21272 21440
rect 21324 21468 21330 21480
rect 21560 21468 21588 21576
rect 21637 21539 21695 21545
rect 21637 21505 21649 21539
rect 21683 21505 21695 21539
rect 21744 21536 21772 21576
rect 21818 21564 21824 21616
rect 21876 21604 21882 21616
rect 22278 21604 22284 21616
rect 21876 21576 22284 21604
rect 21876 21564 21882 21576
rect 22278 21564 22284 21576
rect 22336 21564 22342 21616
rect 22388 21545 22416 21644
rect 22006 21539 22064 21545
rect 22006 21536 22018 21539
rect 21744 21508 22018 21536
rect 21637 21499 21695 21505
rect 22006 21505 22018 21508
rect 22052 21505 22064 21539
rect 22006 21499 22064 21505
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21505 22431 21539
rect 22554 21536 22560 21548
rect 22515 21508 22560 21536
rect 22373 21499 22431 21505
rect 21324 21440 21588 21468
rect 21652 21468 21680 21499
rect 22554 21496 22560 21508
rect 22612 21496 22618 21548
rect 23075 21539 23133 21545
rect 23075 21536 23087 21539
rect 22756 21508 23087 21536
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 21652 21440 22477 21468
rect 21324 21428 21330 21440
rect 22465 21437 22477 21440
rect 22511 21468 22523 21471
rect 22756 21468 22784 21508
rect 23075 21505 23087 21508
rect 23121 21536 23133 21539
rect 23198 21536 23204 21548
rect 23121 21508 23204 21536
rect 23121 21505 23133 21508
rect 23075 21499 23133 21505
rect 23198 21496 23204 21508
rect 23256 21496 23262 21548
rect 23474 21536 23480 21548
rect 23435 21508 23480 21536
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 22511 21440 22784 21468
rect 22511 21437 22523 21440
rect 22465 21431 22523 21437
rect 23290 21428 23296 21480
rect 23348 21468 23354 21480
rect 23385 21471 23443 21477
rect 23385 21468 23397 21471
rect 23348 21440 23397 21468
rect 23348 21428 23354 21440
rect 23385 21437 23397 21440
rect 23431 21437 23443 21471
rect 23385 21431 23443 21437
rect 19061 21363 19119 21369
rect 19168 21372 19748 21400
rect 19812 21372 20484 21400
rect 3142 21332 3148 21344
rect 3103 21304 3148 21332
rect 3142 21292 3148 21304
rect 3200 21292 3206 21344
rect 3326 21332 3332 21344
rect 3287 21304 3332 21332
rect 3326 21292 3332 21304
rect 3384 21292 3390 21344
rect 7377 21335 7435 21341
rect 7377 21301 7389 21335
rect 7423 21332 7435 21335
rect 7650 21332 7656 21344
rect 7423 21304 7656 21332
rect 7423 21301 7435 21304
rect 7377 21295 7435 21301
rect 7650 21292 7656 21304
rect 7708 21292 7714 21344
rect 8938 21332 8944 21344
rect 8899 21304 8944 21332
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 16022 21292 16028 21344
rect 16080 21332 16086 21344
rect 16393 21335 16451 21341
rect 16393 21332 16405 21335
rect 16080 21304 16405 21332
rect 16080 21292 16086 21304
rect 16393 21301 16405 21304
rect 16439 21332 16451 21335
rect 19168 21332 19196 21372
rect 19334 21332 19340 21344
rect 16439 21304 19196 21332
rect 19295 21304 19340 21332
rect 16439 21301 16451 21304
rect 16393 21295 16451 21301
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 19610 21332 19616 21344
rect 19571 21304 19616 21332
rect 19610 21292 19616 21304
rect 19668 21292 19674 21344
rect 19720 21332 19748 21372
rect 21450 21360 21456 21412
rect 21508 21400 21514 21412
rect 21821 21403 21879 21409
rect 21821 21400 21833 21403
rect 21508 21372 21833 21400
rect 21508 21360 21514 21372
rect 21821 21369 21833 21372
rect 21867 21369 21879 21403
rect 21821 21363 21879 21369
rect 21634 21332 21640 21344
rect 19720 21304 21640 21332
rect 21634 21292 21640 21304
rect 21692 21292 21698 21344
rect 22741 21335 22799 21341
rect 22741 21301 22753 21335
rect 22787 21332 22799 21335
rect 22830 21332 22836 21344
rect 22787 21304 22836 21332
rect 22787 21301 22799 21304
rect 22741 21295 22799 21301
rect 22830 21292 22836 21304
rect 22888 21292 22894 21344
rect 22922 21292 22928 21344
rect 22980 21332 22986 21344
rect 22980 21304 23025 21332
rect 22980 21292 22986 21304
rect 1104 21242 26220 21264
rect 1104 21190 5136 21242
rect 5188 21190 5200 21242
rect 5252 21190 5264 21242
rect 5316 21190 5328 21242
rect 5380 21190 5392 21242
rect 5444 21190 13508 21242
rect 13560 21190 13572 21242
rect 13624 21190 13636 21242
rect 13688 21190 13700 21242
rect 13752 21190 13764 21242
rect 13816 21190 21880 21242
rect 21932 21190 21944 21242
rect 21996 21190 22008 21242
rect 22060 21190 22072 21242
rect 22124 21190 22136 21242
rect 22188 21190 26220 21242
rect 1104 21168 26220 21190
rect 2866 21088 2872 21140
rect 2924 21128 2930 21140
rect 3789 21131 3847 21137
rect 3789 21128 3801 21131
rect 2924 21100 3801 21128
rect 2924 21088 2930 21100
rect 3789 21097 3801 21100
rect 3835 21097 3847 21131
rect 3789 21091 3847 21097
rect 4154 21088 4160 21140
rect 4212 21128 4218 21140
rect 4798 21128 4804 21140
rect 4212 21100 4804 21128
rect 4212 21088 4218 21100
rect 4798 21088 4804 21100
rect 4856 21128 4862 21140
rect 4985 21131 5043 21137
rect 4985 21128 4997 21131
rect 4856 21100 4997 21128
rect 4856 21088 4862 21100
rect 4985 21097 4997 21100
rect 5031 21097 5043 21131
rect 4985 21091 5043 21097
rect 9030 21088 9036 21140
rect 9088 21128 9094 21140
rect 9861 21131 9919 21137
rect 9861 21128 9873 21131
rect 9088 21100 9873 21128
rect 9088 21088 9094 21100
rect 9861 21097 9873 21100
rect 9907 21097 9919 21131
rect 10042 21128 10048 21140
rect 10003 21100 10048 21128
rect 9861 21091 9919 21097
rect 10042 21088 10048 21100
rect 10100 21088 10106 21140
rect 12434 21128 12440 21140
rect 11808 21100 12440 21128
rect 9214 21060 9220 21072
rect 7944 21032 9220 21060
rect 1486 20992 1492 21004
rect 1447 20964 1492 20992
rect 1486 20952 1492 20964
rect 1544 20952 1550 21004
rect 3142 20952 3148 21004
rect 3200 20992 3206 21004
rect 3329 20995 3387 21001
rect 3329 20992 3341 20995
rect 3200 20964 3341 20992
rect 3200 20952 3206 20964
rect 3329 20961 3341 20964
rect 3375 20992 3387 20995
rect 4430 20992 4436 21004
rect 3375 20964 3648 20992
rect 4391 20964 4436 20992
rect 3375 20961 3387 20964
rect 3329 20955 3387 20961
rect 3418 20924 3424 20936
rect 3379 20896 3424 20924
rect 3418 20884 3424 20896
rect 3476 20884 3482 20936
rect 3620 20924 3648 20964
rect 4430 20952 4436 20964
rect 4488 20952 4494 21004
rect 7944 21001 7972 21032
rect 9214 21020 9220 21032
rect 9272 21020 9278 21072
rect 7929 20995 7987 21001
rect 7929 20961 7941 20995
rect 7975 20961 7987 20995
rect 8294 20992 8300 21004
rect 8255 20964 8300 20992
rect 7929 20955 7987 20961
rect 8294 20952 8300 20964
rect 8352 20952 8358 21004
rect 8665 20995 8723 21001
rect 8665 20961 8677 20995
rect 8711 20992 8723 20995
rect 8938 20992 8944 21004
rect 8711 20964 8944 20992
rect 8711 20961 8723 20964
rect 8665 20955 8723 20961
rect 8938 20952 8944 20964
rect 8996 20952 9002 21004
rect 4617 20927 4675 20933
rect 4617 20924 4629 20927
rect 3620 20896 4629 20924
rect 4617 20893 4629 20896
rect 4663 20893 4675 20927
rect 4617 20887 4675 20893
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 6365 20927 6423 20933
rect 6365 20924 6377 20927
rect 5592 20896 6377 20924
rect 5592 20884 5598 20896
rect 6365 20893 6377 20896
rect 6411 20924 6423 20927
rect 6822 20924 6828 20936
rect 6411 20896 6828 20924
rect 6411 20893 6423 20896
rect 6365 20887 6423 20893
rect 6822 20884 6828 20896
rect 6880 20884 6886 20936
rect 6914 20884 6920 20936
rect 6972 20924 6978 20936
rect 7834 20924 7840 20936
rect 6972 20896 7840 20924
rect 6972 20884 6978 20896
rect 7834 20884 7840 20896
rect 7892 20924 7898 20936
rect 8021 20927 8079 20933
rect 8021 20924 8033 20927
rect 7892 20896 8033 20924
rect 7892 20884 7898 20896
rect 8021 20893 8033 20896
rect 8067 20893 8079 20927
rect 8021 20887 8079 20893
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20924 8631 20927
rect 8846 20924 8852 20936
rect 8619 20896 8852 20924
rect 8619 20893 8631 20896
rect 8573 20887 8631 20893
rect 8846 20884 8852 20896
rect 8904 20884 8910 20936
rect 9953 20927 10011 20933
rect 9953 20893 9965 20927
rect 9999 20924 10011 20927
rect 10226 20924 10232 20936
rect 9999 20896 10232 20924
rect 9999 20893 10011 20896
rect 9953 20887 10011 20893
rect 10226 20884 10232 20896
rect 10284 20884 10290 20936
rect 11422 20884 11428 20936
rect 11480 20924 11486 20936
rect 11808 20933 11836 21100
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 17494 21128 17500 21140
rect 17455 21100 17500 21128
rect 17494 21088 17500 21100
rect 17552 21128 17558 21140
rect 17957 21131 18015 21137
rect 17957 21128 17969 21131
rect 17552 21100 17969 21128
rect 17552 21088 17558 21100
rect 17957 21097 17969 21100
rect 18003 21097 18015 21131
rect 19245 21131 19303 21137
rect 19245 21128 19257 21131
rect 17957 21091 18015 21097
rect 18616 21100 19257 21128
rect 18616 21069 18644 21100
rect 19245 21097 19257 21100
rect 19291 21097 19303 21131
rect 19245 21091 19303 21097
rect 20533 21131 20591 21137
rect 20533 21097 20545 21131
rect 20579 21128 20591 21131
rect 20579 21100 22324 21128
rect 20579 21097 20591 21100
rect 20533 21091 20591 21097
rect 18601 21063 18659 21069
rect 18601 21029 18613 21063
rect 18647 21029 18659 21063
rect 18601 21023 18659 21029
rect 18693 21063 18751 21069
rect 18693 21029 18705 21063
rect 18739 21029 18751 21063
rect 18693 21023 18751 21029
rect 11974 20992 11980 21004
rect 11935 20964 11980 20992
rect 11974 20952 11980 20964
rect 12032 20952 12038 21004
rect 16206 20952 16212 21004
rect 16264 20992 16270 21004
rect 18233 20995 18291 21001
rect 18233 20992 18245 20995
rect 16264 20964 18245 20992
rect 16264 20952 16270 20964
rect 18233 20961 18245 20964
rect 18279 20961 18291 20995
rect 18233 20955 18291 20961
rect 11609 20927 11667 20933
rect 11609 20924 11621 20927
rect 11480 20896 11621 20924
rect 11480 20884 11486 20896
rect 11609 20893 11621 20896
rect 11655 20893 11667 20927
rect 11609 20887 11667 20893
rect 11792 20927 11850 20933
rect 11792 20893 11804 20927
rect 11838 20893 11850 20927
rect 11792 20887 11850 20893
rect 11885 20927 11943 20933
rect 11885 20893 11897 20927
rect 11931 20893 11943 20927
rect 12158 20924 12164 20936
rect 12119 20896 12164 20924
rect 11885 20887 11943 20893
rect 1756 20859 1814 20865
rect 1756 20825 1768 20859
rect 1802 20856 1814 20859
rect 2498 20856 2504 20868
rect 1802 20828 2504 20856
rect 1802 20825 1814 20828
rect 1756 20819 1814 20825
rect 2498 20816 2504 20828
rect 2556 20816 2562 20868
rect 3050 20856 3056 20868
rect 2884 20828 3056 20856
rect 2884 20797 2912 20828
rect 3050 20816 3056 20828
rect 3108 20856 3114 20868
rect 4157 20859 4215 20865
rect 4157 20856 4169 20859
rect 3108 20828 4169 20856
rect 3108 20816 3114 20828
rect 4157 20825 4169 20828
rect 4203 20825 4215 20859
rect 4157 20819 4215 20825
rect 4249 20859 4307 20865
rect 4249 20825 4261 20859
rect 4295 20856 4307 20859
rect 5994 20856 6000 20868
rect 4295 20828 6000 20856
rect 4295 20825 4307 20828
rect 4249 20819 4307 20825
rect 5994 20816 6000 20828
rect 6052 20816 6058 20868
rect 6086 20816 6092 20868
rect 6144 20865 6150 20868
rect 6144 20856 6156 20865
rect 6144 20828 6189 20856
rect 6144 20819 6156 20828
rect 6144 20816 6150 20819
rect 6270 20816 6276 20868
rect 6328 20856 6334 20868
rect 7662 20859 7720 20865
rect 7662 20856 7674 20859
rect 6328 20828 7674 20856
rect 6328 20816 6334 20828
rect 7662 20825 7674 20828
rect 7708 20825 7720 20859
rect 7662 20819 7720 20825
rect 9858 20816 9864 20868
rect 9916 20856 9922 20868
rect 10962 20856 10968 20868
rect 9916 20828 10968 20856
rect 9916 20816 9922 20828
rect 10962 20816 10968 20828
rect 11020 20816 11026 20868
rect 2869 20791 2927 20797
rect 2869 20757 2881 20791
rect 2915 20757 2927 20791
rect 2869 20751 2927 20757
rect 4430 20748 4436 20800
rect 4488 20788 4494 20800
rect 4801 20791 4859 20797
rect 4801 20788 4813 20791
rect 4488 20760 4813 20788
rect 4488 20748 4494 20760
rect 4801 20757 4813 20760
rect 4847 20757 4859 20791
rect 6012 20788 6040 20816
rect 6549 20791 6607 20797
rect 6549 20788 6561 20791
rect 6012 20760 6561 20788
rect 4801 20751 4859 20757
rect 6549 20757 6561 20760
rect 6595 20757 6607 20791
rect 9674 20788 9680 20800
rect 9635 20760 9680 20788
rect 6549 20751 6607 20757
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 11900 20788 11928 20887
rect 12158 20884 12164 20896
rect 12216 20884 12222 20936
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20924 12495 20927
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 12483 20896 14473 20924
rect 12483 20893 12495 20896
rect 12437 20887 12495 20893
rect 14461 20893 14473 20896
rect 14507 20924 14519 20927
rect 15010 20924 15016 20936
rect 14507 20896 15016 20924
rect 14507 20893 14519 20896
rect 14461 20887 14519 20893
rect 15010 20884 15016 20896
rect 15068 20924 15074 20936
rect 15470 20924 15476 20936
rect 15068 20896 15476 20924
rect 15068 20884 15074 20896
rect 15470 20884 15476 20896
rect 15528 20884 15534 20936
rect 18708 20924 18736 21023
rect 18874 21020 18880 21072
rect 18932 21020 18938 21072
rect 19058 21060 19064 21072
rect 19019 21032 19064 21060
rect 19058 21020 19064 21032
rect 19116 21020 19122 21072
rect 20441 21063 20499 21069
rect 19536 21032 19840 21060
rect 18892 20992 18920 21020
rect 19536 20992 19564 21032
rect 18892 20964 19564 20992
rect 19610 20952 19616 21004
rect 19668 20992 19674 21004
rect 19812 21001 19840 21032
rect 20441 21029 20453 21063
rect 20487 21060 20499 21063
rect 20898 21060 20904 21072
rect 20487 21032 20904 21060
rect 20487 21029 20499 21032
rect 20441 21023 20499 21029
rect 20898 21020 20904 21032
rect 20956 21020 20962 21072
rect 19705 20995 19763 21001
rect 19705 20992 19717 20995
rect 19668 20964 19717 20992
rect 19668 20952 19674 20964
rect 19705 20961 19717 20964
rect 19751 20961 19763 20995
rect 19705 20955 19763 20961
rect 19797 20995 19855 21001
rect 19797 20961 19809 20995
rect 19843 20992 19855 20995
rect 20530 20992 20536 21004
rect 19843 20964 20536 20992
rect 19843 20961 19855 20964
rect 19797 20955 19855 20961
rect 20530 20952 20536 20964
rect 20588 20952 20594 21004
rect 18877 20927 18935 20933
rect 18877 20924 18889 20927
rect 18708 20896 18889 20924
rect 18877 20893 18889 20896
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 18984 20896 20760 20924
rect 12345 20859 12403 20865
rect 12345 20825 12357 20859
rect 12391 20856 12403 20859
rect 12526 20856 12532 20868
rect 12391 20828 12532 20856
rect 12391 20825 12403 20828
rect 12345 20819 12403 20825
rect 12526 20816 12532 20828
rect 12584 20816 12590 20868
rect 12704 20859 12762 20865
rect 12704 20825 12716 20859
rect 12750 20856 12762 20859
rect 14366 20856 14372 20868
rect 12750 20828 14372 20856
rect 12750 20825 12762 20828
rect 12704 20819 12762 20825
rect 14366 20816 14372 20828
rect 14424 20816 14430 20868
rect 14728 20859 14786 20865
rect 14728 20825 14740 20859
rect 14774 20856 14786 20859
rect 15286 20856 15292 20868
rect 14774 20828 15292 20856
rect 14774 20825 14786 20828
rect 14728 20819 14786 20825
rect 15286 20816 15292 20828
rect 15344 20816 15350 20868
rect 18984 20856 19012 20896
rect 15856 20828 19012 20856
rect 20073 20859 20131 20865
rect 13630 20788 13636 20800
rect 11900 20760 13636 20788
rect 13630 20748 13636 20760
rect 13688 20748 13694 20800
rect 13817 20791 13875 20797
rect 13817 20757 13829 20791
rect 13863 20788 13875 20791
rect 14090 20788 14096 20800
rect 13863 20760 14096 20788
rect 13863 20757 13875 20760
rect 13817 20751 13875 20757
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 15856 20797 15884 20828
rect 20073 20825 20085 20859
rect 20119 20856 20131 20859
rect 20162 20856 20168 20868
rect 20119 20828 20168 20856
rect 20119 20825 20131 20828
rect 20073 20819 20131 20825
rect 20162 20816 20168 20828
rect 20220 20856 20226 20868
rect 20622 20856 20628 20868
rect 20220 20828 20628 20856
rect 20220 20816 20226 20828
rect 20622 20816 20628 20828
rect 20680 20816 20686 20868
rect 20732 20856 20760 20896
rect 21634 20884 21640 20936
rect 21692 20924 21698 20936
rect 22189 20927 22247 20933
rect 22189 20924 22201 20927
rect 21692 20896 22201 20924
rect 21692 20884 21698 20896
rect 22189 20893 22201 20896
rect 22235 20893 22247 20927
rect 22296 20924 22324 21100
rect 23290 21088 23296 21140
rect 23348 21128 23354 21140
rect 23937 21131 23995 21137
rect 23937 21128 23949 21131
rect 23348 21100 23949 21128
rect 23348 21088 23354 21100
rect 23937 21097 23949 21100
rect 23983 21097 23995 21131
rect 23937 21091 23995 21097
rect 22830 20933 22836 20936
rect 22465 20927 22523 20933
rect 22465 20924 22477 20927
rect 22296 20896 22477 20924
rect 22189 20887 22247 20893
rect 22465 20893 22477 20896
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20893 22615 20927
rect 22824 20924 22836 20933
rect 22791 20896 22836 20924
rect 22557 20887 22615 20893
rect 22824 20887 22836 20896
rect 21726 20856 21732 20868
rect 20732 20828 21732 20856
rect 21726 20816 21732 20828
rect 21784 20816 21790 20868
rect 21944 20859 22002 20865
rect 21944 20825 21956 20859
rect 21990 20856 22002 20859
rect 22204 20856 22232 20887
rect 22572 20856 22600 20887
rect 22830 20884 22836 20887
rect 22888 20884 22894 20936
rect 21990 20828 22094 20856
rect 22204 20828 22600 20856
rect 21990 20825 22002 20828
rect 21944 20819 22002 20825
rect 15841 20791 15899 20797
rect 15841 20788 15853 20791
rect 15252 20760 15853 20788
rect 15252 20748 15258 20760
rect 15841 20757 15853 20760
rect 15887 20757 15899 20791
rect 19610 20788 19616 20800
rect 19571 20760 19616 20788
rect 15841 20751 15899 20757
rect 19610 20748 19616 20760
rect 19668 20748 19674 20800
rect 20809 20791 20867 20797
rect 20809 20757 20821 20791
rect 20855 20788 20867 20791
rect 21358 20788 21364 20800
rect 20855 20760 21364 20788
rect 20855 20757 20867 20760
rect 20809 20751 20867 20757
rect 21358 20748 21364 20760
rect 21416 20748 21422 20800
rect 22066 20788 22094 20828
rect 22281 20791 22339 20797
rect 22281 20788 22293 20791
rect 22066 20760 22293 20788
rect 22281 20757 22293 20760
rect 22327 20757 22339 20791
rect 22281 20751 22339 20757
rect 1104 20698 26220 20720
rect 1104 20646 9322 20698
rect 9374 20646 9386 20698
rect 9438 20646 9450 20698
rect 9502 20646 9514 20698
rect 9566 20646 9578 20698
rect 9630 20646 17694 20698
rect 17746 20646 17758 20698
rect 17810 20646 17822 20698
rect 17874 20646 17886 20698
rect 17938 20646 17950 20698
rect 18002 20646 26220 20698
rect 1104 20624 26220 20646
rect 2498 20584 2504 20596
rect 2459 20556 2504 20584
rect 2498 20544 2504 20556
rect 2556 20544 2562 20596
rect 3145 20587 3203 20593
rect 3145 20584 3157 20587
rect 2746 20556 3157 20584
rect 2746 20516 2774 20556
rect 3145 20553 3157 20556
rect 3191 20553 3203 20587
rect 3145 20547 3203 20553
rect 4157 20587 4215 20593
rect 4157 20553 4169 20587
rect 4203 20553 4215 20587
rect 4338 20584 4344 20596
rect 4299 20556 4344 20584
rect 4157 20547 4215 20553
rect 2958 20516 2964 20528
rect 2700 20488 2774 20516
rect 2884 20488 2964 20516
rect 2700 20457 2728 20488
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20417 2743 20451
rect 2685 20411 2743 20417
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20448 2835 20451
rect 2884 20448 2912 20488
rect 2958 20476 2964 20488
rect 3016 20516 3022 20528
rect 4062 20516 4068 20528
rect 3016 20488 4068 20516
rect 3016 20476 3022 20488
rect 4062 20476 4068 20488
rect 4120 20516 4126 20528
rect 4172 20516 4200 20547
rect 4338 20544 4344 20556
rect 4396 20584 4402 20596
rect 4522 20584 4528 20596
rect 4396 20556 4528 20584
rect 4396 20544 4402 20556
rect 4522 20544 4528 20556
rect 4580 20544 4586 20596
rect 4709 20587 4767 20593
rect 4709 20553 4721 20587
rect 4755 20584 4767 20587
rect 6086 20584 6092 20596
rect 4755 20556 6092 20584
rect 4755 20553 4767 20556
rect 4709 20547 4767 20553
rect 6086 20544 6092 20556
rect 6144 20544 6150 20596
rect 6362 20544 6368 20596
rect 6420 20584 6426 20596
rect 7377 20587 7435 20593
rect 7377 20584 7389 20587
rect 6420 20556 7389 20584
rect 6420 20544 6426 20556
rect 7377 20553 7389 20556
rect 7423 20553 7435 20587
rect 7377 20547 7435 20553
rect 8570 20544 8576 20596
rect 8628 20544 8634 20596
rect 8846 20544 8852 20596
rect 8904 20584 8910 20596
rect 9125 20587 9183 20593
rect 9125 20584 9137 20587
rect 8904 20556 9137 20584
rect 8904 20544 8910 20556
rect 9125 20553 9137 20556
rect 9171 20553 9183 20587
rect 9125 20547 9183 20553
rect 9585 20587 9643 20593
rect 9585 20553 9597 20587
rect 9631 20584 9643 20587
rect 9950 20584 9956 20596
rect 9631 20556 9956 20584
rect 9631 20553 9643 20556
rect 9585 20547 9643 20553
rect 9950 20544 9956 20556
rect 10008 20584 10014 20596
rect 10410 20584 10416 20596
rect 10008 20556 10416 20584
rect 10008 20544 10014 20556
rect 10410 20544 10416 20556
rect 10468 20544 10474 20596
rect 10594 20584 10600 20596
rect 10507 20556 10600 20584
rect 10594 20544 10600 20556
rect 10652 20584 10658 20596
rect 13262 20584 13268 20596
rect 10652 20556 13268 20584
rect 10652 20544 10658 20556
rect 13262 20544 13268 20556
rect 13320 20544 13326 20596
rect 13630 20584 13636 20596
rect 13591 20556 13636 20584
rect 13630 20544 13636 20556
rect 13688 20584 13694 20596
rect 13688 20556 14320 20584
rect 13688 20544 13694 20556
rect 6181 20519 6239 20525
rect 4120 20488 4200 20516
rect 5736 20488 6132 20516
rect 4120 20476 4126 20488
rect 3050 20448 3056 20460
rect 2823 20420 2912 20448
rect 3011 20420 3056 20448
rect 2823 20417 2835 20420
rect 2777 20411 2835 20417
rect 3050 20408 3056 20420
rect 3108 20408 3114 20460
rect 3510 20448 3516 20460
rect 3471 20420 3516 20448
rect 3510 20408 3516 20420
rect 3568 20408 3574 20460
rect 3970 20448 3976 20460
rect 3931 20420 3976 20448
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 4246 20408 4252 20460
rect 4304 20448 4310 20460
rect 4798 20448 4804 20460
rect 4304 20420 4568 20448
rect 4759 20420 4804 20448
rect 4304 20408 4310 20420
rect 3602 20380 3608 20392
rect 3563 20352 3608 20380
rect 3602 20340 3608 20352
rect 3660 20340 3666 20392
rect 3789 20383 3847 20389
rect 3789 20349 3801 20383
rect 3835 20380 3847 20383
rect 4338 20380 4344 20392
rect 3835 20352 4344 20380
rect 3835 20349 3847 20352
rect 3789 20343 3847 20349
rect 4338 20340 4344 20352
rect 4396 20340 4402 20392
rect 4430 20340 4436 20392
rect 4488 20340 4494 20392
rect 4540 20389 4568 20420
rect 4798 20408 4804 20420
rect 4856 20408 4862 20460
rect 5170 20451 5228 20457
rect 5170 20448 5182 20451
rect 4908 20420 5182 20448
rect 4525 20383 4583 20389
rect 4525 20349 4537 20383
rect 4571 20380 4583 20383
rect 4908 20380 4936 20420
rect 5170 20417 5182 20420
rect 5216 20448 5228 20451
rect 5258 20448 5264 20460
rect 5216 20420 5264 20448
rect 5216 20417 5228 20420
rect 5170 20411 5228 20417
rect 5258 20408 5264 20420
rect 5316 20408 5322 20460
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20448 5411 20451
rect 5442 20448 5448 20460
rect 5399 20420 5448 20448
rect 5399 20417 5411 20420
rect 5353 20411 5411 20417
rect 5442 20408 5448 20420
rect 5500 20408 5506 20460
rect 5626 20448 5632 20460
rect 5587 20420 5632 20448
rect 5626 20408 5632 20420
rect 5684 20408 5690 20460
rect 5736 20389 5764 20488
rect 5994 20448 6000 20460
rect 5955 20420 6000 20448
rect 5994 20408 6000 20420
rect 6052 20408 6058 20460
rect 6104 20448 6132 20488
rect 6181 20485 6193 20519
rect 6227 20516 6239 20519
rect 6270 20516 6276 20528
rect 6227 20488 6276 20516
rect 6227 20485 6239 20488
rect 6181 20479 6239 20485
rect 6270 20476 6276 20488
rect 6328 20476 6334 20528
rect 6638 20516 6644 20528
rect 6472 20488 6644 20516
rect 6472 20448 6500 20488
rect 6638 20476 6644 20488
rect 6696 20516 6702 20528
rect 7285 20519 7343 20525
rect 6696 20488 6868 20516
rect 6696 20476 6702 20488
rect 6104 20420 6500 20448
rect 6546 20408 6552 20460
rect 6604 20448 6610 20460
rect 6840 20457 6868 20488
rect 7285 20485 7297 20519
rect 7331 20516 7343 20519
rect 8588 20516 8616 20544
rect 7331 20488 8616 20516
rect 7331 20485 7343 20488
rect 7285 20479 7343 20485
rect 6825 20451 6883 20457
rect 6604 20420 6649 20448
rect 6604 20408 6610 20420
rect 6825 20417 6837 20451
rect 6871 20417 6883 20451
rect 6825 20411 6883 20417
rect 6918 20451 6976 20457
rect 6918 20417 6930 20451
rect 6964 20417 6976 20451
rect 7098 20448 7104 20460
rect 7059 20420 7104 20448
rect 6918 20411 6976 20417
rect 4571 20352 4936 20380
rect 4985 20383 5043 20389
rect 4571 20349 4583 20352
rect 4525 20343 4583 20349
rect 4985 20349 4997 20383
rect 5031 20349 5043 20383
rect 4985 20343 5043 20349
rect 5077 20383 5135 20389
rect 5077 20349 5089 20383
rect 5123 20380 5135 20383
rect 5721 20383 5779 20389
rect 5721 20380 5733 20383
rect 5123 20352 5733 20380
rect 5123 20349 5135 20352
rect 5077 20343 5135 20349
rect 5721 20349 5733 20352
rect 5767 20349 5779 20383
rect 5721 20343 5779 20349
rect 5813 20383 5871 20389
rect 5813 20349 5825 20383
rect 5859 20380 5871 20383
rect 6730 20380 6736 20392
rect 5859 20352 6736 20380
rect 5859 20349 5871 20352
rect 5813 20343 5871 20349
rect 2961 20315 3019 20321
rect 2961 20281 2973 20315
rect 3007 20312 3019 20315
rect 4448 20312 4476 20340
rect 3007 20284 4476 20312
rect 5000 20312 5028 20343
rect 5828 20312 5856 20343
rect 6730 20340 6736 20352
rect 6788 20340 6794 20392
rect 6933 20380 6961 20411
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 7300 20380 7328 20479
rect 9214 20476 9220 20528
rect 9272 20516 9278 20528
rect 14292 20516 14320 20556
rect 14366 20544 14372 20596
rect 14424 20584 14430 20596
rect 14461 20587 14519 20593
rect 14461 20584 14473 20587
rect 14424 20556 14473 20584
rect 14424 20544 14430 20556
rect 14461 20553 14473 20556
rect 14507 20553 14519 20587
rect 15286 20584 15292 20596
rect 15247 20556 15292 20584
rect 14461 20547 14519 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 16114 20584 16120 20596
rect 15436 20556 15792 20584
rect 16075 20556 16120 20584
rect 15436 20544 15442 20556
rect 9272 20488 12296 20516
rect 9272 20476 9278 20488
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20448 8631 20451
rect 9033 20451 9091 20457
rect 8619 20420 8708 20448
rect 8619 20417 8631 20420
rect 8573 20411 8631 20417
rect 6933 20352 7328 20380
rect 8386 20340 8392 20392
rect 8444 20380 8450 20392
rect 8481 20383 8539 20389
rect 8481 20380 8493 20383
rect 8444 20352 8493 20380
rect 8444 20340 8450 20352
rect 8481 20349 8493 20352
rect 8527 20349 8539 20383
rect 8481 20343 8539 20349
rect 7098 20312 7104 20324
rect 5000 20284 5856 20312
rect 5920 20284 7104 20312
rect 3007 20281 3019 20284
rect 2961 20275 3019 20281
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 5920 20244 5948 20284
rect 7098 20272 7104 20284
rect 7156 20272 7162 20324
rect 7282 20272 7288 20324
rect 7340 20312 7346 20324
rect 8680 20321 8708 20420
rect 9033 20417 9045 20451
rect 9079 20448 9091 20451
rect 9674 20448 9680 20460
rect 9079 20420 9680 20448
rect 9079 20417 9091 20420
rect 9033 20411 9091 20417
rect 9674 20408 9680 20420
rect 9732 20408 9738 20460
rect 9858 20408 9864 20460
rect 9916 20448 9922 20460
rect 10045 20451 10103 20457
rect 10045 20448 10057 20451
rect 9916 20420 10057 20448
rect 9916 20408 9922 20420
rect 10045 20417 10057 20420
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 10137 20451 10195 20457
rect 10137 20417 10149 20451
rect 10183 20448 10195 20451
rect 10502 20448 10508 20460
rect 10183 20420 10508 20448
rect 10183 20417 10195 20420
rect 10137 20411 10195 20417
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 12268 20457 12296 20488
rect 12360 20488 13860 20516
rect 14292 20488 15608 20516
rect 12253 20451 12311 20457
rect 12253 20417 12265 20451
rect 12299 20417 12311 20451
rect 12253 20411 12311 20417
rect 9122 20340 9128 20392
rect 9180 20380 9186 20392
rect 9217 20383 9275 20389
rect 9217 20380 9229 20383
rect 9180 20352 9229 20380
rect 9180 20340 9186 20352
rect 9217 20349 9229 20352
rect 9263 20349 9275 20383
rect 9217 20343 9275 20349
rect 9769 20383 9827 20389
rect 9769 20349 9781 20383
rect 9815 20380 9827 20383
rect 10226 20380 10232 20392
rect 9815 20352 10232 20380
rect 9815 20349 9827 20352
rect 9769 20343 9827 20349
rect 10226 20340 10232 20352
rect 10284 20340 10290 20392
rect 11422 20340 11428 20392
rect 11480 20380 11486 20392
rect 12360 20380 12388 20488
rect 12526 20457 12532 20460
rect 12520 20411 12532 20457
rect 12584 20448 12590 20460
rect 12584 20420 12620 20448
rect 12526 20408 12532 20411
rect 12584 20408 12590 20420
rect 12894 20408 12900 20460
rect 12952 20448 12958 20460
rect 13832 20457 13860 20488
rect 13817 20451 13875 20457
rect 12952 20420 13768 20448
rect 12952 20408 12958 20420
rect 11480 20352 12388 20380
rect 13740 20380 13768 20420
rect 13817 20417 13829 20451
rect 13863 20417 13875 20451
rect 13982 20451 14040 20457
rect 13982 20448 13994 20451
rect 13817 20411 13875 20417
rect 13924 20420 13994 20448
rect 13924 20380 13952 20420
rect 13982 20417 13994 20420
rect 14028 20417 14040 20451
rect 13982 20411 14040 20417
rect 14090 20408 14096 20460
rect 14148 20448 14154 20460
rect 14369 20451 14427 20457
rect 14369 20448 14381 20451
rect 14148 20420 14193 20448
rect 14292 20420 14381 20448
rect 14148 20408 14154 20420
rect 14182 20380 14188 20392
rect 13740 20352 13952 20380
rect 14143 20352 14188 20380
rect 11480 20340 11486 20352
rect 14182 20340 14188 20352
rect 14240 20340 14246 20392
rect 8205 20315 8263 20321
rect 8205 20312 8217 20315
rect 7340 20284 8217 20312
rect 7340 20272 7346 20284
rect 8205 20281 8217 20284
rect 8251 20281 8263 20315
rect 8205 20275 8263 20281
rect 8665 20315 8723 20321
rect 8665 20281 8677 20315
rect 8711 20281 8723 20315
rect 8665 20275 8723 20281
rect 9674 20272 9680 20324
rect 9732 20312 9738 20324
rect 9861 20315 9919 20321
rect 9861 20312 9873 20315
rect 9732 20284 9873 20312
rect 9732 20272 9738 20284
rect 9861 20281 9873 20284
rect 9907 20312 9919 20315
rect 10594 20312 10600 20324
rect 9907 20284 10600 20312
rect 9907 20281 9919 20284
rect 9861 20275 9919 20281
rect 10594 20272 10600 20284
rect 10652 20272 10658 20324
rect 14292 20312 14320 20420
rect 14369 20417 14381 20420
rect 14415 20417 14427 20451
rect 14642 20448 14648 20460
rect 14603 20420 14648 20448
rect 14369 20411 14427 20417
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 14826 20408 14832 20460
rect 14884 20448 14890 20460
rect 15194 20448 15200 20460
rect 14884 20420 14928 20448
rect 15155 20420 15200 20448
rect 14884 20408 14890 20420
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20417 15531 20451
rect 15580 20448 15608 20488
rect 15638 20451 15696 20457
rect 15638 20448 15650 20451
rect 15580 20420 15650 20448
rect 15473 20411 15531 20417
rect 15638 20417 15650 20420
rect 15684 20417 15696 20451
rect 15764 20448 15792 20556
rect 16114 20544 16120 20556
rect 16172 20544 16178 20596
rect 18874 20544 18880 20596
rect 18932 20584 18938 20596
rect 19061 20587 19119 20593
rect 19061 20584 19073 20587
rect 18932 20556 19073 20584
rect 18932 20544 18938 20556
rect 19061 20553 19073 20556
rect 19107 20553 19119 20587
rect 20070 20584 20076 20596
rect 19061 20547 19119 20553
rect 19904 20556 20076 20584
rect 19702 20516 19708 20528
rect 19663 20488 19708 20516
rect 19702 20476 19708 20488
rect 19760 20476 19766 20528
rect 19904 20525 19932 20556
rect 20070 20544 20076 20556
rect 20128 20544 20134 20596
rect 20530 20544 20536 20596
rect 20588 20584 20594 20596
rect 20717 20587 20775 20593
rect 20717 20584 20729 20587
rect 20588 20556 20729 20584
rect 20588 20544 20594 20556
rect 20717 20553 20729 20556
rect 20763 20553 20775 20587
rect 20898 20584 20904 20596
rect 20859 20556 20904 20584
rect 20717 20547 20775 20553
rect 19889 20519 19947 20525
rect 19889 20485 19901 20519
rect 19935 20485 19947 20519
rect 19889 20479 19947 20485
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 15764 20420 15853 20448
rect 15638 20411 15696 20417
rect 15841 20417 15853 20420
rect 15887 20417 15899 20451
rect 16022 20448 16028 20460
rect 15983 20420 16028 20448
rect 15841 20411 15899 20417
rect 14921 20383 14979 20389
rect 14921 20349 14933 20383
rect 14967 20349 14979 20383
rect 14921 20343 14979 20349
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20380 15071 20383
rect 15286 20380 15292 20392
rect 15059 20352 15292 20380
rect 15059 20349 15071 20352
rect 15013 20343 15071 20349
rect 13556 20284 14320 20312
rect 14936 20312 14964 20343
rect 15286 20340 15292 20352
rect 15344 20340 15350 20392
rect 15194 20312 15200 20324
rect 14936 20284 15200 20312
rect 5592 20216 5948 20244
rect 6457 20247 6515 20253
rect 5592 20204 5598 20216
rect 6457 20213 6469 20247
rect 6503 20244 6515 20247
rect 6546 20244 6552 20256
rect 6503 20216 6552 20244
rect 6503 20213 6515 20216
rect 6457 20207 6515 20213
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 8573 20247 8631 20253
rect 8573 20213 8585 20247
rect 8619 20244 8631 20247
rect 9950 20244 9956 20256
rect 8619 20216 9956 20244
rect 8619 20213 8631 20216
rect 8573 20207 8631 20213
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 10318 20244 10324 20256
rect 10279 20216 10324 20244
rect 10318 20204 10324 20216
rect 10376 20204 10382 20256
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 12158 20244 12164 20256
rect 11940 20216 12164 20244
rect 11940 20204 11946 20216
rect 12158 20204 12164 20216
rect 12216 20244 12222 20256
rect 13556 20244 13584 20284
rect 15194 20272 15200 20284
rect 15252 20272 15258 20324
rect 15488 20312 15516 20411
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 20073 20451 20131 20457
rect 20073 20417 20085 20451
rect 20119 20448 20131 20451
rect 20254 20448 20260 20460
rect 20119 20420 20260 20448
rect 20119 20417 20131 20420
rect 20073 20411 20131 20417
rect 20254 20408 20260 20420
rect 20312 20408 20318 20460
rect 15746 20380 15752 20392
rect 15707 20352 15752 20380
rect 15746 20340 15752 20352
rect 15804 20340 15810 20392
rect 20732 20380 20760 20547
rect 20898 20544 20904 20556
rect 20956 20544 20962 20596
rect 21361 20587 21419 20593
rect 21361 20553 21373 20587
rect 21407 20584 21419 20587
rect 21450 20584 21456 20596
rect 21407 20556 21456 20584
rect 21407 20553 21419 20556
rect 21361 20547 21419 20553
rect 21450 20544 21456 20556
rect 21508 20544 21514 20596
rect 22557 20587 22615 20593
rect 22557 20553 22569 20587
rect 22603 20584 22615 20587
rect 22922 20584 22928 20596
rect 22603 20556 22928 20584
rect 22603 20553 22615 20556
rect 22557 20547 22615 20553
rect 22922 20544 22928 20556
rect 22980 20544 22986 20596
rect 23198 20516 23204 20528
rect 23159 20488 23204 20516
rect 23198 20476 23204 20488
rect 23256 20476 23262 20528
rect 23290 20476 23296 20528
rect 23348 20516 23354 20528
rect 23385 20519 23443 20525
rect 23385 20516 23397 20519
rect 23348 20488 23397 20516
rect 23348 20476 23354 20488
rect 23385 20485 23397 20488
rect 23431 20485 23443 20519
rect 23385 20479 23443 20485
rect 23474 20476 23480 20528
rect 23532 20516 23538 20528
rect 23569 20519 23627 20525
rect 23569 20516 23581 20519
rect 23532 20488 23581 20516
rect 23532 20476 23538 20488
rect 23569 20485 23581 20488
rect 23615 20485 23627 20519
rect 23569 20479 23627 20485
rect 21266 20448 21272 20460
rect 21227 20420 21272 20448
rect 21266 20408 21272 20420
rect 21324 20408 21330 20460
rect 22370 20408 22376 20460
rect 22428 20448 22434 20460
rect 22465 20451 22523 20457
rect 22465 20448 22477 20451
rect 22428 20420 22477 20448
rect 22428 20408 22434 20420
rect 22465 20417 22477 20420
rect 22511 20417 22523 20451
rect 22465 20411 22523 20417
rect 21453 20383 21511 20389
rect 21453 20380 21465 20383
rect 20732 20352 21465 20380
rect 21453 20349 21465 20352
rect 21499 20380 21511 20383
rect 21913 20383 21971 20389
rect 21913 20380 21925 20383
rect 21499 20352 21925 20380
rect 21499 20349 21511 20352
rect 21453 20343 21511 20349
rect 21913 20349 21925 20352
rect 21959 20380 21971 20383
rect 22738 20380 22744 20392
rect 21959 20352 22744 20380
rect 21959 20349 21971 20352
rect 21913 20343 21971 20349
rect 22738 20340 22744 20352
rect 22796 20340 22802 20392
rect 17310 20312 17316 20324
rect 15488 20284 17316 20312
rect 12216 20216 13584 20244
rect 12216 20204 12222 20216
rect 14918 20204 14924 20256
rect 14976 20244 14982 20256
rect 15488 20244 15516 20284
rect 17310 20272 17316 20284
rect 17368 20272 17374 20324
rect 14976 20216 15516 20244
rect 22097 20247 22155 20253
rect 14976 20204 14982 20216
rect 22097 20213 22109 20247
rect 22143 20244 22155 20247
rect 22278 20244 22284 20256
rect 22143 20216 22284 20244
rect 22143 20213 22155 20216
rect 22097 20207 22155 20213
rect 22278 20204 22284 20216
rect 22336 20204 22342 20256
rect 1104 20154 26220 20176
rect 1104 20102 5136 20154
rect 5188 20102 5200 20154
rect 5252 20102 5264 20154
rect 5316 20102 5328 20154
rect 5380 20102 5392 20154
rect 5444 20102 13508 20154
rect 13560 20102 13572 20154
rect 13624 20102 13636 20154
rect 13688 20102 13700 20154
rect 13752 20102 13764 20154
rect 13816 20102 21880 20154
rect 21932 20102 21944 20154
rect 21996 20102 22008 20154
rect 22060 20102 22072 20154
rect 22124 20102 22136 20154
rect 22188 20102 26220 20154
rect 1104 20080 26220 20102
rect 3602 20000 3608 20052
rect 3660 20040 3666 20052
rect 5445 20043 5503 20049
rect 5445 20040 5457 20043
rect 3660 20012 5457 20040
rect 3660 20000 3666 20012
rect 5445 20009 5457 20012
rect 5491 20040 5503 20043
rect 6454 20040 6460 20052
rect 5491 20012 6460 20040
rect 5491 20009 5503 20012
rect 5445 20003 5503 20009
rect 6454 20000 6460 20012
rect 6512 20000 6518 20052
rect 7098 20000 7104 20052
rect 7156 20040 7162 20052
rect 7156 20012 8432 20040
rect 7156 20000 7162 20012
rect 3145 19975 3203 19981
rect 3145 19941 3157 19975
rect 3191 19972 3203 19975
rect 3510 19972 3516 19984
rect 3191 19944 3516 19972
rect 3191 19941 3203 19944
rect 3145 19935 3203 19941
rect 3510 19932 3516 19944
rect 3568 19972 3574 19984
rect 3568 19944 3832 19972
rect 3568 19932 3574 19944
rect 3804 19913 3832 19944
rect 3970 19932 3976 19984
rect 4028 19972 4034 19984
rect 7745 19975 7803 19981
rect 4028 19944 4568 19972
rect 4028 19932 4034 19944
rect 3789 19907 3847 19913
rect 3789 19873 3801 19907
rect 3835 19873 3847 19907
rect 3789 19867 3847 19873
rect 3881 19907 3939 19913
rect 3881 19873 3893 19907
rect 3927 19904 3939 19907
rect 4430 19904 4436 19916
rect 3927 19876 4436 19904
rect 3927 19873 3939 19876
rect 3881 19867 3939 19873
rect 4430 19864 4436 19876
rect 4488 19864 4494 19916
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19836 1823 19839
rect 1811 19808 2176 19836
rect 1811 19805 1823 19808
rect 1765 19799 1823 19805
rect 2148 19780 2176 19808
rect 3418 19796 3424 19848
rect 3476 19836 3482 19848
rect 3513 19839 3571 19845
rect 3513 19836 3525 19839
rect 3476 19808 3525 19836
rect 3476 19796 3482 19808
rect 3513 19805 3525 19808
rect 3559 19836 3571 19839
rect 3694 19836 3700 19848
rect 3559 19808 3700 19836
rect 3559 19805 3571 19808
rect 3513 19799 3571 19805
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 4062 19836 4068 19848
rect 4023 19808 4068 19836
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19836 4215 19839
rect 4338 19836 4344 19848
rect 4203 19808 4344 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4338 19796 4344 19808
rect 4396 19796 4402 19848
rect 2032 19771 2090 19777
rect 2032 19737 2044 19771
rect 2078 19737 2090 19771
rect 2032 19731 2090 19737
rect 2056 19700 2084 19731
rect 2130 19728 2136 19780
rect 2188 19728 2194 19780
rect 4540 19768 4568 19944
rect 7745 19941 7757 19975
rect 7791 19972 7803 19975
rect 7791 19944 8340 19972
rect 7791 19941 7803 19944
rect 7745 19935 7803 19941
rect 6822 19904 6828 19916
rect 6783 19876 6828 19904
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 7834 19864 7840 19916
rect 7892 19904 7898 19916
rect 7929 19907 7987 19913
rect 7929 19904 7941 19907
rect 7892 19876 7941 19904
rect 7892 19864 7898 19876
rect 7929 19873 7941 19876
rect 7975 19873 7987 19907
rect 7929 19867 7987 19873
rect 6546 19796 6552 19848
rect 6604 19845 6610 19848
rect 8312 19845 8340 19944
rect 8404 19904 8432 20012
rect 9122 20000 9128 20052
rect 9180 20040 9186 20052
rect 9401 20043 9459 20049
rect 9401 20040 9413 20043
rect 9180 20012 9413 20040
rect 9180 20000 9186 20012
rect 9401 20009 9413 20012
rect 9447 20009 9459 20043
rect 9674 20040 9680 20052
rect 9635 20012 9680 20040
rect 9401 20003 9459 20009
rect 8938 19972 8944 19984
rect 8899 19944 8944 19972
rect 8938 19932 8944 19944
rect 8996 19932 9002 19984
rect 9416 19904 9444 20003
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 10686 20040 10692 20052
rect 10647 20012 10692 20040
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 11698 20000 11704 20052
rect 11756 20040 11762 20052
rect 13173 20043 13231 20049
rect 13173 20040 13185 20043
rect 11756 20012 13185 20040
rect 11756 20000 11762 20012
rect 13173 20009 13185 20012
rect 13219 20040 13231 20043
rect 14826 20040 14832 20052
rect 13219 20012 14832 20040
rect 13219 20009 13231 20012
rect 13173 20003 13231 20009
rect 14826 20000 14832 20012
rect 14884 20000 14890 20052
rect 15194 20040 15200 20052
rect 14936 20012 15200 20040
rect 10045 19907 10103 19913
rect 10045 19904 10057 19907
rect 8404 19876 9260 19904
rect 9416 19876 10057 19904
rect 6604 19836 6616 19845
rect 7561 19839 7619 19845
rect 7561 19836 7573 19839
rect 6604 19808 6649 19836
rect 7484 19808 7573 19836
rect 6604 19799 6616 19808
rect 6604 19796 6610 19799
rect 7282 19768 7288 19780
rect 2240 19740 4384 19768
rect 4540 19740 7288 19768
rect 2240 19700 2268 19740
rect 2056 19672 2268 19700
rect 3329 19703 3387 19709
rect 3329 19669 3341 19703
rect 3375 19700 3387 19703
rect 3786 19700 3792 19712
rect 3375 19672 3792 19700
rect 3375 19669 3387 19672
rect 3329 19663 3387 19669
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 4356 19709 4384 19740
rect 7282 19728 7288 19740
rect 7340 19728 7346 19780
rect 7484 19712 7512 19808
rect 7561 19805 7573 19808
rect 7607 19805 7619 19839
rect 7561 19799 7619 19805
rect 8113 19839 8171 19845
rect 8113 19805 8125 19839
rect 8159 19805 8171 19839
rect 8113 19799 8171 19805
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19836 8355 19839
rect 8386 19836 8392 19848
rect 8343 19808 8392 19836
rect 8343 19805 8355 19808
rect 8297 19799 8355 19805
rect 8128 19768 8156 19799
rect 8386 19796 8392 19808
rect 8444 19796 8450 19848
rect 9030 19796 9036 19848
rect 9088 19836 9094 19848
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 9088 19808 9137 19836
rect 9088 19796 9094 19808
rect 9125 19805 9137 19808
rect 9171 19805 9183 19839
rect 9232 19836 9260 19876
rect 10045 19873 10057 19876
rect 10091 19904 10103 19907
rect 10091 19876 11928 19904
rect 10091 19873 10103 19876
rect 10045 19867 10103 19873
rect 9766 19836 9772 19848
rect 9232 19808 9444 19836
rect 9727 19808 9772 19836
rect 9125 19799 9183 19805
rect 8846 19768 8852 19780
rect 8128 19740 8852 19768
rect 8846 19728 8852 19740
rect 8904 19728 8910 19780
rect 9214 19728 9220 19780
rect 9272 19768 9278 19780
rect 9309 19771 9367 19777
rect 9309 19768 9321 19771
rect 9272 19740 9321 19768
rect 9272 19728 9278 19740
rect 9309 19737 9321 19740
rect 9355 19737 9367 19771
rect 9416 19768 9444 19808
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 10318 19836 10324 19848
rect 10279 19808 10324 19836
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 11790 19836 11796 19848
rect 11751 19808 11796 19836
rect 11790 19796 11796 19808
rect 11848 19796 11854 19848
rect 11900 19836 11928 19876
rect 14090 19864 14096 19916
rect 14148 19904 14154 19916
rect 14936 19913 14964 20012
rect 15194 20000 15200 20012
rect 15252 20040 15258 20052
rect 15746 20040 15752 20052
rect 15252 20012 15752 20040
rect 15252 20000 15258 20012
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 22370 20040 22376 20052
rect 22331 20012 22376 20040
rect 22370 20000 22376 20012
rect 22428 20000 22434 20052
rect 25317 20043 25375 20049
rect 25317 20009 25329 20043
rect 25363 20040 25375 20043
rect 26329 20043 26387 20049
rect 26329 20040 26341 20043
rect 25363 20012 26341 20040
rect 25363 20009 25375 20012
rect 25317 20003 25375 20009
rect 26329 20009 26341 20012
rect 26375 20009 26387 20043
rect 26329 20003 26387 20009
rect 22097 19975 22155 19981
rect 22097 19941 22109 19975
rect 22143 19972 22155 19975
rect 22278 19972 22284 19984
rect 22143 19944 22284 19972
rect 22143 19941 22155 19944
rect 22097 19935 22155 19941
rect 22278 19932 22284 19944
rect 22336 19932 22342 19984
rect 14921 19907 14979 19913
rect 14148 19876 14780 19904
rect 14148 19864 14154 19876
rect 12986 19836 12992 19848
rect 11900 19808 12992 19836
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19805 14703 19839
rect 14752 19836 14780 19876
rect 14921 19873 14933 19907
rect 14967 19873 14979 19907
rect 14921 19867 14979 19873
rect 15013 19907 15071 19913
rect 15013 19873 15025 19907
rect 15059 19904 15071 19907
rect 15286 19904 15292 19916
rect 15059 19876 15292 19904
rect 15059 19873 15071 19876
rect 15013 19867 15071 19873
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 15470 19904 15476 19916
rect 15431 19876 15476 19904
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 16666 19864 16672 19916
rect 16724 19904 16730 19916
rect 17589 19907 17647 19913
rect 17589 19904 17601 19907
rect 16724 19876 17601 19904
rect 16724 19864 16730 19876
rect 17589 19873 17601 19876
rect 17635 19873 17647 19907
rect 17589 19867 17647 19873
rect 20162 19864 20168 19916
rect 20220 19904 20226 19916
rect 21729 19907 21787 19913
rect 21729 19904 21741 19907
rect 20220 19876 21741 19904
rect 20220 19864 20226 19876
rect 21729 19873 21741 19876
rect 21775 19873 21787 19907
rect 21729 19867 21787 19873
rect 22370 19864 22376 19916
rect 22428 19904 22434 19916
rect 22925 19907 22983 19913
rect 22925 19904 22937 19907
rect 22428 19876 22937 19904
rect 22428 19864 22434 19876
rect 22925 19873 22937 19876
rect 22971 19873 22983 19907
rect 22925 19867 22983 19873
rect 14810 19839 14868 19845
rect 14810 19836 14822 19839
rect 14752 19808 14822 19836
rect 14645 19799 14703 19805
rect 14810 19805 14822 19808
rect 14856 19805 14868 19839
rect 15194 19836 15200 19848
rect 15155 19808 15200 19836
rect 14810 19799 14868 19805
rect 12060 19771 12118 19777
rect 9416 19740 10456 19768
rect 9309 19731 9367 19737
rect 4341 19703 4399 19709
rect 4341 19669 4353 19703
rect 4387 19669 4399 19703
rect 7466 19700 7472 19712
rect 7427 19672 7472 19700
rect 4341 19663 4399 19669
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 8573 19703 8631 19709
rect 8573 19669 8585 19703
rect 8619 19700 8631 19703
rect 8662 19700 8668 19712
rect 8619 19672 8668 19700
rect 8619 19669 8631 19672
rect 8573 19663 8631 19669
rect 8662 19660 8668 19672
rect 8720 19660 8726 19712
rect 10229 19703 10287 19709
rect 10229 19669 10241 19703
rect 10275 19700 10287 19703
rect 10318 19700 10324 19712
rect 10275 19672 10324 19700
rect 10275 19669 10287 19672
rect 10229 19663 10287 19669
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 10428 19700 10456 19740
rect 12060 19737 12072 19771
rect 12106 19768 12118 19771
rect 12158 19768 12164 19780
rect 12106 19740 12164 19768
rect 12106 19737 12118 19740
rect 12060 19731 12118 19737
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 13998 19728 14004 19780
rect 14056 19768 14062 19780
rect 14660 19768 14688 19799
rect 15194 19796 15200 19808
rect 15252 19796 15258 19848
rect 25133 19839 25191 19845
rect 25133 19805 25145 19839
rect 25179 19836 25191 19839
rect 25332 19836 25360 20003
rect 25179 19808 25360 19836
rect 25179 19805 25191 19808
rect 25133 19799 25191 19805
rect 14918 19768 14924 19780
rect 14056 19740 14924 19768
rect 14056 19728 14062 19740
rect 14918 19728 14924 19740
rect 14976 19728 14982 19780
rect 15381 19771 15439 19777
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 15718 19771 15776 19777
rect 15718 19768 15730 19771
rect 15427 19740 15730 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 15718 19737 15730 19740
rect 15764 19737 15776 19771
rect 15718 19731 15776 19737
rect 16758 19728 16764 19780
rect 16816 19768 16822 19780
rect 17497 19771 17555 19777
rect 17497 19768 17509 19771
rect 16816 19740 17509 19768
rect 16816 19728 16822 19740
rect 17497 19737 17509 19740
rect 17543 19737 17555 19771
rect 18325 19771 18383 19777
rect 18325 19768 18337 19771
rect 17497 19731 17555 19737
rect 18064 19740 18337 19768
rect 18064 19712 18092 19740
rect 18325 19737 18337 19740
rect 18371 19737 18383 19771
rect 18325 19731 18383 19737
rect 12618 19700 12624 19712
rect 10428 19672 12624 19700
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 13262 19660 13268 19712
rect 13320 19700 13326 19712
rect 16666 19700 16672 19712
rect 13320 19672 16672 19700
rect 13320 19660 13326 19672
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 16850 19700 16856 19712
rect 16811 19672 16856 19700
rect 16850 19660 16856 19672
rect 16908 19660 16914 19712
rect 17034 19700 17040 19712
rect 16995 19672 17040 19700
rect 17034 19660 17040 19672
rect 17092 19660 17098 19712
rect 17402 19700 17408 19712
rect 17363 19672 17408 19700
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 18046 19700 18052 19712
rect 18007 19672 18052 19700
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 18414 19700 18420 19712
rect 18375 19672 18420 19700
rect 18414 19660 18420 19672
rect 18472 19660 18478 19712
rect 22189 19703 22247 19709
rect 22189 19669 22201 19703
rect 22235 19700 22247 19703
rect 22462 19700 22468 19712
rect 22235 19672 22468 19700
rect 22235 19669 22247 19672
rect 22189 19663 22247 19669
rect 22462 19660 22468 19672
rect 22520 19660 22526 19712
rect 22554 19660 22560 19712
rect 22612 19700 22618 19712
rect 22741 19703 22799 19709
rect 22741 19700 22753 19703
rect 22612 19672 22753 19700
rect 22612 19660 22618 19672
rect 22741 19669 22753 19672
rect 22787 19669 22799 19703
rect 22741 19663 22799 19669
rect 22830 19660 22836 19712
rect 22888 19700 22894 19712
rect 25038 19700 25044 19712
rect 22888 19672 22933 19700
rect 24999 19672 25044 19700
rect 22888 19660 22894 19672
rect 25038 19660 25044 19672
rect 25096 19660 25102 19712
rect 1104 19610 26220 19632
rect 1104 19558 9322 19610
rect 9374 19558 9386 19610
rect 9438 19558 9450 19610
rect 9502 19558 9514 19610
rect 9566 19558 9578 19610
rect 9630 19558 17694 19610
rect 17746 19558 17758 19610
rect 17810 19558 17822 19610
rect 17874 19558 17886 19610
rect 17938 19558 17950 19610
rect 18002 19558 26220 19610
rect 1104 19536 26220 19558
rect 4338 19496 4344 19508
rect 4299 19468 4344 19496
rect 4338 19456 4344 19468
rect 4396 19456 4402 19508
rect 4522 19496 4528 19508
rect 4483 19468 4528 19496
rect 4522 19456 4528 19468
rect 4580 19456 4586 19508
rect 6089 19499 6147 19505
rect 6089 19465 6101 19499
rect 6135 19465 6147 19499
rect 6089 19459 6147 19465
rect 3881 19431 3939 19437
rect 3881 19397 3893 19431
rect 3927 19428 3939 19431
rect 6104 19428 6132 19459
rect 7098 19456 7104 19508
rect 7156 19496 7162 19508
rect 7469 19499 7527 19505
rect 7469 19496 7481 19499
rect 7156 19468 7481 19496
rect 7156 19456 7162 19468
rect 7469 19465 7481 19468
rect 7515 19465 7527 19499
rect 7469 19459 7527 19465
rect 10505 19499 10563 19505
rect 10505 19465 10517 19499
rect 10551 19465 10563 19499
rect 12158 19496 12164 19508
rect 12119 19468 12164 19496
rect 10505 19459 10563 19465
rect 8386 19428 8392 19440
rect 3927 19400 6592 19428
rect 3927 19397 3939 19400
rect 3881 19391 3939 19397
rect 2958 19360 2964 19372
rect 2919 19332 2964 19360
rect 2958 19320 2964 19332
rect 3016 19320 3022 19372
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19360 3111 19363
rect 3234 19360 3240 19372
rect 3099 19332 3240 19360
rect 3099 19329 3111 19332
rect 3053 19323 3111 19329
rect 3234 19320 3240 19332
rect 3292 19320 3298 19372
rect 3970 19360 3976 19372
rect 3931 19332 3976 19360
rect 3970 19320 3976 19332
rect 4028 19320 4034 19372
rect 6564 19369 6592 19400
rect 7668 19400 8392 19428
rect 7377 19387 7435 19393
rect 4976 19363 5034 19369
rect 4976 19329 4988 19363
rect 5022 19360 5034 19363
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 5022 19332 6377 19360
rect 5022 19329 5034 19332
rect 4976 19323 5034 19329
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 6549 19363 6607 19369
rect 6549 19329 6561 19363
rect 6595 19329 6607 19363
rect 6730 19360 6736 19372
rect 6691 19332 6736 19360
rect 6549 19323 6607 19329
rect 6730 19320 6736 19332
rect 6788 19320 6794 19372
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7101 19363 7159 19369
rect 6972 19332 7017 19360
rect 6972 19320 6978 19332
rect 7101 19329 7113 19363
rect 7147 19360 7159 19363
rect 7282 19360 7288 19372
rect 7147 19332 7288 19360
rect 7147 19329 7159 19332
rect 7101 19323 7159 19329
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7377 19353 7389 19387
rect 7423 19353 7435 19387
rect 7668 19369 7696 19400
rect 8386 19388 8392 19400
rect 8444 19388 8450 19440
rect 8481 19431 8539 19437
rect 8481 19397 8493 19431
rect 8527 19428 8539 19431
rect 8938 19428 8944 19440
rect 8527 19400 8944 19428
rect 8527 19397 8539 19400
rect 8481 19391 8539 19397
rect 8938 19388 8944 19400
rect 8996 19388 9002 19440
rect 9033 19431 9091 19437
rect 9033 19397 9045 19431
rect 9079 19428 9091 19431
rect 9370 19431 9428 19437
rect 9370 19428 9382 19431
rect 9079 19400 9382 19428
rect 9079 19397 9091 19400
rect 9033 19391 9091 19397
rect 9370 19397 9382 19400
rect 9416 19397 9428 19431
rect 9370 19391 9428 19397
rect 7377 19347 7435 19353
rect 7653 19363 7711 19369
rect 7392 19304 7420 19347
rect 7653 19329 7665 19363
rect 7699 19329 7711 19363
rect 7653 19323 7711 19329
rect 8297 19363 8355 19369
rect 8297 19329 8309 19363
rect 8343 19329 8355 19363
rect 8662 19360 8668 19372
rect 8623 19332 8668 19360
rect 8297 19323 8355 19329
rect 3329 19295 3387 19301
rect 3329 19261 3341 19295
rect 3375 19292 3387 19295
rect 3513 19295 3571 19301
rect 3513 19292 3525 19295
rect 3375 19264 3525 19292
rect 3375 19261 3387 19264
rect 3329 19255 3387 19261
rect 3513 19261 3525 19264
rect 3559 19292 3571 19295
rect 3789 19295 3847 19301
rect 3789 19292 3801 19295
rect 3559 19264 3801 19292
rect 3559 19261 3571 19264
rect 3513 19255 3571 19261
rect 3789 19261 3801 19264
rect 3835 19292 3847 19295
rect 4522 19292 4528 19304
rect 3835 19264 4528 19292
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 4706 19292 4712 19304
rect 4667 19264 4712 19292
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 6638 19252 6644 19304
rect 6696 19292 6702 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6696 19264 6837 19292
rect 6696 19252 6702 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 7374 19292 7380 19304
rect 7287 19264 7380 19292
rect 6825 19255 6883 19261
rect 3237 19227 3295 19233
rect 3237 19193 3249 19227
rect 3283 19224 3295 19227
rect 4062 19224 4068 19236
rect 3283 19196 4068 19224
rect 3283 19193 3295 19196
rect 3237 19187 3295 19193
rect 4062 19184 4068 19196
rect 4120 19184 4126 19236
rect 6840 19224 6868 19255
rect 7374 19252 7380 19264
rect 7432 19292 7438 19304
rect 8113 19295 8171 19301
rect 8113 19292 8125 19295
rect 7432 19264 8125 19292
rect 7432 19252 7438 19264
rect 8113 19261 8125 19264
rect 8159 19261 8171 19295
rect 8312 19292 8340 19323
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 8849 19363 8907 19369
rect 8849 19329 8861 19363
rect 8895 19360 8907 19363
rect 10226 19360 10232 19372
rect 8895 19332 10232 19360
rect 8895 19329 8907 19332
rect 8849 19323 8907 19329
rect 10226 19320 10232 19332
rect 10284 19320 10290 19372
rect 10520 19360 10548 19459
rect 12158 19456 12164 19468
rect 12216 19456 12222 19508
rect 12618 19496 12624 19508
rect 12531 19468 12624 19496
rect 12618 19456 12624 19468
rect 12676 19496 12682 19508
rect 14642 19496 14648 19508
rect 12676 19468 14648 19496
rect 12676 19456 12682 19468
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 15565 19499 15623 19505
rect 15565 19496 15577 19499
rect 15252 19468 15577 19496
rect 15252 19456 15258 19468
rect 15565 19465 15577 19468
rect 15611 19496 15623 19499
rect 16850 19496 16856 19508
rect 15611 19468 16856 19496
rect 15611 19465 15623 19468
rect 15565 19459 15623 19465
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 17497 19499 17555 19505
rect 17497 19465 17509 19499
rect 17543 19496 17555 19499
rect 18230 19496 18236 19508
rect 17543 19468 18236 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 18230 19456 18236 19468
rect 18288 19496 18294 19508
rect 18598 19496 18604 19508
rect 18288 19468 18604 19496
rect 18288 19456 18294 19468
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 20346 19496 20352 19508
rect 19392 19468 20352 19496
rect 19392 19456 19398 19468
rect 20346 19456 20352 19468
rect 20404 19456 20410 19508
rect 22281 19499 22339 19505
rect 22281 19465 22293 19499
rect 22327 19496 22339 19499
rect 22370 19496 22376 19508
rect 22327 19468 22376 19496
rect 22327 19465 22339 19468
rect 22281 19459 22339 19465
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 22554 19496 22560 19508
rect 22515 19468 22560 19496
rect 22554 19456 22560 19468
rect 22612 19456 22618 19508
rect 12434 19428 12440 19440
rect 11808 19400 12440 19428
rect 10689 19363 10747 19369
rect 10689 19360 10701 19363
rect 10520 19332 10701 19360
rect 10689 19329 10701 19332
rect 10735 19329 10747 19363
rect 10689 19323 10747 19329
rect 11422 19320 11428 19372
rect 11480 19360 11486 19372
rect 11517 19363 11575 19369
rect 11517 19360 11529 19363
rect 11480 19332 11529 19360
rect 11480 19320 11486 19332
rect 11517 19329 11529 19332
rect 11563 19329 11575 19363
rect 11698 19360 11704 19372
rect 11659 19332 11704 19360
rect 11517 19323 11575 19329
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 11808 19369 11836 19400
rect 12434 19388 12440 19400
rect 12492 19388 12498 19440
rect 15746 19428 15752 19440
rect 14108 19400 15752 19428
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19329 11851 19363
rect 12066 19360 12072 19372
rect 12027 19332 12072 19360
rect 11793 19323 11851 19329
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 12345 19363 12403 19369
rect 12345 19329 12357 19363
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 8938 19292 8944 19304
rect 8312 19264 8944 19292
rect 8113 19255 8171 19261
rect 8938 19252 8944 19264
rect 8996 19252 9002 19304
rect 9122 19292 9128 19304
rect 9083 19264 9128 19292
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 11882 19252 11888 19304
rect 11940 19292 11946 19304
rect 11940 19264 11985 19292
rect 11940 19252 11946 19264
rect 7193 19227 7251 19233
rect 7193 19224 7205 19227
rect 6840 19196 7205 19224
rect 7193 19193 7205 19196
rect 7239 19193 7251 19227
rect 12158 19224 12164 19236
rect 7193 19187 7251 19193
rect 10612 19196 12164 19224
rect 2774 19116 2780 19168
rect 2832 19156 2838 19168
rect 2832 19128 2877 19156
rect 2832 19116 2838 19128
rect 7834 19116 7840 19168
rect 7892 19156 7898 19168
rect 7929 19159 7987 19165
rect 7929 19156 7941 19159
rect 7892 19128 7941 19156
rect 7892 19116 7898 19128
rect 7929 19125 7941 19128
rect 7975 19156 7987 19159
rect 8662 19156 8668 19168
rect 7975 19128 8668 19156
rect 7975 19125 7987 19128
rect 7929 19119 7987 19125
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 8846 19116 8852 19168
rect 8904 19156 8910 19168
rect 10612 19156 10640 19196
rect 12158 19184 12164 19196
rect 12216 19224 12222 19236
rect 12360 19224 12388 19323
rect 12618 19320 12624 19372
rect 12676 19360 12682 19372
rect 12805 19363 12863 19369
rect 12805 19360 12817 19363
rect 12676 19332 12817 19360
rect 12676 19320 12682 19332
rect 12805 19329 12817 19332
rect 12851 19360 12863 19363
rect 13357 19363 13415 19369
rect 13357 19360 13369 19363
rect 12851 19332 13369 19360
rect 12851 19329 12863 19332
rect 12805 19323 12863 19329
rect 13357 19329 13369 19332
rect 13403 19329 13415 19363
rect 13998 19360 14004 19372
rect 13357 19323 13415 19329
rect 13740 19332 14004 19360
rect 13740 19292 13768 19332
rect 13998 19320 14004 19332
rect 14056 19320 14062 19372
rect 13556 19264 13768 19292
rect 14108 19292 14136 19400
rect 15746 19388 15752 19400
rect 15804 19388 15810 19440
rect 17954 19388 17960 19440
rect 18012 19428 18018 19440
rect 19214 19431 19272 19437
rect 19214 19428 19226 19431
rect 18012 19400 19226 19428
rect 18012 19388 18018 19400
rect 19214 19397 19226 19400
rect 19260 19397 19272 19431
rect 19214 19391 19272 19397
rect 23017 19431 23075 19437
rect 23017 19397 23029 19431
rect 23063 19428 23075 19431
rect 23106 19428 23112 19440
rect 23063 19400 23112 19428
rect 23063 19397 23075 19400
rect 23017 19391 23075 19397
rect 23106 19388 23112 19400
rect 23164 19388 23170 19440
rect 14182 19320 14188 19372
rect 14240 19360 14246 19372
rect 14240 19332 14284 19360
rect 14240 19320 14246 19332
rect 14458 19320 14464 19372
rect 14516 19360 14522 19372
rect 14553 19363 14611 19369
rect 14553 19360 14565 19363
rect 14516 19332 14565 19360
rect 14516 19320 14522 19332
rect 14553 19329 14565 19332
rect 14599 19329 14611 19363
rect 14553 19323 14611 19329
rect 16666 19320 16672 19372
rect 16724 19360 16730 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16724 19332 16865 19360
rect 16724 19320 16730 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 18230 19320 18236 19372
rect 18288 19360 18294 19372
rect 18610 19363 18668 19369
rect 18610 19360 18622 19363
rect 18288 19332 18622 19360
rect 18288 19320 18294 19332
rect 18610 19329 18622 19332
rect 18656 19329 18668 19363
rect 18610 19323 18668 19329
rect 22462 19320 22468 19372
rect 22520 19360 22526 19372
rect 22830 19360 22836 19372
rect 22520 19332 22836 19360
rect 22520 19320 22526 19332
rect 22830 19320 22836 19332
rect 22888 19360 22894 19372
rect 22925 19363 22983 19369
rect 22925 19360 22937 19363
rect 22888 19332 22937 19360
rect 22888 19320 22894 19332
rect 22925 19329 22937 19332
rect 22971 19329 22983 19363
rect 22925 19323 22983 19329
rect 14277 19295 14335 19301
rect 14277 19292 14289 19295
rect 14108 19264 14289 19292
rect 13556 19233 13584 19264
rect 14277 19261 14289 19264
rect 14323 19261 14335 19295
rect 14277 19255 14335 19261
rect 14369 19295 14427 19301
rect 14369 19261 14381 19295
rect 14415 19292 14427 19295
rect 15286 19292 15292 19304
rect 14415 19264 15292 19292
rect 14415 19261 14427 19264
rect 14369 19255 14427 19261
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 18877 19295 18935 19301
rect 18877 19261 18889 19295
rect 18923 19292 18935 19295
rect 18966 19292 18972 19304
rect 18923 19264 18972 19292
rect 18923 19261 18935 19264
rect 18877 19255 18935 19261
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 22373 19295 22431 19301
rect 22373 19261 22385 19295
rect 22419 19292 22431 19295
rect 23109 19295 23167 19301
rect 23109 19292 23121 19295
rect 22419 19264 23121 19292
rect 22419 19261 22431 19264
rect 22373 19255 22431 19261
rect 23109 19261 23121 19264
rect 23155 19292 23167 19295
rect 23290 19292 23296 19304
rect 23155 19264 23296 19292
rect 23155 19261 23167 19264
rect 23109 19255 23167 19261
rect 23290 19252 23296 19264
rect 23348 19252 23354 19304
rect 12216 19196 12388 19224
rect 13541 19227 13599 19233
rect 12216 19184 12222 19196
rect 13541 19193 13553 19227
rect 13587 19193 13599 19227
rect 25038 19224 25044 19236
rect 13541 19187 13599 19193
rect 22066 19196 25044 19224
rect 10778 19156 10784 19168
rect 8904 19128 10640 19156
rect 10739 19128 10784 19156
rect 8904 19116 8910 19128
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12529 19159 12587 19165
rect 12529 19156 12541 19159
rect 12492 19128 12541 19156
rect 12492 19116 12498 19128
rect 12529 19125 12541 19128
rect 12575 19156 12587 19159
rect 12894 19156 12900 19168
rect 12575 19128 12900 19156
rect 12575 19125 12587 19128
rect 12529 19119 12587 19125
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 14642 19156 14648 19168
rect 14603 19128 14648 19156
rect 14642 19116 14648 19128
rect 14700 19116 14706 19168
rect 14826 19116 14832 19168
rect 14884 19156 14890 19168
rect 22066 19156 22094 19196
rect 25038 19184 25044 19196
rect 25096 19184 25102 19236
rect 14884 19128 22094 19156
rect 14884 19116 14890 19128
rect 22370 19116 22376 19168
rect 22428 19156 22434 19168
rect 23198 19156 23204 19168
rect 22428 19128 23204 19156
rect 22428 19116 22434 19128
rect 23198 19116 23204 19128
rect 23256 19116 23262 19168
rect 1104 19066 26220 19088
rect 1104 19014 5136 19066
rect 5188 19014 5200 19066
rect 5252 19014 5264 19066
rect 5316 19014 5328 19066
rect 5380 19014 5392 19066
rect 5444 19014 13508 19066
rect 13560 19014 13572 19066
rect 13624 19014 13636 19066
rect 13688 19014 13700 19066
rect 13752 19014 13764 19066
rect 13816 19014 21880 19066
rect 21932 19014 21944 19066
rect 21996 19014 22008 19066
rect 22060 19014 22072 19066
rect 22124 19014 22136 19066
rect 22188 19014 26220 19066
rect 1104 18992 26220 19014
rect 3513 18955 3571 18961
rect 3513 18921 3525 18955
rect 3559 18952 3571 18955
rect 3970 18952 3976 18964
rect 3559 18924 3976 18952
rect 3559 18921 3571 18924
rect 3513 18915 3571 18921
rect 3970 18912 3976 18924
rect 4028 18912 4034 18964
rect 6181 18955 6239 18961
rect 6181 18921 6193 18955
rect 6227 18952 6239 18955
rect 6730 18952 6736 18964
rect 6227 18924 6736 18952
rect 6227 18921 6239 18924
rect 6181 18915 6239 18921
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 7653 18955 7711 18961
rect 7653 18921 7665 18955
rect 7699 18952 7711 18955
rect 7742 18952 7748 18964
rect 7699 18924 7748 18952
rect 7699 18921 7711 18924
rect 7653 18915 7711 18921
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 8846 18912 8852 18964
rect 8904 18952 8910 18964
rect 9125 18955 9183 18961
rect 9125 18952 9137 18955
rect 8904 18924 9137 18952
rect 8904 18912 8910 18924
rect 9125 18921 9137 18924
rect 9171 18921 9183 18955
rect 10226 18952 10232 18964
rect 10187 18924 10232 18952
rect 9125 18915 9183 18921
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 11701 18955 11759 18961
rect 11701 18921 11713 18955
rect 11747 18952 11759 18955
rect 12066 18952 12072 18964
rect 11747 18924 12072 18952
rect 11747 18921 11759 18924
rect 11701 18915 11759 18921
rect 12066 18912 12072 18924
rect 12124 18912 12130 18964
rect 15286 18912 15292 18964
rect 15344 18952 15350 18964
rect 15657 18955 15715 18961
rect 15657 18952 15669 18955
rect 15344 18924 15669 18952
rect 15344 18912 15350 18924
rect 15657 18921 15669 18924
rect 15703 18921 15715 18955
rect 15657 18915 15715 18921
rect 15746 18912 15752 18964
rect 15804 18952 15810 18964
rect 15933 18955 15991 18961
rect 15933 18952 15945 18955
rect 15804 18924 15945 18952
rect 15804 18912 15810 18924
rect 15933 18921 15945 18924
rect 15979 18921 15991 18955
rect 15933 18915 15991 18921
rect 17126 18912 17132 18964
rect 17184 18952 17190 18964
rect 17221 18955 17279 18961
rect 17221 18952 17233 18955
rect 17184 18924 17233 18952
rect 17184 18912 17190 18924
rect 17221 18921 17233 18924
rect 17267 18921 17279 18955
rect 17221 18915 17279 18921
rect 17862 18912 17868 18964
rect 17920 18952 17926 18964
rect 18049 18955 18107 18961
rect 18049 18952 18061 18955
rect 17920 18924 18061 18952
rect 17920 18912 17926 18924
rect 18049 18921 18061 18924
rect 18095 18921 18107 18955
rect 18506 18952 18512 18964
rect 18049 18915 18107 18921
rect 18156 18924 18512 18952
rect 7190 18844 7196 18896
rect 7248 18884 7254 18896
rect 8021 18887 8079 18893
rect 8021 18884 8033 18887
rect 7248 18856 8033 18884
rect 7248 18844 7254 18856
rect 8021 18853 8033 18856
rect 8067 18884 8079 18887
rect 8386 18884 8392 18896
rect 8067 18856 8392 18884
rect 8067 18853 8079 18856
rect 8021 18847 8079 18853
rect 8386 18844 8392 18856
rect 8444 18884 8450 18896
rect 9674 18884 9680 18896
rect 8444 18856 9352 18884
rect 8444 18844 8450 18856
rect 6914 18816 6920 18828
rect 6827 18788 6920 18816
rect 6914 18776 6920 18788
rect 6972 18816 6978 18828
rect 8757 18819 8815 18825
rect 6972 18788 8708 18816
rect 6972 18776 6978 18788
rect 2130 18748 2136 18760
rect 2043 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18748 2194 18760
rect 4706 18748 4712 18760
rect 2188 18720 4712 18748
rect 2188 18708 2194 18720
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 6365 18751 6423 18757
rect 6365 18717 6377 18751
rect 6411 18748 6423 18751
rect 6546 18748 6552 18760
rect 6411 18720 6552 18748
rect 6411 18717 6423 18720
rect 6365 18711 6423 18717
rect 6546 18708 6552 18720
rect 6604 18748 6610 18760
rect 6641 18751 6699 18757
rect 6641 18748 6653 18751
rect 6604 18720 6653 18748
rect 6604 18708 6610 18720
rect 6641 18717 6653 18720
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 6733 18751 6791 18757
rect 6733 18717 6745 18751
rect 6779 18748 6791 18751
rect 7006 18748 7012 18760
rect 6779 18720 7012 18748
rect 6779 18717 6791 18720
rect 6733 18711 6791 18717
rect 7006 18708 7012 18720
rect 7064 18748 7070 18760
rect 7374 18748 7380 18760
rect 7064 18720 7380 18748
rect 7064 18708 7070 18720
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18748 7527 18751
rect 7650 18748 7656 18760
rect 7515 18720 7656 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 7650 18708 7656 18720
rect 7708 18708 7714 18760
rect 7837 18751 7895 18757
rect 7837 18717 7849 18751
rect 7883 18748 7895 18751
rect 8018 18748 8024 18760
rect 7883 18720 8024 18748
rect 7883 18717 7895 18720
rect 7837 18711 7895 18717
rect 8018 18708 8024 18720
rect 8076 18708 8082 18760
rect 8386 18748 8392 18760
rect 8347 18720 8392 18748
rect 8386 18708 8392 18720
rect 8444 18708 8450 18760
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18717 8631 18751
rect 8680 18748 8708 18788
rect 8757 18785 8769 18819
rect 8803 18816 8815 18819
rect 8803 18788 9260 18816
rect 8803 18785 8815 18788
rect 8757 18779 8815 18785
rect 9232 18760 9260 18788
rect 8938 18748 8944 18760
rect 8680 18720 8800 18748
rect 8899 18720 8944 18748
rect 8573 18711 8631 18717
rect 2400 18683 2458 18689
rect 2400 18649 2412 18683
rect 2446 18680 2458 18683
rect 3418 18680 3424 18692
rect 2446 18652 3424 18680
rect 2446 18649 2458 18652
rect 2400 18643 2458 18649
rect 3418 18640 3424 18652
rect 3476 18640 3482 18692
rect 8297 18683 8355 18689
rect 8297 18680 8309 18683
rect 6748 18652 8309 18680
rect 2498 18572 2504 18624
rect 2556 18612 2562 18624
rect 6748 18612 6776 18652
rect 8297 18649 8309 18652
rect 8343 18680 8355 18683
rect 8588 18680 8616 18711
rect 8662 18680 8668 18692
rect 8343 18652 8668 18680
rect 8343 18649 8355 18652
rect 8297 18643 8355 18649
rect 8662 18640 8668 18652
rect 8720 18640 8726 18692
rect 8772 18680 8800 18720
rect 8938 18708 8944 18720
rect 8996 18708 9002 18760
rect 9214 18748 9220 18760
rect 9175 18720 9220 18748
rect 9214 18708 9220 18720
rect 9272 18708 9278 18760
rect 8846 18680 8852 18692
rect 8772 18652 8852 18680
rect 8846 18640 8852 18652
rect 8904 18640 8910 18692
rect 9324 18680 9352 18856
rect 9416 18856 9680 18884
rect 9416 18757 9444 18856
rect 9674 18844 9680 18856
rect 9732 18844 9738 18896
rect 18156 18884 18184 18924
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 19061 18955 19119 18961
rect 19061 18921 19073 18955
rect 19107 18952 19119 18955
rect 20625 18955 20683 18961
rect 20625 18952 20637 18955
rect 19107 18924 20637 18952
rect 19107 18921 19119 18924
rect 19061 18915 19119 18921
rect 20625 18921 20637 18924
rect 20671 18921 20683 18955
rect 20625 18915 20683 18921
rect 18874 18884 18880 18896
rect 17696 18856 18184 18884
rect 18248 18856 18880 18884
rect 9861 18819 9919 18825
rect 9861 18785 9873 18819
rect 9907 18816 9919 18819
rect 10226 18816 10232 18828
rect 9907 18788 10232 18816
rect 9907 18785 9919 18788
rect 9861 18779 9919 18785
rect 10226 18776 10232 18788
rect 10284 18816 10290 18828
rect 10689 18819 10747 18825
rect 10689 18816 10701 18819
rect 10284 18788 10701 18816
rect 10284 18776 10290 18788
rect 10689 18785 10701 18788
rect 10735 18785 10747 18819
rect 10689 18779 10747 18785
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 11149 18819 11207 18825
rect 10836 18788 10881 18816
rect 10836 18776 10842 18788
rect 11149 18785 11161 18819
rect 11195 18816 11207 18819
rect 11698 18816 11704 18828
rect 11195 18788 11704 18816
rect 11195 18785 11207 18788
rect 11149 18779 11207 18785
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 11882 18776 11888 18828
rect 11940 18816 11946 18828
rect 12713 18819 12771 18825
rect 12713 18816 12725 18819
rect 11940 18788 12725 18816
rect 11940 18776 11946 18788
rect 12713 18785 12725 18788
rect 12759 18785 12771 18819
rect 12713 18779 12771 18785
rect 12805 18819 12863 18825
rect 12805 18785 12817 18819
rect 12851 18816 12863 18819
rect 14182 18816 14188 18828
rect 12851 18788 14188 18816
rect 12851 18785 12863 18788
rect 12805 18779 12863 18785
rect 14182 18776 14188 18788
rect 14240 18776 14246 18828
rect 17696 18825 17724 18856
rect 16577 18819 16635 18825
rect 16577 18816 16589 18819
rect 16316 18788 16589 18816
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18717 9459 18751
rect 9401 18711 9459 18717
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18717 9551 18751
rect 9493 18711 9551 18717
rect 9619 18748 9677 18751
rect 9766 18748 9772 18760
rect 9619 18745 9772 18748
rect 9619 18711 9631 18745
rect 9665 18720 9772 18745
rect 9665 18711 9677 18720
rect 9508 18680 9536 18711
rect 9619 18705 9677 18711
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 10134 18708 10140 18760
rect 10192 18748 10198 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 10192 18720 10425 18748
rect 10192 18708 10198 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18717 10563 18751
rect 10796 18748 10824 18776
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 10796 18720 11253 18748
rect 10505 18711 10563 18717
rect 11241 18717 11253 18720
rect 11287 18717 11299 18751
rect 12526 18748 12532 18760
rect 12487 18720 12532 18748
rect 11241 18711 11299 18717
rect 9324 18652 9536 18680
rect 7374 18612 7380 18624
rect 2556 18584 6776 18612
rect 7335 18584 7380 18612
rect 2556 18572 2562 18584
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 9508 18612 9536 18652
rect 9950 18612 9956 18624
rect 9508 18584 9956 18612
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 10520 18612 10548 18711
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 12894 18708 12900 18760
rect 12952 18748 12958 18760
rect 12952 18720 12997 18748
rect 12952 18708 12958 18720
rect 13078 18708 13084 18760
rect 13136 18748 13142 18760
rect 13136 18720 13181 18748
rect 13136 18708 13142 18720
rect 14090 18708 14096 18760
rect 14148 18748 14154 18760
rect 15565 18751 15623 18757
rect 15565 18748 15577 18751
rect 14148 18720 15577 18748
rect 14148 18708 14154 18720
rect 15565 18717 15577 18720
rect 15611 18717 15623 18751
rect 15838 18748 15844 18760
rect 15799 18720 15844 18748
rect 15565 18711 15623 18717
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18717 16175 18751
rect 16117 18711 16175 18717
rect 12342 18640 12348 18692
rect 12400 18680 12406 18692
rect 12400 18652 12848 18680
rect 12400 18640 12406 18652
rect 11054 18612 11060 18624
rect 10520 18584 11060 18612
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 11333 18615 11391 18621
rect 11333 18581 11345 18615
rect 11379 18612 11391 18615
rect 11606 18612 11612 18624
rect 11379 18584 11612 18612
rect 11379 18581 11391 18584
rect 11333 18575 11391 18581
rect 11606 18572 11612 18584
rect 11664 18572 11670 18624
rect 12434 18572 12440 18624
rect 12492 18612 12498 18624
rect 12820 18612 12848 18652
rect 12986 18640 12992 18692
rect 13044 18680 13050 18692
rect 13044 18652 14601 18680
rect 13044 18640 13050 18652
rect 14185 18615 14243 18621
rect 14185 18612 14197 18615
rect 12492 18584 12537 18612
rect 12820 18584 14197 18612
rect 12492 18572 12498 18584
rect 14185 18581 14197 18584
rect 14231 18612 14243 18615
rect 14458 18612 14464 18624
rect 14231 18584 14464 18612
rect 14231 18581 14243 18584
rect 14185 18575 14243 18581
rect 14458 18572 14464 18584
rect 14516 18572 14522 18624
rect 14573 18612 14601 18652
rect 14642 18640 14648 18692
rect 14700 18680 14706 18692
rect 15298 18683 15356 18689
rect 15298 18680 15310 18683
rect 14700 18652 15310 18680
rect 14700 18640 14706 18652
rect 15298 18649 15310 18652
rect 15344 18649 15356 18683
rect 15298 18643 15356 18649
rect 15654 18640 15660 18692
rect 15712 18680 15718 18692
rect 16132 18680 16160 18711
rect 15712 18652 16160 18680
rect 15712 18640 15718 18652
rect 16316 18621 16344 18788
rect 16577 18785 16589 18788
rect 16623 18785 16635 18819
rect 16577 18779 16635 18785
rect 17681 18819 17739 18825
rect 17681 18785 17693 18819
rect 17727 18785 17739 18819
rect 17681 18779 17739 18785
rect 17773 18819 17831 18825
rect 17773 18785 17785 18819
rect 17819 18816 17831 18819
rect 18138 18816 18144 18828
rect 17819 18788 18144 18816
rect 17819 18785 17831 18788
rect 17773 18779 17831 18785
rect 18138 18776 18144 18788
rect 18196 18776 18202 18828
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 17034 18748 17040 18760
rect 16899 18720 17040 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 17034 18708 17040 18720
rect 17092 18708 17098 18760
rect 17310 18708 17316 18760
rect 17368 18748 17374 18760
rect 17405 18751 17463 18757
rect 17405 18748 17417 18751
rect 17368 18720 17417 18748
rect 17368 18708 17374 18720
rect 17405 18717 17417 18720
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 17586 18708 17592 18760
rect 17644 18748 17650 18760
rect 17954 18748 17960 18760
rect 17644 18720 17688 18748
rect 17915 18720 17960 18748
rect 17644 18708 17650 18720
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 18248 18757 18276 18856
rect 18874 18844 18880 18856
rect 18932 18844 18938 18896
rect 18601 18819 18659 18825
rect 18601 18816 18613 18819
rect 18340 18788 18613 18816
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18717 18291 18751
rect 18233 18711 18291 18717
rect 18138 18640 18144 18692
rect 18196 18680 18202 18692
rect 18340 18680 18368 18788
rect 18601 18785 18613 18788
rect 18647 18785 18659 18819
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 18601 18779 18659 18785
rect 18800 18788 19073 18816
rect 18398 18745 18456 18751
rect 18398 18711 18410 18745
rect 18444 18711 18456 18745
rect 18398 18705 18456 18711
rect 18506 18708 18512 18760
rect 18564 18748 18570 18760
rect 18800 18757 18828 18788
rect 19061 18785 19073 18788
rect 19107 18785 19119 18819
rect 20640 18816 20668 18915
rect 21174 18912 21180 18964
rect 21232 18952 21238 18964
rect 21269 18955 21327 18961
rect 21269 18952 21281 18955
rect 21232 18924 21281 18952
rect 21232 18912 21238 18924
rect 21269 18921 21281 18924
rect 21315 18921 21327 18955
rect 21269 18915 21327 18921
rect 21726 18912 21732 18964
rect 21784 18952 21790 18964
rect 22922 18952 22928 18964
rect 21784 18924 22928 18952
rect 21784 18912 21790 18924
rect 22922 18912 22928 18924
rect 22980 18912 22986 18964
rect 20714 18844 20720 18896
rect 20772 18884 20778 18896
rect 21085 18887 21143 18893
rect 21085 18884 21097 18887
rect 20772 18856 21097 18884
rect 20772 18844 20778 18856
rect 21085 18853 21097 18856
rect 21131 18884 21143 18887
rect 21634 18884 21640 18896
rect 21131 18856 21640 18884
rect 21131 18853 21143 18856
rect 21085 18847 21143 18853
rect 21634 18844 21640 18856
rect 21692 18844 21698 18896
rect 20640 18788 21128 18816
rect 19061 18779 19119 18785
rect 18785 18751 18843 18757
rect 18564 18720 18609 18748
rect 18564 18708 18570 18720
rect 18785 18717 18797 18751
rect 18831 18717 18843 18751
rect 18785 18711 18843 18717
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 19024 18720 19257 18748
rect 19024 18708 19030 18720
rect 19245 18717 19257 18720
rect 19291 18748 19303 18751
rect 20714 18748 20720 18760
rect 19291 18720 20720 18748
rect 19291 18717 19303 18720
rect 19245 18711 19303 18717
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 18196 18652 18368 18680
rect 18196 18640 18202 18652
rect 16301 18615 16359 18621
rect 16301 18612 16313 18615
rect 14573 18584 16313 18612
rect 16301 18581 16313 18584
rect 16347 18581 16359 18615
rect 16301 18575 16359 18581
rect 16761 18615 16819 18621
rect 16761 18581 16773 18615
rect 16807 18612 16819 18615
rect 17126 18612 17132 18624
rect 16807 18584 17132 18612
rect 16807 18581 16819 18584
rect 16761 18575 16819 18581
rect 17126 18572 17132 18584
rect 17184 18612 17190 18624
rect 17402 18612 17408 18624
rect 17184 18584 17408 18612
rect 17184 18572 17190 18584
rect 17402 18572 17408 18584
rect 17460 18572 17466 18624
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 18412 18612 18440 18705
rect 19501 18683 19559 18689
rect 19501 18680 19513 18683
rect 19444 18652 19513 18680
rect 17552 18584 18440 18612
rect 18877 18615 18935 18621
rect 17552 18572 17558 18584
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 19444 18612 19472 18652
rect 19501 18649 19513 18652
rect 19547 18649 19559 18683
rect 19501 18643 19559 18649
rect 19886 18640 19892 18692
rect 19944 18680 19950 18692
rect 20901 18683 20959 18689
rect 20901 18680 20913 18683
rect 19944 18652 20913 18680
rect 19944 18640 19950 18652
rect 20901 18649 20913 18652
rect 20947 18649 20959 18683
rect 21100 18680 21128 18788
rect 21634 18708 21640 18760
rect 21692 18748 21698 18760
rect 22649 18751 22707 18757
rect 22649 18748 22661 18751
rect 21692 18720 22661 18748
rect 21692 18708 21698 18720
rect 22649 18717 22661 18720
rect 22695 18748 22707 18751
rect 24210 18748 24216 18760
rect 22695 18720 24216 18748
rect 22695 18717 22707 18720
rect 22649 18711 22707 18717
rect 24210 18708 24216 18720
rect 24268 18708 24274 18760
rect 21100 18652 22094 18680
rect 20901 18643 20959 18649
rect 18923 18584 19472 18612
rect 22066 18612 22094 18652
rect 22370 18640 22376 18692
rect 22428 18689 22434 18692
rect 22428 18680 22440 18689
rect 22428 18652 22473 18680
rect 22428 18643 22440 18652
rect 22428 18640 22434 18643
rect 23382 18640 23388 18692
rect 23440 18680 23446 18692
rect 23946 18683 24004 18689
rect 23946 18680 23958 18683
rect 23440 18652 23958 18680
rect 23440 18640 23446 18652
rect 23946 18649 23958 18652
rect 23992 18649 24004 18683
rect 23946 18643 24004 18649
rect 22554 18612 22560 18624
rect 22066 18584 22560 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 22554 18572 22560 18584
rect 22612 18572 22618 18624
rect 22830 18612 22836 18624
rect 22791 18584 22836 18612
rect 22830 18572 22836 18584
rect 22888 18572 22894 18624
rect 1104 18522 26220 18544
rect 1104 18470 9322 18522
rect 9374 18470 9386 18522
rect 9438 18470 9450 18522
rect 9502 18470 9514 18522
rect 9566 18470 9578 18522
rect 9630 18470 17694 18522
rect 17746 18470 17758 18522
rect 17810 18470 17822 18522
rect 17874 18470 17886 18522
rect 17938 18470 17950 18522
rect 18002 18470 26220 18522
rect 1104 18448 26220 18470
rect 2958 18368 2964 18420
rect 3016 18408 3022 18420
rect 3237 18411 3295 18417
rect 3237 18408 3249 18411
rect 3016 18380 3249 18408
rect 3016 18368 3022 18380
rect 3237 18377 3249 18380
rect 3283 18377 3295 18411
rect 3237 18371 3295 18377
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 3513 18411 3571 18417
rect 3513 18408 3525 18411
rect 3476 18380 3525 18408
rect 3476 18368 3482 18380
rect 3513 18377 3525 18380
rect 3559 18377 3571 18411
rect 8662 18408 8668 18420
rect 8623 18380 8668 18408
rect 3513 18371 3571 18377
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 9585 18411 9643 18417
rect 9585 18377 9597 18411
rect 9631 18408 9643 18411
rect 9674 18408 9680 18420
rect 9631 18380 9680 18408
rect 9631 18377 9643 18380
rect 9585 18371 9643 18377
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 11882 18368 11888 18420
rect 11940 18408 11946 18420
rect 12069 18411 12127 18417
rect 12069 18408 12081 18411
rect 11940 18380 12081 18408
rect 11940 18368 11946 18380
rect 12069 18377 12081 18380
rect 12115 18377 12127 18411
rect 12069 18371 12127 18377
rect 13541 18411 13599 18417
rect 13541 18377 13553 18411
rect 13587 18408 13599 18411
rect 14182 18408 14188 18420
rect 13587 18380 14188 18408
rect 13587 18377 13599 18380
rect 13541 18371 13599 18377
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 15562 18408 15568 18420
rect 15475 18380 15568 18408
rect 15562 18368 15568 18380
rect 15620 18408 15626 18420
rect 17494 18408 17500 18420
rect 15620 18380 17500 18408
rect 15620 18368 15626 18380
rect 17494 18368 17500 18380
rect 17552 18368 17558 18420
rect 18506 18408 18512 18420
rect 17972 18380 18512 18408
rect 2124 18343 2182 18349
rect 2124 18309 2136 18343
rect 2170 18340 2182 18343
rect 2774 18340 2780 18352
rect 2170 18312 2780 18340
rect 2170 18309 2182 18312
rect 2124 18303 2182 18309
rect 2774 18300 2780 18312
rect 2832 18300 2838 18352
rect 4706 18300 4712 18352
rect 4764 18340 4770 18352
rect 4985 18343 5043 18349
rect 4985 18340 4997 18343
rect 4764 18312 4997 18340
rect 4764 18300 4770 18312
rect 4985 18309 4997 18312
rect 5031 18309 5043 18343
rect 4985 18303 5043 18309
rect 5169 18343 5227 18349
rect 5169 18309 5181 18343
rect 5215 18340 5227 18343
rect 7374 18340 7380 18352
rect 5215 18312 7380 18340
rect 5215 18309 5227 18312
rect 5169 18303 5227 18309
rect 7374 18300 7380 18312
rect 7432 18340 7438 18352
rect 12434 18349 12440 18352
rect 9217 18343 9275 18349
rect 9217 18340 9229 18343
rect 7432 18312 9229 18340
rect 7432 18300 7438 18312
rect 9217 18309 9229 18312
rect 9263 18309 9275 18343
rect 9217 18303 9275 18309
rect 12428 18303 12440 18349
rect 12492 18340 12498 18352
rect 12492 18312 12528 18340
rect 12434 18300 12440 18303
rect 12492 18300 12498 18312
rect 16758 18300 16764 18352
rect 16816 18340 16822 18352
rect 16816 18312 17705 18340
rect 16816 18300 16822 18312
rect 17677 18284 17705 18312
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18272 1915 18275
rect 1946 18272 1952 18284
rect 1903 18244 1952 18272
rect 1903 18241 1915 18244
rect 1857 18235 1915 18241
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 3694 18272 3700 18284
rect 3655 18244 3700 18272
rect 3694 18232 3700 18244
rect 3752 18232 3758 18284
rect 3786 18232 3792 18284
rect 3844 18272 3850 18284
rect 3844 18244 3937 18272
rect 3844 18232 3850 18244
rect 3970 18232 3976 18284
rect 4028 18272 4034 18284
rect 4065 18275 4123 18281
rect 4065 18272 4077 18275
rect 4028 18244 4077 18272
rect 4028 18232 4034 18244
rect 4065 18241 4077 18244
rect 4111 18241 4123 18275
rect 6546 18272 6552 18284
rect 6507 18244 6552 18272
rect 4065 18235 4123 18241
rect 6546 18232 6552 18244
rect 6604 18232 6610 18284
rect 7006 18272 7012 18284
rect 6967 18244 7012 18272
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 8662 18232 8668 18284
rect 8720 18272 8726 18284
rect 8849 18275 8907 18281
rect 8849 18272 8861 18275
rect 8720 18244 8861 18272
rect 8720 18232 8726 18244
rect 8849 18241 8861 18244
rect 8895 18241 8907 18275
rect 9674 18272 9680 18284
rect 9635 18244 9680 18272
rect 8849 18235 8907 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 9766 18232 9772 18284
rect 9824 18272 9830 18284
rect 9953 18275 10011 18281
rect 9953 18272 9965 18275
rect 9824 18244 9965 18272
rect 9824 18232 9830 18244
rect 9953 18241 9965 18244
rect 9999 18241 10011 18275
rect 10226 18272 10232 18284
rect 10187 18244 10232 18272
rect 9953 18235 10011 18241
rect 10226 18232 10232 18244
rect 10284 18232 10290 18284
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 10502 18272 10508 18284
rect 10367 18244 10508 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 10502 18232 10508 18244
rect 10560 18232 10566 18284
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18272 11759 18275
rect 11885 18275 11943 18281
rect 11885 18272 11897 18275
rect 11747 18244 11897 18272
rect 11747 18241 11759 18244
rect 11701 18235 11759 18241
rect 11885 18241 11897 18244
rect 11931 18272 11943 18275
rect 12986 18272 12992 18284
rect 11931 18244 12992 18272
rect 11931 18241 11943 18244
rect 11885 18235 11943 18241
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 14274 18232 14280 18284
rect 14332 18272 14338 18284
rect 14441 18275 14499 18281
rect 14441 18272 14453 18275
rect 14332 18244 14453 18272
rect 14332 18232 14338 18244
rect 14441 18241 14453 18244
rect 14487 18241 14499 18275
rect 17494 18272 17500 18284
rect 17455 18244 17500 18272
rect 14441 18235 14499 18241
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 17662 18278 17720 18284
rect 17662 18244 17674 18278
rect 17708 18244 17720 18278
rect 17662 18238 17720 18244
rect 17780 18275 17838 18281
rect 17780 18241 17792 18275
rect 17826 18272 17838 18275
rect 17972 18272 18000 18380
rect 18506 18368 18512 18380
rect 18564 18368 18570 18420
rect 19610 18368 19616 18420
rect 19668 18408 19674 18420
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 19668 18380 19809 18408
rect 19668 18368 19674 18380
rect 19797 18377 19809 18380
rect 19843 18377 19855 18411
rect 20990 18408 20996 18420
rect 19797 18371 19855 18377
rect 19904 18380 20996 18408
rect 18598 18340 18604 18352
rect 18110 18312 18604 18340
rect 18110 18296 18138 18312
rect 18598 18300 18604 18312
rect 18656 18300 18662 18352
rect 19904 18340 19932 18380
rect 20990 18368 20996 18380
rect 21048 18408 21054 18420
rect 21177 18411 21235 18417
rect 21177 18408 21189 18411
rect 21048 18380 21189 18408
rect 21048 18368 21054 18380
rect 21177 18377 21189 18380
rect 21223 18377 21235 18411
rect 21177 18371 21235 18377
rect 21358 18368 21364 18420
rect 21416 18408 21422 18420
rect 21416 18380 22416 18408
rect 21416 18368 21422 18380
rect 18800 18312 19932 18340
rect 18063 18281 18138 18296
rect 18800 18284 18828 18312
rect 17826 18244 18000 18272
rect 18049 18275 18138 18281
rect 17826 18241 17838 18244
rect 17780 18235 17838 18241
rect 18049 18241 18061 18275
rect 18095 18268 18138 18275
rect 18325 18275 18383 18281
rect 18095 18241 18107 18268
rect 18049 18235 18107 18241
rect 18325 18241 18337 18275
rect 18371 18272 18383 18275
rect 18371 18244 18644 18272
rect 18371 18241 18383 18244
rect 18325 18235 18383 18241
rect 3142 18164 3148 18216
rect 3200 18204 3206 18216
rect 3803 18204 3831 18232
rect 3200 18176 3831 18204
rect 3200 18164 3206 18176
rect 7650 18164 7656 18216
rect 7708 18204 7714 18216
rect 7708 18176 11744 18204
rect 7708 18164 7714 18176
rect 9122 18096 9128 18148
rect 9180 18136 9186 18148
rect 9398 18136 9404 18148
rect 9180 18108 9404 18136
rect 9180 18096 9186 18108
rect 9398 18096 9404 18108
rect 9456 18096 9462 18148
rect 10137 18139 10195 18145
rect 10137 18105 10149 18139
rect 10183 18136 10195 18139
rect 10594 18136 10600 18148
rect 10183 18108 10600 18136
rect 10183 18105 10195 18108
rect 10137 18099 10195 18105
rect 10594 18096 10600 18108
rect 10652 18096 10658 18148
rect 11716 18136 11744 18176
rect 11790 18164 11796 18216
rect 11848 18204 11854 18216
rect 12161 18207 12219 18213
rect 12161 18204 12173 18207
rect 11848 18176 12173 18204
rect 11848 18164 11854 18176
rect 12161 18173 12173 18176
rect 12207 18173 12219 18207
rect 12161 18167 12219 18173
rect 14090 18164 14096 18216
rect 14148 18204 14154 18216
rect 14185 18207 14243 18213
rect 14185 18204 14197 18207
rect 14148 18176 14197 18204
rect 14148 18164 14154 18176
rect 14185 18173 14197 18176
rect 14231 18173 14243 18207
rect 17862 18204 17868 18216
rect 17823 18176 17868 18204
rect 14185 18167 14243 18173
rect 17862 18164 17868 18176
rect 17920 18164 17926 18216
rect 18138 18164 18144 18216
rect 18196 18204 18202 18216
rect 18616 18204 18644 18244
rect 18782 18232 18788 18284
rect 18840 18272 18846 18284
rect 18840 18244 18885 18272
rect 18840 18232 18846 18244
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 19886 18272 19892 18284
rect 19300 18244 19892 18272
rect 19300 18232 19306 18244
rect 19886 18232 19892 18244
rect 19944 18232 19950 18284
rect 20162 18272 20168 18284
rect 20123 18244 20168 18272
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18272 20315 18275
rect 20346 18272 20352 18284
rect 20303 18244 20352 18272
rect 20303 18241 20315 18244
rect 20257 18235 20315 18241
rect 20346 18232 20352 18244
rect 20404 18232 20410 18284
rect 21082 18232 21088 18284
rect 21140 18272 21146 18284
rect 21361 18275 21419 18281
rect 21361 18272 21373 18275
rect 21140 18244 21373 18272
rect 21140 18232 21146 18244
rect 21361 18241 21373 18244
rect 21407 18272 21419 18275
rect 21453 18275 21511 18281
rect 21453 18272 21465 18275
rect 21407 18244 21465 18272
rect 21407 18241 21419 18244
rect 21361 18235 21419 18241
rect 21453 18241 21465 18244
rect 21499 18241 21511 18275
rect 21453 18235 21511 18241
rect 21545 18275 21603 18281
rect 21545 18241 21557 18275
rect 21591 18272 21603 18275
rect 22005 18275 22063 18281
rect 22005 18272 22017 18275
rect 21591 18244 22017 18272
rect 21591 18241 21603 18244
rect 21545 18235 21603 18241
rect 22005 18241 22017 18244
rect 22051 18272 22063 18275
rect 22278 18272 22284 18284
rect 22051 18244 22284 18272
rect 22051 18241 22063 18244
rect 22005 18235 22063 18241
rect 22278 18232 22284 18244
rect 22336 18232 22342 18284
rect 22388 18281 22416 18380
rect 22554 18368 22560 18420
rect 22612 18368 22618 18420
rect 22572 18340 22600 18368
rect 22480 18312 22600 18340
rect 22373 18275 22431 18281
rect 22373 18241 22385 18275
rect 22419 18241 22431 18275
rect 22373 18235 22431 18241
rect 19705 18207 19763 18213
rect 18196 18176 18552 18204
rect 18616 18176 18828 18204
rect 18196 18164 18202 18176
rect 13998 18136 14004 18148
rect 11716 18108 12204 18136
rect 3973 18071 4031 18077
rect 3973 18037 3985 18071
rect 4019 18068 4031 18071
rect 4430 18068 4436 18080
rect 4019 18040 4436 18068
rect 4019 18037 4031 18040
rect 3973 18031 4031 18037
rect 4430 18028 4436 18040
rect 4488 18028 4494 18080
rect 5810 18028 5816 18080
rect 5868 18068 5874 18080
rect 6730 18068 6736 18080
rect 5868 18040 6736 18068
rect 5868 18028 5874 18040
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 6822 18028 6828 18080
rect 6880 18068 6886 18080
rect 7650 18068 7656 18080
rect 6880 18040 6925 18068
rect 7611 18040 7656 18068
rect 6880 18028 6886 18040
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 9033 18071 9091 18077
rect 9033 18037 9045 18071
rect 9079 18068 9091 18071
rect 9306 18068 9312 18080
rect 9079 18040 9312 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 9306 18028 9312 18040
rect 9364 18068 9370 18080
rect 9769 18071 9827 18077
rect 9769 18068 9781 18071
rect 9364 18040 9781 18068
rect 9364 18028 9370 18040
rect 9769 18037 9781 18040
rect 9815 18037 9827 18071
rect 9769 18031 9827 18037
rect 10318 18028 10324 18080
rect 10376 18068 10382 18080
rect 10413 18071 10471 18077
rect 10413 18068 10425 18071
rect 10376 18040 10425 18068
rect 10376 18028 10382 18040
rect 10413 18037 10425 18040
rect 10459 18068 10471 18071
rect 11698 18068 11704 18080
rect 10459 18040 11704 18068
rect 10459 18037 10471 18040
rect 10413 18031 10471 18037
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 12176 18068 12204 18108
rect 13464 18108 14004 18136
rect 13464 18068 13492 18108
rect 13998 18096 14004 18108
rect 14056 18096 14062 18148
rect 18230 18136 18236 18148
rect 18191 18108 18236 18136
rect 18230 18096 18236 18108
rect 18288 18096 18294 18148
rect 18524 18145 18552 18176
rect 18800 18148 18828 18176
rect 19705 18173 19717 18207
rect 19751 18204 19763 18207
rect 20441 18207 20499 18213
rect 20441 18204 20453 18207
rect 19751 18176 20453 18204
rect 19751 18173 19763 18176
rect 19705 18167 19763 18173
rect 20441 18173 20453 18176
rect 20487 18204 20499 18207
rect 20898 18204 20904 18216
rect 20487 18176 20904 18204
rect 20487 18173 20499 18176
rect 20441 18167 20499 18173
rect 20898 18164 20904 18176
rect 20956 18164 20962 18216
rect 20990 18164 20996 18216
rect 21048 18204 21054 18216
rect 22480 18204 22508 18312
rect 22738 18300 22744 18352
rect 22796 18300 22802 18352
rect 23109 18343 23167 18349
rect 23109 18309 23121 18343
rect 23155 18340 23167 18343
rect 23382 18340 23388 18352
rect 23155 18312 23388 18340
rect 23155 18309 23167 18312
rect 23109 18303 23167 18309
rect 23382 18300 23388 18312
rect 23440 18300 23446 18352
rect 22556 18275 22614 18281
rect 22556 18241 22568 18275
rect 22602 18241 22614 18275
rect 22556 18235 22614 18241
rect 22649 18275 22707 18281
rect 22649 18241 22661 18275
rect 22695 18272 22707 18275
rect 22756 18272 22784 18300
rect 22695 18244 22784 18272
rect 22695 18241 22707 18244
rect 22649 18235 22707 18241
rect 21048 18176 22508 18204
rect 21048 18164 21054 18176
rect 18509 18139 18567 18145
rect 18509 18105 18521 18139
rect 18555 18105 18567 18139
rect 18509 18099 18567 18105
rect 18598 18096 18604 18148
rect 18656 18136 18662 18148
rect 18656 18108 18701 18136
rect 18656 18096 18662 18108
rect 18782 18096 18788 18148
rect 18840 18136 18846 18148
rect 21726 18136 21732 18148
rect 18840 18108 21732 18136
rect 18840 18096 18846 18108
rect 21726 18096 21732 18108
rect 21784 18136 21790 18148
rect 21821 18139 21879 18145
rect 21821 18136 21833 18139
rect 21784 18108 21833 18136
rect 21784 18096 21790 18108
rect 21821 18105 21833 18108
rect 21867 18105 21879 18139
rect 21821 18099 21879 18105
rect 22186 18096 22192 18148
rect 22244 18136 22250 18148
rect 22571 18136 22599 18235
rect 22830 18232 22836 18284
rect 22888 18275 22894 18284
rect 22925 18275 22983 18281
rect 22888 18247 22937 18275
rect 22888 18232 22894 18247
rect 22925 18241 22937 18247
rect 22971 18241 22983 18275
rect 22925 18235 22983 18241
rect 22738 18204 22744 18216
rect 22699 18176 22744 18204
rect 22738 18164 22744 18176
rect 22796 18164 22802 18216
rect 22830 18136 22836 18148
rect 22244 18108 22599 18136
rect 22628 18108 22836 18136
rect 22244 18096 22250 18108
rect 12176 18040 13492 18068
rect 15102 18028 15108 18080
rect 15160 18068 15166 18080
rect 22628 18068 22656 18108
rect 22830 18096 22836 18108
rect 22888 18136 22894 18148
rect 23201 18139 23259 18145
rect 23201 18136 23213 18139
rect 22888 18108 23213 18136
rect 22888 18096 22894 18108
rect 23201 18105 23213 18108
rect 23247 18105 23259 18139
rect 23201 18099 23259 18105
rect 15160 18040 22656 18068
rect 15160 18028 15166 18040
rect 1104 17978 26220 18000
rect 1104 17926 5136 17978
rect 5188 17926 5200 17978
rect 5252 17926 5264 17978
rect 5316 17926 5328 17978
rect 5380 17926 5392 17978
rect 5444 17926 13508 17978
rect 13560 17926 13572 17978
rect 13624 17926 13636 17978
rect 13688 17926 13700 17978
rect 13752 17926 13764 17978
rect 13816 17926 21880 17978
rect 21932 17926 21944 17978
rect 21996 17926 22008 17978
rect 22060 17926 22072 17978
rect 22124 17926 22136 17978
rect 22188 17926 26220 17978
rect 1104 17904 26220 17926
rect 4522 17824 4528 17876
rect 4580 17864 4586 17876
rect 4617 17867 4675 17873
rect 4617 17864 4629 17867
rect 4580 17836 4629 17864
rect 4580 17824 4586 17836
rect 4617 17833 4629 17836
rect 4663 17864 4675 17867
rect 4801 17867 4859 17873
rect 4801 17864 4813 17867
rect 4663 17836 4813 17864
rect 4663 17833 4675 17836
rect 4617 17827 4675 17833
rect 4801 17833 4813 17836
rect 4847 17833 4859 17867
rect 4801 17827 4859 17833
rect 6181 17867 6239 17873
rect 6181 17833 6193 17867
rect 6227 17864 6239 17867
rect 8386 17864 8392 17876
rect 6227 17836 8392 17864
rect 6227 17833 6239 17836
rect 6181 17827 6239 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 9950 17864 9956 17876
rect 9911 17836 9956 17864
rect 9950 17824 9956 17836
rect 10008 17864 10014 17876
rect 10321 17867 10379 17873
rect 10321 17864 10333 17867
rect 10008 17836 10333 17864
rect 10008 17824 10014 17836
rect 10321 17833 10333 17836
rect 10367 17833 10379 17867
rect 11790 17864 11796 17876
rect 10321 17827 10379 17833
rect 11624 17836 11796 17864
rect 3789 17799 3847 17805
rect 3789 17796 3801 17799
rect 3068 17768 3801 17796
rect 3068 17669 3096 17768
rect 3789 17765 3801 17768
rect 3835 17765 3847 17799
rect 3789 17759 3847 17765
rect 3326 17728 3332 17740
rect 3287 17700 3332 17728
rect 3326 17688 3332 17700
rect 3384 17688 3390 17740
rect 4338 17688 4344 17740
rect 4396 17728 4402 17740
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 4396 17700 4445 17728
rect 4396 17688 4402 17700
rect 4433 17697 4445 17700
rect 4479 17728 4491 17731
rect 4540 17728 4568 17824
rect 9398 17756 9404 17808
rect 9456 17796 9462 17808
rect 11624 17796 11652 17836
rect 11790 17824 11796 17836
rect 11848 17824 11854 17876
rect 12250 17824 12256 17876
rect 12308 17864 12314 17876
rect 12710 17864 12716 17876
rect 12308 17836 12716 17864
rect 12308 17824 12314 17836
rect 12710 17824 12716 17836
rect 12768 17824 12774 17876
rect 15473 17867 15531 17873
rect 15473 17864 15485 17867
rect 13924 17836 15485 17864
rect 9456 17768 11652 17796
rect 9456 17756 9462 17768
rect 4479 17700 4568 17728
rect 8205 17731 8263 17737
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 8205 17697 8217 17731
rect 8251 17728 8263 17731
rect 8294 17728 8300 17740
rect 8251 17700 8300 17728
rect 8251 17697 8263 17700
rect 8205 17691 8263 17697
rect 8294 17688 8300 17700
rect 8352 17728 8358 17740
rect 9416 17728 9444 17756
rect 11624 17737 11652 17768
rect 12989 17799 13047 17805
rect 12989 17765 13001 17799
rect 13035 17796 13047 17799
rect 13035 17768 13584 17796
rect 13035 17765 13047 17768
rect 12989 17759 13047 17765
rect 13556 17737 13584 17768
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 8352 17700 9444 17728
rect 9600 17700 9873 17728
rect 8352 17688 8358 17700
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17629 3111 17663
rect 3053 17623 3111 17629
rect 3142 17620 3148 17672
rect 3200 17660 3206 17672
rect 3421 17663 3479 17669
rect 3200 17632 3245 17660
rect 3200 17620 3206 17632
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 4154 17660 4160 17672
rect 3467 17632 4160 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 4154 17620 4160 17632
rect 4212 17620 4218 17672
rect 6362 17620 6368 17672
rect 6420 17660 6426 17672
rect 8754 17660 8760 17672
rect 6420 17632 8760 17660
rect 6420 17620 6426 17632
rect 8754 17620 8760 17632
rect 8812 17620 8818 17672
rect 9306 17660 9312 17672
rect 9267 17632 9312 17660
rect 9306 17620 9312 17632
rect 9364 17660 9370 17672
rect 9600 17660 9628 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 11609 17731 11667 17737
rect 11609 17697 11621 17731
rect 11655 17697 11667 17731
rect 11609 17691 11667 17697
rect 13541 17731 13599 17737
rect 13541 17697 13553 17731
rect 13587 17697 13599 17731
rect 13924 17728 13952 17836
rect 15473 17833 15485 17836
rect 15519 17864 15531 17867
rect 17586 17864 17592 17876
rect 15519 17836 17592 17864
rect 15519 17833 15531 17836
rect 15473 17827 15531 17833
rect 17586 17824 17592 17836
rect 17644 17824 17650 17876
rect 17862 17824 17868 17876
rect 17920 17864 17926 17876
rect 18138 17864 18144 17876
rect 17920 17836 18144 17864
rect 17920 17824 17926 17836
rect 18138 17824 18144 17836
rect 18196 17824 18202 17876
rect 18414 17824 18420 17876
rect 18472 17864 18478 17876
rect 19242 17864 19248 17876
rect 18472 17836 19248 17864
rect 18472 17824 18478 17836
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 20162 17864 20168 17876
rect 20123 17836 20168 17864
rect 20162 17824 20168 17836
rect 20220 17824 20226 17876
rect 20254 17824 20260 17876
rect 20312 17864 20318 17876
rect 22005 17867 22063 17873
rect 20312 17836 21404 17864
rect 20312 17824 20318 17836
rect 15378 17756 15384 17808
rect 15436 17796 15442 17808
rect 17402 17796 17408 17808
rect 15436 17768 17408 17796
rect 15436 17756 15442 17768
rect 17402 17756 17408 17768
rect 17460 17796 17466 17808
rect 17681 17799 17739 17805
rect 17681 17796 17693 17799
rect 17460 17768 17693 17796
rect 17460 17756 17466 17768
rect 17681 17765 17693 17768
rect 17727 17765 17739 17799
rect 17681 17759 17739 17765
rect 21269 17799 21327 17805
rect 21269 17765 21281 17799
rect 21315 17765 21327 17799
rect 21376 17796 21404 17836
rect 22005 17833 22017 17867
rect 22051 17864 22063 17867
rect 22370 17864 22376 17876
rect 22051 17836 22376 17864
rect 22051 17833 22063 17836
rect 22005 17827 22063 17833
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 23014 17796 23020 17808
rect 21376 17768 22508 17796
rect 21269 17759 21327 17765
rect 14090 17728 14096 17740
rect 13541 17691 13599 17697
rect 13648 17700 13952 17728
rect 14051 17700 14096 17728
rect 9364 17632 9628 17660
rect 9769 17663 9827 17669
rect 9364 17620 9370 17632
rect 9769 17629 9781 17663
rect 9815 17629 9827 17663
rect 10594 17660 10600 17672
rect 10555 17632 10600 17660
rect 9769 17623 9827 17629
rect 4249 17595 4307 17601
rect 4249 17561 4261 17595
rect 4295 17592 4307 17595
rect 7926 17592 7932 17604
rect 7984 17601 7990 17604
rect 4295 17564 6868 17592
rect 7896 17564 7932 17592
rect 4295 17561 4307 17564
rect 4249 17555 4307 17561
rect 2866 17524 2872 17536
rect 2827 17496 2872 17524
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 2958 17484 2964 17536
rect 3016 17524 3022 17536
rect 4157 17527 4215 17533
rect 4157 17524 4169 17527
rect 3016 17496 4169 17524
rect 3016 17484 3022 17496
rect 4157 17493 4169 17496
rect 4203 17493 4215 17527
rect 4157 17487 4215 17493
rect 6086 17484 6092 17536
rect 6144 17524 6150 17536
rect 6840 17533 6868 17564
rect 7926 17552 7932 17564
rect 7984 17555 7996 17601
rect 7984 17552 7990 17555
rect 9030 17552 9036 17604
rect 9088 17592 9094 17604
rect 9125 17595 9183 17601
rect 9125 17592 9137 17595
rect 9088 17564 9137 17592
rect 9088 17552 9094 17564
rect 9125 17561 9137 17564
rect 9171 17561 9183 17595
rect 9125 17555 9183 17561
rect 9493 17595 9551 17601
rect 9493 17561 9505 17595
rect 9539 17592 9551 17595
rect 9674 17592 9680 17604
rect 9539 17564 9680 17592
rect 9539 17561 9551 17564
rect 9493 17555 9551 17561
rect 6181 17527 6239 17533
rect 6181 17524 6193 17527
rect 6144 17496 6193 17524
rect 6144 17484 6150 17496
rect 6181 17493 6193 17496
rect 6227 17524 6239 17527
rect 6273 17527 6331 17533
rect 6273 17524 6285 17527
rect 6227 17496 6285 17524
rect 6227 17493 6239 17496
rect 6181 17487 6239 17493
rect 6273 17493 6285 17496
rect 6319 17493 6331 17527
rect 6273 17487 6331 17493
rect 6825 17527 6883 17533
rect 6825 17493 6837 17527
rect 6871 17524 6883 17527
rect 8110 17524 8116 17536
rect 6871 17496 8116 17524
rect 6871 17493 6883 17496
rect 6825 17487 6883 17493
rect 8110 17484 8116 17496
rect 8168 17484 8174 17536
rect 8938 17484 8944 17536
rect 8996 17524 9002 17536
rect 9508 17524 9536 17555
rect 9674 17552 9680 17564
rect 9732 17592 9738 17604
rect 9784 17592 9812 17623
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 12250 17660 12256 17672
rect 11164 17632 12256 17660
rect 11164 17592 11192 17632
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 13078 17620 13084 17672
rect 13136 17660 13142 17672
rect 13173 17663 13231 17669
rect 13173 17660 13185 17663
rect 13136 17632 13185 17660
rect 13136 17620 13142 17632
rect 13173 17629 13185 17632
rect 13219 17629 13231 17663
rect 13173 17623 13231 17629
rect 13321 17660 13379 17666
rect 13321 17626 13333 17660
rect 13367 17626 13379 17660
rect 13321 17620 13379 17626
rect 13449 17663 13507 17669
rect 13449 17629 13461 17663
rect 13495 17660 13507 17663
rect 13648 17660 13676 17700
rect 14090 17688 14096 17700
rect 14148 17688 14154 17740
rect 20073 17731 20131 17737
rect 20073 17697 20085 17731
rect 20119 17728 20131 17731
rect 20717 17731 20775 17737
rect 20717 17728 20729 17731
rect 20119 17700 20729 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 20717 17697 20729 17700
rect 20763 17728 20775 17731
rect 20898 17728 20904 17740
rect 20763 17700 20904 17728
rect 20763 17697 20775 17700
rect 20717 17691 20775 17697
rect 20898 17688 20904 17700
rect 20956 17688 20962 17740
rect 21284 17728 21312 17759
rect 21634 17728 21640 17740
rect 21284 17700 21640 17728
rect 21634 17688 21640 17700
rect 21692 17688 21698 17740
rect 21729 17731 21787 17737
rect 21729 17697 21741 17731
rect 21775 17728 21787 17731
rect 22370 17728 22376 17740
rect 21775 17700 22376 17728
rect 21775 17697 21787 17700
rect 21729 17691 21787 17697
rect 22370 17688 22376 17700
rect 22428 17688 22434 17740
rect 13495 17632 13676 17660
rect 13495 17629 13507 17632
rect 13449 17623 13507 17629
rect 13722 17620 13728 17672
rect 13780 17660 13786 17672
rect 14108 17660 14136 17688
rect 16666 17660 16672 17672
rect 13780 17632 13825 17660
rect 14108 17632 16672 17660
rect 13780 17620 13786 17632
rect 16666 17620 16672 17632
rect 16724 17660 16730 17672
rect 17037 17663 17095 17669
rect 17037 17660 17049 17663
rect 16724 17632 17049 17660
rect 16724 17620 16730 17632
rect 17037 17629 17049 17632
rect 17083 17629 17095 17663
rect 17037 17623 17095 17629
rect 17221 17663 17279 17669
rect 17221 17629 17233 17663
rect 17267 17660 17279 17663
rect 18414 17660 18420 17672
rect 17267 17632 18420 17660
rect 17267 17629 17279 17632
rect 17221 17623 17279 17629
rect 9732 17564 9812 17592
rect 10152 17564 11192 17592
rect 9732 17552 9738 17564
rect 8996 17496 9536 17524
rect 9585 17527 9643 17533
rect 8996 17484 9002 17496
rect 9585 17493 9597 17527
rect 9631 17524 9643 17527
rect 9950 17524 9956 17536
rect 9631 17496 9956 17524
rect 9631 17493 9643 17496
rect 9585 17487 9643 17493
rect 9950 17484 9956 17496
rect 10008 17484 10014 17536
rect 10152 17533 10180 17564
rect 11238 17552 11244 17604
rect 11296 17592 11302 17604
rect 11854 17595 11912 17601
rect 11854 17592 11866 17595
rect 11296 17564 11866 17592
rect 11296 17552 11302 17564
rect 11854 17561 11866 17564
rect 11900 17561 11912 17595
rect 11854 17555 11912 17561
rect 12158 17552 12164 17604
rect 12216 17592 12222 17604
rect 13336 17592 13364 17620
rect 13538 17592 13544 17604
rect 12216 17564 13544 17592
rect 12216 17552 12222 17564
rect 13538 17552 13544 17564
rect 13596 17552 13602 17604
rect 13909 17595 13967 17601
rect 13909 17561 13921 17595
rect 13955 17592 13967 17595
rect 14338 17595 14396 17601
rect 14338 17592 14350 17595
rect 13955 17564 14350 17592
rect 13955 17561 13967 17564
rect 13909 17555 13967 17561
rect 14338 17561 14350 17564
rect 14384 17561 14396 17595
rect 17052 17592 17080 17623
rect 18414 17620 18420 17632
rect 18472 17620 18478 17672
rect 19058 17660 19064 17672
rect 18524 17632 19064 17660
rect 18524 17592 18552 17632
rect 19058 17620 19064 17632
rect 19116 17620 19122 17672
rect 21082 17660 21088 17672
rect 19168 17632 21088 17660
rect 17052 17564 18552 17592
rect 14338 17555 14396 17561
rect 18598 17552 18604 17604
rect 18656 17592 18662 17604
rect 18794 17595 18852 17601
rect 18794 17592 18806 17595
rect 18656 17564 18806 17592
rect 18656 17552 18662 17564
rect 18794 17561 18806 17564
rect 18840 17561 18852 17595
rect 18794 17555 18852 17561
rect 10137 17527 10195 17533
rect 10137 17493 10149 17527
rect 10183 17493 10195 17527
rect 10137 17487 10195 17493
rect 10781 17527 10839 17533
rect 10781 17493 10793 17527
rect 10827 17524 10839 17527
rect 11054 17524 11060 17536
rect 10827 17496 11060 17524
rect 10827 17493 10839 17496
rect 10781 17487 10839 17493
rect 11054 17484 11060 17496
rect 11112 17524 11118 17536
rect 12250 17524 12256 17536
rect 11112 17496 12256 17524
rect 11112 17484 11118 17496
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 19168 17524 19196 17632
rect 21082 17620 21088 17632
rect 21140 17620 21146 17672
rect 21358 17660 21364 17672
rect 21319 17632 21364 17660
rect 21358 17620 21364 17632
rect 21416 17620 21422 17672
rect 21509 17657 21567 17663
rect 21910 17660 21916 17672
rect 21509 17634 21521 17657
rect 21468 17623 21521 17634
rect 21555 17623 21567 17657
rect 21871 17632 21916 17660
rect 21468 17617 21567 17623
rect 21910 17620 21916 17632
rect 21968 17620 21974 17672
rect 22189 17663 22247 17669
rect 22189 17629 22201 17663
rect 22235 17660 22247 17663
rect 22278 17660 22284 17672
rect 22235 17632 22284 17660
rect 22235 17629 22247 17632
rect 22189 17623 22247 17629
rect 22278 17620 22284 17632
rect 22336 17620 22342 17672
rect 22480 17669 22508 17768
rect 22756 17768 23020 17796
rect 22756 17672 22784 17768
rect 23014 17756 23020 17768
rect 23072 17756 23078 17808
rect 24210 17688 24216 17740
rect 24268 17728 24274 17740
rect 24397 17731 24455 17737
rect 24397 17728 24409 17731
rect 24268 17700 24409 17728
rect 24268 17688 24274 17700
rect 24397 17697 24409 17700
rect 24443 17697 24455 17731
rect 24397 17691 24455 17697
rect 22465 17663 22523 17669
rect 22465 17629 22477 17663
rect 22511 17629 22523 17663
rect 22465 17623 22523 17629
rect 22613 17660 22671 17666
rect 22738 17660 22744 17672
rect 22613 17626 22625 17660
rect 22659 17626 22671 17660
rect 22699 17632 22744 17660
rect 22613 17620 22671 17626
rect 22738 17620 22744 17632
rect 22796 17620 22802 17672
rect 22830 17620 22836 17672
rect 22888 17660 22894 17672
rect 23017 17663 23075 17669
rect 22888 17632 22933 17660
rect 22888 17620 22894 17632
rect 23017 17629 23029 17663
rect 23063 17629 23075 17663
rect 23017 17623 23075 17629
rect 21468 17606 21552 17617
rect 20714 17552 20720 17604
rect 20772 17592 20778 17604
rect 21468 17592 21496 17606
rect 22628 17592 22656 17620
rect 20772 17564 21496 17592
rect 22296 17564 22656 17592
rect 20772 17552 20778 17564
rect 22296 17536 22324 17564
rect 20530 17524 20536 17536
rect 12768 17496 19196 17524
rect 20491 17496 20536 17524
rect 12768 17484 12774 17496
rect 20530 17484 20536 17496
rect 20588 17484 20594 17536
rect 20622 17484 20628 17536
rect 20680 17524 20686 17536
rect 20680 17496 20725 17524
rect 20680 17484 20686 17496
rect 21174 17484 21180 17536
rect 21232 17524 21238 17536
rect 21910 17524 21916 17536
rect 21232 17496 21916 17524
rect 21232 17484 21238 17496
rect 21910 17484 21916 17496
rect 21968 17484 21974 17536
rect 22278 17484 22284 17536
rect 22336 17484 22342 17536
rect 22370 17484 22376 17536
rect 22428 17524 22434 17536
rect 22830 17524 22836 17536
rect 22428 17496 22836 17524
rect 22428 17484 22434 17496
rect 22830 17484 22836 17496
rect 22888 17484 22894 17536
rect 23032 17524 23060 17623
rect 23201 17595 23259 17601
rect 23201 17561 23213 17595
rect 23247 17592 23259 17595
rect 24642 17595 24700 17601
rect 24642 17592 24654 17595
rect 23247 17564 24654 17592
rect 23247 17561 23259 17564
rect 23201 17555 23259 17561
rect 24642 17561 24654 17564
rect 24688 17561 24700 17595
rect 24642 17555 24700 17561
rect 25774 17524 25780 17536
rect 23032 17496 25780 17524
rect 25774 17484 25780 17496
rect 25832 17484 25838 17536
rect 1104 17434 26220 17456
rect 1104 17382 9322 17434
rect 9374 17382 9386 17434
rect 9438 17382 9450 17434
rect 9502 17382 9514 17434
rect 9566 17382 9578 17434
rect 9630 17382 17694 17434
rect 17746 17382 17758 17434
rect 17810 17382 17822 17434
rect 17874 17382 17886 17434
rect 17938 17382 17950 17434
rect 18002 17382 26220 17434
rect 1104 17360 26220 17382
rect 3694 17280 3700 17332
rect 3752 17320 3758 17332
rect 3789 17323 3847 17329
rect 3789 17320 3801 17323
rect 3752 17292 3801 17320
rect 3752 17280 3758 17292
rect 3789 17289 3801 17292
rect 3835 17289 3847 17323
rect 5537 17323 5595 17329
rect 3789 17283 3847 17289
rect 4172 17292 4936 17320
rect 2124 17255 2182 17261
rect 2124 17221 2136 17255
rect 2170 17252 2182 17255
rect 2866 17252 2872 17264
rect 2170 17224 2872 17252
rect 2170 17221 2182 17224
rect 2124 17215 2182 17221
rect 2866 17212 2872 17224
rect 2924 17212 2930 17264
rect 3142 17212 3148 17264
rect 3200 17252 3206 17264
rect 4172 17252 4200 17292
rect 3200 17224 4200 17252
rect 4249 17255 4307 17261
rect 3200 17212 3206 17224
rect 4249 17221 4261 17255
rect 4295 17252 4307 17255
rect 4295 17224 4844 17252
rect 4295 17221 4307 17224
rect 4249 17215 4307 17221
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 1946 17184 1952 17196
rect 1903 17156 1952 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 4157 17187 4215 17193
rect 4157 17184 4169 17187
rect 3568 17156 4169 17184
rect 3568 17144 3574 17156
rect 4157 17153 4169 17156
rect 4203 17184 4215 17187
rect 4617 17187 4675 17193
rect 4617 17184 4629 17187
rect 4203 17156 4629 17184
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 4617 17153 4629 17156
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 4338 17116 4344 17128
rect 4299 17088 4344 17116
rect 4338 17076 4344 17088
rect 4396 17076 4402 17128
rect 4430 17076 4436 17128
rect 4488 17116 4494 17128
rect 4709 17119 4767 17125
rect 4709 17116 4721 17119
rect 4488 17088 4721 17116
rect 4488 17076 4494 17088
rect 4709 17085 4721 17088
rect 4755 17085 4767 17119
rect 4816 17116 4844 17224
rect 4908 17193 4936 17292
rect 5537 17289 5549 17323
rect 5583 17320 5595 17323
rect 6178 17320 6184 17332
rect 5583 17292 6184 17320
rect 5583 17289 5595 17292
rect 5537 17283 5595 17289
rect 6178 17280 6184 17292
rect 6236 17280 6242 17332
rect 8294 17320 8300 17332
rect 8036 17292 8300 17320
rect 7570 17255 7628 17261
rect 7570 17252 7582 17255
rect 6380 17224 7582 17252
rect 6380 17196 6408 17224
rect 7570 17221 7582 17224
rect 7616 17221 7628 17255
rect 7926 17252 7932 17264
rect 7887 17224 7932 17252
rect 7570 17215 7628 17221
rect 7926 17212 7932 17224
rect 7984 17212 7990 17264
rect 4893 17187 4951 17193
rect 4893 17153 4905 17187
rect 4939 17153 4951 17187
rect 4893 17147 4951 17153
rect 4982 17144 4988 17196
rect 5040 17184 5046 17196
rect 5629 17187 5687 17193
rect 5040 17156 5085 17184
rect 5040 17144 5046 17156
rect 5629 17153 5641 17187
rect 5675 17153 5687 17187
rect 5810 17184 5816 17196
rect 5771 17156 5816 17184
rect 5629 17147 5687 17153
rect 5644 17116 5672 17147
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 5998 17187 6056 17193
rect 5998 17153 6010 17187
rect 6044 17184 6056 17187
rect 6086 17184 6092 17196
rect 6044 17156 6092 17184
rect 6044 17153 6056 17156
rect 5998 17147 6056 17153
rect 6086 17144 6092 17156
rect 6144 17144 6150 17196
rect 6178 17144 6184 17196
rect 6236 17184 6242 17196
rect 6236 17156 6281 17184
rect 6236 17144 6242 17156
rect 6362 17144 6368 17196
rect 6420 17144 6426 17196
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 7837 17187 7895 17193
rect 6788 17156 7788 17184
rect 6788 17144 6794 17156
rect 4816 17088 5672 17116
rect 4709 17079 4767 17085
rect 4062 17008 4068 17060
rect 4120 17048 4126 17060
rect 5644 17048 5672 17088
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 6822 17116 6828 17128
rect 5951 17088 6828 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 7760 17116 7788 17156
rect 7837 17153 7849 17187
rect 7883 17184 7895 17187
rect 8036 17184 8064 17292
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 9122 17320 9128 17332
rect 8588 17292 9128 17320
rect 7883 17156 8064 17184
rect 7883 17153 7895 17156
rect 7837 17147 7895 17153
rect 8110 17144 8116 17196
rect 8168 17184 8174 17196
rect 8499 17187 8557 17193
rect 8168 17156 8213 17184
rect 8168 17144 8174 17156
rect 8499 17153 8511 17187
rect 8545 17184 8557 17187
rect 8588 17184 8616 17292
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 11238 17320 11244 17332
rect 9324 17292 10088 17320
rect 11199 17292 11244 17320
rect 8545 17156 8616 17184
rect 8545 17153 8557 17156
rect 8499 17147 8557 17153
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 8849 17187 8907 17193
rect 8849 17184 8861 17187
rect 8720 17156 8861 17184
rect 8720 17144 8726 17156
rect 8849 17153 8861 17156
rect 8895 17153 8907 17187
rect 9014 17187 9072 17193
rect 9014 17184 9026 17187
rect 8849 17147 8907 17153
rect 8956 17156 9026 17184
rect 8297 17119 8355 17125
rect 8297 17116 8309 17119
rect 7760 17088 8309 17116
rect 8297 17085 8309 17088
rect 8343 17085 8355 17119
rect 8297 17079 8355 17085
rect 8389 17119 8447 17125
rect 8389 17085 8401 17119
rect 8435 17085 8447 17119
rect 8389 17079 8447 17085
rect 6457 17051 6515 17057
rect 6457 17048 6469 17051
rect 4120 17020 5304 17048
rect 5644 17020 6469 17048
rect 4120 17008 4126 17020
rect 3237 16983 3295 16989
rect 3237 16949 3249 16983
rect 3283 16980 3295 16983
rect 4154 16980 4160 16992
rect 3283 16952 4160 16980
rect 3283 16949 3295 16952
rect 3237 16943 3295 16949
rect 4154 16940 4160 16952
rect 4212 16940 4218 16992
rect 4798 16940 4804 16992
rect 4856 16980 4862 16992
rect 5169 16983 5227 16989
rect 5169 16980 5181 16983
rect 4856 16952 5181 16980
rect 4856 16940 4862 16952
rect 5169 16949 5181 16952
rect 5215 16949 5227 16983
rect 5276 16980 5304 17020
rect 6457 17017 6469 17020
rect 6503 17017 6515 17051
rect 6457 17011 6515 17017
rect 7926 17008 7932 17060
rect 7984 17048 7990 17060
rect 8404 17048 8432 17079
rect 8754 17076 8760 17128
rect 8812 17116 8818 17128
rect 8956 17116 8984 17156
rect 9014 17153 9026 17156
rect 9060 17153 9072 17187
rect 9014 17147 9072 17153
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17184 9275 17187
rect 9324 17184 9352 17292
rect 9490 17212 9496 17264
rect 9548 17252 9554 17264
rect 9548 17224 9720 17252
rect 9548 17212 9554 17224
rect 9263 17156 9352 17184
rect 9263 17153 9275 17156
rect 9217 17147 9275 17153
rect 9398 17144 9404 17196
rect 9456 17184 9462 17196
rect 9692 17193 9720 17224
rect 9950 17212 9956 17264
rect 10008 17212 10014 17264
rect 9677 17187 9735 17193
rect 9456 17156 9501 17184
rect 9456 17144 9462 17156
rect 9677 17153 9689 17187
rect 9723 17153 9735 17187
rect 9677 17147 9735 17153
rect 9860 17187 9918 17193
rect 9860 17153 9872 17187
rect 9906 17184 9918 17187
rect 9968 17184 9996 17212
rect 9906 17156 9996 17184
rect 9906 17153 9918 17156
rect 9860 17147 9918 17153
rect 9122 17116 9128 17128
rect 8812 17088 8984 17116
rect 9083 17088 9128 17116
rect 8812 17076 8818 17088
rect 9122 17076 9128 17088
rect 9180 17076 9186 17128
rect 10060 17125 10088 17292
rect 11238 17280 11244 17292
rect 11296 17280 11302 17332
rect 15562 17320 15568 17332
rect 13740 17292 15568 17320
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17184 10287 17187
rect 10502 17184 10508 17196
rect 10275 17156 10508 17184
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 11054 17184 11060 17196
rect 11015 17156 11060 17184
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 13078 17144 13084 17196
rect 13136 17184 13142 17196
rect 13449 17187 13507 17193
rect 13449 17184 13461 17187
rect 13136 17156 13461 17184
rect 13136 17144 13142 17156
rect 13449 17153 13461 17156
rect 13495 17153 13507 17187
rect 13449 17147 13507 17153
rect 9953 17119 10011 17125
rect 9953 17116 9965 17119
rect 9508 17088 9965 17116
rect 7984 17020 8432 17048
rect 9140 17048 9168 17076
rect 9508 17048 9536 17088
rect 9953 17085 9965 17088
rect 9999 17085 10011 17119
rect 9953 17079 10011 17085
rect 10045 17119 10103 17125
rect 10045 17085 10057 17119
rect 10091 17116 10103 17119
rect 10134 17116 10140 17128
rect 10091 17088 10140 17116
rect 10091 17085 10103 17088
rect 10045 17079 10103 17085
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 12710 17076 12716 17128
rect 12768 17116 12774 17128
rect 13262 17116 13268 17128
rect 12768 17088 13268 17116
rect 12768 17076 12774 17088
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 13464 17116 13492 17147
rect 13538 17144 13544 17196
rect 13596 17190 13655 17196
rect 13740 17193 13768 17292
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 17218 17280 17224 17332
rect 17276 17320 17282 17332
rect 17313 17323 17371 17329
rect 17313 17320 17325 17323
rect 17276 17292 17325 17320
rect 17276 17280 17282 17292
rect 17313 17289 17325 17292
rect 17359 17320 17371 17323
rect 17586 17320 17592 17332
rect 17359 17292 17592 17320
rect 17359 17289 17371 17292
rect 17313 17283 17371 17289
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 18325 17323 18383 17329
rect 17695 17292 17816 17320
rect 14185 17255 14243 17261
rect 14185 17221 14197 17255
rect 14231 17252 14243 17255
rect 14274 17252 14280 17264
rect 14231 17224 14280 17252
rect 14231 17221 14243 17224
rect 14185 17215 14243 17221
rect 14274 17212 14280 17224
rect 14332 17212 14338 17264
rect 16942 17212 16948 17264
rect 17000 17252 17006 17264
rect 17497 17255 17555 17261
rect 17497 17252 17509 17255
rect 17000 17224 17509 17252
rect 17000 17212 17006 17224
rect 17497 17221 17509 17224
rect 17543 17221 17555 17255
rect 17497 17215 17555 17221
rect 17695 17219 17723 17292
rect 17788 17252 17816 17292
rect 18325 17289 18337 17323
rect 18371 17320 18383 17323
rect 18598 17320 18604 17332
rect 18371 17292 18604 17320
rect 18371 17289 18383 17292
rect 18325 17283 18383 17289
rect 18598 17280 18604 17292
rect 18656 17280 18662 17332
rect 20533 17323 20591 17329
rect 20533 17289 20545 17323
rect 20579 17320 20591 17323
rect 20714 17320 20720 17332
rect 20579 17292 20720 17320
rect 20579 17289 20591 17292
rect 20533 17283 20591 17289
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 21174 17320 21180 17332
rect 21135 17292 21180 17320
rect 21174 17280 21180 17292
rect 21232 17280 21238 17332
rect 21266 17280 21272 17332
rect 21324 17320 21330 17332
rect 21821 17323 21879 17329
rect 21821 17320 21833 17323
rect 21324 17292 21833 17320
rect 21324 17280 21330 17292
rect 21821 17289 21833 17292
rect 21867 17289 21879 17323
rect 22646 17320 22652 17332
rect 22607 17292 22652 17320
rect 21821 17283 21879 17289
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 20990 17252 20996 17264
rect 17788 17224 18368 17252
rect 17681 17213 17739 17219
rect 13596 17156 13609 17190
rect 13643 17156 13655 17190
rect 13596 17150 13655 17156
rect 13725 17187 13783 17193
rect 13725 17153 13737 17187
rect 13771 17153 13783 17187
rect 13596 17144 13602 17150
rect 13725 17147 13783 17153
rect 13906 17144 13912 17196
rect 13964 17184 13970 17196
rect 14001 17187 14059 17193
rect 14001 17184 14013 17187
rect 13964 17156 14013 17184
rect 13964 17144 13970 17156
rect 14001 17153 14013 17156
rect 14047 17153 14059 17187
rect 17681 17179 17693 17213
rect 17727 17179 17739 17213
rect 17681 17173 17739 17179
rect 14001 17147 14059 17153
rect 13817 17119 13875 17125
rect 13464 17088 13584 17116
rect 9140 17020 9536 17048
rect 9585 17051 9643 17057
rect 7984 17008 7990 17020
rect 9585 17017 9597 17051
rect 9631 17048 9643 17051
rect 9674 17048 9680 17060
rect 9631 17020 9680 17048
rect 9631 17017 9643 17020
rect 9585 17011 9643 17017
rect 9674 17008 9680 17020
rect 9732 17008 9738 17060
rect 12342 17048 12348 17060
rect 10161 17020 12348 17048
rect 10161 16980 10189 17020
rect 12342 17008 12348 17020
rect 12400 17008 12406 17060
rect 13556 17048 13584 17088
rect 13817 17085 13829 17119
rect 13863 17116 13875 17119
rect 14090 17116 14096 17128
rect 13863 17088 14096 17116
rect 13863 17085 13875 17088
rect 13817 17079 13875 17085
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 17494 17076 17500 17128
rect 17552 17116 17558 17128
rect 17695 17116 17723 17173
rect 17770 17144 17776 17196
rect 17828 17184 17834 17196
rect 17864 17187 17922 17193
rect 17864 17184 17876 17187
rect 17828 17156 17876 17184
rect 17828 17144 17834 17156
rect 17864 17153 17876 17156
rect 17910 17153 17922 17187
rect 17864 17147 17922 17153
rect 18049 17187 18107 17193
rect 18049 17153 18061 17187
rect 18095 17184 18107 17187
rect 18138 17184 18144 17196
rect 18095 17156 18144 17184
rect 18095 17153 18107 17156
rect 18049 17147 18107 17153
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 18233 17187 18291 17193
rect 18233 17153 18245 17187
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 17954 17116 17960 17128
rect 17552 17088 17723 17116
rect 17915 17088 17960 17116
rect 17552 17076 17558 17088
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 14366 17048 14372 17060
rect 13556 17020 14372 17048
rect 14366 17008 14372 17020
rect 14424 17008 14430 17060
rect 17402 17008 17408 17060
rect 17460 17048 17466 17060
rect 18248 17048 18276 17147
rect 18340 17116 18368 17224
rect 19306 17224 20996 17252
rect 18506 17144 18512 17196
rect 18564 17184 18570 17196
rect 18693 17187 18751 17193
rect 18693 17184 18705 17187
rect 18564 17156 18705 17184
rect 18564 17144 18570 17156
rect 18693 17153 18705 17156
rect 18739 17184 18751 17187
rect 19306 17184 19334 17224
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 22189 17255 22247 17261
rect 22189 17221 22201 17255
rect 22235 17252 22247 17255
rect 22278 17252 22284 17264
rect 22235 17224 22284 17252
rect 22235 17221 22247 17224
rect 22189 17215 22247 17221
rect 22278 17212 22284 17224
rect 22336 17212 22342 17264
rect 23109 17255 23167 17261
rect 23109 17221 23121 17255
rect 23155 17252 23167 17255
rect 23198 17252 23204 17264
rect 23155 17224 23204 17252
rect 23155 17221 23167 17224
rect 23109 17215 23167 17221
rect 23198 17212 23204 17224
rect 23256 17212 23262 17264
rect 20714 17184 20720 17196
rect 18739 17156 19334 17184
rect 20675 17156 20720 17184
rect 18739 17153 18751 17156
rect 18693 17147 18751 17153
rect 20714 17144 20720 17156
rect 20772 17144 20778 17196
rect 23014 17184 23020 17196
rect 22975 17156 23020 17184
rect 23014 17144 23020 17156
rect 23072 17144 23078 17196
rect 18874 17116 18880 17128
rect 18340 17088 18880 17116
rect 18874 17076 18880 17088
rect 18932 17116 18938 17128
rect 20254 17116 20260 17128
rect 18932 17088 20260 17116
rect 18932 17076 18938 17088
rect 20254 17076 20260 17088
rect 20312 17076 20318 17128
rect 21542 17076 21548 17128
rect 21600 17116 21606 17128
rect 22281 17119 22339 17125
rect 22281 17116 22293 17119
rect 21600 17088 22293 17116
rect 21600 17076 21606 17088
rect 22281 17085 22293 17088
rect 22327 17085 22339 17119
rect 22281 17079 22339 17085
rect 22370 17076 22376 17128
rect 22428 17116 22434 17128
rect 22465 17119 22523 17125
rect 22465 17116 22477 17119
rect 22428 17088 22477 17116
rect 22428 17076 22434 17088
rect 22465 17085 22477 17088
rect 22511 17116 22523 17119
rect 23106 17116 23112 17128
rect 22511 17088 23112 17116
rect 22511 17085 22523 17088
rect 22465 17079 22523 17085
rect 23106 17076 23112 17088
rect 23164 17116 23170 17128
rect 23201 17119 23259 17125
rect 23201 17116 23213 17119
rect 23164 17088 23213 17116
rect 23164 17076 23170 17088
rect 23201 17085 23213 17088
rect 23247 17085 23259 17119
rect 23201 17079 23259 17085
rect 18509 17051 18567 17057
rect 18509 17048 18521 17051
rect 17460 17020 18521 17048
rect 17460 17008 17466 17020
rect 18509 17017 18521 17020
rect 18555 17017 18567 17051
rect 18509 17011 18567 17017
rect 20990 17008 20996 17060
rect 21048 17048 21054 17060
rect 21637 17051 21695 17057
rect 21637 17048 21649 17051
rect 21048 17020 21649 17048
rect 21048 17008 21054 17020
rect 21637 17017 21649 17020
rect 21683 17048 21695 17051
rect 22388 17048 22416 17076
rect 21683 17020 22416 17048
rect 21683 17017 21695 17020
rect 21637 17011 21695 17017
rect 10318 16980 10324 16992
rect 5276 16952 10189 16980
rect 10279 16952 10324 16980
rect 5169 16943 5227 16949
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 12986 16980 12992 16992
rect 12947 16952 12992 16980
rect 12986 16940 12992 16952
rect 13044 16980 13050 16992
rect 13265 16983 13323 16989
rect 13265 16980 13277 16983
rect 13044 16952 13277 16980
rect 13044 16940 13050 16952
rect 13265 16949 13277 16952
rect 13311 16980 13323 16983
rect 13906 16980 13912 16992
rect 13311 16952 13912 16980
rect 13311 16949 13323 16952
rect 13265 16943 13323 16949
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 17218 16940 17224 16992
rect 17276 16980 17282 16992
rect 17770 16980 17776 16992
rect 17276 16952 17776 16980
rect 17276 16940 17282 16952
rect 17770 16940 17776 16952
rect 17828 16980 17834 16992
rect 18874 16980 18880 16992
rect 17828 16952 18880 16980
rect 17828 16940 17834 16952
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 1104 16890 26220 16912
rect 1104 16838 5136 16890
rect 5188 16838 5200 16890
rect 5252 16838 5264 16890
rect 5316 16838 5328 16890
rect 5380 16838 5392 16890
rect 5444 16838 13508 16890
rect 13560 16838 13572 16890
rect 13624 16838 13636 16890
rect 13688 16838 13700 16890
rect 13752 16838 13764 16890
rect 13816 16838 21880 16890
rect 21932 16838 21944 16890
rect 21996 16838 22008 16890
rect 22060 16838 22072 16890
rect 22124 16838 22136 16890
rect 22188 16838 26220 16890
rect 1104 16816 26220 16838
rect 3510 16776 3516 16788
rect 3471 16748 3516 16776
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 6181 16779 6239 16785
rect 6181 16776 6193 16779
rect 4264 16748 6193 16776
rect 2130 16640 2136 16652
rect 2091 16612 2136 16640
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 4264 16649 4292 16748
rect 6181 16745 6193 16748
rect 6227 16776 6239 16779
rect 6546 16776 6552 16788
rect 6227 16748 6552 16776
rect 6227 16745 6239 16748
rect 6181 16739 6239 16745
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 7926 16776 7932 16788
rect 6880 16748 7932 16776
rect 6880 16736 6886 16748
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8389 16779 8447 16785
rect 8389 16745 8401 16779
rect 8435 16776 8447 16779
rect 8662 16776 8668 16788
rect 8435 16748 8668 16776
rect 8435 16745 8447 16748
rect 8389 16739 8447 16745
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 8754 16736 8760 16788
rect 8812 16776 8818 16788
rect 9033 16779 9091 16785
rect 8812 16748 8857 16776
rect 8812 16736 8818 16748
rect 9033 16745 9045 16779
rect 9079 16776 9091 16779
rect 9306 16776 9312 16788
rect 9079 16748 9312 16776
rect 9079 16745 9091 16748
rect 9033 16739 9091 16745
rect 9306 16736 9312 16748
rect 9364 16776 9370 16788
rect 11514 16776 11520 16788
rect 9364 16748 11520 16776
rect 9364 16736 9370 16748
rect 11514 16736 11520 16748
rect 11572 16776 11578 16788
rect 11882 16776 11888 16788
rect 11572 16748 11888 16776
rect 11572 16736 11578 16748
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12621 16779 12679 16785
rect 12621 16745 12633 16779
rect 12667 16776 12679 16779
rect 12894 16776 12900 16788
rect 12667 16748 12900 16776
rect 12667 16745 12679 16748
rect 12621 16739 12679 16745
rect 12894 16736 12900 16748
rect 12952 16736 12958 16788
rect 13262 16736 13268 16788
rect 13320 16776 13326 16788
rect 13541 16779 13599 16785
rect 13541 16776 13553 16779
rect 13320 16748 13553 16776
rect 13320 16736 13326 16748
rect 13541 16745 13553 16748
rect 13587 16745 13599 16779
rect 13541 16739 13599 16745
rect 16206 16736 16212 16788
rect 16264 16776 16270 16788
rect 17034 16776 17040 16788
rect 16264 16748 17040 16776
rect 16264 16736 16270 16748
rect 17034 16736 17040 16748
rect 17092 16776 17098 16788
rect 20898 16776 20904 16788
rect 17092 16748 17908 16776
rect 20859 16748 20904 16776
rect 17092 16736 17098 16748
rect 4338 16668 4344 16720
rect 4396 16708 4402 16720
rect 4617 16711 4675 16717
rect 4617 16708 4629 16711
rect 4396 16680 4629 16708
rect 4396 16668 4402 16680
rect 4448 16649 4476 16680
rect 4617 16677 4629 16680
rect 4663 16677 4675 16711
rect 4617 16671 4675 16677
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16609 4307 16643
rect 4249 16603 4307 16609
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4479 16612 4513 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4706 16600 4712 16652
rect 4764 16640 4770 16652
rect 4801 16643 4859 16649
rect 4801 16640 4813 16643
rect 4764 16612 4813 16640
rect 4764 16600 4770 16612
rect 4801 16609 4813 16612
rect 4847 16609 4859 16643
rect 4801 16603 4859 16609
rect 7837 16643 7895 16649
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8294 16640 8300 16652
rect 7883 16612 8300 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8294 16600 8300 16612
rect 8352 16640 8358 16652
rect 9401 16643 9459 16649
rect 9401 16640 9413 16643
rect 8352 16612 9413 16640
rect 8352 16600 8358 16612
rect 9401 16609 9413 16612
rect 9447 16640 9459 16643
rect 12912 16640 12940 16736
rect 15562 16668 15568 16720
rect 15620 16708 15626 16720
rect 15749 16711 15807 16717
rect 15749 16708 15761 16711
rect 15620 16680 15761 16708
rect 15620 16668 15626 16680
rect 15749 16677 15761 16680
rect 15795 16708 15807 16711
rect 16574 16708 16580 16720
rect 15795 16680 16160 16708
rect 16535 16680 16580 16708
rect 15795 16677 15807 16680
rect 15749 16671 15807 16677
rect 13265 16643 13323 16649
rect 13265 16640 13277 16643
rect 9447 16612 9536 16640
rect 12912 16612 13277 16640
rect 9447 16609 9459 16612
rect 9401 16603 9459 16609
rect 4154 16572 4160 16584
rect 4115 16544 4160 16572
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 8018 16532 8024 16584
rect 8076 16572 8082 16584
rect 8202 16572 8208 16584
rect 8076 16544 8208 16572
rect 8076 16532 8082 16544
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 9309 16575 9367 16581
rect 9309 16541 9321 16575
rect 9355 16541 9367 16575
rect 9508 16572 9536 16612
rect 13265 16609 13277 16612
rect 13311 16609 13323 16643
rect 13265 16603 13323 16609
rect 15470 16600 15476 16652
rect 15528 16640 15534 16652
rect 16132 16649 16160 16680
rect 16574 16668 16580 16680
rect 16632 16668 16638 16720
rect 17880 16649 17908 16748
rect 20898 16736 20904 16748
rect 20956 16736 20962 16788
rect 22370 16736 22376 16788
rect 22428 16776 22434 16788
rect 22465 16779 22523 16785
rect 22465 16776 22477 16779
rect 22428 16748 22477 16776
rect 22428 16736 22434 16748
rect 22465 16745 22477 16748
rect 22511 16745 22523 16779
rect 23106 16776 23112 16788
rect 22465 16739 22523 16745
rect 22664 16748 23112 16776
rect 18506 16668 18512 16720
rect 18564 16708 18570 16720
rect 18564 16680 19012 16708
rect 18564 16668 18570 16680
rect 18984 16649 19012 16680
rect 19058 16668 19064 16720
rect 19116 16708 19122 16720
rect 20916 16708 20944 16736
rect 22664 16708 22692 16748
rect 23106 16736 23112 16748
rect 23164 16776 23170 16788
rect 23290 16776 23296 16788
rect 23164 16748 23296 16776
rect 23164 16736 23170 16748
rect 23290 16736 23296 16748
rect 23348 16736 23354 16788
rect 19116 16680 19288 16708
rect 19116 16668 19122 16680
rect 19260 16649 19288 16680
rect 20916 16680 22692 16708
rect 16117 16643 16175 16649
rect 15528 16612 15976 16640
rect 15528 16600 15534 16612
rect 10594 16572 10600 16584
rect 9508 16544 9812 16572
rect 9309 16535 9367 16541
rect 2400 16507 2458 16513
rect 2400 16473 2412 16507
rect 2446 16504 2458 16507
rect 4798 16504 4804 16516
rect 2446 16476 4804 16504
rect 2446 16473 2458 16476
rect 2400 16467 2458 16473
rect 4798 16464 4804 16476
rect 4856 16464 4862 16516
rect 5068 16507 5126 16513
rect 5068 16473 5080 16507
rect 5114 16504 5126 16507
rect 6270 16504 6276 16516
rect 5114 16476 6276 16504
rect 5114 16473 5126 16476
rect 5068 16467 5126 16473
rect 6270 16464 6276 16476
rect 6328 16464 6334 16516
rect 7282 16464 7288 16516
rect 7340 16504 7346 16516
rect 7570 16507 7628 16513
rect 7570 16504 7582 16507
rect 7340 16476 7582 16504
rect 7340 16464 7346 16476
rect 7570 16473 7582 16476
rect 7616 16473 7628 16507
rect 7570 16467 7628 16473
rect 3786 16436 3792 16448
rect 3747 16408 3792 16436
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 6362 16396 6368 16448
rect 6420 16436 6426 16448
rect 6457 16439 6515 16445
rect 6457 16436 6469 16439
rect 6420 16408 6469 16436
rect 6420 16396 6426 16408
rect 6457 16405 6469 16408
rect 6503 16405 6515 16439
rect 6457 16399 6515 16405
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16436 9183 16439
rect 9214 16436 9220 16448
rect 9171 16408 9220 16436
rect 9171 16405 9183 16408
rect 9125 16399 9183 16405
rect 9214 16396 9220 16408
rect 9272 16396 9278 16448
rect 9324 16436 9352 16535
rect 9784 16516 9812 16544
rect 10244 16544 10600 16572
rect 9490 16464 9496 16516
rect 9548 16504 9554 16516
rect 9646 16507 9704 16513
rect 9646 16504 9658 16507
rect 9548 16476 9658 16504
rect 9548 16464 9554 16476
rect 9646 16473 9658 16476
rect 9692 16473 9704 16507
rect 9646 16467 9704 16473
rect 9766 16464 9772 16516
rect 9824 16464 9830 16516
rect 10244 16436 10272 16544
rect 10594 16532 10600 16544
rect 10652 16572 10658 16584
rect 10965 16575 11023 16581
rect 10965 16572 10977 16575
rect 10652 16544 10977 16572
rect 10652 16532 10658 16544
rect 10965 16541 10977 16544
rect 11011 16541 11023 16575
rect 15565 16575 15623 16581
rect 15565 16572 15577 16575
rect 10965 16535 11023 16541
rect 15212 16544 15577 16572
rect 12250 16464 12256 16516
rect 12308 16504 12314 16516
rect 15212 16504 15240 16544
rect 15565 16541 15577 16544
rect 15611 16572 15623 16575
rect 15746 16572 15752 16584
rect 15611 16544 15752 16572
rect 15611 16541 15623 16544
rect 15565 16535 15623 16541
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16541 15899 16575
rect 15948 16572 15976 16612
rect 16117 16609 16129 16643
rect 16163 16640 16175 16643
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 16163 16612 16957 16640
rect 16163 16609 16175 16612
rect 16117 16603 16175 16609
rect 16945 16609 16957 16612
rect 16991 16640 17003 16643
rect 17773 16643 17831 16649
rect 17773 16640 17785 16643
rect 16991 16612 17785 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 17773 16609 17785 16612
rect 17819 16609 17831 16643
rect 17773 16603 17831 16609
rect 17865 16643 17923 16649
rect 17865 16609 17877 16643
rect 17911 16609 17923 16643
rect 17865 16603 17923 16609
rect 18233 16643 18291 16649
rect 18233 16609 18245 16643
rect 18279 16640 18291 16643
rect 18969 16643 19027 16649
rect 18279 16612 18920 16640
rect 18279 16609 18291 16612
rect 18233 16603 18291 16609
rect 16006 16575 16064 16581
rect 16006 16572 16018 16575
rect 15948 16544 16018 16572
rect 15841 16535 15899 16541
rect 16006 16541 16018 16544
rect 16052 16541 16064 16575
rect 16206 16572 16212 16584
rect 16167 16544 16212 16572
rect 16006 16535 16064 16541
rect 12308 16476 15240 16504
rect 12308 16464 12314 16476
rect 15286 16464 15292 16516
rect 15344 16504 15350 16516
rect 15856 16504 15884 16535
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 16390 16572 16396 16584
rect 16351 16544 16396 16572
rect 16390 16532 16396 16544
rect 16448 16532 16454 16584
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 16850 16572 16856 16584
rect 16811 16544 16856 16572
rect 16669 16535 16727 16541
rect 16684 16504 16712 16535
rect 16850 16532 16856 16544
rect 16908 16532 16914 16584
rect 17034 16572 17040 16584
rect 16995 16544 17040 16572
rect 17034 16532 17040 16544
rect 17092 16532 17098 16584
rect 17218 16572 17224 16584
rect 17179 16544 17224 16572
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 17494 16572 17500 16584
rect 17455 16544 17500 16572
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 17586 16532 17592 16584
rect 17644 16572 17650 16584
rect 17680 16575 17738 16581
rect 17680 16572 17692 16575
rect 17644 16544 17692 16572
rect 17644 16532 17650 16544
rect 17680 16541 17692 16544
rect 17726 16541 17738 16575
rect 17680 16535 17738 16541
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16541 18107 16575
rect 18892 16572 18920 16612
rect 18969 16609 18981 16643
rect 19015 16609 19027 16643
rect 18969 16603 19027 16609
rect 19245 16643 19303 16649
rect 19245 16609 19257 16643
rect 19291 16609 19303 16643
rect 20916 16640 20944 16680
rect 22830 16668 22836 16720
rect 22888 16708 22894 16720
rect 22888 16680 23244 16708
rect 22888 16668 22894 16680
rect 21085 16643 21143 16649
rect 21085 16640 21097 16643
rect 20916 16612 21097 16640
rect 19245 16603 19303 16609
rect 21085 16609 21097 16612
rect 21131 16609 21143 16643
rect 21085 16603 21143 16609
rect 22738 16600 22744 16652
rect 22796 16640 22802 16652
rect 23216 16649 23244 16680
rect 23109 16643 23167 16649
rect 23109 16640 23121 16643
rect 22796 16612 23121 16640
rect 22796 16600 22802 16612
rect 23109 16609 23121 16612
rect 23155 16609 23167 16643
rect 23109 16603 23167 16609
rect 23201 16643 23259 16649
rect 23201 16609 23213 16643
rect 23247 16609 23259 16643
rect 23201 16603 23259 16609
rect 19501 16575 19559 16581
rect 19501 16572 19513 16575
rect 18892 16544 19513 16572
rect 18049 16535 18107 16541
rect 19501 16541 19513 16544
rect 19547 16541 19559 16575
rect 19501 16535 19559 16541
rect 17512 16504 17540 16532
rect 15344 16476 17540 16504
rect 18064 16504 18092 16535
rect 19886 16532 19892 16584
rect 19944 16572 19950 16584
rect 20622 16572 20628 16584
rect 19944 16544 20628 16572
rect 19944 16532 19950 16544
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 21358 16532 21364 16584
rect 21416 16572 21422 16584
rect 22830 16572 22836 16584
rect 21416 16544 22836 16572
rect 21416 16532 21422 16544
rect 22830 16532 22836 16544
rect 22888 16532 22894 16584
rect 23016 16575 23074 16581
rect 23016 16541 23028 16575
rect 23062 16572 23074 16575
rect 23382 16572 23388 16584
rect 23062 16544 23244 16572
rect 23343 16544 23388 16572
rect 23062 16541 23074 16544
rect 23016 16535 23074 16541
rect 19904 16504 19932 16532
rect 20714 16504 20720 16516
rect 18064 16476 19932 16504
rect 20627 16476 20720 16504
rect 15344 16464 15350 16476
rect 9324 16408 10272 16436
rect 10594 16396 10600 16448
rect 10652 16436 10658 16448
rect 10781 16439 10839 16445
rect 10781 16436 10793 16439
rect 10652 16408 10793 16436
rect 10652 16396 10658 16408
rect 10781 16405 10793 16408
rect 10827 16405 10839 16439
rect 10781 16399 10839 16405
rect 11057 16439 11115 16445
rect 11057 16405 11069 16439
rect 11103 16436 11115 16439
rect 11698 16436 11704 16448
rect 11103 16408 11704 16436
rect 11103 16405 11115 16408
rect 11057 16399 11115 16405
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 12713 16439 12771 16445
rect 12713 16405 12725 16439
rect 12759 16436 12771 16439
rect 12802 16436 12808 16448
rect 12759 16408 12808 16436
rect 12759 16405 12771 16408
rect 12713 16399 12771 16405
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 13078 16436 13084 16448
rect 13039 16408 13084 16436
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 13173 16439 13231 16445
rect 13173 16405 13185 16439
rect 13219 16436 13231 16439
rect 13262 16436 13268 16448
rect 13219 16408 13268 16436
rect 13219 16405 13231 16408
rect 13173 16399 13231 16405
rect 13262 16396 13268 16408
rect 13320 16396 13326 16448
rect 15470 16436 15476 16448
rect 15431 16408 15476 16436
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15930 16396 15936 16448
rect 15988 16436 15994 16448
rect 16758 16436 16764 16448
rect 15988 16408 16764 16436
rect 15988 16396 15994 16408
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 17218 16396 17224 16448
rect 17276 16436 17282 16448
rect 17313 16439 17371 16445
rect 17313 16436 17325 16439
rect 17276 16408 17325 16436
rect 17276 16396 17282 16408
rect 17313 16405 17325 16408
rect 17359 16405 17371 16439
rect 18322 16436 18328 16448
rect 18283 16408 18328 16436
rect 17313 16399 17371 16405
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 18414 16396 18420 16448
rect 18472 16436 18478 16448
rect 18693 16439 18751 16445
rect 18693 16436 18705 16439
rect 18472 16408 18705 16436
rect 18472 16396 18478 16408
rect 18693 16405 18705 16408
rect 18739 16405 18751 16439
rect 18693 16399 18751 16405
rect 18782 16396 18788 16448
rect 18840 16436 18846 16448
rect 20640 16445 20668 16476
rect 20714 16464 20720 16476
rect 20772 16504 20778 16516
rect 23216 16504 23244 16544
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 23290 16504 23296 16516
rect 20772 16476 21312 16504
rect 23216 16476 23296 16504
rect 20772 16464 20778 16476
rect 21284 16448 21312 16476
rect 23290 16464 23296 16476
rect 23348 16464 23354 16516
rect 23569 16507 23627 16513
rect 23569 16473 23581 16507
rect 23615 16504 23627 16507
rect 24118 16504 24124 16516
rect 23615 16476 24124 16504
rect 23615 16473 23627 16476
rect 23569 16467 23627 16473
rect 24118 16464 24124 16476
rect 24176 16464 24182 16516
rect 20625 16439 20683 16445
rect 18840 16408 18885 16436
rect 18840 16396 18846 16408
rect 20625 16405 20637 16439
rect 20671 16405 20683 16439
rect 21266 16436 21272 16448
rect 21227 16408 21272 16436
rect 20625 16399 20683 16405
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 21361 16439 21419 16445
rect 21361 16405 21373 16439
rect 21407 16436 21419 16439
rect 21542 16436 21548 16448
rect 21407 16408 21548 16436
rect 21407 16405 21419 16408
rect 21361 16399 21419 16405
rect 21542 16396 21548 16408
rect 21600 16396 21606 16448
rect 21729 16439 21787 16445
rect 21729 16405 21741 16439
rect 21775 16436 21787 16439
rect 22278 16436 22284 16448
rect 21775 16408 22284 16436
rect 21775 16405 21787 16408
rect 21729 16399 21787 16405
rect 22278 16396 22284 16408
rect 22336 16396 22342 16448
rect 1104 16346 26220 16368
rect 1104 16294 9322 16346
rect 9374 16294 9386 16346
rect 9438 16294 9450 16346
rect 9502 16294 9514 16346
rect 9566 16294 9578 16346
rect 9630 16294 17694 16346
rect 17746 16294 17758 16346
rect 17810 16294 17822 16346
rect 17874 16294 17886 16346
rect 17938 16294 17950 16346
rect 18002 16294 26220 16346
rect 1104 16272 26220 16294
rect 2130 16232 2136 16244
rect 1872 16204 2136 16232
rect 1872 16105 1900 16204
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 3237 16235 3295 16241
rect 3237 16201 3249 16235
rect 3283 16232 3295 16235
rect 3418 16232 3424 16244
rect 3283 16204 3424 16232
rect 3283 16201 3295 16204
rect 3237 16195 3295 16201
rect 3418 16192 3424 16204
rect 3476 16232 3482 16244
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 3476 16204 3893 16232
rect 3476 16192 3482 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 3881 16195 3939 16201
rect 4249 16235 4307 16241
rect 4249 16201 4261 16235
rect 4295 16232 4307 16235
rect 4982 16232 4988 16244
rect 4295 16204 4988 16232
rect 4295 16201 4307 16204
rect 4249 16195 4307 16201
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 6270 16192 6276 16244
rect 6328 16232 6334 16244
rect 6457 16235 6515 16241
rect 6457 16232 6469 16235
rect 6328 16204 6469 16232
rect 6328 16192 6334 16204
rect 6457 16201 6469 16204
rect 6503 16201 6515 16235
rect 7282 16232 7288 16244
rect 7243 16204 7288 16232
rect 6457 16195 6515 16201
rect 7282 16192 7288 16204
rect 7340 16192 7346 16244
rect 7374 16192 7380 16244
rect 7432 16232 7438 16244
rect 7742 16232 7748 16244
rect 7432 16204 7748 16232
rect 7432 16192 7438 16204
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 10134 16232 10140 16244
rect 9417 16204 10140 16232
rect 3789 16167 3847 16173
rect 3789 16133 3801 16167
rect 3835 16164 3847 16167
rect 6362 16164 6368 16176
rect 3835 16136 6368 16164
rect 3835 16133 3847 16136
rect 3789 16127 3847 16133
rect 6362 16124 6368 16136
rect 6420 16164 6426 16176
rect 7760 16164 7788 16192
rect 6420 16136 7420 16164
rect 7760 16136 7972 16164
rect 6420 16124 6426 16136
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16065 1915 16099
rect 1857 16059 1915 16065
rect 2124 16099 2182 16105
rect 2124 16065 2136 16099
rect 2170 16096 2182 16099
rect 2866 16096 2872 16108
rect 2170 16068 2872 16096
rect 2170 16065 2182 16068
rect 2124 16059 2182 16065
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 4338 16096 4344 16108
rect 3712 16068 4344 16096
rect 3712 16037 3740 16068
rect 4338 16056 4344 16068
rect 4396 16056 4402 16108
rect 6546 16096 6552 16108
rect 6507 16068 6552 16096
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 6822 16096 6828 16108
rect 6783 16068 6828 16096
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 7101 16099 7159 16105
rect 6972 16068 7017 16096
rect 6972 16056 6978 16068
rect 7101 16065 7113 16099
rect 7147 16096 7159 16099
rect 7282 16096 7288 16108
rect 7147 16068 7288 16096
rect 7147 16065 7159 16068
rect 7101 16059 7159 16065
rect 7282 16056 7288 16068
rect 7340 16056 7346 16108
rect 7392 16105 7420 16136
rect 7944 16105 7972 16136
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16065 7435 16099
rect 7653 16099 7711 16105
rect 7653 16096 7665 16099
rect 7377 16059 7435 16065
rect 7484 16068 7665 16096
rect 3697 16031 3755 16037
rect 3697 15997 3709 16031
rect 3743 15997 3755 16031
rect 3697 15991 3755 15997
rect 5810 15988 5816 16040
rect 5868 16028 5874 16040
rect 6733 16031 6791 16037
rect 6733 16028 6745 16031
rect 5868 16000 6745 16028
rect 5868 15988 5874 16000
rect 6733 15997 6745 16000
rect 6779 15997 6791 16031
rect 6840 16028 6868 16056
rect 7484 16028 7512 16068
rect 7653 16065 7665 16068
rect 7699 16065 7711 16099
rect 7653 16059 7711 16065
rect 7763 16099 7821 16105
rect 7763 16065 7775 16099
rect 7809 16065 7821 16099
rect 7763 16059 7821 16065
rect 7929 16099 7987 16105
rect 7929 16065 7941 16099
rect 7975 16065 7987 16099
rect 8294 16096 8300 16108
rect 8255 16068 8300 16096
rect 7929 16059 7987 16065
rect 6840 16000 7512 16028
rect 7561 16031 7619 16037
rect 6733 15991 6791 15997
rect 7561 15997 7573 16031
rect 7607 15997 7619 16031
rect 7778 16028 7806 16059
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 8662 16056 8668 16108
rect 8720 16096 8726 16108
rect 8941 16099 8999 16105
rect 8941 16096 8953 16099
rect 8720 16068 8953 16096
rect 8720 16056 8726 16068
rect 8941 16065 8953 16068
rect 8987 16065 8999 16099
rect 9122 16096 9128 16108
rect 8941 16059 8999 16065
rect 9048 16068 9128 16096
rect 8312 16028 8340 16056
rect 7778 16000 8340 16028
rect 7561 15991 7619 15997
rect 6748 15960 6776 15991
rect 7576 15960 7604 15991
rect 8570 15988 8576 16040
rect 8628 16028 8634 16040
rect 9048 16028 9076 16068
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 9309 16099 9367 16105
rect 9309 16065 9321 16099
rect 9355 16096 9367 16099
rect 9417 16096 9445 16204
rect 10134 16192 10140 16204
rect 10192 16232 10198 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 10192 16204 11529 16232
rect 10192 16192 10198 16204
rect 11517 16201 11529 16204
rect 11563 16201 11575 16235
rect 11517 16195 11575 16201
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 12618 16232 12624 16244
rect 12483 16204 12624 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 9582 16124 9588 16176
rect 9640 16164 9646 16176
rect 10036 16167 10094 16173
rect 9640 16136 9904 16164
rect 9640 16124 9646 16136
rect 9355 16068 9445 16096
rect 9493 16099 9551 16105
rect 9355 16065 9367 16068
rect 9309 16059 9367 16065
rect 9493 16065 9505 16099
rect 9539 16065 9551 16099
rect 9766 16096 9772 16108
rect 9727 16068 9772 16096
rect 9493 16059 9551 16065
rect 9214 16028 9220 16040
rect 8628 16000 9076 16028
rect 9175 16000 9220 16028
rect 8628 15988 8634 16000
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 9508 15972 9536 16059
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 9876 16096 9904 16136
rect 10036 16133 10048 16167
rect 10082 16164 10094 16167
rect 10318 16164 10324 16176
rect 10082 16136 10324 16164
rect 10082 16133 10094 16136
rect 10036 16127 10094 16133
rect 10318 16124 10324 16136
rect 10376 16124 10382 16176
rect 12452 16164 12480 16195
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 13081 16235 13139 16241
rect 13081 16201 13093 16235
rect 13127 16232 13139 16235
rect 13541 16235 13599 16241
rect 13541 16232 13553 16235
rect 13127 16204 13553 16232
rect 13127 16201 13139 16204
rect 13081 16195 13139 16201
rect 13541 16201 13553 16204
rect 13587 16201 13599 16235
rect 14366 16232 14372 16244
rect 14279 16204 14372 16232
rect 13541 16195 13599 16201
rect 14366 16192 14372 16204
rect 14424 16232 14430 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 14424 16204 15025 16232
rect 14424 16192 14430 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 15013 16195 15071 16201
rect 16206 16192 16212 16244
rect 16264 16232 16270 16244
rect 16301 16235 16359 16241
rect 16301 16232 16313 16235
rect 16264 16204 16313 16232
rect 16264 16192 16270 16204
rect 16301 16201 16313 16204
rect 16347 16201 16359 16235
rect 16301 16195 16359 16201
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 16448 16204 18061 16232
rect 16448 16192 16454 16204
rect 18049 16201 18061 16204
rect 18095 16232 18107 16235
rect 18230 16232 18236 16244
rect 18095 16204 18236 16232
rect 18095 16201 18107 16204
rect 18049 16195 18107 16201
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 18414 16232 18420 16244
rect 18375 16204 18420 16232
rect 18414 16192 18420 16204
rect 18472 16192 18478 16244
rect 18874 16232 18880 16244
rect 18835 16204 18880 16232
rect 18874 16192 18880 16204
rect 18932 16192 18938 16244
rect 19521 16235 19579 16241
rect 19521 16201 19533 16235
rect 19567 16232 19579 16235
rect 20254 16232 20260 16244
rect 19567 16204 20260 16232
rect 19567 16201 19579 16204
rect 19521 16195 19579 16201
rect 20254 16192 20260 16204
rect 20312 16192 20318 16244
rect 20993 16235 21051 16241
rect 20993 16201 21005 16235
rect 21039 16201 21051 16235
rect 24210 16232 24216 16244
rect 20993 16195 21051 16201
rect 22296 16204 24216 16232
rect 10888 16136 12480 16164
rect 12544 16136 16160 16164
rect 10778 16096 10784 16108
rect 9876 16068 10784 16096
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 9582 15988 9588 16040
rect 9640 16028 9646 16040
rect 9677 16031 9735 16037
rect 9677 16028 9689 16031
rect 9640 16000 9689 16028
rect 9640 15988 9646 16000
rect 9677 15997 9689 16000
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 6748 15932 7604 15960
rect 8754 15920 8760 15972
rect 8812 15960 8818 15972
rect 9490 15960 9496 15972
rect 8812 15932 9496 15960
rect 8812 15920 8818 15932
rect 9490 15920 9496 15932
rect 9548 15920 9554 15972
rect 6914 15852 6920 15904
rect 6972 15892 6978 15904
rect 8018 15892 8024 15904
rect 6972 15864 8024 15892
rect 6972 15852 6978 15864
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 8202 15852 8208 15904
rect 8260 15892 8266 15904
rect 10888 15892 10916 16136
rect 11698 16096 11704 16108
rect 11659 16068 11704 16096
rect 11698 16056 11704 16068
rect 11756 16096 11762 16108
rect 12158 16096 12164 16108
rect 11756 16068 12164 16096
rect 11756 16056 11762 16068
rect 12158 16056 12164 16068
rect 12216 16096 12222 16108
rect 12544 16096 12572 16136
rect 12216 16068 12572 16096
rect 12621 16099 12679 16105
rect 12216 16056 12222 16068
rect 12621 16065 12633 16099
rect 12667 16096 12679 16099
rect 12989 16099 13047 16105
rect 12667 16068 12940 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 12345 16031 12403 16037
rect 12345 15997 12357 16031
rect 12391 16028 12403 16031
rect 12802 16028 12808 16040
rect 12391 16000 12808 16028
rect 12391 15997 12403 16000
rect 12345 15991 12403 15997
rect 12802 15988 12808 16000
rect 12860 15988 12866 16040
rect 12912 15904 12940 16068
rect 12989 16065 13001 16099
rect 13035 16096 13047 16099
rect 13909 16099 13967 16105
rect 13909 16096 13921 16099
rect 13035 16068 13921 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 13909 16065 13921 16068
rect 13955 16096 13967 16099
rect 14182 16096 14188 16108
rect 13955 16068 14188 16096
rect 13955 16065 13967 16068
rect 13909 16059 13967 16065
rect 14182 16056 14188 16068
rect 14240 16056 14246 16108
rect 14274 16056 14280 16108
rect 14332 16096 14338 16108
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 14332 16068 14565 16096
rect 14332 16056 14338 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 15289 16099 15347 16105
rect 15289 16096 15301 16099
rect 15059 16068 15301 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 15289 16065 15301 16068
rect 15335 16065 15347 16099
rect 15454 16099 15512 16105
rect 15454 16096 15466 16099
rect 15289 16059 15347 16065
rect 15396 16068 15466 16096
rect 13354 15988 13360 16040
rect 13412 16028 13418 16040
rect 14001 16031 14059 16037
rect 14001 16028 14013 16031
rect 13412 16000 14013 16028
rect 13412 15988 13418 16000
rect 14001 15997 14013 16000
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 14093 16031 14151 16037
rect 14093 15997 14105 16031
rect 14139 16028 14151 16031
rect 14366 16028 14372 16040
rect 14139 16000 14372 16028
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 15194 15988 15200 16040
rect 15252 16028 15258 16040
rect 15396 16028 15424 16068
rect 15454 16065 15466 16068
rect 15500 16065 15512 16099
rect 15454 16059 15512 16065
rect 15562 16056 15568 16108
rect 15620 16096 15626 16108
rect 15841 16099 15899 16105
rect 15620 16068 15665 16096
rect 15620 16056 15626 16068
rect 15841 16065 15853 16099
rect 15887 16096 15899 16099
rect 15930 16096 15936 16108
rect 15887 16068 15936 16096
rect 15887 16065 15899 16068
rect 15841 16059 15899 16065
rect 15930 16056 15936 16068
rect 15988 16056 15994 16108
rect 16132 16105 16160 16136
rect 16574 16124 16580 16176
rect 16632 16164 16638 16176
rect 16914 16167 16972 16173
rect 16914 16164 16926 16167
rect 16632 16136 16926 16164
rect 16632 16124 16638 16136
rect 16914 16133 16926 16136
rect 16960 16133 16972 16167
rect 16914 16127 16972 16133
rect 19058 16124 19064 16176
rect 19116 16164 19122 16176
rect 20809 16167 20867 16173
rect 20809 16164 20821 16167
rect 19116 16136 20821 16164
rect 19116 16124 19122 16136
rect 20809 16133 20821 16136
rect 20855 16164 20867 16167
rect 21008 16164 21036 16195
rect 20855 16136 21036 16164
rect 20855 16133 20867 16136
rect 20809 16127 20867 16133
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16666 16096 16672 16108
rect 16163 16068 16528 16096
rect 16627 16068 16672 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 15252 16000 15424 16028
rect 15657 16031 15715 16037
rect 15252 15988 15258 16000
rect 15657 15997 15669 16031
rect 15703 16028 15715 16031
rect 16206 16028 16212 16040
rect 15703 16000 16212 16028
rect 15703 15997 15715 16000
rect 15657 15991 15715 15997
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 16500 16028 16528 16068
rect 16666 16056 16672 16068
rect 16724 16056 16730 16108
rect 18598 16056 18604 16108
rect 18656 16096 18662 16108
rect 18782 16096 18788 16108
rect 18656 16068 18788 16096
rect 18656 16056 18662 16068
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19392 16068 19717 16096
rect 19392 16056 19398 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19886 16096 19892 16108
rect 19847 16068 19892 16096
rect 19705 16059 19763 16065
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 20165 16099 20223 16105
rect 20165 16065 20177 16099
rect 20211 16096 20223 16099
rect 20441 16099 20499 16105
rect 20441 16096 20453 16099
rect 20211 16068 20453 16096
rect 20211 16065 20223 16068
rect 20165 16059 20223 16065
rect 20441 16065 20453 16068
rect 20487 16096 20499 16099
rect 20622 16096 20628 16108
rect 20487 16068 20628 16096
rect 20487 16065 20499 16068
rect 20441 16059 20499 16065
rect 16574 16028 16580 16040
rect 16500 16000 16580 16028
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 15997 19027 16031
rect 18969 15991 19027 15997
rect 13170 15920 13176 15972
rect 13228 15960 13234 15972
rect 13449 15963 13507 15969
rect 13449 15960 13461 15963
rect 13228 15932 13461 15960
rect 13228 15920 13234 15932
rect 13449 15929 13461 15932
rect 13495 15929 13507 15963
rect 18782 15960 18788 15972
rect 13449 15923 13507 15929
rect 13556 15932 16068 15960
rect 11146 15892 11152 15904
rect 8260 15864 10916 15892
rect 11107 15864 11152 15892
rect 8260 15852 8266 15864
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 12894 15892 12900 15904
rect 12807 15864 12900 15892
rect 12894 15852 12900 15864
rect 12952 15892 12958 15904
rect 13556 15892 13584 15932
rect 15194 15892 15200 15904
rect 12952 15864 13584 15892
rect 15155 15864 15200 15892
rect 12952 15852 12958 15864
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 15930 15892 15936 15904
rect 15891 15864 15936 15892
rect 15930 15852 15936 15864
rect 15988 15852 15994 15904
rect 16040 15892 16068 15932
rect 17604 15932 18788 15960
rect 17604 15892 17632 15932
rect 18782 15920 18788 15932
rect 18840 15920 18846 15972
rect 16040 15864 17632 15892
rect 18138 15852 18144 15904
rect 18196 15892 18202 15904
rect 18233 15895 18291 15901
rect 18233 15892 18245 15895
rect 18196 15864 18245 15892
rect 18196 15852 18202 15864
rect 18233 15861 18245 15864
rect 18279 15892 18291 15895
rect 18984 15892 19012 15991
rect 18279 15864 19012 15892
rect 19996 15892 20024 16059
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 21361 16099 21419 16105
rect 21361 16096 21373 16099
rect 21100 16068 21373 16096
rect 20346 16028 20352 16040
rect 20307 16000 20352 16028
rect 20346 15988 20352 16000
rect 20404 15988 20410 16040
rect 20070 15920 20076 15972
rect 20128 15960 20134 15972
rect 20441 15963 20499 15969
rect 20441 15960 20453 15963
rect 20128 15932 20453 15960
rect 20128 15920 20134 15932
rect 20441 15929 20453 15932
rect 20487 15960 20499 15963
rect 20530 15960 20536 15972
rect 20487 15932 20536 15960
rect 20487 15929 20499 15932
rect 20441 15923 20499 15929
rect 20530 15920 20536 15932
rect 20588 15920 20594 15972
rect 21100 15904 21128 16068
rect 21361 16065 21373 16068
rect 21407 16065 21419 16099
rect 21361 16059 21419 16065
rect 21726 16056 21732 16108
rect 21784 16096 21790 16108
rect 22296 16096 22324 16204
rect 22370 16105 22376 16108
rect 21784 16068 22324 16096
rect 21784 16056 21790 16068
rect 21269 16031 21327 16037
rect 21269 15997 21281 16031
rect 21315 16028 21327 16031
rect 21450 16028 21456 16040
rect 21315 16000 21456 16028
rect 21315 15997 21327 16000
rect 21269 15991 21327 15997
rect 21450 15988 21456 16000
rect 21508 15988 21514 16040
rect 22112 16037 22140 16068
rect 22364 16059 22376 16105
rect 22428 16096 22434 16108
rect 24044 16105 24072 16204
rect 24210 16192 24216 16204
rect 24268 16192 24274 16244
rect 24118 16124 24124 16176
rect 24176 16164 24182 16176
rect 24296 16167 24354 16173
rect 24296 16164 24308 16167
rect 24176 16136 24308 16164
rect 24176 16124 24182 16136
rect 24296 16133 24308 16136
rect 24342 16133 24354 16167
rect 24296 16127 24354 16133
rect 24029 16099 24087 16105
rect 22428 16068 22464 16096
rect 22370 16056 22376 16059
rect 22428 16056 22434 16068
rect 24029 16065 24041 16099
rect 24075 16065 24087 16099
rect 24029 16059 24087 16065
rect 22097 16031 22155 16037
rect 22097 15997 22109 16031
rect 22143 16028 22155 16031
rect 22143 16000 22177 16028
rect 22143 15997 22155 16000
rect 22097 15991 22155 15997
rect 23382 15920 23388 15972
rect 23440 15960 23446 15972
rect 23440 15932 23612 15960
rect 23440 15920 23446 15932
rect 21082 15892 21088 15904
rect 19996 15864 21088 15892
rect 18279 15861 18291 15864
rect 18233 15855 18291 15861
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 21266 15892 21272 15904
rect 21227 15864 21272 15892
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 23474 15892 23480 15904
rect 23435 15864 23480 15892
rect 23474 15852 23480 15864
rect 23532 15852 23538 15904
rect 23584 15892 23612 15932
rect 25409 15895 25467 15901
rect 25409 15892 25421 15895
rect 23584 15864 25421 15892
rect 25409 15861 25421 15864
rect 25455 15892 25467 15895
rect 26329 15895 26387 15901
rect 26329 15892 26341 15895
rect 25455 15864 26341 15892
rect 25455 15861 25467 15864
rect 25409 15855 25467 15861
rect 26329 15861 26341 15864
rect 26375 15861 26387 15895
rect 26329 15855 26387 15861
rect 1104 15802 26220 15824
rect 1104 15750 5136 15802
rect 5188 15750 5200 15802
rect 5252 15750 5264 15802
rect 5316 15750 5328 15802
rect 5380 15750 5392 15802
rect 5444 15750 13508 15802
rect 13560 15750 13572 15802
rect 13624 15750 13636 15802
rect 13688 15750 13700 15802
rect 13752 15750 13764 15802
rect 13816 15750 21880 15802
rect 21932 15750 21944 15802
rect 21996 15750 22008 15802
rect 22060 15750 22072 15802
rect 22124 15750 22136 15802
rect 22188 15750 26220 15802
rect 1104 15728 26220 15750
rect 2866 15688 2872 15700
rect 2827 15660 2872 15688
rect 2866 15648 2872 15660
rect 2924 15648 2930 15700
rect 3326 15688 3332 15700
rect 3287 15660 3332 15688
rect 3326 15648 3332 15660
rect 3384 15648 3390 15700
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 7742 15688 7748 15700
rect 7248 15660 7748 15688
rect 7248 15648 7254 15660
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 9548 15660 11345 15688
rect 9548 15648 9554 15660
rect 11333 15657 11345 15660
rect 11379 15688 11391 15691
rect 11379 15660 13032 15688
rect 11379 15657 11391 15660
rect 11333 15651 11391 15657
rect 3786 15620 3792 15632
rect 3068 15592 3792 15620
rect 3068 15493 3096 15592
rect 3786 15580 3792 15592
rect 3844 15580 3850 15632
rect 3418 15512 3424 15564
rect 3476 15552 3482 15564
rect 7101 15555 7159 15561
rect 3476 15524 3521 15552
rect 3476 15512 3482 15524
rect 7101 15521 7113 15555
rect 7147 15552 7159 15555
rect 7208 15552 7236 15648
rect 7653 15623 7711 15629
rect 7653 15589 7665 15623
rect 7699 15620 7711 15623
rect 8570 15620 8576 15632
rect 7699 15592 8576 15620
rect 7699 15589 7711 15592
rect 7653 15583 7711 15589
rect 8570 15580 8576 15592
rect 8628 15580 8634 15632
rect 12345 15623 12403 15629
rect 12345 15589 12357 15623
rect 12391 15620 12403 15623
rect 12710 15620 12716 15632
rect 12391 15592 12716 15620
rect 12391 15589 12403 15592
rect 12345 15583 12403 15589
rect 12710 15580 12716 15592
rect 12768 15620 12774 15632
rect 13004 15620 13032 15660
rect 13078 15648 13084 15700
rect 13136 15688 13142 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 13136 15660 13461 15688
rect 13136 15648 13142 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 13449 15651 13507 15657
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 15286 15688 15292 15700
rect 14783 15660 15292 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 16758 15648 16764 15700
rect 16816 15688 16822 15700
rect 16945 15691 17003 15697
rect 16945 15688 16957 15691
rect 16816 15660 16957 15688
rect 16816 15648 16822 15660
rect 16945 15657 16957 15660
rect 16991 15688 17003 15691
rect 17310 15688 17316 15700
rect 16991 15660 17316 15688
rect 16991 15657 17003 15660
rect 16945 15651 17003 15657
rect 17310 15648 17316 15660
rect 17368 15648 17374 15700
rect 17494 15648 17500 15700
rect 17552 15688 17558 15700
rect 18506 15688 18512 15700
rect 17552 15660 18091 15688
rect 18419 15660 18512 15688
rect 17552 15648 17558 15660
rect 13354 15620 13360 15632
rect 12768 15592 12848 15620
rect 13004 15592 13360 15620
rect 12768 15580 12774 15592
rect 7147 15524 7236 15552
rect 7147 15521 7159 15524
rect 7101 15515 7159 15521
rect 8018 15512 8024 15564
rect 8076 15552 8082 15564
rect 9674 15552 9680 15564
rect 8076 15524 9680 15552
rect 8076 15512 8082 15524
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 12820 15561 12848 15592
rect 13354 15580 13360 15592
rect 13412 15580 13418 15632
rect 18063 15620 18091 15660
rect 18506 15648 18512 15660
rect 18564 15688 18570 15700
rect 18874 15688 18880 15700
rect 18564 15660 18880 15688
rect 18564 15648 18570 15660
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 20346 15648 20352 15700
rect 20404 15688 20410 15700
rect 20441 15691 20499 15697
rect 20441 15688 20453 15691
rect 20404 15660 20453 15688
rect 20404 15648 20410 15660
rect 20441 15657 20453 15660
rect 20487 15657 20499 15691
rect 20441 15651 20499 15657
rect 20530 15648 20536 15700
rect 20588 15688 20594 15700
rect 21450 15688 21456 15700
rect 20588 15660 21456 15688
rect 20588 15648 20594 15660
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 22005 15691 22063 15697
rect 22005 15657 22017 15691
rect 22051 15688 22063 15691
rect 22370 15688 22376 15700
rect 22051 15660 22376 15688
rect 22051 15657 22063 15660
rect 22005 15651 22063 15657
rect 22370 15648 22376 15660
rect 22428 15648 22434 15700
rect 22833 15691 22891 15697
rect 22833 15657 22845 15691
rect 22879 15688 22891 15691
rect 23014 15688 23020 15700
rect 22879 15660 23020 15688
rect 22879 15657 22891 15660
rect 22833 15651 22891 15657
rect 23014 15648 23020 15660
rect 23072 15648 23078 15700
rect 22278 15620 22284 15632
rect 18063 15592 21404 15620
rect 9953 15555 10011 15561
rect 9953 15552 9965 15555
rect 9824 15524 9965 15552
rect 9824 15512 9830 15524
rect 9953 15521 9965 15524
rect 9999 15521 10011 15555
rect 9953 15515 10011 15521
rect 12805 15555 12863 15561
rect 12805 15521 12817 15555
rect 12851 15552 12863 15555
rect 14366 15552 14372 15564
rect 12851 15524 14372 15552
rect 12851 15521 12863 15524
rect 12805 15515 12863 15521
rect 14366 15512 14372 15524
rect 14424 15552 14430 15564
rect 14826 15552 14832 15564
rect 14424 15524 14832 15552
rect 14424 15512 14430 15524
rect 14826 15512 14832 15524
rect 14884 15512 14890 15564
rect 18230 15512 18236 15564
rect 18288 15552 18294 15564
rect 20622 15552 20628 15564
rect 18288 15524 20484 15552
rect 20583 15524 20628 15552
rect 18288 15512 18294 15524
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15453 3111 15487
rect 3053 15447 3111 15453
rect 3142 15444 3148 15496
rect 3200 15484 3206 15496
rect 3200 15456 3245 15484
rect 3200 15444 3206 15456
rect 9582 15444 9588 15496
rect 9640 15484 9646 15496
rect 10209 15487 10267 15493
rect 10209 15484 10221 15487
rect 9640 15456 10221 15484
rect 9640 15444 9646 15456
rect 10209 15453 10221 15456
rect 10255 15453 10267 15487
rect 12618 15484 12624 15496
rect 12579 15456 12624 15484
rect 10209 15447 10267 15453
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 13906 15484 13912 15496
rect 13771 15456 13912 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 14274 15444 14280 15496
rect 14332 15484 14338 15496
rect 14553 15487 14611 15493
rect 14553 15484 14565 15487
rect 14332 15456 14565 15484
rect 14332 15444 14338 15456
rect 14553 15453 14565 15456
rect 14599 15453 14611 15487
rect 14553 15447 14611 15453
rect 15565 15487 15623 15493
rect 15565 15453 15577 15487
rect 15611 15484 15623 15487
rect 16666 15484 16672 15496
rect 15611 15456 16672 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 16666 15444 16672 15456
rect 16724 15484 16730 15496
rect 17129 15487 17187 15493
rect 17129 15484 17141 15487
rect 16724 15456 17141 15484
rect 16724 15444 16730 15456
rect 17129 15453 17141 15456
rect 17175 15453 17187 15487
rect 17129 15447 17187 15453
rect 17218 15444 17224 15496
rect 17276 15484 17282 15496
rect 17385 15487 17443 15493
rect 17385 15484 17397 15487
rect 17276 15456 17397 15484
rect 17276 15444 17282 15456
rect 17385 15453 17397 15456
rect 17431 15453 17443 15487
rect 18874 15484 18880 15496
rect 18835 15456 18880 15484
rect 17385 15447 17443 15453
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 18966 15444 18972 15496
rect 19024 15484 19030 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 19024 15456 19257 15484
rect 19024 15444 19030 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 20456 15484 20484 15524
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 21177 15555 21235 15561
rect 21177 15552 21189 15555
rect 21140 15524 21189 15552
rect 21140 15512 21146 15524
rect 21177 15521 21189 15524
rect 21223 15521 21235 15555
rect 21177 15515 21235 15521
rect 20530 15484 20536 15496
rect 20456 15456 20536 15484
rect 19245 15447 19303 15453
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 20714 15444 20720 15496
rect 20772 15484 20778 15496
rect 21376 15493 21404 15592
rect 22066 15592 22284 15620
rect 22066 15552 22094 15592
rect 22278 15580 22284 15592
rect 22336 15580 22342 15632
rect 22741 15623 22799 15629
rect 22741 15589 22753 15623
rect 22787 15620 22799 15623
rect 23106 15620 23112 15632
rect 22787 15592 23112 15620
rect 22787 15589 22799 15592
rect 22741 15583 22799 15589
rect 23106 15580 23112 15592
rect 23164 15580 23170 15632
rect 21560 15524 22094 15552
rect 23124 15552 23152 15580
rect 23385 15555 23443 15561
rect 23385 15552 23397 15555
rect 23124 15524 23397 15552
rect 21560 15493 21588 15524
rect 23385 15521 23397 15524
rect 23431 15521 23443 15555
rect 23385 15515 23443 15521
rect 20993 15487 21051 15493
rect 20993 15484 21005 15487
rect 20772 15456 21005 15484
rect 20772 15444 20778 15456
rect 20993 15453 21005 15456
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 21361 15487 21419 15493
rect 21361 15453 21373 15487
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 21544 15487 21602 15493
rect 21544 15453 21556 15487
rect 21590 15453 21602 15487
rect 21544 15447 21602 15453
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15453 21695 15487
rect 21637 15447 21695 15453
rect 21729 15487 21787 15493
rect 21729 15453 21741 15487
rect 21775 15484 21787 15487
rect 21818 15484 21824 15496
rect 21775 15456 21824 15484
rect 21775 15453 21787 15456
rect 21729 15447 21787 15453
rect 7285 15419 7343 15425
rect 7285 15385 7297 15419
rect 7331 15416 7343 15419
rect 10686 15416 10692 15428
rect 7331 15388 10692 15416
rect 7331 15385 7343 15388
rect 7285 15379 7343 15385
rect 10686 15376 10692 15388
rect 10744 15416 10750 15428
rect 11146 15416 11152 15428
rect 10744 15388 11152 15416
rect 10744 15376 10750 15388
rect 11146 15376 11152 15388
rect 11204 15376 11210 15428
rect 12452 15388 13124 15416
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 7193 15351 7251 15357
rect 7193 15348 7205 15351
rect 5592 15320 7205 15348
rect 5592 15308 5598 15320
rect 7193 15317 7205 15320
rect 7239 15317 7251 15351
rect 7193 15311 7251 15317
rect 9122 15308 9128 15360
rect 9180 15348 9186 15360
rect 9861 15351 9919 15357
rect 9861 15348 9873 15351
rect 9180 15320 9873 15348
rect 9180 15308 9186 15320
rect 9861 15317 9873 15320
rect 9907 15348 9919 15351
rect 10042 15348 10048 15360
rect 9907 15320 10048 15348
rect 9907 15317 9919 15320
rect 9861 15311 9919 15317
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 12452 15357 12480 15388
rect 12437 15351 12495 15357
rect 12437 15317 12449 15351
rect 12483 15317 12495 15351
rect 12437 15311 12495 15317
rect 12802 15308 12808 15360
rect 12860 15348 12866 15360
rect 13096 15357 13124 15388
rect 13262 15376 13268 15428
rect 13320 15416 13326 15428
rect 15378 15416 15384 15428
rect 13320 15388 15384 15416
rect 13320 15376 13326 15388
rect 15378 15376 15384 15388
rect 15436 15376 15442 15428
rect 15832 15419 15890 15425
rect 15832 15385 15844 15419
rect 15878 15416 15890 15419
rect 15930 15416 15936 15428
rect 15878 15388 15936 15416
rect 15878 15385 15890 15388
rect 15832 15379 15890 15385
rect 15930 15376 15936 15388
rect 15988 15376 15994 15428
rect 18322 15376 18328 15428
rect 18380 15416 18386 15428
rect 18693 15419 18751 15425
rect 18693 15416 18705 15419
rect 18380 15388 18705 15416
rect 18380 15376 18386 15388
rect 18693 15385 18705 15388
rect 18739 15385 18751 15419
rect 19058 15416 19064 15428
rect 19019 15388 19064 15416
rect 18693 15379 18751 15385
rect 19058 15376 19064 15388
rect 19116 15376 19122 15428
rect 21266 15376 21272 15428
rect 21324 15416 21330 15428
rect 21450 15416 21456 15428
rect 21324 15388 21456 15416
rect 21324 15376 21330 15388
rect 21450 15376 21456 15388
rect 21508 15416 21514 15428
rect 21652 15416 21680 15447
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 21913 15487 21971 15493
rect 21913 15453 21925 15487
rect 21959 15484 21971 15487
rect 23474 15484 23480 15496
rect 21959 15456 23480 15484
rect 21959 15453 21971 15456
rect 21913 15447 21971 15453
rect 23474 15444 23480 15456
rect 23532 15444 23538 15496
rect 21508 15388 21680 15416
rect 21508 15376 21514 15388
rect 12989 15351 13047 15357
rect 12989 15348 13001 15351
rect 12860 15320 13001 15348
rect 12860 15308 12866 15320
rect 12989 15317 13001 15320
rect 13035 15317 13047 15351
rect 12989 15311 13047 15317
rect 13081 15351 13139 15357
rect 13081 15317 13093 15351
rect 13127 15348 13139 15351
rect 13170 15348 13176 15360
rect 13127 15320 13176 15348
rect 13127 15317 13139 15320
rect 13081 15311 13139 15317
rect 13170 15308 13176 15320
rect 13228 15308 13234 15360
rect 13541 15351 13599 15357
rect 13541 15317 13553 15351
rect 13587 15348 13599 15351
rect 14182 15348 14188 15360
rect 13587 15320 14188 15348
rect 13587 15317 13599 15320
rect 13541 15311 13599 15317
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 18598 15308 18604 15360
rect 18656 15348 18662 15360
rect 19429 15351 19487 15357
rect 19429 15348 19441 15351
rect 18656 15320 19441 15348
rect 18656 15308 18662 15320
rect 19429 15317 19441 15320
rect 19475 15317 19487 15351
rect 19429 15311 19487 15317
rect 20993 15351 21051 15357
rect 20993 15317 21005 15351
rect 21039 15348 21051 15351
rect 21358 15348 21364 15360
rect 21039 15320 21364 15348
rect 21039 15317 21051 15320
rect 20993 15311 21051 15317
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 23198 15348 23204 15360
rect 23159 15320 23204 15348
rect 23198 15308 23204 15320
rect 23256 15308 23262 15360
rect 23290 15308 23296 15360
rect 23348 15348 23354 15360
rect 23348 15320 23393 15348
rect 23348 15308 23354 15320
rect 1104 15258 26220 15280
rect 1104 15206 9322 15258
rect 9374 15206 9386 15258
rect 9438 15206 9450 15258
rect 9502 15206 9514 15258
rect 9566 15206 9578 15258
rect 9630 15206 17694 15258
rect 17746 15206 17758 15258
rect 17810 15206 17822 15258
rect 17874 15206 17886 15258
rect 17938 15206 17950 15258
rect 18002 15206 26220 15258
rect 26326 15212 26332 15224
rect 1104 15184 26220 15206
rect 26287 15184 26332 15212
rect 26326 15172 26332 15184
rect 26384 15172 26390 15224
rect 4890 15104 4896 15156
rect 4948 15144 4954 15156
rect 7285 15147 7343 15153
rect 4948 15116 6316 15144
rect 4948 15104 4954 15116
rect 5534 15076 5540 15088
rect 4264 15048 5540 15076
rect 4264 15017 4292 15048
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 14977 4307 15011
rect 4618 15011 4676 15017
rect 4618 15008 4630 15011
rect 4249 14971 4307 14977
rect 4356 14980 4630 15008
rect 2866 14900 2872 14952
rect 2924 14940 2930 14952
rect 4356 14940 4384 14980
rect 4618 14977 4630 14980
rect 4664 14977 4676 15011
rect 4618 14971 4676 14977
rect 4706 14968 4712 15020
rect 4764 15008 4770 15020
rect 4801 15011 4859 15017
rect 4801 15008 4813 15011
rect 4764 14980 4813 15008
rect 4764 14968 4770 14980
rect 4801 14977 4813 14980
rect 4847 14977 4859 15011
rect 4801 14971 4859 14977
rect 5077 15011 5135 15017
rect 5077 14977 5089 15011
rect 5123 15008 5135 15011
rect 5626 15008 5632 15020
rect 5123 14980 5632 15008
rect 5123 14977 5135 14980
rect 5077 14971 5135 14977
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 6288 15008 6316 15116
rect 7285 15113 7297 15147
rect 7331 15113 7343 15147
rect 7285 15107 7343 15113
rect 7653 15147 7711 15153
rect 7653 15113 7665 15147
rect 7699 15144 7711 15147
rect 9858 15144 9864 15156
rect 7699 15116 9864 15144
rect 7699 15113 7711 15116
rect 7653 15107 7711 15113
rect 7300 15076 7328 15107
rect 9858 15104 9864 15116
rect 9916 15144 9922 15156
rect 10594 15144 10600 15156
rect 9916 15116 10600 15144
rect 9916 15104 9922 15116
rect 10594 15104 10600 15116
rect 10652 15104 10658 15156
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12713 15147 12771 15153
rect 12713 15144 12725 15147
rect 12676 15116 12725 15144
rect 12676 15104 12682 15116
rect 12713 15113 12725 15116
rect 12759 15113 12771 15147
rect 12713 15107 12771 15113
rect 18141 15147 18199 15153
rect 18141 15113 18153 15147
rect 18187 15144 18199 15147
rect 18874 15144 18880 15156
rect 18187 15116 18880 15144
rect 18187 15113 18199 15116
rect 18141 15107 18199 15113
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 18969 15147 19027 15153
rect 18969 15113 18981 15147
rect 19015 15144 19027 15147
rect 19334 15144 19340 15156
rect 19015 15116 19340 15144
rect 19015 15113 19027 15116
rect 18969 15107 19027 15113
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 23290 15144 23296 15156
rect 23251 15116 23296 15144
rect 23290 15104 23296 15116
rect 23348 15104 23354 15156
rect 23382 15104 23388 15156
rect 23440 15144 23446 15156
rect 23661 15147 23719 15153
rect 23661 15144 23673 15147
rect 23440 15116 23673 15144
rect 23440 15104 23446 15116
rect 23661 15113 23673 15116
rect 23707 15113 23719 15147
rect 23661 15107 23719 15113
rect 7116 15048 7328 15076
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 6288 14980 6653 15008
rect 6641 14977 6653 14980
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 7027 15011 7085 15017
rect 7027 14977 7039 15011
rect 7073 15008 7085 15011
rect 7116 15008 7144 15048
rect 7742 15036 7748 15088
rect 7800 15076 7806 15088
rect 8113 15079 8171 15085
rect 8113 15076 8125 15079
rect 7800 15048 8125 15076
rect 7800 15036 7806 15048
rect 7073 14980 7144 15008
rect 7193 15011 7251 15017
rect 7073 14977 7085 14980
rect 7027 14971 7085 14977
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7374 15008 7380 15020
rect 7239 14980 7380 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 2924 14912 4384 14940
rect 4433 14943 4491 14949
rect 2924 14900 2930 14912
rect 4433 14909 4445 14943
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 5810 14940 5816 14952
rect 4571 14912 5816 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 4338 14832 4344 14884
rect 4396 14872 4402 14884
rect 4448 14872 4476 14903
rect 5810 14900 5816 14912
rect 5868 14900 5874 14952
rect 6457 14943 6515 14949
rect 6457 14909 6469 14943
rect 6503 14940 6515 14943
rect 6546 14940 6552 14952
rect 6503 14912 6552 14940
rect 6503 14909 6515 14912
rect 6457 14903 6515 14909
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14940 6975 14943
rect 7282 14940 7288 14952
rect 6963 14912 7288 14940
rect 6963 14909 6975 14912
rect 6917 14903 6975 14909
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 7944 14949 7972 15048
rect 8113 15045 8125 15048
rect 8159 15076 8171 15079
rect 8662 15076 8668 15088
rect 8159 15048 8668 15076
rect 8159 15045 8171 15048
rect 8113 15039 8171 15045
rect 8662 15036 8668 15048
rect 8720 15036 8726 15088
rect 8846 15036 8852 15088
rect 8904 15076 8910 15088
rect 9490 15076 9496 15088
rect 8904 15048 9496 15076
rect 8904 15036 8910 15048
rect 9490 15036 9496 15048
rect 9548 15076 9554 15088
rect 18046 15076 18052 15088
rect 9548 15048 9812 15076
rect 9548 15036 9554 15048
rect 9674 15008 9680 15020
rect 9635 14980 9680 15008
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 9784 15008 9812 15048
rect 14936 15048 18052 15076
rect 9842 15011 9900 15017
rect 9842 15008 9854 15011
rect 9784 14980 9854 15008
rect 9842 14977 9854 14980
rect 9888 14977 9900 15011
rect 9842 14971 9900 14977
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 10134 15008 10140 15020
rect 10091 14980 10140 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 10134 14968 10140 14980
rect 10192 14968 10198 15020
rect 10226 14968 10232 15020
rect 10284 15008 10290 15020
rect 10686 15008 10692 15020
rect 10284 14980 10329 15008
rect 10647 14980 10692 15008
rect 10284 14968 10290 14980
rect 10686 14968 10692 14980
rect 10744 15008 10750 15020
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 10744 14980 12173 15008
rect 10744 14968 10750 14980
rect 12161 14977 12173 14980
rect 12207 15008 12219 15011
rect 12342 15008 12348 15020
rect 12207 14980 12348 15008
rect 12207 14977 12219 14980
rect 12161 14971 12219 14977
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 12620 15011 12678 15017
rect 12620 14977 12632 15011
rect 12666 15008 12678 15011
rect 12710 15008 12716 15020
rect 12666 14980 12716 15008
rect 12666 14977 12678 14980
rect 12620 14971 12678 14977
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 12897 15011 12955 15017
rect 12897 14977 12909 15011
rect 12943 14977 12955 15011
rect 12897 14971 12955 14977
rect 7745 14943 7803 14949
rect 7745 14909 7757 14943
rect 7791 14909 7803 14943
rect 7745 14903 7803 14909
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14909 7987 14943
rect 7929 14903 7987 14909
rect 4396 14844 4476 14872
rect 4396 14832 4402 14844
rect 4798 14832 4804 14884
rect 4856 14872 4862 14884
rect 7760 14872 7788 14903
rect 9214 14900 9220 14952
rect 9272 14940 9278 14952
rect 9953 14943 10011 14949
rect 9953 14940 9965 14943
rect 9272 14912 9965 14940
rect 9272 14900 9278 14912
rect 9953 14909 9965 14912
rect 9999 14909 10011 14943
rect 9953 14903 10011 14909
rect 10594 14900 10600 14952
rect 10652 14940 10658 14952
rect 12253 14943 12311 14949
rect 12253 14940 12265 14943
rect 10652 14912 12265 14940
rect 10652 14900 10658 14912
rect 12253 14909 12265 14912
rect 12299 14940 12311 14943
rect 12802 14940 12808 14952
rect 12299 14912 12808 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 11422 14872 11428 14884
rect 4856 14844 7788 14872
rect 8128 14844 11428 14872
rect 4856 14832 4862 14844
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 4157 14807 4215 14813
rect 4157 14804 4169 14807
rect 4120 14776 4169 14804
rect 4120 14764 4126 14776
rect 4157 14773 4169 14776
rect 4203 14773 4215 14807
rect 4157 14767 4215 14773
rect 4706 14764 4712 14816
rect 4764 14804 4770 14816
rect 4893 14807 4951 14813
rect 4893 14804 4905 14807
rect 4764 14776 4905 14804
rect 4764 14764 4770 14776
rect 4893 14773 4905 14776
rect 4939 14804 4951 14807
rect 8128 14804 8156 14844
rect 11422 14832 11428 14844
rect 11480 14832 11486 14884
rect 12912 14872 12940 14971
rect 14936 14952 14964 15048
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 21266 15076 21272 15088
rect 19812 15048 21272 15076
rect 15102 15008 15108 15020
rect 15063 14980 15108 15008
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 18322 15017 18328 15020
rect 16761 15011 16819 15017
rect 16761 15008 16773 15011
rect 16632 14980 16773 15008
rect 16632 14968 16638 14980
rect 16761 14977 16773 14980
rect 16807 14977 16819 15011
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 16761 14971 16819 14977
rect 16868 14980 17049 15008
rect 13998 14900 14004 14952
rect 14056 14940 14062 14952
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 14056 14912 14657 14940
rect 14056 14900 14062 14912
rect 14645 14909 14657 14912
rect 14691 14940 14703 14943
rect 14918 14940 14924 14952
rect 14691 14912 14924 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 14918 14900 14924 14912
rect 14976 14900 14982 14952
rect 15194 14940 15200 14952
rect 15155 14912 15200 14940
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14909 15347 14943
rect 15289 14903 15347 14909
rect 12084 14844 12940 14872
rect 12084 14816 12112 14844
rect 9490 14804 9496 14816
rect 4939 14776 8156 14804
rect 9451 14776 9496 14804
rect 4939 14773 4951 14776
rect 4893 14767 4951 14773
rect 9490 14764 9496 14776
rect 9548 14764 9554 14816
rect 10318 14804 10324 14816
rect 10279 14776 10324 14804
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 10505 14807 10563 14813
rect 10505 14773 10517 14807
rect 10551 14804 10563 14807
rect 10594 14804 10600 14816
rect 10551 14776 10600 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 12066 14804 12072 14816
rect 12027 14776 12072 14804
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 14458 14764 14464 14816
rect 14516 14804 14522 14816
rect 14737 14807 14795 14813
rect 14737 14804 14749 14807
rect 14516 14776 14749 14804
rect 14516 14764 14522 14776
rect 14737 14773 14749 14776
rect 14783 14773 14795 14807
rect 14737 14767 14795 14773
rect 14826 14764 14832 14816
rect 14884 14804 14890 14816
rect 15304 14804 15332 14903
rect 15746 14900 15752 14952
rect 15804 14940 15810 14952
rect 16868 14940 16896 14980
rect 17037 14977 17049 14980
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 18291 15011 18328 15017
rect 18291 14977 18303 15011
rect 18291 14971 18328 14977
rect 18322 14968 18328 14971
rect 18380 14968 18386 15020
rect 18506 14968 18512 15020
rect 18564 15008 18570 15020
rect 18601 15011 18659 15017
rect 18601 15008 18613 15011
rect 18564 14980 18613 15008
rect 18564 14968 18570 14980
rect 18601 14977 18613 14980
rect 18647 14977 18659 15011
rect 18782 15008 18788 15020
rect 18743 14980 18788 15008
rect 18601 14971 18659 14977
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 17494 14940 17500 14952
rect 15804 14912 16896 14940
rect 16960 14912 17500 14940
rect 15804 14900 15810 14912
rect 16960 14881 16988 14912
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14940 18751 14943
rect 19058 14940 19064 14952
rect 18739 14912 19064 14940
rect 18739 14909 18751 14912
rect 18693 14903 18751 14909
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 16945 14875 17003 14881
rect 16945 14841 16957 14875
rect 16991 14841 17003 14875
rect 19812 14872 19840 15048
rect 20898 15008 20904 15020
rect 20859 14980 20904 15008
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 21192 15017 21220 15048
rect 21266 15036 21272 15048
rect 21324 15036 21330 15088
rect 21637 15079 21695 15085
rect 21637 15045 21649 15079
rect 21683 15076 21695 15079
rect 22158 15079 22216 15085
rect 22158 15076 22170 15079
rect 21683 15048 22170 15076
rect 21683 15045 21695 15048
rect 21637 15039 21695 15045
rect 22158 15045 22170 15048
rect 22204 15045 22216 15079
rect 22158 15039 22216 15045
rect 21066 15011 21124 15017
rect 21066 15008 21078 15011
rect 21008 14980 21078 15008
rect 16945 14835 17003 14841
rect 17420 14844 19840 14872
rect 17420 14816 17448 14844
rect 14884 14776 15332 14804
rect 17221 14807 17279 14813
rect 14884 14764 14890 14776
rect 17221 14773 17233 14807
rect 17267 14804 17279 14807
rect 17402 14804 17408 14816
rect 17267 14776 17408 14804
rect 17267 14773 17279 14776
rect 17221 14767 17279 14773
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 19150 14764 19156 14816
rect 19208 14804 19214 14816
rect 20717 14807 20775 14813
rect 20717 14804 20729 14807
rect 19208 14776 20729 14804
rect 19208 14764 19214 14776
rect 20717 14773 20729 14776
rect 20763 14804 20775 14807
rect 21008 14804 21036 14980
rect 21066 14977 21078 14980
rect 21112 14977 21124 15011
rect 21066 14971 21124 14977
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 14977 21235 15011
rect 21177 14971 21235 14977
rect 21453 15011 21511 15017
rect 21453 14977 21465 15011
rect 21499 14977 21511 15011
rect 21453 14971 21511 14977
rect 21266 14900 21272 14952
rect 21324 14940 21330 14952
rect 21324 14912 21369 14940
rect 21324 14900 21330 14912
rect 21468 14872 21496 14971
rect 21726 14968 21732 15020
rect 21784 15008 21790 15020
rect 21913 15011 21971 15017
rect 21913 15008 21925 15011
rect 21784 14980 21925 15008
rect 21784 14968 21790 14980
rect 21913 14977 21925 14980
rect 21959 14977 21971 15011
rect 23308 15008 23336 15104
rect 23477 15011 23535 15017
rect 23477 15008 23489 15011
rect 23308 14980 23489 15008
rect 21913 14971 21971 14977
rect 23477 14977 23489 14980
rect 23523 14977 23535 15011
rect 23477 14971 23535 14977
rect 21468 14844 21772 14872
rect 20763 14776 21036 14804
rect 21744 14804 21772 14844
rect 23382 14804 23388 14816
rect 21744 14776 23388 14804
rect 20763 14773 20775 14776
rect 20717 14767 20775 14773
rect 23382 14764 23388 14776
rect 23440 14764 23446 14816
rect 1104 14714 26220 14736
rect 1104 14662 5136 14714
rect 5188 14662 5200 14714
rect 5252 14662 5264 14714
rect 5316 14662 5328 14714
rect 5380 14662 5392 14714
rect 5444 14662 13508 14714
rect 13560 14662 13572 14714
rect 13624 14662 13636 14714
rect 13688 14662 13700 14714
rect 13752 14662 13764 14714
rect 13816 14662 21880 14714
rect 21932 14662 21944 14714
rect 21996 14662 22008 14714
rect 22060 14662 22072 14714
rect 22124 14662 22136 14714
rect 22188 14662 26220 14714
rect 1104 14640 26220 14662
rect 5169 14603 5227 14609
rect 5169 14569 5181 14603
rect 5215 14600 5227 14603
rect 5534 14600 5540 14612
rect 5215 14572 5540 14600
rect 5215 14569 5227 14572
rect 5169 14563 5227 14569
rect 5534 14560 5540 14572
rect 5592 14560 5598 14612
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 8478 14600 8484 14612
rect 7423 14572 8484 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 9732 14572 12265 14600
rect 9732 14560 9738 14572
rect 12253 14569 12265 14572
rect 12299 14569 12311 14603
rect 12253 14563 12311 14569
rect 12710 14560 12716 14612
rect 12768 14600 12774 14612
rect 12897 14603 12955 14609
rect 12897 14600 12909 14603
rect 12768 14572 12909 14600
rect 12768 14560 12774 14572
rect 12897 14569 12909 14572
rect 12943 14569 12955 14603
rect 13078 14600 13084 14612
rect 13039 14572 13084 14600
rect 12897 14563 12955 14569
rect 4890 14492 4896 14544
rect 4948 14532 4954 14544
rect 5445 14535 5503 14541
rect 5445 14532 5457 14535
rect 4948 14504 5457 14532
rect 4948 14492 4954 14504
rect 5445 14501 5457 14504
rect 5491 14501 5503 14535
rect 5445 14495 5503 14501
rect 10318 14424 10324 14476
rect 10376 14464 10382 14476
rect 12912 14464 12940 14563
rect 13078 14560 13084 14572
rect 13136 14600 13142 14612
rect 14366 14600 14372 14612
rect 13136 14572 14372 14600
rect 13136 14560 13142 14572
rect 13906 14532 13912 14544
rect 13867 14504 13912 14532
rect 13906 14492 13912 14504
rect 13964 14492 13970 14544
rect 13265 14467 13323 14473
rect 13265 14464 13277 14467
rect 10376 14436 10548 14464
rect 12912 14436 13277 14464
rect 10376 14424 10382 14436
rect 3418 14356 3424 14408
rect 3476 14396 3482 14408
rect 4062 14405 4068 14408
rect 3789 14399 3847 14405
rect 3789 14396 3801 14399
rect 3476 14368 3801 14396
rect 3476 14356 3482 14368
rect 3789 14365 3801 14368
rect 3835 14365 3847 14399
rect 4056 14396 4068 14405
rect 4023 14368 4068 14396
rect 3789 14359 3847 14365
rect 4056 14359 4068 14368
rect 4062 14356 4068 14359
rect 4120 14356 4126 14408
rect 6546 14356 6552 14408
rect 6604 14405 6610 14408
rect 6604 14396 6616 14405
rect 6825 14399 6883 14405
rect 6604 14368 6649 14396
rect 6604 14359 6616 14368
rect 6825 14365 6837 14399
rect 6871 14396 6883 14399
rect 7926 14396 7932 14408
rect 6871 14368 7932 14396
rect 6871 14365 6883 14368
rect 6825 14359 6883 14365
rect 6604 14356 6610 14359
rect 7926 14356 7932 14368
rect 7984 14396 7990 14408
rect 8757 14399 8815 14405
rect 8757 14396 8769 14399
rect 7984 14368 8769 14396
rect 7984 14356 7990 14368
rect 8757 14365 8769 14368
rect 8803 14396 8815 14399
rect 9214 14396 9220 14408
rect 8803 14368 9220 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 9214 14356 9220 14368
rect 9272 14396 9278 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 9272 14368 10425 14396
rect 9272 14356 9278 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10520 14396 10548 14436
rect 13265 14433 13277 14436
rect 13311 14464 13323 14467
rect 13814 14464 13820 14476
rect 13311 14436 13820 14464
rect 13311 14433 13323 14436
rect 13265 14427 13323 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 14199 14473 14227 14572
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 14734 14560 14740 14612
rect 14792 14600 14798 14612
rect 14829 14603 14887 14609
rect 14829 14600 14841 14603
rect 14792 14572 14841 14600
rect 14792 14560 14798 14572
rect 14829 14569 14841 14572
rect 14875 14569 14887 14603
rect 14829 14563 14887 14569
rect 17494 14560 17500 14612
rect 17552 14600 17558 14612
rect 21266 14600 21272 14612
rect 17552 14572 21272 14600
rect 17552 14560 17558 14572
rect 21266 14560 21272 14572
rect 21324 14600 21330 14612
rect 21726 14600 21732 14612
rect 21324 14572 21732 14600
rect 21324 14560 21330 14572
rect 21726 14560 21732 14572
rect 21784 14560 21790 14612
rect 14642 14492 14648 14544
rect 14700 14532 14706 14544
rect 19334 14532 19340 14544
rect 14700 14504 19340 14532
rect 14700 14492 14706 14504
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 20625 14535 20683 14541
rect 20625 14501 20637 14535
rect 20671 14532 20683 14535
rect 22370 14532 22376 14544
rect 20671 14504 22376 14532
rect 20671 14501 20683 14504
rect 20625 14495 20683 14501
rect 22370 14492 22376 14504
rect 22428 14532 22434 14544
rect 22830 14532 22836 14544
rect 22428 14504 22836 14532
rect 22428 14492 22434 14504
rect 22830 14492 22836 14504
rect 22888 14492 22894 14544
rect 14185 14467 14243 14473
rect 14185 14433 14197 14467
rect 14231 14433 14243 14467
rect 14369 14467 14427 14473
rect 14369 14464 14381 14467
rect 14185 14427 14243 14433
rect 14292 14436 14381 14464
rect 10669 14399 10727 14405
rect 10669 14396 10681 14399
rect 10520 14368 10681 14396
rect 10413 14359 10471 14365
rect 10669 14365 10681 14368
rect 10715 14365 10727 14399
rect 12158 14396 12164 14408
rect 12119 14368 12164 14396
rect 10669 14359 10727 14365
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 12437 14399 12495 14405
rect 12437 14365 12449 14399
rect 12483 14396 12495 14399
rect 12526 14396 12532 14408
rect 12483 14368 12532 14396
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 12802 14396 12808 14408
rect 12763 14368 12808 14396
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 13354 14396 13360 14408
rect 13315 14368 13360 14396
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 13446 14356 13452 14408
rect 13504 14396 13510 14408
rect 13667 14399 13725 14405
rect 13667 14396 13679 14399
rect 13504 14368 13679 14396
rect 13504 14356 13510 14368
rect 13667 14365 13679 14368
rect 13713 14365 13725 14399
rect 13667 14359 13725 14365
rect 13998 14356 14004 14408
rect 14056 14396 14062 14408
rect 14292 14396 14320 14436
rect 14369 14433 14381 14436
rect 14415 14464 14427 14467
rect 15102 14464 15108 14476
rect 14415 14436 15108 14464
rect 14415 14433 14427 14436
rect 14369 14427 14427 14433
rect 15102 14424 15108 14436
rect 15160 14424 15166 14476
rect 14458 14396 14464 14408
rect 14056 14368 14320 14396
rect 14419 14368 14464 14396
rect 14056 14356 14062 14368
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 14826 14356 14832 14408
rect 14884 14396 14890 14408
rect 18138 14396 18144 14408
rect 14884 14368 18144 14396
rect 14884 14356 14890 14368
rect 15120 14340 15148 14368
rect 18138 14356 18144 14368
rect 18196 14356 18202 14408
rect 19352 14396 19380 14492
rect 23106 14464 23112 14476
rect 22572 14436 23112 14464
rect 20441 14399 20499 14405
rect 20441 14396 20453 14399
rect 19352 14368 20453 14396
rect 20441 14365 20453 14368
rect 20487 14365 20499 14399
rect 20441 14359 20499 14365
rect 21082 14356 21088 14408
rect 21140 14396 21146 14408
rect 21910 14396 21916 14408
rect 21140 14368 21916 14396
rect 21140 14356 21146 14368
rect 21910 14356 21916 14368
rect 21968 14396 21974 14408
rect 22572 14405 22600 14436
rect 23106 14424 23112 14436
rect 23164 14424 23170 14476
rect 22189 14399 22247 14405
rect 22189 14396 22201 14399
rect 21968 14368 22201 14396
rect 21968 14356 21974 14368
rect 22189 14365 22201 14368
rect 22235 14365 22247 14399
rect 22189 14359 22247 14365
rect 22557 14399 22615 14405
rect 22557 14365 22569 14399
rect 22603 14365 22615 14399
rect 22557 14359 22615 14365
rect 22741 14399 22799 14405
rect 22741 14365 22753 14399
rect 22787 14396 22799 14399
rect 23385 14399 23443 14405
rect 23385 14396 23397 14399
rect 22787 14368 23397 14396
rect 22787 14365 22799 14368
rect 22741 14359 22799 14365
rect 23385 14365 23397 14368
rect 23431 14365 23443 14399
rect 23385 14359 23443 14365
rect 23474 14356 23480 14408
rect 23532 14396 23538 14408
rect 23532 14368 23577 14396
rect 23532 14356 23538 14368
rect 7282 14288 7288 14340
rect 7340 14328 7346 14340
rect 8202 14328 8208 14340
rect 7340 14300 8208 14328
rect 7340 14288 7346 14300
rect 8202 14288 8208 14300
rect 8260 14288 8266 14340
rect 8294 14288 8300 14340
rect 8352 14328 8358 14340
rect 8490 14331 8548 14337
rect 8490 14328 8502 14331
rect 8352 14300 8502 14328
rect 8352 14288 8358 14300
rect 8490 14297 8502 14300
rect 8536 14297 8548 14331
rect 8490 14291 8548 14297
rect 11808 14300 12296 14328
rect 10226 14220 10232 14272
rect 10284 14260 10290 14272
rect 11808 14269 11836 14300
rect 11793 14263 11851 14269
rect 11793 14260 11805 14263
rect 10284 14232 11805 14260
rect 10284 14220 10290 14232
rect 11793 14229 11805 14232
rect 11839 14229 11851 14263
rect 11793 14223 11851 14229
rect 11977 14263 12035 14269
rect 11977 14229 11989 14263
rect 12023 14260 12035 14263
rect 12066 14260 12072 14272
rect 12023 14232 12072 14260
rect 12023 14229 12035 14232
rect 11977 14223 12035 14229
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 12268 14260 12296 14300
rect 12342 14288 12348 14340
rect 12400 14328 12406 14340
rect 12621 14331 12679 14337
rect 12621 14328 12633 14331
rect 12400 14300 12633 14328
rect 12400 14288 12406 14300
rect 12621 14297 12633 14300
rect 12667 14297 12679 14331
rect 12621 14291 12679 14297
rect 15102 14288 15108 14340
rect 15160 14288 15166 14340
rect 22281 14331 22339 14337
rect 22281 14297 22293 14331
rect 22327 14328 22339 14331
rect 22462 14328 22468 14340
rect 22327 14300 22468 14328
rect 22327 14297 22339 14300
rect 22281 14291 22339 14297
rect 22462 14288 22468 14300
rect 22520 14288 22526 14340
rect 22833 14331 22891 14337
rect 22833 14297 22845 14331
rect 22879 14297 22891 14331
rect 22833 14291 22891 14297
rect 23017 14331 23075 14337
rect 23017 14297 23029 14331
rect 23063 14297 23075 14331
rect 23017 14291 23075 14297
rect 23201 14331 23259 14337
rect 23201 14297 23213 14331
rect 23247 14328 23259 14331
rect 23290 14328 23296 14340
rect 23247 14300 23296 14328
rect 23247 14297 23259 14300
rect 23201 14291 23259 14297
rect 14458 14260 14464 14272
rect 12268 14232 14464 14260
rect 14458 14220 14464 14232
rect 14516 14260 14522 14272
rect 14826 14260 14832 14272
rect 14516 14232 14832 14260
rect 14516 14220 14522 14232
rect 14826 14220 14832 14232
rect 14884 14260 14890 14272
rect 15194 14260 15200 14272
rect 14884 14232 15200 14260
rect 14884 14220 14890 14232
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 19981 14263 20039 14269
rect 19981 14229 19993 14263
rect 20027 14260 20039 14263
rect 20162 14260 20168 14272
rect 20027 14232 20168 14260
rect 20027 14229 20039 14232
rect 19981 14223 20039 14229
rect 20162 14220 20168 14232
rect 20220 14220 20226 14272
rect 22002 14220 22008 14272
rect 22060 14260 22066 14272
rect 22848 14260 22876 14291
rect 22060 14232 22876 14260
rect 23032 14260 23060 14291
rect 23290 14288 23296 14300
rect 23348 14288 23354 14340
rect 23492 14260 23520 14356
rect 23032 14232 23520 14260
rect 22060 14220 22066 14232
rect 1104 14170 26220 14192
rect 1104 14118 9322 14170
rect 9374 14118 9386 14170
rect 9438 14118 9450 14170
rect 9502 14118 9514 14170
rect 9566 14118 9578 14170
rect 9630 14118 17694 14170
rect 17746 14118 17758 14170
rect 17810 14118 17822 14170
rect 17874 14118 17886 14170
rect 17938 14118 17950 14170
rect 18002 14118 26220 14170
rect 1104 14096 26220 14118
rect 2866 14056 2872 14068
rect 2827 14028 2872 14056
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 4798 14056 4804 14068
rect 4759 14028 4804 14056
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 8389 14059 8447 14065
rect 8389 14056 8401 14059
rect 7336 14028 8401 14056
rect 1504 13960 3464 13988
rect 1504 13864 1532 13960
rect 3436 13932 3464 13960
rect 6822 13948 6828 14000
rect 6880 13988 6886 14000
rect 6880 13960 7144 13988
rect 6880 13948 6886 13960
rect 1756 13923 1814 13929
rect 1756 13889 1768 13923
rect 1802 13920 1814 13923
rect 2314 13920 2320 13932
rect 1802 13892 2320 13920
rect 1802 13889 1814 13892
rect 1756 13883 1814 13889
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 3418 13920 3424 13932
rect 3331 13892 3424 13920
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 3688 13923 3746 13929
rect 3688 13889 3700 13923
rect 3734 13920 3746 13923
rect 4430 13920 4436 13932
rect 3734 13892 4436 13920
rect 3734 13889 3746 13892
rect 3688 13883 3746 13889
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 6914 13920 6920 13932
rect 6875 13892 6920 13920
rect 6914 13880 6920 13892
rect 6972 13880 6978 13932
rect 7116 13929 7144 13960
rect 7336 13932 7364 14028
rect 8389 14025 8401 14028
rect 8435 14025 8447 14059
rect 8389 14019 8447 14025
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 9493 14059 9551 14065
rect 9493 14056 9505 14059
rect 8720 14028 9505 14056
rect 8720 14016 8726 14028
rect 8294 13988 8300 14000
rect 8255 13960 8300 13988
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 8478 13948 8484 14000
rect 8536 13948 8542 14000
rect 8754 13988 8760 14000
rect 8715 13960 8760 13988
rect 8754 13948 8760 13960
rect 8812 13948 8818 14000
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7321 13926 7379 13932
rect 7248 13892 7293 13920
rect 7321 13892 7333 13926
rect 7367 13892 7379 13926
rect 7248 13880 7254 13892
rect 7321 13886 7379 13892
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 7561 13923 7619 13929
rect 7561 13920 7573 13923
rect 7515 13892 7573 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7561 13889 7573 13892
rect 7607 13889 7619 13923
rect 7561 13883 7619 13889
rect 1486 13852 1492 13864
rect 1447 13824 1492 13852
rect 1486 13812 1492 13824
rect 1544 13812 1550 13864
rect 6733 13855 6791 13861
rect 6733 13821 6745 13855
rect 6779 13852 6791 13855
rect 7006 13852 7012 13864
rect 6779 13824 7012 13852
rect 6779 13821 6791 13824
rect 6733 13815 6791 13821
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7374 13676 7380 13728
rect 7432 13716 7438 13728
rect 7484 13716 7512 13883
rect 7742 13880 7748 13932
rect 7800 13920 7806 13932
rect 7929 13923 7987 13929
rect 7800 13892 7844 13920
rect 7800 13880 7806 13892
rect 7929 13889 7941 13923
rect 7975 13920 7987 13923
rect 8018 13920 8024 13932
rect 7975 13892 8024 13920
rect 7975 13889 7987 13892
rect 7929 13883 7987 13889
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 8113 13923 8171 13929
rect 8113 13889 8125 13923
rect 8159 13920 8171 13923
rect 8496 13920 8524 13948
rect 8159 13892 8524 13920
rect 8159 13889 8171 13892
rect 8113 13883 8171 13889
rect 8956 13864 8984 14028
rect 9493 14025 9505 14028
rect 9539 14025 9551 14059
rect 13173 14059 13231 14065
rect 13173 14056 13185 14059
rect 9493 14019 9551 14025
rect 12406 14028 13185 14056
rect 9306 13948 9312 14000
rect 9364 13988 9370 14000
rect 12406 13988 12434 14028
rect 13173 14025 13185 14028
rect 13219 14025 13231 14059
rect 14274 14056 14280 14068
rect 13173 14019 13231 14025
rect 13280 14028 14280 14056
rect 13280 13988 13308 14028
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 16117 14059 16175 14065
rect 16117 14056 16129 14059
rect 14424 14028 16129 14056
rect 14424 14016 14430 14028
rect 16117 14025 16129 14028
rect 16163 14056 16175 14059
rect 16850 14056 16856 14068
rect 16163 14028 16856 14056
rect 16163 14025 16175 14028
rect 16117 14019 16175 14025
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 17221 14059 17279 14065
rect 17221 14025 17233 14059
rect 17267 14056 17279 14059
rect 18138 14056 18144 14068
rect 17267 14028 18144 14056
rect 17267 14025 17279 14028
rect 17221 14019 17279 14025
rect 18138 14016 18144 14028
rect 18196 14056 18202 14068
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 18196 14028 19073 14056
rect 18196 14016 18202 14028
rect 19061 14025 19073 14028
rect 19107 14056 19119 14059
rect 19242 14056 19248 14068
rect 19107 14028 19248 14056
rect 19107 14025 19119 14028
rect 19061 14019 19119 14025
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 19610 14056 19616 14068
rect 19571 14028 19616 14056
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 19978 14056 19984 14068
rect 19939 14028 19984 14056
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20806 14056 20812 14068
rect 20767 14028 20812 14056
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 21910 14016 21916 14068
rect 21968 14056 21974 14068
rect 22281 14059 22339 14065
rect 22281 14056 22293 14059
rect 21968 14028 22293 14056
rect 21968 14016 21974 14028
rect 22281 14025 22293 14028
rect 22327 14025 22339 14059
rect 22281 14019 22339 14025
rect 13446 13988 13452 14000
rect 9364 13960 12434 13988
rect 12728 13960 13308 13988
rect 13407 13960 13452 13988
rect 9364 13948 9370 13960
rect 9030 13880 9036 13932
rect 9088 13920 9094 13932
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 9088 13892 9413 13920
rect 9088 13880 9094 13892
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13920 11759 13923
rect 12250 13920 12256 13932
rect 11747 13892 12256 13920
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 12250 13880 12256 13892
rect 12308 13880 12314 13932
rect 12618 13880 12624 13932
rect 12676 13920 12682 13932
rect 12728 13929 12756 13960
rect 13446 13948 13452 13960
rect 13504 13988 13510 14000
rect 14645 13991 14703 13997
rect 14645 13988 14657 13991
rect 13504 13960 14657 13988
rect 13504 13948 13510 13960
rect 12713 13923 12771 13929
rect 12713 13920 12725 13923
rect 12676 13892 12725 13920
rect 12676 13880 12682 13892
rect 12713 13889 12725 13892
rect 12759 13889 12771 13923
rect 12713 13883 12771 13889
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8202 13852 8208 13864
rect 7883 13824 8208 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8536 13824 8861 13852
rect 8536 13812 8542 13824
rect 8849 13821 8861 13824
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 8938 13812 8944 13864
rect 8996 13852 9002 13864
rect 13372 13852 13400 13883
rect 13538 13880 13544 13932
rect 13596 13920 13602 13932
rect 13633 13923 13691 13929
rect 13633 13920 13645 13923
rect 13596 13892 13645 13920
rect 13596 13880 13602 13892
rect 13633 13889 13645 13892
rect 13679 13889 13691 13923
rect 13814 13920 13820 13932
rect 13775 13892 13820 13920
rect 13633 13883 13691 13889
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 14151 13923 14209 13929
rect 14151 13889 14163 13923
rect 14197 13920 14209 13923
rect 14458 13920 14464 13932
rect 14197 13892 14320 13920
rect 14419 13892 14464 13920
rect 14197 13889 14209 13892
rect 14151 13883 14209 13889
rect 8996 13824 9089 13852
rect 13372 13824 13676 13852
rect 8996 13812 9002 13824
rect 8294 13744 8300 13796
rect 8352 13784 8358 13796
rect 13262 13784 13268 13796
rect 8352 13756 13268 13784
rect 8352 13744 8358 13756
rect 13262 13744 13268 13756
rect 13320 13744 13326 13796
rect 13648 13784 13676 13824
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13780 13824 13921 13852
rect 13780 13812 13786 13824
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 14292 13852 14320 13892
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 14573 13929 14601 13960
rect 14645 13957 14657 13960
rect 14691 13957 14703 13991
rect 14826 13988 14832 14000
rect 14787 13960 14832 13988
rect 14645 13951 14703 13957
rect 14826 13948 14832 13960
rect 14884 13948 14890 14000
rect 16868 13988 16896 14016
rect 17773 13991 17831 13997
rect 17773 13988 17785 13991
rect 16868 13960 17785 13988
rect 17773 13957 17785 13960
rect 17819 13988 17831 13991
rect 18506 13988 18512 14000
rect 17819 13960 18512 13988
rect 17819 13957 17831 13960
rect 17773 13951 17831 13957
rect 18506 13948 18512 13960
rect 18564 13988 18570 14000
rect 18877 13991 18935 13997
rect 18877 13988 18889 13991
rect 18564 13960 18889 13988
rect 18564 13948 18570 13960
rect 18877 13957 18889 13960
rect 18923 13988 18935 13991
rect 23109 13991 23167 13997
rect 23109 13988 23121 13991
rect 18923 13960 19334 13988
rect 18923 13957 18935 13960
rect 18877 13951 18935 13957
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13889 14611 13923
rect 19306 13920 19334 13960
rect 22296 13960 23121 13988
rect 22296 13932 22324 13960
rect 23109 13957 23121 13960
rect 23155 13957 23167 13991
rect 23109 13951 23167 13957
rect 20438 13920 20444 13932
rect 19306 13892 20208 13920
rect 20399 13892 20444 13920
rect 14553 13883 14611 13889
rect 14734 13852 14740 13864
rect 14292 13824 14740 13852
rect 13909 13815 13967 13821
rect 14734 13812 14740 13824
rect 14792 13852 14798 13864
rect 19444 13861 19472 13892
rect 20180 13864 20208 13892
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 20806 13880 20812 13932
rect 20864 13920 20870 13932
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 20864 13892 21833 13920
rect 20864 13880 20870 13892
rect 21821 13889 21833 13892
rect 21867 13889 21879 13923
rect 22002 13920 22008 13932
rect 21963 13892 22008 13920
rect 21821 13883 21879 13889
rect 22002 13880 22008 13892
rect 22060 13880 22066 13932
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13920 22155 13923
rect 22278 13920 22284 13932
rect 22143 13892 22284 13920
rect 22143 13889 22155 13892
rect 22097 13883 22155 13889
rect 22278 13880 22284 13892
rect 22336 13880 22342 13932
rect 22830 13880 22836 13932
rect 22888 13920 22894 13932
rect 23017 13923 23075 13929
rect 23017 13920 23029 13923
rect 22888 13892 23029 13920
rect 22888 13880 22894 13892
rect 23017 13889 23029 13892
rect 23063 13889 23075 13923
rect 23017 13883 23075 13889
rect 15013 13855 15071 13861
rect 15013 13852 15025 13855
rect 14792 13824 15025 13852
rect 14792 13812 14798 13824
rect 15013 13821 15025 13824
rect 15059 13821 15071 13855
rect 15013 13815 15071 13821
rect 19429 13855 19487 13861
rect 19429 13821 19441 13855
rect 19475 13821 19487 13855
rect 19429 13815 19487 13821
rect 19521 13855 19579 13861
rect 19521 13821 19533 13855
rect 19567 13852 19579 13855
rect 19886 13852 19892 13864
rect 19567 13824 19892 13852
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 19886 13812 19892 13824
rect 19944 13812 19950 13864
rect 20162 13852 20168 13864
rect 20123 13824 20168 13852
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20346 13852 20352 13864
rect 20307 13824 20352 13852
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 22554 13852 22560 13864
rect 22515 13824 22560 13852
rect 22554 13812 22560 13824
rect 22612 13812 22618 13864
rect 23201 13855 23259 13861
rect 23201 13852 23213 13855
rect 23032 13824 23213 13852
rect 23032 13796 23060 13824
rect 23201 13821 23213 13824
rect 23247 13821 23259 13855
rect 23201 13815 23259 13821
rect 14458 13784 14464 13796
rect 13648 13756 14464 13784
rect 14458 13744 14464 13756
rect 14516 13784 14522 13796
rect 14642 13784 14648 13796
rect 14516 13756 14648 13784
rect 14516 13744 14522 13756
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 17037 13787 17095 13793
rect 17037 13753 17049 13787
rect 17083 13784 17095 13787
rect 17218 13784 17224 13796
rect 17083 13756 17224 13784
rect 17083 13753 17095 13756
rect 17037 13747 17095 13753
rect 17218 13744 17224 13756
rect 17276 13744 17282 13796
rect 23014 13784 23020 13796
rect 21560 13756 23020 13784
rect 7432 13688 7512 13716
rect 7432 13676 7438 13688
rect 8202 13676 8208 13728
rect 8260 13716 8266 13728
rect 9217 13719 9275 13725
rect 9217 13716 9229 13719
rect 8260 13688 9229 13716
rect 8260 13676 8266 13688
rect 9217 13685 9229 13688
rect 9263 13685 9275 13719
rect 11514 13716 11520 13728
rect 11427 13688 11520 13716
rect 9217 13679 9275 13685
rect 11514 13676 11520 13688
rect 11572 13716 11578 13728
rect 11974 13716 11980 13728
rect 11572 13688 11980 13716
rect 11572 13676 11578 13688
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 12894 13716 12900 13728
rect 12807 13688 12900 13716
rect 12894 13676 12900 13688
rect 12952 13716 12958 13728
rect 17494 13716 17500 13728
rect 12952 13688 17500 13716
rect 12952 13676 12958 13688
rect 17494 13676 17500 13688
rect 17552 13716 17558 13728
rect 20898 13716 20904 13728
rect 17552 13688 20904 13716
rect 17552 13676 17558 13688
rect 20898 13676 20904 13688
rect 20956 13676 20962 13728
rect 20990 13676 20996 13728
rect 21048 13716 21054 13728
rect 21560 13725 21588 13756
rect 23014 13744 23020 13756
rect 23072 13744 23078 13796
rect 21545 13719 21603 13725
rect 21545 13716 21557 13719
rect 21048 13688 21557 13716
rect 21048 13676 21054 13688
rect 21545 13685 21557 13688
rect 21591 13685 21603 13719
rect 21545 13679 21603 13685
rect 21634 13676 21640 13728
rect 21692 13716 21698 13728
rect 21821 13719 21879 13725
rect 21821 13716 21833 13719
rect 21692 13688 21833 13716
rect 21692 13676 21698 13688
rect 21821 13685 21833 13688
rect 21867 13685 21879 13719
rect 22646 13716 22652 13728
rect 22607 13688 22652 13716
rect 21821 13679 21879 13685
rect 22646 13676 22652 13688
rect 22704 13676 22710 13728
rect 1104 13626 26220 13648
rect 1104 13574 5136 13626
rect 5188 13574 5200 13626
rect 5252 13574 5264 13626
rect 5316 13574 5328 13626
rect 5380 13574 5392 13626
rect 5444 13574 13508 13626
rect 13560 13574 13572 13626
rect 13624 13574 13636 13626
rect 13688 13574 13700 13626
rect 13752 13574 13764 13626
rect 13816 13574 21880 13626
rect 21932 13574 21944 13626
rect 21996 13574 22008 13626
rect 22060 13574 22072 13626
rect 22124 13574 22136 13626
rect 22188 13574 26220 13626
rect 1104 13552 26220 13574
rect 3326 13472 3332 13524
rect 3384 13512 3390 13524
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 3384 13484 5181 13512
rect 3384 13472 3390 13484
rect 5169 13481 5181 13484
rect 5215 13512 5227 13515
rect 8478 13512 8484 13524
rect 5215 13484 8484 13512
rect 5215 13481 5227 13484
rect 5169 13475 5227 13481
rect 8478 13472 8484 13484
rect 8536 13472 8542 13524
rect 8662 13472 8668 13524
rect 8720 13512 8726 13524
rect 8938 13512 8944 13524
rect 8720 13484 8944 13512
rect 8720 13472 8726 13484
rect 8938 13472 8944 13484
rect 8996 13472 9002 13524
rect 9324 13484 10364 13512
rect 2498 13404 2504 13456
rect 2556 13444 2562 13456
rect 2869 13447 2927 13453
rect 2869 13444 2881 13447
rect 2556 13416 2881 13444
rect 2556 13404 2562 13416
rect 2869 13413 2881 13416
rect 2915 13444 2927 13447
rect 3605 13447 3663 13453
rect 3605 13444 3617 13447
rect 2915 13416 3617 13444
rect 2915 13413 2927 13416
rect 2869 13407 2927 13413
rect 3605 13413 3617 13416
rect 3651 13413 3663 13447
rect 3605 13407 3663 13413
rect 8110 13404 8116 13456
rect 8168 13444 8174 13456
rect 9324 13453 9352 13484
rect 9309 13447 9367 13453
rect 9309 13444 9321 13447
rect 8168 13416 9321 13444
rect 8168 13404 8174 13416
rect 3418 13336 3424 13388
rect 3476 13376 3482 13388
rect 3789 13379 3847 13385
rect 3789 13376 3801 13379
rect 3476 13348 3801 13376
rect 3476 13336 3482 13348
rect 3789 13345 3801 13348
rect 3835 13345 3847 13379
rect 7926 13376 7932 13388
rect 7887 13348 7932 13376
rect 3789 13339 3847 13345
rect 7926 13336 7932 13348
rect 7984 13336 7990 13388
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 8352 13348 8493 13376
rect 8352 13336 8358 13348
rect 8481 13345 8493 13348
rect 8527 13345 8539 13379
rect 8481 13339 8539 13345
rect 1486 13308 1492 13320
rect 1447 13280 1492 13308
rect 1486 13268 1492 13280
rect 1544 13268 1550 13320
rect 3234 13268 3240 13320
rect 3292 13308 3298 13320
rect 3329 13311 3387 13317
rect 3329 13308 3341 13311
rect 3292 13280 3341 13308
rect 3292 13268 3298 13280
rect 3329 13277 3341 13280
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13308 3571 13311
rect 3605 13311 3663 13317
rect 3605 13308 3617 13311
rect 3559 13280 3617 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 3605 13277 3617 13280
rect 3651 13308 3663 13311
rect 4982 13308 4988 13320
rect 3651 13280 4988 13308
rect 3651 13277 3663 13280
rect 3605 13271 3663 13277
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 8205 13311 8263 13317
rect 8205 13308 8217 13311
rect 6512 13280 8217 13308
rect 6512 13268 6518 13280
rect 8205 13277 8217 13280
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 1756 13243 1814 13249
rect 1756 13209 1768 13243
rect 1802 13240 1814 13243
rect 2130 13240 2136 13252
rect 1802 13212 2136 13240
rect 1802 13209 1814 13212
rect 1756 13203 1814 13209
rect 2130 13200 2136 13212
rect 2188 13200 2194 13252
rect 3418 13200 3424 13252
rect 3476 13240 3482 13252
rect 4034 13243 4092 13249
rect 4034 13240 4046 13243
rect 3476 13212 4046 13240
rect 3476 13200 3482 13212
rect 4034 13209 4046 13212
rect 4080 13209 4092 13243
rect 4034 13203 4092 13209
rect 7006 13200 7012 13252
rect 7064 13240 7070 13252
rect 7662 13243 7720 13249
rect 7662 13240 7674 13243
rect 7064 13212 7674 13240
rect 7064 13200 7070 13212
rect 7662 13209 7674 13212
rect 7708 13209 7720 13243
rect 7662 13203 7720 13209
rect 8018 13200 8024 13252
rect 8076 13240 8082 13252
rect 8404 13240 8432 13271
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 8772 13317 8800 13416
rect 9309 13413 9321 13416
rect 9355 13413 9367 13447
rect 10336 13444 10364 13484
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 10781 13515 10839 13521
rect 10781 13512 10793 13515
rect 10468 13484 10793 13512
rect 10468 13472 10474 13484
rect 10781 13481 10793 13484
rect 10827 13481 10839 13515
rect 12158 13512 12164 13524
rect 10781 13475 10839 13481
rect 11624 13484 12164 13512
rect 11624 13444 11652 13484
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 13998 13512 14004 13524
rect 13587 13484 14004 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 14185 13515 14243 13521
rect 14185 13481 14197 13515
rect 14231 13512 14243 13515
rect 14366 13512 14372 13524
rect 14231 13484 14372 13512
rect 14231 13481 14243 13484
rect 14185 13475 14243 13481
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 14550 13512 14556 13524
rect 14511 13484 14556 13512
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 16301 13515 16359 13521
rect 16301 13481 16313 13515
rect 16347 13512 16359 13515
rect 16482 13512 16488 13524
rect 16347 13484 16488 13512
rect 16347 13481 16359 13484
rect 16301 13475 16359 13481
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 17494 13512 17500 13524
rect 17144 13484 17500 13512
rect 12894 13444 12900 13456
rect 10336 13416 11652 13444
rect 11716 13416 12900 13444
rect 9309 13407 9367 13413
rect 9214 13336 9220 13388
rect 9272 13376 9278 13388
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 9272 13348 9413 13376
rect 9272 13336 9278 13348
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 8757 13311 8815 13317
rect 8628 13280 8673 13308
rect 8628 13268 8634 13280
rect 8757 13277 8769 13311
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 11716 13317 11744 13416
rect 12894 13404 12900 13416
rect 12952 13404 12958 13456
rect 13078 13404 13084 13456
rect 13136 13444 13142 13456
rect 14277 13447 14335 13453
rect 14277 13444 14289 13447
rect 13136 13416 14289 13444
rect 13136 13404 13142 13416
rect 14277 13413 14289 13416
rect 14323 13444 14335 13447
rect 14323 13416 15424 13444
rect 14323 13413 14335 13416
rect 14277 13407 14335 13413
rect 11974 13376 11980 13388
rect 11935 13348 11980 13376
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 12066 13336 12072 13388
rect 12124 13376 12130 13388
rect 12529 13379 12587 13385
rect 12529 13376 12541 13379
rect 12124 13348 12169 13376
rect 12360 13348 12541 13376
rect 12124 13336 12130 13348
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 9088 13280 9137 13308
rect 9088 13268 9094 13280
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13277 11759 13311
rect 11882 13308 11888 13320
rect 11843 13280 11888 13308
rect 11701 13271 11759 13277
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 9674 13249 9680 13252
rect 8076 13212 8432 13240
rect 8076 13200 8082 13212
rect 9668 13203 9680 13249
rect 9732 13240 9738 13252
rect 9732 13212 9768 13240
rect 9674 13200 9680 13203
rect 9732 13200 9738 13212
rect 11238 13200 11244 13252
rect 11296 13240 11302 13252
rect 12084 13240 12112 13336
rect 12250 13308 12256 13320
rect 12211 13280 12256 13308
rect 12250 13268 12256 13280
rect 12308 13268 12314 13320
rect 11296 13212 12112 13240
rect 11296 13200 11302 13212
rect 3142 13172 3148 13184
rect 3103 13144 3148 13172
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 6549 13175 6607 13181
rect 6549 13141 6561 13175
rect 6595 13172 6607 13175
rect 6914 13172 6920 13184
rect 6595 13144 6920 13172
rect 6595 13141 6607 13144
rect 6549 13135 6607 13141
rect 6914 13132 6920 13144
rect 6972 13172 6978 13184
rect 7190 13172 7196 13184
rect 6972 13144 7196 13172
rect 6972 13132 6978 13144
rect 7190 13132 7196 13144
rect 7248 13132 7254 13184
rect 8110 13172 8116 13184
rect 8071 13144 8116 13172
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8996 13144 9045 13172
rect 8996 13132 9002 13144
rect 9033 13141 9045 13144
rect 9079 13141 9091 13175
rect 9033 13135 9091 13141
rect 9858 13132 9864 13184
rect 9916 13172 9922 13184
rect 10686 13172 10692 13184
rect 9916 13144 10692 13172
rect 9916 13132 9922 13144
rect 10686 13132 10692 13144
rect 10744 13172 10750 13184
rect 11422 13172 11428 13184
rect 10744 13144 11428 13172
rect 10744 13132 10750 13144
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 12360 13172 12388 13348
rect 12529 13345 12541 13348
rect 12575 13345 12587 13379
rect 12529 13339 12587 13345
rect 14366 13336 14372 13388
rect 14424 13376 14430 13388
rect 15105 13379 15163 13385
rect 15105 13376 15117 13379
rect 14424 13348 15117 13376
rect 14424 13336 14430 13348
rect 15105 13345 15117 13348
rect 15151 13345 15163 13379
rect 15105 13339 15163 13345
rect 13354 13308 13360 13320
rect 13315 13280 13360 13308
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 14274 13308 14280 13320
rect 14056 13280 14280 13308
rect 14056 13268 14062 13280
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 14458 13308 14464 13320
rect 14419 13280 14464 13308
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 15396 13317 15424 13416
rect 15469 13416 17080 13444
rect 15381 13311 15439 13317
rect 15381 13277 15393 13311
rect 15427 13277 15439 13311
rect 15469 13308 15497 13416
rect 15654 13376 15660 13388
rect 15615 13348 15660 13376
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 15749 13379 15807 13385
rect 15749 13345 15761 13379
rect 15795 13376 15807 13379
rect 15838 13376 15844 13388
rect 15795 13348 15844 13376
rect 15795 13345 15807 13348
rect 15749 13339 15807 13345
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 16850 13376 16856 13388
rect 16811 13348 16856 13376
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 15529 13311 15587 13317
rect 15529 13308 15541 13311
rect 15469 13280 15541 13308
rect 15381 13271 15439 13277
rect 15529 13277 15541 13280
rect 15575 13277 15587 13311
rect 15529 13271 15587 13277
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 12437 13243 12495 13249
rect 12437 13209 12449 13243
rect 12483 13240 12495 13243
rect 13262 13240 13268 13252
rect 12483 13212 13268 13240
rect 12483 13209 12495 13212
rect 12437 13203 12495 13209
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 15102 13200 15108 13252
rect 15160 13240 15166 13252
rect 15948 13240 15976 13271
rect 15160 13212 15976 13240
rect 15160 13200 15166 13212
rect 16574 13200 16580 13252
rect 16632 13240 16638 13252
rect 16761 13243 16819 13249
rect 16761 13240 16773 13243
rect 16632 13212 16773 13240
rect 16632 13200 16638 13212
rect 16761 13209 16773 13212
rect 16807 13209 16819 13243
rect 17052 13240 17080 13416
rect 17144 13317 17172 13484
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 17586 13472 17592 13524
rect 17644 13472 17650 13524
rect 17957 13515 18015 13521
rect 17957 13481 17969 13515
rect 18003 13512 18015 13515
rect 18690 13512 18696 13524
rect 18003 13484 18696 13512
rect 18003 13481 18015 13484
rect 17957 13475 18015 13481
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 19337 13515 19395 13521
rect 19337 13481 19349 13515
rect 19383 13512 19395 13515
rect 19610 13512 19616 13524
rect 19383 13484 19616 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 20165 13515 20223 13521
rect 20165 13481 20177 13515
rect 20211 13512 20223 13515
rect 20438 13512 20444 13524
rect 20211 13484 20444 13512
rect 20211 13481 20223 13484
rect 20165 13475 20223 13481
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 20990 13512 20996 13524
rect 20732 13484 20996 13512
rect 17604 13444 17632 13472
rect 18877 13447 18935 13453
rect 18877 13444 18889 13447
rect 17512 13416 17632 13444
rect 18708 13416 18889 13444
rect 17402 13376 17408 13388
rect 17363 13348 17408 13376
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 17512 13385 17540 13416
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13345 17555 13379
rect 17497 13339 17555 13345
rect 17586 13336 17592 13388
rect 17644 13376 17650 13388
rect 18417 13379 18475 13385
rect 18417 13376 18429 13379
rect 17644 13348 18429 13376
rect 17644 13336 17650 13348
rect 18417 13345 18429 13348
rect 18463 13345 18475 13379
rect 18417 13339 18475 13345
rect 18506 13336 18512 13388
rect 18564 13376 18570 13388
rect 18564 13348 18609 13376
rect 18564 13336 18570 13348
rect 17129 13311 17187 13317
rect 17129 13277 17141 13311
rect 17175 13277 17187 13311
rect 17129 13271 17187 13277
rect 17218 13268 17224 13320
rect 17276 13308 17282 13320
rect 17312 13311 17370 13317
rect 17312 13308 17324 13311
rect 17276 13280 17324 13308
rect 17276 13268 17282 13280
rect 17312 13277 17324 13280
rect 17358 13277 17370 13311
rect 17312 13271 17370 13277
rect 17681 13311 17739 13317
rect 17681 13277 17693 13311
rect 17727 13308 17739 13311
rect 18708 13308 18736 13416
rect 18877 13413 18889 13416
rect 18923 13444 18935 13447
rect 19518 13444 19524 13456
rect 18923 13416 19524 13444
rect 18923 13413 18935 13416
rect 18877 13407 18935 13413
rect 19518 13404 19524 13416
rect 19576 13404 19582 13456
rect 19242 13336 19248 13388
rect 19300 13376 19306 13388
rect 20732 13385 20760 13484
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 22278 13472 22284 13524
rect 22336 13512 22342 13524
rect 23385 13515 23443 13521
rect 23385 13512 23397 13515
rect 22336 13484 23397 13512
rect 22336 13472 22342 13484
rect 23385 13481 23397 13484
rect 23431 13481 23443 13515
rect 23385 13475 23443 13481
rect 21266 13444 21272 13456
rect 20824 13416 21272 13444
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 19300 13348 19901 13376
rect 19300 13336 19306 13348
rect 19889 13345 19901 13348
rect 19935 13376 19947 13379
rect 20717 13379 20775 13385
rect 20717 13376 20729 13379
rect 19935 13348 20729 13376
rect 19935 13345 19947 13348
rect 19889 13339 19947 13345
rect 20717 13345 20729 13348
rect 20763 13345 20775 13379
rect 20717 13339 20775 13345
rect 17727 13280 18736 13308
rect 19061 13311 19119 13317
rect 17727 13277 17739 13280
rect 17681 13271 17739 13277
rect 19061 13277 19073 13311
rect 19107 13308 19119 13311
rect 19107 13280 20300 13308
rect 19107 13277 19119 13280
rect 19061 13271 19119 13277
rect 17696 13240 17724 13271
rect 17052 13212 17724 13240
rect 17865 13243 17923 13249
rect 16761 13203 16819 13209
rect 17865 13209 17877 13243
rect 17911 13240 17923 13243
rect 18230 13240 18236 13252
rect 17911 13212 18236 13240
rect 17911 13209 17923 13212
rect 17865 13203 17923 13209
rect 18230 13200 18236 13212
rect 18288 13200 18294 13252
rect 19705 13243 19763 13249
rect 19705 13209 19717 13243
rect 19751 13240 19763 13243
rect 19886 13240 19892 13252
rect 19751 13212 19892 13240
rect 19751 13209 19763 13212
rect 19705 13203 19763 13209
rect 19886 13200 19892 13212
rect 19944 13200 19950 13252
rect 20272 13240 20300 13280
rect 20346 13268 20352 13320
rect 20404 13308 20410 13320
rect 20533 13311 20591 13317
rect 20533 13308 20545 13311
rect 20404 13280 20545 13308
rect 20404 13268 20410 13280
rect 20533 13277 20545 13280
rect 20579 13308 20591 13311
rect 20622 13308 20628 13320
rect 20579 13280 20628 13308
rect 20579 13277 20591 13280
rect 20533 13271 20591 13277
rect 20622 13268 20628 13280
rect 20680 13268 20686 13320
rect 20824 13240 20852 13416
rect 21266 13404 21272 13416
rect 21324 13444 21330 13456
rect 21634 13444 21640 13456
rect 21324 13416 21640 13444
rect 21324 13404 21330 13416
rect 21634 13404 21640 13416
rect 21692 13404 21698 13456
rect 21376 13348 22140 13376
rect 20898 13268 20904 13320
rect 20956 13308 20962 13320
rect 21376 13317 21404 13348
rect 21177 13311 21235 13317
rect 21177 13308 21189 13311
rect 20956 13280 21189 13308
rect 20956 13268 20962 13280
rect 21177 13277 21189 13280
rect 21223 13277 21235 13311
rect 21177 13271 21235 13277
rect 21360 13311 21418 13317
rect 21360 13277 21372 13311
rect 21406 13277 21418 13311
rect 21360 13271 21418 13277
rect 21450 13311 21508 13317
rect 21450 13296 21462 13311
rect 21496 13296 21508 13311
rect 21545 13311 21603 13317
rect 21450 13244 21456 13296
rect 21508 13244 21514 13296
rect 21545 13277 21557 13311
rect 21591 13277 21603 13311
rect 21726 13308 21732 13320
rect 21687 13280 21732 13308
rect 21545 13271 21603 13277
rect 20272 13212 20852 13240
rect 21560 13240 21588 13271
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 22002 13308 22008 13320
rect 21963 13280 22008 13308
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 22112 13308 22140 13348
rect 22554 13308 22560 13320
rect 22112 13280 22560 13308
rect 22554 13268 22560 13280
rect 22612 13308 22618 13320
rect 23382 13308 23388 13320
rect 22612 13280 23388 13308
rect 22612 13268 22618 13280
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 23474 13268 23480 13320
rect 23532 13308 23538 13320
rect 23569 13311 23627 13317
rect 23569 13308 23581 13311
rect 23532 13280 23581 13308
rect 23532 13268 23538 13280
rect 23569 13277 23581 13280
rect 23615 13277 23627 13311
rect 23569 13271 23627 13277
rect 23658 13268 23664 13320
rect 23716 13308 23722 13320
rect 23753 13311 23811 13317
rect 23753 13308 23765 13311
rect 23716 13280 23765 13308
rect 23716 13268 23722 13280
rect 23753 13277 23765 13280
rect 23799 13277 23811 13311
rect 23753 13271 23811 13277
rect 21818 13240 21824 13252
rect 21560 13212 21824 13240
rect 11940 13144 12388 13172
rect 11940 13132 11946 13144
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 14884 13144 14933 13172
rect 14884 13132 14890 13144
rect 14921 13141 14933 13144
rect 14967 13141 14979 13175
rect 14921 13135 14979 13141
rect 15013 13175 15071 13181
rect 15013 13141 15025 13175
rect 15059 13172 15071 13175
rect 15286 13172 15292 13184
rect 15059 13144 15292 13172
rect 15059 13141 15071 13144
rect 15013 13135 15071 13141
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 16022 13172 16028 13184
rect 15983 13144 16028 13172
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 16669 13175 16727 13181
rect 16669 13141 16681 13175
rect 16715 13172 16727 13175
rect 16942 13172 16948 13184
rect 16715 13144 16948 13172
rect 16715 13141 16727 13144
rect 16669 13135 16727 13141
rect 16942 13132 16948 13144
rect 17000 13132 17006 13184
rect 18046 13132 18052 13184
rect 18104 13172 18110 13184
rect 18325 13175 18383 13181
rect 18325 13172 18337 13175
rect 18104 13144 18337 13172
rect 18104 13132 18110 13144
rect 18325 13141 18337 13144
rect 18371 13141 18383 13175
rect 19794 13172 19800 13184
rect 19755 13144 19800 13172
rect 18325 13135 18383 13141
rect 19794 13132 19800 13144
rect 19852 13132 19858 13184
rect 20625 13175 20683 13181
rect 20625 13141 20637 13175
rect 20671 13172 20683 13175
rect 20824 13172 20852 13212
rect 21818 13200 21824 13212
rect 21876 13200 21882 13252
rect 21913 13243 21971 13249
rect 21913 13209 21925 13243
rect 21959 13240 21971 13243
rect 22250 13243 22308 13249
rect 22250 13240 22262 13243
rect 21959 13212 22262 13240
rect 21959 13209 21971 13212
rect 21913 13203 21971 13209
rect 22250 13209 22262 13212
rect 22296 13209 22308 13243
rect 23768 13240 23796 13271
rect 22250 13203 22308 13209
rect 23032 13212 23796 13240
rect 20671 13144 20852 13172
rect 20671 13141 20683 13144
rect 20625 13135 20683 13141
rect 21634 13132 21640 13184
rect 21692 13172 21698 13184
rect 23032 13172 23060 13212
rect 21692 13144 23060 13172
rect 21692 13132 21698 13144
rect 23106 13132 23112 13184
rect 23164 13172 23170 13184
rect 23290 13172 23296 13184
rect 23164 13144 23296 13172
rect 23164 13132 23170 13144
rect 23290 13132 23296 13144
rect 23348 13172 23354 13184
rect 23661 13175 23719 13181
rect 23661 13172 23673 13175
rect 23348 13144 23673 13172
rect 23348 13132 23354 13144
rect 23661 13141 23673 13144
rect 23707 13141 23719 13175
rect 23661 13135 23719 13141
rect 1104 13082 26220 13104
rect 1104 13030 9322 13082
rect 9374 13030 9386 13082
rect 9438 13030 9450 13082
rect 9502 13030 9514 13082
rect 9566 13030 9578 13082
rect 9630 13030 17694 13082
rect 17746 13030 17758 13082
rect 17810 13030 17822 13082
rect 17874 13030 17886 13082
rect 17938 13030 17950 13082
rect 18002 13030 26220 13082
rect 1104 13008 26220 13030
rect 2130 12968 2136 12980
rect 2091 12940 2136 12968
rect 2130 12928 2136 12940
rect 2188 12928 2194 12980
rect 2958 12968 2964 12980
rect 2792 12940 2964 12968
rect 2498 12900 2504 12912
rect 2332 12872 2504 12900
rect 2332 12841 2360 12872
rect 2498 12860 2504 12872
rect 2556 12860 2562 12912
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12801 2375 12835
rect 2317 12795 2375 12801
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12832 2467 12835
rect 2590 12832 2596 12844
rect 2455 12804 2596 12832
rect 2455 12801 2467 12804
rect 2409 12795 2467 12801
rect 2590 12792 2596 12804
rect 2648 12792 2654 12844
rect 2792 12841 2820 12940
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 3418 12968 3424 12980
rect 3160 12940 3326 12968
rect 3379 12940 3424 12968
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 2960 12835 3018 12841
rect 2960 12801 2972 12835
rect 3006 12801 3018 12835
rect 3160 12832 3188 12940
rect 3298 12900 3326 12940
rect 3418 12928 3424 12940
rect 3476 12928 3482 12980
rect 3970 12968 3976 12980
rect 3528 12940 3976 12968
rect 3528 12900 3556 12940
rect 3298 12872 3556 12900
rect 2960 12795 3018 12801
rect 3068 12804 3188 12832
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12733 2743 12767
rect 2685 12727 2743 12733
rect 2700 12696 2728 12727
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 2976 12764 3004 12795
rect 3068 12773 3096 12804
rect 3326 12792 3332 12844
rect 3384 12832 3390 12844
rect 3384 12804 3429 12832
rect 3384 12792 3390 12804
rect 3510 12792 3516 12844
rect 3568 12832 3574 12844
rect 3602 12835 3660 12841
rect 3602 12832 3614 12835
rect 3568 12804 3614 12832
rect 3568 12792 3574 12804
rect 3602 12801 3614 12804
rect 3648 12801 3660 12835
rect 3786 12832 3792 12844
rect 3747 12804 3792 12832
rect 3602 12795 3660 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 3896 12841 3924 12940
rect 3970 12928 3976 12940
rect 4028 12968 4034 12980
rect 4890 12968 4896 12980
rect 4028 12940 4896 12968
rect 4028 12928 4034 12940
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 6454 12968 6460 12980
rect 6415 12940 6460 12968
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 7800 12940 7941 12968
rect 7800 12928 7806 12940
rect 7929 12937 7941 12940
rect 7975 12937 7987 12971
rect 7929 12931 7987 12937
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8444 12940 8769 12968
rect 8444 12928 8450 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 8757 12931 8815 12937
rect 9585 12971 9643 12977
rect 9585 12937 9597 12971
rect 9631 12968 9643 12971
rect 9674 12968 9680 12980
rect 9631 12940 9680 12968
rect 9631 12937 9643 12940
rect 9585 12931 9643 12937
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 10502 12968 10508 12980
rect 9824 12940 10508 12968
rect 9824 12928 9830 12940
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 11146 12928 11152 12980
rect 11204 12928 11210 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 12250 12968 12256 12980
rect 11756 12940 12256 12968
rect 11756 12928 11762 12940
rect 12250 12928 12256 12940
rect 12308 12968 12314 12980
rect 12308 12940 13584 12968
rect 12308 12928 12314 12940
rect 4430 12900 4436 12912
rect 4391 12872 4436 12900
rect 4430 12860 4436 12872
rect 4488 12860 4494 12912
rect 4798 12900 4804 12912
rect 4632 12872 4804 12900
rect 3881 12835 3939 12841
rect 3881 12801 3893 12835
rect 3927 12801 3939 12835
rect 3881 12795 3939 12801
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12832 4215 12835
rect 4522 12832 4528 12844
rect 4203 12804 4528 12832
rect 4203 12801 4215 12804
rect 4157 12795 4215 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 4632 12841 4660 12872
rect 4798 12860 4804 12872
rect 4856 12860 4862 12912
rect 7592 12903 7650 12909
rect 7592 12869 7604 12903
rect 7638 12900 7650 12903
rect 8110 12900 8116 12912
rect 7638 12872 8116 12900
rect 7638 12869 7650 12872
rect 7592 12863 7650 12869
rect 8110 12860 8116 12872
rect 8168 12860 8174 12912
rect 8297 12903 8355 12909
rect 8297 12869 8309 12903
rect 8343 12900 8355 12903
rect 11164 12900 11192 12928
rect 11514 12900 11520 12912
rect 8343 12872 9628 12900
rect 8343 12869 8355 12872
rect 8297 12863 8355 12869
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12801 4675 12835
rect 4982 12832 4988 12844
rect 4944 12804 4988 12832
rect 4617 12795 4675 12801
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 5166 12832 5172 12844
rect 5127 12804 5172 12832
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 5718 12832 5724 12844
rect 5491 12804 5724 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 5810 12792 5816 12844
rect 5868 12832 5874 12844
rect 7837 12835 7895 12841
rect 5868 12804 5913 12832
rect 5868 12792 5874 12804
rect 7837 12801 7849 12835
rect 7883 12832 7895 12835
rect 7926 12832 7932 12844
rect 7883 12804 7932 12832
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 8754 12792 8760 12844
rect 8812 12832 8818 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8812 12804 8953 12832
rect 8812 12792 8818 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9124 12835 9182 12841
rect 9124 12801 9136 12835
rect 9170 12832 9182 12835
rect 9398 12832 9404 12844
rect 9170 12804 9404 12832
rect 9170 12801 9182 12804
rect 9124 12795 9182 12801
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 2924 12736 3004 12764
rect 3053 12767 3111 12773
rect 2924 12724 2930 12736
rect 3053 12733 3065 12767
rect 3099 12733 3111 12767
rect 3053 12727 3111 12733
rect 3145 12767 3203 12773
rect 3145 12733 3157 12767
rect 3191 12764 3203 12767
rect 3973 12767 4031 12773
rect 3191 12736 3740 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 2958 12696 2964 12708
rect 2700 12668 2964 12696
rect 2958 12656 2964 12668
rect 3016 12656 3022 12708
rect 3712 12696 3740 12736
rect 3973 12733 3985 12767
rect 4019 12764 4031 12767
rect 4338 12764 4344 12776
rect 4019 12736 4344 12764
rect 4019 12733 4031 12736
rect 3973 12727 4031 12733
rect 3988 12696 4016 12727
rect 4338 12724 4344 12736
rect 4396 12764 4402 12776
rect 4798 12764 4804 12776
rect 4396 12736 4804 12764
rect 4396 12724 4402 12736
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 4890 12724 4896 12776
rect 4948 12764 4954 12776
rect 8389 12767 8447 12773
rect 4948 12736 5672 12764
rect 4948 12724 4954 12736
rect 3712 12668 4016 12696
rect 4706 12656 4712 12708
rect 4764 12696 4770 12708
rect 5644 12705 5672 12736
rect 8389 12733 8401 12767
rect 8435 12733 8447 12767
rect 8389 12727 8447 12733
rect 5261 12699 5319 12705
rect 5261 12696 5273 12699
rect 4764 12668 5273 12696
rect 4764 12656 4770 12668
rect 5261 12665 5273 12668
rect 5307 12665 5319 12699
rect 5261 12659 5319 12665
rect 5629 12699 5687 12705
rect 5629 12665 5641 12699
rect 5675 12665 5687 12699
rect 5629 12659 5687 12665
rect 2593 12631 2651 12637
rect 2593 12597 2605 12631
rect 2639 12628 2651 12631
rect 3326 12628 3332 12640
rect 2639 12600 3332 12628
rect 2639 12597 2651 12600
rect 2593 12591 2651 12597
rect 3326 12588 3332 12600
rect 3384 12588 3390 12640
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4249 12631 4307 12637
rect 4249 12628 4261 12631
rect 4212 12600 4261 12628
rect 4212 12588 4218 12600
rect 4249 12597 4261 12600
rect 4295 12597 4307 12631
rect 4249 12591 4307 12597
rect 4522 12588 4528 12640
rect 4580 12628 4586 12640
rect 4982 12628 4988 12640
rect 4580 12600 4988 12628
rect 4580 12588 4586 12600
rect 4982 12588 4988 12600
rect 5040 12628 5046 12640
rect 8404 12628 8432 12727
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 8536 12736 8585 12764
rect 8536 12724 8542 12736
rect 8573 12733 8585 12736
rect 8619 12764 8631 12767
rect 8662 12764 8668 12776
rect 8619 12736 8668 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 9214 12764 9220 12776
rect 9175 12736 9220 12764
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9030 12656 9036 12708
rect 9088 12696 9094 12708
rect 9324 12696 9352 12727
rect 9088 12668 9352 12696
rect 9088 12656 9094 12668
rect 5040 12600 8432 12628
rect 9508 12628 9536 12795
rect 9600 12696 9628 12872
rect 10060 12872 11520 12900
rect 9766 12832 9772 12844
rect 9727 12804 9772 12832
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 9950 12832 9956 12844
rect 9911 12804 9956 12832
rect 9950 12792 9956 12804
rect 10008 12792 10014 12844
rect 10060 12841 10088 12872
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12801 10103 12835
rect 10318 12832 10324 12844
rect 10279 12804 10324 12832
rect 10045 12795 10103 12801
rect 10318 12792 10324 12804
rect 10376 12792 10382 12844
rect 10502 12792 10508 12844
rect 10560 12832 10566 12844
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 10560 12804 10609 12832
rect 10560 12792 10566 12804
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 10888 12841 10916 12872
rect 11514 12860 11520 12872
rect 11572 12860 11578 12912
rect 11624 12872 12434 12900
rect 10780 12835 10838 12841
rect 10780 12832 10792 12835
rect 10744 12804 10792 12832
rect 10744 12792 10750 12804
rect 10780 12801 10792 12804
rect 10826 12801 10838 12835
rect 10780 12795 10838 12801
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12801 10931 12835
rect 10873 12795 10931 12801
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 11330 12832 11336 12844
rect 11195 12804 11336 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 11624 12841 11652 12872
rect 12406 12844 12434 12872
rect 13262 12860 13268 12912
rect 13320 12900 13326 12912
rect 13418 12903 13476 12909
rect 13418 12900 13430 12903
rect 13320 12872 13430 12900
rect 13320 12860 13326 12872
rect 13418 12869 13430 12872
rect 13464 12869 13476 12903
rect 13556 12900 13584 12940
rect 14550 12928 14556 12980
rect 14608 12968 14614 12980
rect 15102 12968 15108 12980
rect 14608 12940 15108 12968
rect 14608 12928 14614 12940
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 16390 12928 16396 12980
rect 16448 12968 16454 12980
rect 17221 12971 17279 12977
rect 17221 12968 17233 12971
rect 16448 12940 17233 12968
rect 16448 12928 16454 12940
rect 17221 12937 17233 12940
rect 17267 12937 17279 12971
rect 17221 12931 17279 12937
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 17681 12971 17739 12977
rect 17681 12968 17693 12971
rect 17552 12940 17693 12968
rect 17552 12928 17558 12940
rect 17681 12937 17693 12940
rect 17727 12937 17739 12971
rect 18046 12968 18052 12980
rect 18007 12940 18052 12968
rect 17681 12931 17739 12937
rect 18046 12928 18052 12940
rect 18104 12928 18110 12980
rect 19521 12971 19579 12977
rect 19521 12937 19533 12971
rect 19567 12968 19579 12971
rect 21266 12968 21272 12980
rect 19567 12940 21272 12968
rect 19567 12937 19579 12940
rect 19521 12931 19579 12937
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 22925 12971 22983 12977
rect 22204 12940 22508 12968
rect 13556 12872 14601 12900
rect 13418 12863 13476 12869
rect 11609 12835 11667 12841
rect 11609 12801 11621 12835
rect 11655 12801 11667 12835
rect 11865 12835 11923 12841
rect 11865 12832 11877 12835
rect 11609 12795 11667 12801
rect 11716 12804 11877 12832
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12764 10195 12767
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 10183 12736 10977 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 10965 12733 10977 12736
rect 11011 12764 11023 12767
rect 11238 12764 11244 12776
rect 11011 12736 11244 12764
rect 11011 12733 11023 12736
rect 10965 12727 11023 12733
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 11716 12764 11744 12804
rect 11865 12801 11877 12804
rect 11911 12801 11923 12835
rect 12406 12804 12440 12844
rect 11865 12795 11923 12801
rect 12434 12792 12440 12804
rect 12492 12832 12498 12844
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 12492 12804 13185 12832
rect 12492 12792 12498 12804
rect 13173 12801 13185 12804
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 14573 12832 14601 12872
rect 16022 12860 16028 12912
rect 16080 12900 16086 12912
rect 16218 12903 16276 12909
rect 16218 12900 16230 12903
rect 16080 12872 16230 12900
rect 16080 12860 16086 12872
rect 16218 12869 16230 12872
rect 16264 12869 16276 12903
rect 17586 12900 17592 12912
rect 16218 12863 16276 12869
rect 16500 12872 17592 12900
rect 16500 12841 16528 12872
rect 17586 12860 17592 12872
rect 17644 12900 17650 12912
rect 22002 12900 22008 12912
rect 17644 12872 22008 12900
rect 17644 12860 17650 12872
rect 16485 12835 16543 12841
rect 14573 12804 16436 12832
rect 11624 12736 11744 12764
rect 10226 12696 10232 12708
rect 9600 12668 10232 12696
rect 10226 12656 10232 12668
rect 10284 12656 10290 12708
rect 10505 12699 10563 12705
rect 10505 12665 10517 12699
rect 10551 12696 10563 12699
rect 11624 12696 11652 12736
rect 14573 12705 14601 12804
rect 16408 12764 16436 12804
rect 16485 12801 16497 12835
rect 16531 12801 16543 12835
rect 16666 12832 16672 12844
rect 16627 12804 16672 12832
rect 16485 12795 16543 12801
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 18046 12832 18052 12844
rect 17267 12804 18052 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 16758 12764 16764 12776
rect 16408 12736 16528 12764
rect 16719 12736 16764 12764
rect 10551 12668 11652 12696
rect 14553 12699 14611 12705
rect 10551 12665 10563 12668
rect 10505 12659 10563 12665
rect 14553 12665 14565 12699
rect 14599 12665 14611 12699
rect 16500 12696 16528 12736
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 17420 12773 17448 12804
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 18156 12841 18184 12872
rect 22002 12860 22008 12872
rect 22060 12900 22066 12912
rect 22204 12900 22232 12940
rect 22060 12872 22232 12900
rect 22480 12900 22508 12940
rect 22925 12937 22937 12971
rect 22971 12968 22983 12971
rect 22971 12940 23888 12968
rect 22971 12937 22983 12940
rect 22925 12931 22983 12937
rect 23860 12900 23888 12940
rect 23998 12903 24056 12909
rect 23998 12900 24010 12903
rect 22480 12872 23796 12900
rect 23860 12872 24010 12900
rect 22060 12860 22066 12872
rect 18141 12835 18199 12841
rect 18141 12801 18153 12835
rect 18187 12801 18199 12835
rect 18141 12795 18199 12801
rect 18230 12792 18236 12844
rect 18288 12832 18294 12844
rect 19978 12841 19984 12844
rect 18397 12835 18455 12841
rect 18397 12832 18409 12835
rect 18288 12804 18409 12832
rect 18288 12792 18294 12804
rect 18397 12801 18409 12804
rect 18443 12801 18455 12835
rect 18397 12795 18455 12801
rect 19947 12835 19984 12841
rect 19947 12801 19959 12835
rect 19947 12795 19984 12801
rect 19978 12792 19984 12795
rect 20036 12792 20042 12844
rect 20441 12835 20499 12841
rect 20441 12801 20453 12835
rect 20487 12801 20499 12835
rect 20441 12795 20499 12801
rect 20625 12835 20683 12841
rect 20625 12801 20637 12835
rect 20671 12801 20683 12835
rect 20806 12832 20812 12844
rect 20767 12804 20812 12832
rect 20625 12795 20683 12801
rect 17405 12767 17463 12773
rect 17405 12733 17417 12767
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 17589 12767 17647 12773
rect 17589 12764 17601 12767
rect 17552 12736 17601 12764
rect 17552 12724 17558 12736
rect 17589 12733 17601 12736
rect 17635 12733 17647 12767
rect 17589 12727 17647 12733
rect 20257 12767 20315 12773
rect 20257 12733 20269 12767
rect 20303 12733 20315 12767
rect 20257 12727 20315 12733
rect 19702 12696 19708 12708
rect 16500 12668 17172 12696
rect 19663 12668 19708 12696
rect 14553 12659 14611 12665
rect 10410 12628 10416 12640
rect 9508 12600 10416 12628
rect 5040 12588 5046 12600
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 11241 12631 11299 12637
rect 11241 12597 11253 12631
rect 11287 12628 11299 12631
rect 12250 12628 12256 12640
rect 11287 12600 12256 12628
rect 11287 12597 11299 12600
rect 11241 12591 11299 12597
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 12342 12588 12348 12640
rect 12400 12628 12406 12640
rect 12989 12631 13047 12637
rect 12989 12628 13001 12631
rect 12400 12600 13001 12628
rect 12400 12588 12406 12600
rect 12989 12597 13001 12600
rect 13035 12628 13047 12631
rect 15378 12628 15384 12640
rect 13035 12600 15384 12628
rect 13035 12597 13047 12600
rect 12989 12591 13047 12597
rect 15378 12588 15384 12600
rect 15436 12628 15442 12640
rect 16669 12631 16727 12637
rect 16669 12628 16681 12631
rect 15436 12600 16681 12628
rect 15436 12588 15442 12600
rect 16669 12597 16681 12600
rect 16715 12597 16727 12631
rect 16669 12591 16727 12597
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 17037 12631 17095 12637
rect 17037 12628 17049 12631
rect 16908 12600 17049 12628
rect 16908 12588 16914 12600
rect 17037 12597 17049 12600
rect 17083 12597 17095 12631
rect 17144 12628 17172 12668
rect 19702 12656 19708 12668
rect 19760 12656 19766 12708
rect 20272 12696 20300 12727
rect 20346 12724 20352 12776
rect 20404 12764 20410 12776
rect 20456 12764 20484 12795
rect 20404 12736 20484 12764
rect 20404 12724 20410 12736
rect 20640 12696 20668 12795
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 20990 12792 20996 12844
rect 21048 12832 21054 12844
rect 21269 12835 21327 12841
rect 21269 12832 21281 12835
rect 21048 12804 21281 12832
rect 21048 12792 21054 12804
rect 21269 12801 21281 12804
rect 21315 12801 21327 12835
rect 21634 12832 21640 12844
rect 21595 12804 21640 12832
rect 21269 12795 21327 12801
rect 21634 12792 21640 12804
rect 21692 12792 21698 12844
rect 22186 12832 22192 12844
rect 22147 12804 22192 12832
rect 22186 12792 22192 12804
rect 22244 12792 22250 12844
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12832 22339 12835
rect 22370 12832 22376 12844
rect 22327 12804 22376 12832
rect 22327 12801 22339 12804
rect 22281 12795 22339 12801
rect 22370 12792 22376 12804
rect 22428 12792 22434 12844
rect 22464 12835 22522 12841
rect 22464 12801 22476 12835
rect 22510 12801 22522 12835
rect 22464 12795 22522 12801
rect 22557 12835 22615 12841
rect 22557 12801 22569 12835
rect 22603 12832 22615 12835
rect 22738 12832 22744 12844
rect 22603 12804 22744 12832
rect 22603 12801 22615 12804
rect 22557 12795 22615 12801
rect 21450 12764 21456 12776
rect 21411 12736 21456 12764
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 21726 12724 21732 12776
rect 21784 12764 21790 12776
rect 21913 12767 21971 12773
rect 21913 12764 21925 12767
rect 21784 12736 21925 12764
rect 21784 12724 21790 12736
rect 21913 12733 21925 12736
rect 21959 12764 21971 12767
rect 22480 12764 22508 12795
rect 22738 12792 22744 12804
rect 22796 12792 22802 12844
rect 22833 12835 22891 12841
rect 22833 12801 22845 12835
rect 22879 12832 22891 12835
rect 23130 12835 23188 12841
rect 22879 12804 23060 12832
rect 22879 12801 22891 12804
rect 22833 12795 22891 12801
rect 21959 12736 22508 12764
rect 22649 12767 22707 12773
rect 21959 12733 21971 12736
rect 21913 12727 21971 12733
rect 22649 12733 22661 12767
rect 22695 12764 22707 12767
rect 22922 12764 22928 12776
rect 22695 12736 22928 12764
rect 22695 12733 22707 12736
rect 22649 12727 22707 12733
rect 22922 12724 22928 12736
rect 22980 12724 22986 12776
rect 23032 12764 23060 12804
rect 23130 12801 23142 12835
rect 23176 12832 23188 12835
rect 23290 12832 23296 12844
rect 23176 12804 23296 12832
rect 23176 12801 23188 12804
rect 23130 12795 23188 12801
rect 23290 12792 23296 12804
rect 23348 12792 23354 12844
rect 23474 12832 23480 12844
rect 23435 12804 23480 12832
rect 23474 12792 23480 12804
rect 23532 12792 23538 12844
rect 23658 12832 23664 12844
rect 23619 12804 23664 12832
rect 23658 12792 23664 12804
rect 23716 12792 23722 12844
rect 23768 12841 23796 12872
rect 23998 12869 24010 12872
rect 24044 12869 24056 12903
rect 23998 12863 24056 12869
rect 23753 12835 23811 12841
rect 23753 12801 23765 12835
rect 23799 12801 23811 12835
rect 23753 12795 23811 12801
rect 23032 12736 23796 12764
rect 20272 12668 20668 12696
rect 21545 12699 21603 12705
rect 19794 12628 19800 12640
rect 17144 12600 19800 12628
rect 17037 12591 17095 12597
rect 19794 12588 19800 12600
rect 19852 12628 19858 12640
rect 20272 12628 20300 12668
rect 21545 12665 21557 12699
rect 21591 12696 21603 12699
rect 22738 12696 22744 12708
rect 21591 12668 22744 12696
rect 21591 12665 21603 12668
rect 21545 12659 21603 12665
rect 22738 12656 22744 12668
rect 22796 12656 22802 12708
rect 23014 12656 23020 12708
rect 23072 12696 23078 12708
rect 23201 12699 23259 12705
rect 23201 12696 23213 12699
rect 23072 12668 23213 12696
rect 23072 12656 23078 12668
rect 23201 12665 23213 12668
rect 23247 12665 23259 12699
rect 23201 12659 23259 12665
rect 19852 12600 20300 12628
rect 21913 12631 21971 12637
rect 19852 12588 19858 12600
rect 21913 12597 21925 12631
rect 21959 12628 21971 12631
rect 22005 12631 22063 12637
rect 22005 12628 22017 12631
rect 21959 12600 22017 12628
rect 21959 12597 21971 12600
rect 21913 12591 21971 12597
rect 22005 12597 22017 12600
rect 22051 12597 22063 12631
rect 23768 12628 23796 12736
rect 25130 12628 25136 12640
rect 23768 12600 25136 12628
rect 22005 12591 22063 12597
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 1104 12538 26220 12560
rect 1104 12486 5136 12538
rect 5188 12486 5200 12538
rect 5252 12486 5264 12538
rect 5316 12486 5328 12538
rect 5380 12486 5392 12538
rect 5444 12486 13508 12538
rect 13560 12486 13572 12538
rect 13624 12486 13636 12538
rect 13688 12486 13700 12538
rect 13752 12486 13764 12538
rect 13816 12486 21880 12538
rect 21932 12486 21944 12538
rect 21996 12486 22008 12538
rect 22060 12486 22072 12538
rect 22124 12486 22136 12538
rect 22188 12486 26220 12538
rect 1104 12464 26220 12486
rect 2314 12424 2320 12436
rect 2275 12396 2320 12424
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 3142 12424 3148 12436
rect 2823 12396 3148 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 3326 12424 3332 12436
rect 3287 12396 3332 12424
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 4798 12384 4804 12436
rect 4856 12384 4862 12436
rect 4982 12384 4988 12436
rect 5040 12424 5046 12436
rect 5261 12427 5319 12433
rect 5261 12424 5273 12427
rect 5040 12396 5273 12424
rect 5040 12384 5046 12396
rect 5261 12393 5273 12396
rect 5307 12393 5319 12427
rect 5261 12387 5319 12393
rect 5445 12427 5503 12433
rect 5445 12393 5457 12427
rect 5491 12424 5503 12427
rect 5534 12424 5540 12436
rect 5491 12396 5540 12424
rect 5491 12393 5503 12396
rect 5445 12387 5503 12393
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 5902 12384 5908 12436
rect 5960 12424 5966 12436
rect 6549 12427 6607 12433
rect 6549 12424 6561 12427
rect 5960 12396 6561 12424
rect 5960 12384 5966 12396
rect 6549 12393 6561 12396
rect 6595 12424 6607 12427
rect 7650 12424 7656 12436
rect 6595 12396 7656 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 7926 12424 7932 12436
rect 7887 12396 7932 12424
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 8205 12427 8263 12433
rect 8205 12424 8217 12427
rect 8076 12396 8217 12424
rect 8076 12384 8082 12396
rect 8205 12393 8217 12396
rect 8251 12393 8263 12427
rect 8478 12424 8484 12436
rect 8439 12396 8484 12424
rect 8205 12387 8263 12393
rect 8478 12384 8484 12396
rect 8536 12424 8542 12436
rect 8665 12427 8723 12433
rect 8665 12424 8677 12427
rect 8536 12396 8677 12424
rect 8536 12384 8542 12396
rect 8665 12393 8677 12396
rect 8711 12393 8723 12427
rect 8665 12387 8723 12393
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 9493 12427 9551 12433
rect 9493 12424 9505 12427
rect 9456 12396 9505 12424
rect 9456 12384 9462 12396
rect 9493 12393 9505 12396
rect 9539 12393 9551 12427
rect 9493 12387 9551 12393
rect 10318 12384 10324 12436
rect 10376 12424 10382 12436
rect 12342 12424 12348 12436
rect 10376 12396 12348 12424
rect 10376 12384 10382 12396
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 14826 12384 14832 12436
rect 14884 12424 14890 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 14884 12396 14933 12424
rect 14884 12384 14890 12396
rect 14921 12393 14933 12396
rect 14967 12393 14979 12427
rect 16942 12424 16948 12436
rect 16903 12396 16948 12424
rect 14921 12387 14979 12393
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 18601 12427 18659 12433
rect 18601 12393 18613 12427
rect 18647 12424 18659 12427
rect 20346 12424 20352 12436
rect 18647 12396 20352 12424
rect 18647 12393 18659 12396
rect 18601 12387 18659 12393
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 4816 12356 4844 12384
rect 6181 12359 6239 12365
rect 6181 12356 6193 12359
rect 2924 12328 3004 12356
rect 4816 12328 6193 12356
rect 2924 12316 2930 12328
rect 2682 12288 2688 12300
rect 2516 12260 2688 12288
rect 2516 12229 2544 12260
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 2976 12297 3004 12328
rect 6181 12325 6193 12328
rect 6227 12325 6239 12359
rect 6181 12319 6239 12325
rect 6270 12316 6276 12368
rect 6328 12356 6334 12368
rect 10962 12356 10968 12368
rect 6328 12328 10968 12356
rect 6328 12316 6334 12328
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 14734 12316 14740 12368
rect 14792 12356 14798 12368
rect 16666 12356 16672 12368
rect 14792 12328 16672 12356
rect 14792 12316 14798 12328
rect 2961 12291 3019 12297
rect 2961 12257 2973 12291
rect 3007 12257 3019 12291
rect 2961 12251 3019 12257
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 7558 12288 7564 12300
rect 4948 12260 7564 12288
rect 4948 12248 4954 12260
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 10137 12291 10195 12297
rect 10137 12288 10149 12291
rect 8536 12260 10149 12288
rect 8536 12248 8542 12260
rect 10137 12257 10149 12260
rect 10183 12288 10195 12291
rect 10413 12291 10471 12297
rect 10413 12288 10425 12291
rect 10183 12260 10425 12288
rect 10183 12257 10195 12260
rect 10137 12251 10195 12257
rect 10413 12257 10425 12260
rect 10459 12257 10471 12291
rect 11238 12288 11244 12300
rect 11199 12260 11244 12288
rect 10413 12251 10471 12257
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 14829 12291 14887 12297
rect 14829 12257 14841 12291
rect 14875 12288 14887 12291
rect 15010 12288 15016 12300
rect 14875 12260 15016 12288
rect 14875 12257 14887 12260
rect 14829 12251 14887 12257
rect 15010 12248 15016 12260
rect 15068 12288 15074 12300
rect 15473 12291 15531 12297
rect 15473 12288 15485 12291
rect 15068 12260 15485 12288
rect 15068 12248 15074 12260
rect 15473 12257 15485 12260
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12189 2559 12223
rect 2501 12183 2559 12189
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12189 2651 12223
rect 2593 12183 2651 12189
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 3050 12220 3056 12232
rect 2915 12192 3056 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 2608 12152 2636 12183
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12220 3203 12223
rect 3234 12220 3240 12232
rect 3191 12192 3240 12220
rect 3191 12189 3203 12192
rect 3145 12183 3203 12189
rect 3234 12180 3240 12192
rect 3292 12220 3298 12232
rect 3418 12220 3424 12232
rect 3292 12192 3424 12220
rect 3292 12180 3298 12192
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3878 12220 3884 12232
rect 3839 12192 3884 12220
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 4154 12229 4160 12232
rect 4148 12183 4160 12229
rect 4212 12220 4218 12232
rect 5626 12220 5632 12232
rect 4212 12192 4248 12220
rect 5539 12192 5632 12220
rect 4154 12180 4160 12183
rect 4212 12180 4218 12192
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 5718 12180 5724 12232
rect 5776 12220 5782 12232
rect 5776 12192 6132 12220
rect 5776 12180 5782 12192
rect 2682 12152 2688 12164
rect 2608 12124 2688 12152
rect 2682 12112 2688 12124
rect 2740 12112 2746 12164
rect 3896 12152 3924 12180
rect 4706 12152 4712 12164
rect 3896 12124 4712 12152
rect 4706 12112 4712 12124
rect 4764 12112 4770 12164
rect 5644 12084 5672 12180
rect 5902 12152 5908 12164
rect 5863 12124 5908 12152
rect 5902 12112 5908 12124
rect 5960 12112 5966 12164
rect 6104 12161 6132 12192
rect 6178 12180 6184 12232
rect 6236 12220 6242 12232
rect 6365 12223 6423 12229
rect 6365 12220 6377 12223
rect 6236 12192 6377 12220
rect 6236 12180 6242 12192
rect 6365 12189 6377 12192
rect 6411 12220 6423 12223
rect 8389 12223 8447 12229
rect 6411 12192 7972 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6089 12155 6147 12161
rect 6089 12121 6101 12155
rect 6135 12152 6147 12155
rect 7837 12155 7895 12161
rect 7837 12152 7849 12155
rect 6135 12124 7849 12152
rect 6135 12121 6147 12124
rect 6089 12115 6147 12121
rect 7837 12121 7849 12124
rect 7883 12121 7895 12155
rect 7944 12152 7972 12192
rect 8389 12189 8401 12223
rect 8435 12220 8447 12223
rect 8938 12220 8944 12232
rect 8435 12192 8944 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 9180 12192 9413 12220
rect 9180 12180 9186 12192
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12220 9919 12223
rect 10318 12220 10324 12232
rect 9907 12192 10324 12220
rect 9907 12189 9919 12192
rect 9861 12183 9919 12189
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10502 12180 10508 12232
rect 10560 12220 10566 12232
rect 10873 12223 10931 12229
rect 10873 12220 10885 12223
rect 10560 12192 10885 12220
rect 10560 12180 10566 12192
rect 10873 12189 10885 12192
rect 10919 12189 10931 12223
rect 11038 12223 11096 12229
rect 11038 12220 11050 12223
rect 10873 12183 10931 12189
rect 10980 12192 11050 12220
rect 10226 12152 10232 12164
rect 7944 12124 10232 12152
rect 7837 12115 7895 12121
rect 10226 12112 10232 12124
rect 10284 12112 10290 12164
rect 10980 12152 11008 12192
rect 11038 12189 11050 12192
rect 11084 12189 11096 12223
rect 11038 12183 11096 12189
rect 11146 12180 11152 12232
rect 11204 12220 11210 12232
rect 11425 12223 11483 12229
rect 11204 12192 11249 12220
rect 11204 12180 11210 12192
rect 11425 12189 11437 12223
rect 11471 12220 11483 12223
rect 11701 12223 11759 12229
rect 11471 12192 11560 12220
rect 11471 12189 11483 12192
rect 11425 12183 11483 12189
rect 10704 12124 11008 12152
rect 10704 12096 10732 12124
rect 6270 12084 6276 12096
rect 5644 12056 6276 12084
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 9122 12084 9128 12096
rect 9083 12056 9128 12084
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 9950 12084 9956 12096
rect 9272 12056 9317 12084
rect 9911 12056 9956 12084
rect 9272 12044 9278 12056
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 10686 12084 10692 12096
rect 10647 12056 10692 12084
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 11532 12084 11560 12192
rect 11701 12189 11713 12223
rect 11747 12220 11759 12223
rect 12434 12220 12440 12232
rect 11747 12192 12440 12220
rect 11747 12189 11759 12192
rect 11701 12183 11759 12189
rect 12434 12180 12440 12192
rect 12492 12180 12498 12232
rect 15286 12220 15292 12232
rect 15247 12192 15292 12220
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 15378 12180 15384 12232
rect 15436 12220 15442 12232
rect 15948 12229 15976 12328
rect 16666 12316 16672 12328
rect 16724 12316 16730 12368
rect 17494 12316 17500 12368
rect 17552 12356 17558 12368
rect 17678 12356 17684 12368
rect 17552 12328 17684 12356
rect 17552 12316 17558 12328
rect 17678 12316 17684 12328
rect 17736 12356 17742 12368
rect 18230 12356 18236 12368
rect 17736 12328 18236 12356
rect 17736 12316 17742 12328
rect 18230 12316 18236 12328
rect 18288 12316 18294 12368
rect 16390 12288 16396 12300
rect 16351 12260 16396 12288
rect 16390 12248 16396 12260
rect 16448 12248 16454 12300
rect 18322 12288 18328 12300
rect 17144 12260 18328 12288
rect 15933 12223 15991 12229
rect 15436 12192 15481 12220
rect 15436 12180 15442 12192
rect 15933 12189 15945 12223
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 16485 12223 16543 12229
rect 16485 12189 16497 12223
rect 16531 12220 16543 12223
rect 16574 12220 16580 12232
rect 16531 12192 16580 12220
rect 16531 12189 16543 12192
rect 16485 12183 16543 12189
rect 11609 12155 11667 12161
rect 11609 12121 11621 12155
rect 11655 12152 11667 12155
rect 11946 12155 12004 12161
rect 11946 12152 11958 12155
rect 11655 12124 11958 12152
rect 11655 12121 11667 12124
rect 11609 12115 11667 12121
rect 11946 12121 11958 12124
rect 11992 12121 12004 12155
rect 15396 12152 15424 12180
rect 16040 12152 16068 12183
rect 16574 12180 16580 12192
rect 16632 12220 16638 12232
rect 16758 12220 16764 12232
rect 16632 12192 16764 12220
rect 16632 12180 16638 12192
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17144 12229 17172 12260
rect 18322 12248 18328 12260
rect 18380 12248 18386 12300
rect 17129 12223 17187 12229
rect 17129 12189 17141 12223
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 17313 12223 17371 12229
rect 17313 12220 17325 12223
rect 17276 12192 17325 12220
rect 17276 12180 17282 12192
rect 17313 12189 17325 12192
rect 17359 12189 17371 12223
rect 17313 12183 17371 12189
rect 17494 12180 17500 12232
rect 17552 12220 17558 12232
rect 17589 12223 17647 12229
rect 17589 12220 17601 12223
rect 17552 12192 17601 12220
rect 17552 12180 17558 12192
rect 17589 12189 17601 12192
rect 17635 12189 17647 12223
rect 17589 12183 17647 12189
rect 17034 12152 17040 12164
rect 15396 12124 16068 12152
rect 16995 12124 17040 12152
rect 11946 12115 12004 12121
rect 17034 12112 17040 12124
rect 17092 12112 17098 12164
rect 17604 12152 17632 12183
rect 17678 12180 17684 12232
rect 17736 12220 17742 12232
rect 18048 12223 18106 12229
rect 17736 12192 17781 12220
rect 17736 12180 17742 12192
rect 18048 12189 18060 12223
rect 18094 12220 18106 12223
rect 18616 12220 18644 12387
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 21266 12424 21272 12436
rect 21227 12396 21272 12424
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 21634 12424 21640 12436
rect 21595 12396 21640 12424
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 22373 12427 22431 12433
rect 22373 12424 22385 12427
rect 22020 12396 22385 12424
rect 19518 12316 19524 12368
rect 19576 12316 19582 12368
rect 20162 12316 20168 12368
rect 20220 12356 20226 12368
rect 20220 12328 21128 12356
rect 20220 12316 20226 12328
rect 19536 12288 19564 12316
rect 20533 12291 20591 12297
rect 19536 12260 20208 12288
rect 18094 12192 18644 12220
rect 19521 12223 19579 12229
rect 18094 12189 18106 12192
rect 18048 12183 18106 12189
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 19702 12220 19708 12232
rect 19567 12192 19708 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 19702 12180 19708 12192
rect 19760 12180 19766 12232
rect 19978 12220 19984 12232
rect 19939 12192 19984 12220
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 20180 12229 20208 12260
rect 20533 12257 20545 12291
rect 20579 12288 20591 12291
rect 20990 12288 20996 12300
rect 20579 12260 20996 12288
rect 20579 12257 20591 12260
rect 20533 12251 20591 12257
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 21100 12288 21128 12328
rect 21450 12316 21456 12368
rect 21508 12356 21514 12368
rect 21913 12359 21971 12365
rect 21913 12356 21925 12359
rect 21508 12328 21925 12356
rect 21508 12316 21514 12328
rect 21913 12325 21925 12328
rect 21959 12325 21971 12359
rect 21913 12319 21971 12325
rect 22020 12288 22048 12396
rect 22373 12393 22385 12396
rect 22419 12424 22431 12427
rect 22419 12396 23060 12424
rect 22419 12393 22431 12396
rect 22373 12387 22431 12393
rect 22462 12356 22468 12368
rect 22423 12328 22468 12356
rect 22462 12316 22468 12328
rect 22520 12316 22526 12368
rect 22830 12316 22836 12368
rect 22888 12356 22894 12368
rect 22888 12328 22968 12356
rect 22888 12316 22894 12328
rect 22940 12297 22968 12328
rect 23032 12297 23060 12396
rect 21100 12260 22048 12288
rect 22925 12291 22983 12297
rect 22925 12257 22937 12291
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 23017 12291 23075 12297
rect 23017 12257 23029 12291
rect 23063 12257 23075 12291
rect 23017 12251 23075 12257
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12220 20223 12223
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 20211 12192 20637 12220
rect 20211 12189 20223 12192
rect 20165 12183 20223 12189
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 20809 12223 20867 12229
rect 20809 12189 20821 12223
rect 20855 12220 20867 12223
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 20855 12192 21281 12220
rect 20855 12189 20867 12192
rect 20809 12183 20867 12189
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 21269 12183 21327 12189
rect 21453 12223 21511 12229
rect 21453 12189 21465 12223
rect 21499 12220 21511 12223
rect 21726 12220 21732 12232
rect 21499 12192 21732 12220
rect 21499 12189 21511 12192
rect 21453 12183 21511 12189
rect 18325 12155 18383 12161
rect 18325 12152 18337 12155
rect 17604 12124 18337 12152
rect 18325 12121 18337 12124
rect 18371 12121 18383 12155
rect 18325 12115 18383 12121
rect 18509 12155 18567 12161
rect 18509 12121 18521 12155
rect 18555 12121 18567 12155
rect 19996 12152 20024 12180
rect 20824 12152 20852 12183
rect 21726 12180 21732 12192
rect 21784 12220 21790 12232
rect 22005 12223 22063 12229
rect 22005 12220 22017 12223
rect 21784 12192 22017 12220
rect 21784 12180 21790 12192
rect 22005 12189 22017 12192
rect 22051 12189 22063 12223
rect 22005 12183 22063 12189
rect 22646 12180 22652 12232
rect 22704 12220 22710 12232
rect 22833 12223 22891 12229
rect 22833 12220 22845 12223
rect 22704 12192 22845 12220
rect 22704 12180 22710 12192
rect 22833 12189 22845 12192
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 19996 12124 20852 12152
rect 18509 12115 18567 12121
rect 12342 12084 12348 12096
rect 11532 12056 12348 12084
rect 12342 12044 12348 12056
rect 12400 12084 12406 12096
rect 13081 12087 13139 12093
rect 13081 12084 13093 12087
rect 12400 12056 13093 12084
rect 12400 12044 12406 12056
rect 13081 12053 13093 12056
rect 13127 12053 13139 12087
rect 13081 12047 13139 12053
rect 15841 12087 15899 12093
rect 15841 12053 15853 12087
rect 15887 12084 15899 12087
rect 15930 12084 15936 12096
rect 15887 12056 15936 12084
rect 15887 12053 15899 12056
rect 15841 12047 15899 12053
rect 15930 12044 15936 12056
rect 15988 12044 15994 12096
rect 16482 12044 16488 12096
rect 16540 12084 16546 12096
rect 16577 12087 16635 12093
rect 16577 12084 16589 12087
rect 16540 12056 16589 12084
rect 16540 12044 16546 12056
rect 16577 12053 16589 12056
rect 16623 12084 16635 12087
rect 16758 12084 16764 12096
rect 16623 12056 16764 12084
rect 16623 12053 16635 12056
rect 16577 12047 16635 12053
rect 16758 12044 16764 12056
rect 16816 12044 16822 12096
rect 18046 12044 18052 12096
rect 18104 12084 18110 12096
rect 18141 12087 18199 12093
rect 18141 12084 18153 12087
rect 18104 12056 18153 12084
rect 18104 12044 18110 12056
rect 18141 12053 18153 12056
rect 18187 12053 18199 12087
rect 18141 12047 18199 12053
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 18524 12084 18552 12115
rect 18288 12056 18552 12084
rect 19337 12087 19395 12093
rect 18288 12044 18294 12056
rect 19337 12053 19349 12087
rect 19383 12084 19395 12087
rect 19886 12084 19892 12096
rect 19383 12056 19892 12084
rect 19383 12053 19395 12056
rect 19337 12047 19395 12053
rect 19886 12044 19892 12056
rect 19944 12044 19950 12096
rect 20346 12044 20352 12096
rect 20404 12084 20410 12096
rect 20441 12087 20499 12093
rect 20441 12084 20453 12087
rect 20404 12056 20453 12084
rect 20404 12044 20410 12056
rect 20441 12053 20453 12056
rect 20487 12053 20499 12087
rect 20441 12047 20499 12053
rect 1104 11994 26220 12016
rect 1104 11942 9322 11994
rect 9374 11942 9386 11994
rect 9438 11942 9450 11994
rect 9502 11942 9514 11994
rect 9566 11942 9578 11994
rect 9630 11942 17694 11994
rect 17746 11942 17758 11994
rect 17810 11942 17822 11994
rect 17874 11942 17886 11994
rect 17938 11942 17950 11994
rect 18002 11942 26220 11994
rect 1104 11920 26220 11942
rect 2866 11880 2872 11892
rect 2827 11852 2872 11880
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 5166 11880 5172 11892
rect 4488 11852 5172 11880
rect 4488 11840 4494 11852
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 7098 11880 7104 11892
rect 5316 11852 7104 11880
rect 5316 11840 5322 11852
rect 7098 11840 7104 11852
rect 7156 11880 7162 11892
rect 7193 11883 7251 11889
rect 7193 11880 7205 11883
rect 7156 11852 7205 11880
rect 7156 11840 7162 11852
rect 7193 11849 7205 11852
rect 7239 11849 7251 11883
rect 7193 11843 7251 11849
rect 9401 11883 9459 11889
rect 9401 11849 9413 11883
rect 9447 11880 9459 11883
rect 10413 11883 10471 11889
rect 9447 11852 10364 11880
rect 9447 11849 9459 11852
rect 9401 11843 9459 11849
rect 1486 11772 1492 11824
rect 1544 11812 1550 11824
rect 3878 11812 3884 11824
rect 1544 11784 3884 11812
rect 1544 11772 1550 11784
rect 1756 11747 1814 11753
rect 1756 11713 1768 11747
rect 1802 11744 1814 11747
rect 2314 11744 2320 11756
rect 1802 11716 2320 11744
rect 1802 11713 1814 11716
rect 1756 11707 1814 11713
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 3803 11753 3831 11784
rect 3878 11772 3884 11784
rect 3936 11772 3942 11824
rect 9582 11772 9588 11824
rect 9640 11812 9646 11824
rect 9950 11812 9956 11824
rect 9640 11784 9956 11812
rect 9640 11772 9646 11784
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10045 11815 10103 11821
rect 10045 11781 10057 11815
rect 10091 11781 10103 11815
rect 10045 11775 10103 11781
rect 10229 11815 10287 11821
rect 10229 11781 10241 11815
rect 10275 11781 10287 11815
rect 10336 11812 10364 11852
rect 10413 11849 10425 11883
rect 10459 11880 10471 11883
rect 11054 11880 11060 11892
rect 10459 11852 11060 11880
rect 10459 11849 10471 11852
rect 10413 11843 10471 11849
rect 11054 11840 11060 11852
rect 11112 11840 11118 11892
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 13357 11883 13415 11889
rect 13357 11880 13369 11883
rect 11388 11852 13369 11880
rect 11388 11840 11394 11852
rect 13357 11849 13369 11852
rect 13403 11880 13415 11883
rect 16390 11880 16396 11892
rect 13403 11852 14872 11880
rect 16351 11852 16396 11880
rect 13403 11849 13415 11852
rect 13357 11843 13415 11849
rect 11698 11812 11704 11824
rect 10336 11784 11704 11812
rect 10229 11775 10287 11781
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 4056 11747 4114 11753
rect 4056 11713 4068 11747
rect 4102 11744 4114 11747
rect 4522 11744 4528 11756
rect 4102 11716 4528 11744
rect 4102 11713 4114 11716
rect 4056 11707 4114 11713
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 5350 11744 5356 11756
rect 5311 11716 5356 11744
rect 5350 11704 5356 11716
rect 5408 11704 5414 11756
rect 5445 11747 5503 11753
rect 5445 11713 5457 11747
rect 5491 11744 5503 11747
rect 5813 11747 5871 11753
rect 5813 11744 5825 11747
rect 5491 11716 5825 11744
rect 5491 11713 5503 11716
rect 5445 11707 5503 11713
rect 5813 11713 5825 11716
rect 5859 11744 5871 11747
rect 6178 11744 6184 11756
rect 5859 11716 6184 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 6822 11744 6828 11756
rect 6783 11716 6828 11744
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11713 6975 11747
rect 6917 11707 6975 11713
rect 1486 11676 1492 11688
rect 1447 11648 1492 11676
rect 1486 11636 1492 11648
rect 1544 11636 1550 11688
rect 4798 11636 4804 11688
rect 4856 11676 4862 11688
rect 5258 11676 5264 11688
rect 4856 11648 5264 11676
rect 4856 11636 4862 11648
rect 5258 11636 5264 11648
rect 5316 11636 5322 11688
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 6932 11676 6960 11707
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 9548 11716 9593 11744
rect 9548 11704 9554 11716
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10060 11744 10088 11775
rect 9916 11716 10088 11744
rect 9916 11704 9922 11716
rect 5592 11648 6960 11676
rect 7101 11679 7159 11685
rect 5592 11636 5598 11648
rect 7101 11645 7113 11679
rect 7147 11676 7159 11679
rect 8018 11676 8024 11688
rect 7147 11648 8024 11676
rect 7147 11645 7159 11648
rect 7101 11639 7159 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 9456 11648 9689 11676
rect 9456 11636 9462 11648
rect 9677 11645 9689 11648
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 9766 11636 9772 11688
rect 9824 11676 9830 11688
rect 10244 11676 10272 11775
rect 11698 11772 11704 11784
rect 11756 11772 11762 11824
rect 12434 11812 12440 11824
rect 11992 11784 12440 11812
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11744 10655 11747
rect 10778 11744 10784 11756
rect 10643 11716 10784 11744
rect 10643 11713 10655 11716
rect 10597 11707 10655 11713
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11744 10931 11747
rect 11882 11744 11888 11756
rect 10919 11716 11888 11744
rect 10919 11713 10931 11716
rect 10873 11707 10931 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 11992 11753 12020 11784
rect 12434 11772 12440 11784
rect 12492 11812 12498 11824
rect 13541 11815 13599 11821
rect 13541 11812 13553 11815
rect 12492 11784 13553 11812
rect 12492 11772 12498 11784
rect 13541 11781 13553 11784
rect 13587 11781 13599 11815
rect 13541 11775 13599 11781
rect 12250 11753 12256 11756
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11713 12035 11747
rect 12244 11744 12256 11753
rect 12211 11716 12256 11744
rect 11977 11707 12035 11713
rect 12244 11707 12256 11716
rect 12250 11704 12256 11707
rect 12308 11704 12314 11756
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11744 13783 11747
rect 13906 11744 13912 11756
rect 13771 11716 13912 11744
rect 13771 11713 13783 11716
rect 13725 11707 13783 11713
rect 13906 11704 13912 11716
rect 13964 11704 13970 11756
rect 11606 11676 11612 11688
rect 9824 11648 11612 11676
rect 9824 11636 9830 11648
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 14844 11676 14872 11852
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 16850 11840 16856 11892
rect 16908 11840 16914 11892
rect 17586 11840 17592 11892
rect 17644 11880 17650 11892
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 17644 11852 17693 11880
rect 17644 11840 17650 11852
rect 17681 11849 17693 11852
rect 17727 11849 17739 11883
rect 17681 11843 17739 11849
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 20441 11883 20499 11889
rect 20441 11880 20453 11883
rect 20036 11852 20453 11880
rect 20036 11840 20042 11852
rect 20441 11849 20453 11852
rect 20487 11849 20499 11883
rect 20441 11843 20499 11849
rect 22925 11883 22983 11889
rect 22925 11849 22937 11883
rect 22971 11880 22983 11883
rect 23106 11880 23112 11892
rect 22971 11852 23112 11880
rect 22971 11849 22983 11852
rect 22925 11843 22983 11849
rect 23106 11840 23112 11852
rect 23164 11880 23170 11892
rect 23382 11880 23388 11892
rect 23164 11852 23388 11880
rect 23164 11840 23170 11852
rect 23382 11840 23388 11852
rect 23440 11840 23446 11892
rect 16666 11812 16672 11824
rect 14936 11784 16672 11812
rect 14936 11753 14964 11784
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 16868 11812 16896 11840
rect 17494 11812 17500 11824
rect 16776 11784 17500 11812
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 15105 11747 15163 11753
rect 15105 11713 15117 11747
rect 15151 11744 15163 11747
rect 15378 11744 15384 11756
rect 15151 11716 15384 11744
rect 15151 11713 15163 11716
rect 15105 11707 15163 11713
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11744 15531 11747
rect 15930 11744 15936 11756
rect 15519 11716 15936 11744
rect 15519 11713 15531 11716
rect 15473 11707 15531 11713
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16776 11744 16804 11784
rect 17494 11772 17500 11784
rect 17552 11772 17558 11824
rect 16347 11716 16804 11744
rect 16853 11747 16911 11753
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16853 11713 16865 11747
rect 16899 11744 16911 11747
rect 17034 11744 17040 11756
rect 16899 11716 17040 11744
rect 16899 11713 16911 11716
rect 16853 11707 16911 11713
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 17218 11744 17224 11756
rect 17179 11716 17224 11744
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 17586 11744 17592 11756
rect 17547 11716 17592 11744
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 18046 11744 18052 11756
rect 18007 11716 18052 11744
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 20346 11744 20352 11756
rect 20307 11716 20352 11744
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11744 20683 11747
rect 20806 11744 20812 11756
rect 20671 11716 20812 11744
rect 20671 11713 20683 11716
rect 20625 11707 20683 11713
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 23014 11744 23020 11756
rect 22975 11716 23020 11744
rect 23014 11704 23020 11716
rect 23072 11704 23078 11756
rect 15838 11676 15844 11688
rect 14844 11648 15700 11676
rect 15799 11648 15844 11676
rect 4982 11568 4988 11620
rect 5040 11608 5046 11620
rect 15381 11611 15439 11617
rect 5040 11580 10823 11608
rect 5040 11568 5046 11580
rect 5626 11540 5632 11552
rect 5587 11512 5632 11540
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 8662 11500 8668 11552
rect 8720 11540 8726 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8720 11512 9045 11540
rect 8720 11500 8726 11512
rect 9033 11509 9045 11512
rect 9079 11509 9091 11543
rect 9033 11503 9091 11509
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 9582 11540 9588 11552
rect 9456 11512 9588 11540
rect 9456 11500 9462 11512
rect 9582 11500 9588 11512
rect 9640 11540 9646 11552
rect 9861 11543 9919 11549
rect 9861 11540 9873 11543
rect 9640 11512 9873 11540
rect 9640 11500 9646 11512
rect 9861 11509 9873 11512
rect 9907 11509 9919 11543
rect 10226 11540 10232 11552
rect 10187 11512 10232 11540
rect 9861 11503 9919 11509
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 10597 11543 10655 11549
rect 10597 11509 10609 11543
rect 10643 11540 10655 11543
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 10643 11512 10701 11540
rect 10643 11509 10655 11512
rect 10597 11503 10655 11509
rect 10689 11509 10701 11512
rect 10735 11509 10747 11543
rect 10795 11540 10823 11580
rect 13280 11580 13584 11608
rect 13280 11540 13308 11580
rect 10795 11512 13308 11540
rect 13556 11540 13584 11580
rect 15381 11577 15393 11611
rect 15427 11608 15439 11611
rect 15562 11608 15568 11620
rect 15427 11580 15568 11608
rect 15427 11577 15439 11580
rect 15381 11571 15439 11577
rect 15562 11568 15568 11580
rect 15620 11568 15626 11620
rect 15672 11608 15700 11648
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11676 17463 11679
rect 18322 11676 18328 11688
rect 17451 11648 18328 11676
rect 17451 11645 17463 11648
rect 17405 11639 17463 11645
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 16942 11608 16948 11620
rect 15672 11580 16804 11608
rect 16903 11580 16948 11608
rect 15470 11540 15476 11552
rect 13556 11512 15476 11540
rect 10689 11503 10747 11509
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 16209 11543 16267 11549
rect 16209 11509 16221 11543
rect 16255 11540 16267 11543
rect 16666 11540 16672 11552
rect 16255 11512 16672 11540
rect 16255 11509 16267 11512
rect 16209 11503 16267 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 16776 11540 16804 11580
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 17310 11568 17316 11620
rect 17368 11608 17374 11620
rect 17865 11611 17923 11617
rect 17865 11608 17877 11611
rect 17368 11580 17877 11608
rect 17368 11568 17374 11580
rect 17865 11577 17877 11580
rect 17911 11577 17923 11611
rect 17865 11571 17923 11577
rect 17402 11540 17408 11552
rect 16776 11512 17408 11540
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 20257 11543 20315 11549
rect 20257 11509 20269 11543
rect 20303 11540 20315 11543
rect 20622 11540 20628 11552
rect 20303 11512 20628 11540
rect 20303 11509 20315 11512
rect 20257 11503 20315 11509
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 1104 11450 26220 11472
rect 1104 11398 5136 11450
rect 5188 11398 5200 11450
rect 5252 11398 5264 11450
rect 5316 11398 5328 11450
rect 5380 11398 5392 11450
rect 5444 11398 13508 11450
rect 13560 11398 13572 11450
rect 13624 11398 13636 11450
rect 13688 11398 13700 11450
rect 13752 11398 13764 11450
rect 13816 11398 21880 11450
rect 21932 11398 21944 11450
rect 21996 11398 22008 11450
rect 22060 11398 22072 11450
rect 22124 11398 22136 11450
rect 22188 11398 26220 11450
rect 1104 11376 26220 11398
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 2372 11308 2421 11336
rect 2372 11296 2378 11308
rect 2409 11305 2421 11308
rect 2455 11305 2467 11339
rect 2866 11336 2872 11348
rect 2409 11299 2467 11305
rect 2746 11308 2872 11336
rect 2746 11268 2774 11308
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 4522 11336 4528 11348
rect 4483 11308 4528 11336
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 7466 11336 7472 11348
rect 5828 11308 7052 11336
rect 7379 11308 7472 11336
rect 2608 11240 2774 11268
rect 2608 11141 2636 11240
rect 2866 11200 2872 11212
rect 2827 11172 2872 11200
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 2961 11203 3019 11209
rect 2961 11169 2973 11203
rect 3007 11200 3019 11203
rect 3050 11200 3056 11212
rect 3007 11172 3056 11200
rect 3007 11169 3019 11172
rect 2961 11163 3019 11169
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 3510 11160 3516 11212
rect 3568 11200 3574 11212
rect 3568 11172 3924 11200
rect 3568 11160 3574 11172
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11101 2651 11135
rect 2593 11095 2651 11101
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 2774 11132 2780 11144
rect 2731 11104 2780 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 2774 11092 2780 11104
rect 2832 11132 2838 11144
rect 3694 11132 3700 11144
rect 2832 11104 3700 11132
rect 2832 11092 2838 11104
rect 3694 11092 3700 11104
rect 3752 11092 3758 11144
rect 3896 11141 3924 11172
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4157 11203 4215 11209
rect 4157 11200 4169 11203
rect 4028 11172 4169 11200
rect 4028 11160 4034 11172
rect 4157 11169 4169 11172
rect 4203 11169 4215 11203
rect 4157 11163 4215 11169
rect 4614 11160 4620 11212
rect 4672 11200 4678 11212
rect 5626 11200 5632 11212
rect 4672 11172 5488 11200
rect 5587 11172 5632 11200
rect 4672 11160 4678 11172
rect 3881 11135 3939 11141
rect 3881 11101 3893 11135
rect 3927 11101 3939 11135
rect 3881 11095 3939 11101
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4249 11135 4307 11141
rect 4120 11104 4164 11132
rect 4120 11092 4126 11104
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4430 11132 4436 11144
rect 4391 11104 4436 11132
rect 4249 11095 4307 11101
rect 4264 11064 4292 11095
rect 4430 11092 4436 11104
rect 4488 11092 4494 11144
rect 4890 11092 4896 11144
rect 4948 11132 4954 11144
rect 5258 11132 5264 11144
rect 4948 11104 5264 11132
rect 4948 11092 4954 11104
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5460 11141 5488 11172
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5444 11135 5502 11141
rect 5444 11101 5456 11135
rect 5490 11101 5502 11135
rect 5444 11095 5502 11101
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 5828 11141 5856 11308
rect 7024 11268 7052 11308
rect 7466 11296 7472 11308
rect 7524 11336 7530 11348
rect 9306 11336 9312 11348
rect 7524 11308 9312 11336
rect 7524 11296 7530 11308
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 9858 11336 9864 11348
rect 9416 11308 9864 11336
rect 7742 11268 7748 11280
rect 7024 11240 7748 11268
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 9416 11268 9444 11308
rect 9858 11296 9864 11308
rect 9916 11296 9922 11348
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 15289 11339 15347 11345
rect 15289 11336 15301 11339
rect 13964 11308 15301 11336
rect 13964 11296 13970 11308
rect 15289 11305 15301 11308
rect 15335 11336 15347 11339
rect 17586 11336 17592 11348
rect 15335 11308 17592 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 21453 11339 21511 11345
rect 21453 11305 21465 11339
rect 21499 11336 21511 11339
rect 21542 11336 21548 11348
rect 21499 11308 21548 11336
rect 21499 11305 21511 11308
rect 21453 11299 21511 11305
rect 21542 11296 21548 11308
rect 21600 11336 21606 11348
rect 21600 11308 22094 11336
rect 21600 11296 21606 11308
rect 7852 11240 9444 11268
rect 5813 11135 5871 11141
rect 5592 11104 5637 11132
rect 5592 11092 5598 11104
rect 5813 11101 5825 11135
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6914 11132 6920 11144
rect 6135 11104 6920 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7852 11141 7880 11240
rect 14918 11228 14924 11280
rect 14976 11268 14982 11280
rect 15013 11271 15071 11277
rect 15013 11268 15025 11271
rect 14976 11240 15025 11268
rect 14976 11228 14982 11240
rect 15013 11237 15025 11240
rect 15059 11237 15071 11271
rect 15013 11231 15071 11237
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 9030 11200 9036 11212
rect 8536 11172 9036 11200
rect 8536 11160 8542 11172
rect 9030 11160 9036 11172
rect 9088 11200 9094 11212
rect 9217 11203 9275 11209
rect 9217 11200 9229 11203
rect 9088 11172 9229 11200
rect 9088 11160 9094 11172
rect 9217 11169 9229 11172
rect 9263 11200 9275 11203
rect 9582 11200 9588 11212
rect 9263 11172 9588 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 9582 11160 9588 11172
rect 9640 11200 9646 11212
rect 10137 11203 10195 11209
rect 10137 11200 10149 11203
rect 9640 11172 10149 11200
rect 9640 11160 9646 11172
rect 10137 11169 10149 11172
rect 10183 11200 10195 11203
rect 10781 11203 10839 11209
rect 10781 11200 10793 11203
rect 10183 11172 10793 11200
rect 10183 11169 10195 11172
rect 10137 11163 10195 11169
rect 10781 11169 10793 11172
rect 10827 11169 10839 11203
rect 10781 11163 10839 11169
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 11330 11132 11336 11144
rect 9539 11104 11336 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 15028 11132 15056 11231
rect 15838 11228 15844 11280
rect 15896 11268 15902 11280
rect 15933 11271 15991 11277
rect 15933 11268 15945 11271
rect 15896 11240 15945 11268
rect 15896 11228 15902 11240
rect 15933 11237 15945 11240
rect 15979 11237 15991 11271
rect 15933 11231 15991 11237
rect 17126 11228 17132 11280
rect 17184 11268 17190 11280
rect 17313 11271 17371 11277
rect 17313 11268 17325 11271
rect 17184 11240 17325 11268
rect 17184 11228 17190 11240
rect 17313 11237 17325 11240
rect 17359 11268 17371 11271
rect 17402 11268 17408 11280
rect 17359 11240 17408 11268
rect 17359 11237 17371 11240
rect 17313 11231 17371 11237
rect 17402 11228 17408 11240
rect 17460 11228 17466 11280
rect 20993 11271 21051 11277
rect 20993 11268 21005 11271
rect 19306 11240 21005 11268
rect 15286 11160 15292 11212
rect 15344 11200 15350 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 15344 11172 15669 11200
rect 15344 11160 15350 11172
rect 15657 11169 15669 11172
rect 15703 11200 15715 11203
rect 15746 11200 15752 11212
rect 15703 11172 15752 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 19306 11200 19334 11240
rect 20993 11237 21005 11240
rect 21039 11268 21051 11271
rect 21174 11268 21180 11280
rect 21039 11240 21180 11268
rect 21039 11237 21051 11240
rect 20993 11231 21051 11237
rect 21174 11228 21180 11240
rect 21232 11228 21238 11280
rect 22066 11268 22094 11308
rect 22186 11268 22192 11280
rect 22066 11240 22192 11268
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 20717 11203 20775 11209
rect 20717 11200 20729 11203
rect 16776 11172 19334 11200
rect 20272 11172 20729 11200
rect 16776 11144 16804 11172
rect 15378 11132 15384 11144
rect 15028 11104 15384 11132
rect 15378 11092 15384 11104
rect 15436 11092 15442 11144
rect 15562 11132 15568 11144
rect 15523 11104 15568 11132
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 16025 11135 16083 11141
rect 16025 11101 16037 11135
rect 16071 11132 16083 11135
rect 16574 11132 16580 11144
rect 16071 11104 16580 11132
rect 16071 11101 16083 11104
rect 16025 11095 16083 11101
rect 5626 11064 5632 11076
rect 4264 11036 5632 11064
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 6178 11024 6184 11076
rect 6236 11064 6242 11076
rect 6334 11067 6392 11073
rect 6334 11064 6346 11067
rect 6236 11036 6346 11064
rect 6236 11024 6242 11036
rect 6334 11033 6346 11036
rect 6380 11033 6392 11067
rect 6334 11027 6392 11033
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 7616 11036 7696 11064
rect 7616 11024 7622 11036
rect 5905 10999 5963 11005
rect 5905 10965 5917 10999
rect 5951 10996 5963 10999
rect 6454 10996 6460 11008
rect 5951 10968 6460 10996
rect 5951 10965 5963 10968
rect 5905 10959 5963 10965
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 7668 11005 7696 11036
rect 7742 11024 7748 11076
rect 7800 11064 7806 11076
rect 10229 11067 10287 11073
rect 10229 11064 10241 11067
rect 7800 11036 10241 11064
rect 7800 11024 7806 11036
rect 10229 11033 10241 11036
rect 10275 11033 10287 11067
rect 10229 11027 10287 11033
rect 10321 11067 10379 11073
rect 10321 11033 10333 11067
rect 10367 11064 10379 11067
rect 12342 11064 12348 11076
rect 10367 11036 12348 11064
rect 10367 11033 10379 11036
rect 10321 11027 10379 11033
rect 12342 11024 12348 11036
rect 12400 11064 12406 11076
rect 16040 11064 16068 11095
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 16758 11132 16764 11144
rect 16715 11104 16764 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 16942 11132 16948 11144
rect 16903 11104 16948 11132
rect 16942 11092 16948 11104
rect 17000 11132 17006 11144
rect 17221 11135 17279 11141
rect 17221 11132 17233 11135
rect 17000 11104 17233 11132
rect 17000 11092 17006 11104
rect 17221 11101 17233 11104
rect 17267 11101 17279 11135
rect 17221 11095 17279 11101
rect 19610 11092 19616 11144
rect 19668 11132 19674 11144
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 19668 11104 19717 11132
rect 19668 11092 19674 11104
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 19886 11132 19892 11144
rect 19847 11104 19892 11132
rect 19705 11095 19763 11101
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 20272 11141 20300 11172
rect 20717 11169 20729 11172
rect 20763 11169 20775 11203
rect 23017 11203 23075 11209
rect 23017 11200 23029 11203
rect 20717 11163 20775 11169
rect 22388 11172 23029 11200
rect 20257 11135 20315 11141
rect 20257 11132 20269 11135
rect 19996 11104 20269 11132
rect 17126 11064 17132 11076
rect 12400 11036 16068 11064
rect 17087 11036 17132 11064
rect 12400 11024 12406 11036
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 7653 10999 7711 11005
rect 7653 10965 7665 10999
rect 7699 10965 7711 10999
rect 7653 10959 7711 10965
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 9401 10999 9459 11005
rect 9401 10996 9413 10999
rect 8352 10968 9413 10996
rect 8352 10956 8358 10968
rect 9401 10965 9413 10968
rect 9447 10965 9459 10999
rect 9401 10959 9459 10965
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 9861 10999 9919 11005
rect 9861 10996 9873 10999
rect 9732 10968 9873 10996
rect 9732 10956 9738 10968
rect 9861 10965 9873 10968
rect 9907 10965 9919 10999
rect 9861 10959 9919 10965
rect 10502 10956 10508 11008
rect 10560 10996 10566 11008
rect 10689 10999 10747 11005
rect 10689 10996 10701 10999
rect 10560 10968 10701 10996
rect 10560 10956 10566 10968
rect 10689 10965 10701 10968
rect 10735 10965 10747 10999
rect 10689 10959 10747 10965
rect 15194 10956 15200 11008
rect 15252 10996 15258 11008
rect 19996 10996 20024 11104
rect 20257 11101 20269 11104
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 20346 11092 20352 11144
rect 20404 11132 20410 11144
rect 20441 11135 20499 11141
rect 20441 11132 20453 11135
rect 20404 11104 20453 11132
rect 20404 11092 20410 11104
rect 20441 11101 20453 11104
rect 20487 11101 20499 11135
rect 21358 11132 21364 11144
rect 21319 11104 21364 11132
rect 20441 11095 20499 11101
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 22388 11076 22416 11172
rect 23017 11169 23029 11172
rect 23063 11200 23075 11203
rect 23290 11200 23296 11212
rect 23063 11172 23296 11200
rect 23063 11169 23075 11172
rect 23017 11163 23075 11169
rect 23290 11160 23296 11172
rect 23348 11160 23354 11212
rect 22554 11092 22560 11144
rect 22612 11132 22618 11144
rect 22833 11135 22891 11141
rect 22833 11132 22845 11135
rect 22612 11104 22845 11132
rect 22612 11092 22618 11104
rect 22833 11101 22845 11104
rect 22879 11132 22891 11135
rect 23198 11132 23204 11144
rect 22879 11104 23204 11132
rect 22879 11101 22891 11104
rect 22833 11095 22891 11101
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 20073 11067 20131 11073
rect 20073 11033 20085 11067
rect 20119 11064 20131 11067
rect 21726 11064 21732 11076
rect 20119 11036 21732 11064
rect 20119 11033 20131 11036
rect 20073 11027 20131 11033
rect 21726 11024 21732 11036
rect 21784 11024 21790 11076
rect 22281 11067 22339 11073
rect 22281 11064 22293 11067
rect 22066 11036 22293 11064
rect 20530 10996 20536 11008
rect 15252 10968 20024 10996
rect 20491 10968 20536 10996
rect 15252 10956 15258 10968
rect 20530 10956 20536 10968
rect 20588 10956 20594 11008
rect 21450 10956 21456 11008
rect 21508 10996 21514 11008
rect 21637 10999 21695 11005
rect 21637 10996 21649 10999
rect 21508 10968 21649 10996
rect 21508 10956 21514 10968
rect 21637 10965 21649 10968
rect 21683 10996 21695 10999
rect 22066 10996 22094 11036
rect 22281 11033 22293 11036
rect 22327 11064 22339 11067
rect 22370 11064 22376 11076
rect 22327 11036 22376 11064
rect 22327 11033 22339 11036
rect 22281 11027 22339 11033
rect 22370 11024 22376 11036
rect 22428 11024 22434 11076
rect 22922 11064 22928 11076
rect 22883 11036 22928 11064
rect 22922 11024 22928 11036
rect 22980 11024 22986 11076
rect 22462 10996 22468 11008
rect 21683 10968 22094 10996
rect 22423 10968 22468 10996
rect 21683 10965 21695 10968
rect 21637 10959 21695 10965
rect 22462 10956 22468 10968
rect 22520 10956 22526 11008
rect 1104 10906 26220 10928
rect 1104 10854 9322 10906
rect 9374 10854 9386 10906
rect 9438 10854 9450 10906
rect 9502 10854 9514 10906
rect 9566 10854 9578 10906
rect 9630 10854 17694 10906
rect 17746 10854 17758 10906
rect 17810 10854 17822 10906
rect 17874 10854 17886 10906
rect 17938 10854 17950 10906
rect 18002 10854 26220 10906
rect 1104 10832 26220 10854
rect 2866 10792 2872 10804
rect 2827 10764 2872 10792
rect 2866 10752 2872 10764
rect 2924 10752 2930 10804
rect 4798 10752 4804 10804
rect 4856 10752 4862 10804
rect 5534 10792 5540 10804
rect 4908 10764 5540 10792
rect 4816 10724 4844 10752
rect 4632 10696 4844 10724
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3326 10656 3332 10668
rect 3099 10628 3332 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3326 10616 3332 10628
rect 3384 10616 3390 10668
rect 4632 10665 4660 10696
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10625 4675 10659
rect 4798 10656 4804 10668
rect 4759 10628 4804 10656
rect 4617 10619 4675 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 4908 10665 4936 10764
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 5626 10752 5632 10804
rect 5684 10752 5690 10804
rect 7466 10792 7472 10804
rect 6012 10764 7472 10792
rect 5644 10724 5672 10752
rect 5000 10696 5856 10724
rect 5000 10665 5028 10696
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 2866 10548 2872 10600
rect 2924 10588 2930 10600
rect 3237 10591 3295 10597
rect 3237 10588 3249 10591
rect 2924 10560 3249 10588
rect 2924 10548 2930 10560
rect 3237 10557 3249 10560
rect 3283 10588 3295 10591
rect 3786 10588 3792 10600
rect 3283 10560 3792 10588
rect 3283 10557 3295 10560
rect 3237 10551 3295 10557
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 5184 10588 5212 10619
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 5828 10665 5856 10696
rect 6012 10665 6040 10764
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7742 10792 7748 10804
rect 7703 10764 7748 10792
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 9309 10795 9367 10801
rect 9309 10761 9321 10795
rect 9355 10792 9367 10795
rect 9766 10792 9772 10804
rect 9355 10764 9772 10792
rect 9355 10761 9367 10764
rect 9309 10755 9367 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 12253 10795 12311 10801
rect 12253 10792 12265 10795
rect 9916 10764 12265 10792
rect 9916 10752 9922 10764
rect 12253 10761 12265 10764
rect 12299 10792 12311 10795
rect 12345 10795 12403 10801
rect 12345 10792 12357 10795
rect 12299 10764 12357 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12345 10761 12357 10764
rect 12391 10761 12403 10795
rect 12345 10755 12403 10761
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 14090 10792 14096 10804
rect 13863 10764 14096 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 17034 10752 17040 10804
rect 17092 10792 17098 10804
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 17092 10764 17141 10792
rect 17092 10752 17098 10764
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 19337 10795 19395 10801
rect 19337 10761 19349 10795
rect 19383 10792 19395 10795
rect 19886 10792 19892 10804
rect 19383 10764 19892 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 19886 10752 19892 10764
rect 19944 10752 19950 10804
rect 20530 10792 20536 10804
rect 20491 10764 20536 10792
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 21174 10752 21180 10804
rect 21232 10792 21238 10804
rect 21637 10795 21695 10801
rect 21637 10792 21649 10795
rect 21232 10764 21649 10792
rect 21232 10752 21238 10764
rect 21637 10761 21649 10764
rect 21683 10761 21695 10795
rect 22186 10792 22192 10804
rect 22147 10764 22192 10792
rect 21637 10755 21695 10761
rect 22186 10752 22192 10764
rect 22244 10792 22250 10804
rect 22554 10792 22560 10804
rect 22244 10764 22560 10792
rect 22244 10752 22250 10764
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 23014 10752 23020 10804
rect 23072 10752 23078 10804
rect 6178 10724 6184 10736
rect 6139 10696 6184 10724
rect 6178 10684 6184 10696
rect 6236 10684 6242 10736
rect 6914 10724 6920 10736
rect 6380 10696 6920 10724
rect 6380 10665 6408 10696
rect 6914 10684 6920 10696
rect 6972 10724 6978 10736
rect 13078 10724 13084 10736
rect 6972 10696 7972 10724
rect 6972 10684 6978 10696
rect 7944 10668 7972 10696
rect 9508 10696 13084 10724
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 5316 10628 5457 10656
rect 5316 10616 5322 10628
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 5593 10659 5651 10665
rect 5593 10625 5605 10659
rect 5639 10656 5651 10659
rect 5813 10659 5871 10665
rect 5639 10625 5672 10656
rect 5593 10619 5672 10625
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6365 10659 6423 10665
rect 6365 10625 6377 10659
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 5184 10560 5580 10588
rect 5552 10532 5580 10560
rect 5534 10480 5540 10532
rect 5592 10480 5598 10532
rect 5644 10520 5672 10619
rect 6454 10616 6460 10668
rect 6512 10656 6518 10668
rect 6621 10659 6679 10665
rect 6621 10656 6633 10659
rect 6512 10628 6633 10656
rect 6512 10616 6518 10628
rect 6621 10625 6633 10628
rect 6667 10625 6679 10659
rect 7926 10656 7932 10668
rect 7887 10628 7932 10656
rect 6621 10619 6679 10625
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8018 10616 8024 10668
rect 8076 10656 8082 10668
rect 8185 10659 8243 10665
rect 8185 10656 8197 10659
rect 8076 10628 8197 10656
rect 8076 10616 8082 10628
rect 8185 10625 8197 10628
rect 8231 10625 8243 10659
rect 8185 10619 8243 10625
rect 8754 10616 8760 10668
rect 8812 10656 8818 10668
rect 9508 10665 9536 10696
rect 9493 10659 9551 10665
rect 9493 10656 9505 10659
rect 8812 10628 9505 10656
rect 8812 10616 8818 10628
rect 9493 10625 9505 10628
rect 9539 10625 9551 10659
rect 9674 10656 9680 10668
rect 9635 10628 9680 10656
rect 9493 10619 9551 10625
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 10226 10656 10232 10668
rect 10091 10628 10232 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 10226 10616 10232 10628
rect 10284 10616 10290 10668
rect 10336 10665 10364 10696
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 16390 10684 16396 10736
rect 16448 10724 16454 10736
rect 16448 10696 17540 10724
rect 16448 10684 16454 10696
rect 10321 10659 10379 10665
rect 10321 10625 10333 10659
rect 10367 10625 10379 10659
rect 10502 10656 10508 10668
rect 10463 10628 10508 10656
rect 10321 10619 10379 10625
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10656 10655 10659
rect 10873 10659 10931 10665
rect 10643 10628 10823 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 5718 10548 5724 10600
rect 5776 10588 5782 10600
rect 5776 10560 5821 10588
rect 5776 10548 5782 10560
rect 9398 10548 9404 10600
rect 9456 10588 9462 10600
rect 9769 10591 9827 10597
rect 9769 10588 9781 10591
rect 9456 10560 9781 10588
rect 9456 10548 9462 10560
rect 9769 10557 9781 10560
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 5994 10520 6000 10532
rect 5644 10492 6000 10520
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 9784 10520 9812 10551
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10689 10591 10747 10597
rect 10689 10588 10701 10591
rect 9916 10560 10701 10588
rect 9916 10548 9922 10560
rect 10689 10557 10701 10560
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 10795 10520 10823 10628
rect 10873 10625 10885 10659
rect 10919 10656 10931 10659
rect 11606 10656 11612 10668
rect 10919 10628 11612 10656
rect 10919 10625 10931 10628
rect 10873 10619 10931 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 11882 10616 11888 10668
rect 11940 10656 11946 10668
rect 12710 10665 12716 10668
rect 12069 10659 12127 10665
rect 12069 10656 12081 10659
rect 11940 10628 12081 10656
rect 11940 10616 11946 10628
rect 12069 10625 12081 10628
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 12704 10619 12716 10665
rect 12768 10656 12774 10668
rect 12768 10628 12804 10656
rect 12710 10616 12716 10619
rect 12768 10616 12774 10628
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 15289 10659 15347 10665
rect 15289 10656 15301 10659
rect 15252 10628 15301 10656
rect 15252 10616 15258 10628
rect 15289 10625 15301 10628
rect 15335 10625 15347 10659
rect 15562 10656 15568 10668
rect 15523 10628 15568 10656
rect 15289 10619 15347 10625
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 16485 10659 16543 10665
rect 16485 10656 16497 10659
rect 15979 10628 16497 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 16485 10625 16497 10628
rect 16531 10656 16543 10659
rect 16574 10656 16580 10668
rect 16531 10628 16580 10656
rect 16531 10625 16543 10628
rect 16485 10619 16543 10625
rect 16574 10616 16580 10628
rect 16632 10616 16638 10668
rect 17034 10656 17040 10668
rect 16995 10628 17040 10656
rect 17034 10616 17040 10628
rect 17092 10616 17098 10668
rect 17512 10665 17540 10696
rect 17586 10684 17592 10736
rect 17644 10724 17650 10736
rect 22646 10724 22652 10736
rect 17644 10696 22652 10724
rect 17644 10684 17650 10696
rect 22646 10684 22652 10696
rect 22704 10684 22710 10736
rect 23032 10724 23060 10752
rect 23032 10696 23612 10724
rect 17497 10659 17555 10665
rect 17497 10625 17509 10659
rect 17543 10625 17555 10659
rect 17678 10656 17684 10668
rect 17639 10628 17684 10656
rect 17497 10619 17555 10625
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 17221 10591 17279 10597
rect 17221 10588 17233 10591
rect 12492 10560 12537 10588
rect 16316 10560 17233 10588
rect 12492 10548 12498 10560
rect 15470 10520 15476 10532
rect 9784 10492 10823 10520
rect 15028 10492 15476 10520
rect 5261 10455 5319 10461
rect 5261 10421 5273 10455
rect 5307 10452 5319 10455
rect 6086 10452 6092 10464
rect 5307 10424 6092 10452
rect 5307 10421 5319 10424
rect 5261 10415 5319 10421
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 10134 10452 10140 10464
rect 10095 10424 10140 10452
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 10962 10452 10968 10464
rect 10923 10424 10968 10452
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 12345 10455 12403 10461
rect 12345 10421 12357 10455
rect 12391 10452 12403 10455
rect 15028 10452 15056 10492
rect 15470 10480 15476 10492
rect 15528 10480 15534 10532
rect 15565 10523 15623 10529
rect 15565 10489 15577 10523
rect 15611 10520 15623 10523
rect 15654 10520 15660 10532
rect 15611 10492 15660 10520
rect 15611 10489 15623 10492
rect 15565 10483 15623 10489
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 16316 10464 16344 10560
rect 17221 10557 17233 10560
rect 17267 10557 17279 10591
rect 17512 10588 17540 10619
rect 17678 10616 17684 10628
rect 17736 10616 17742 10668
rect 17770 10616 17776 10668
rect 17828 10656 17834 10668
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 17828 10628 18061 10656
rect 17828 10616 17834 10628
rect 18049 10625 18061 10628
rect 18095 10625 18107 10659
rect 18782 10656 18788 10668
rect 18743 10628 18788 10656
rect 18049 10619 18107 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 19426 10656 19432 10668
rect 19076 10628 19288 10656
rect 19387 10628 19432 10656
rect 19076 10588 19104 10628
rect 17512 10560 19104 10588
rect 19153 10591 19211 10597
rect 17221 10551 17279 10557
rect 19153 10557 19165 10591
rect 19199 10557 19211 10591
rect 19260 10588 19288 10628
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 20622 10656 20628 10668
rect 20583 10628 20628 10656
rect 20622 10616 20628 10628
rect 20680 10616 20686 10668
rect 21174 10656 21180 10668
rect 21135 10628 21180 10656
rect 21174 10616 21180 10628
rect 21232 10616 21238 10668
rect 21358 10656 21364 10668
rect 21319 10628 21364 10656
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 21637 10659 21695 10665
rect 21637 10625 21649 10659
rect 21683 10656 21695 10659
rect 23014 10656 23020 10668
rect 21683 10628 22885 10656
rect 22975 10628 23020 10656
rect 21683 10625 21695 10628
rect 21637 10619 21695 10625
rect 19610 10588 19616 10600
rect 19260 10560 19616 10588
rect 19153 10551 19211 10557
rect 17236 10520 17264 10551
rect 18601 10523 18659 10529
rect 18601 10520 18613 10523
rect 17236 10492 18613 10520
rect 18601 10489 18613 10492
rect 18647 10520 18659 10523
rect 19168 10520 19196 10551
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 20349 10591 20407 10597
rect 20349 10557 20361 10591
rect 20395 10588 20407 10591
rect 21450 10588 21456 10600
rect 20395 10560 21456 10588
rect 20395 10557 20407 10560
rect 20349 10551 20407 10557
rect 18647 10492 19196 10520
rect 18647 10489 18659 10492
rect 18601 10483 18659 10489
rect 15194 10452 15200 10464
rect 12391 10424 15056 10452
rect 15155 10424 15200 10452
rect 12391 10421 12403 10424
rect 12345 10415 12403 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 15749 10455 15807 10461
rect 15749 10452 15761 10455
rect 15344 10424 15761 10452
rect 15344 10412 15350 10424
rect 15749 10421 15761 10424
rect 15795 10452 15807 10455
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 15795 10424 15945 10452
rect 15795 10421 15807 10424
rect 15749 10415 15807 10421
rect 15933 10421 15945 10424
rect 15979 10421 15991 10455
rect 15933 10415 15991 10421
rect 16117 10455 16175 10461
rect 16117 10421 16129 10455
rect 16163 10452 16175 10455
rect 16298 10452 16304 10464
rect 16163 10424 16304 10452
rect 16163 10421 16175 10424
rect 16117 10415 16175 10421
rect 16298 10412 16304 10424
rect 16356 10412 16362 10464
rect 16482 10412 16488 10464
rect 16540 10452 16546 10464
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 16540 10424 16681 10452
rect 16540 10412 16546 10424
rect 16669 10421 16681 10424
rect 16715 10421 16727 10455
rect 17862 10452 17868 10464
rect 17823 10424 17868 10452
rect 16669 10415 16727 10421
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 18966 10452 18972 10464
rect 18927 10424 18972 10452
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 19794 10452 19800 10464
rect 19755 10424 19800 10452
rect 19794 10412 19800 10424
rect 19852 10412 19858 10464
rect 19978 10452 19984 10464
rect 19939 10424 19984 10452
rect 19978 10412 19984 10424
rect 20036 10452 20042 10464
rect 20073 10455 20131 10461
rect 20073 10452 20085 10455
rect 20036 10424 20085 10452
rect 20036 10412 20042 10424
rect 20073 10421 20085 10424
rect 20119 10452 20131 10455
rect 20364 10452 20392 10551
rect 21450 10548 21456 10560
rect 21508 10548 21514 10600
rect 21545 10591 21603 10597
rect 21545 10557 21557 10591
rect 21591 10588 21603 10591
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 21591 10560 22293 10588
rect 21591 10557 21603 10560
rect 21545 10551 21603 10557
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 22370 10548 22376 10600
rect 22428 10588 22434 10600
rect 22428 10560 22473 10588
rect 22428 10548 22434 10560
rect 20993 10523 21051 10529
rect 20993 10489 21005 10523
rect 21039 10520 21051 10523
rect 22857 10520 22885 10628
rect 23014 10616 23020 10628
rect 23072 10616 23078 10668
rect 23584 10665 23612 10696
rect 23109 10659 23167 10665
rect 23109 10625 23121 10659
rect 23155 10656 23167 10659
rect 23477 10659 23535 10665
rect 23477 10656 23489 10659
rect 23155 10628 23489 10656
rect 23155 10625 23167 10628
rect 23109 10619 23167 10625
rect 23477 10625 23489 10628
rect 23523 10625 23535 10659
rect 23477 10619 23535 10625
rect 23569 10659 23627 10665
rect 23569 10625 23581 10659
rect 23615 10625 23627 10659
rect 23569 10619 23627 10625
rect 23753 10659 23811 10665
rect 23753 10625 23765 10659
rect 23799 10625 23811 10659
rect 23753 10619 23811 10625
rect 23290 10588 23296 10600
rect 23251 10560 23296 10588
rect 23290 10548 23296 10560
rect 23348 10548 23354 10600
rect 23768 10520 23796 10619
rect 23937 10523 23995 10529
rect 23937 10520 23949 10523
rect 21039 10492 22324 10520
rect 22857 10492 23949 10520
rect 21039 10489 21051 10492
rect 20993 10483 21051 10489
rect 22296 10464 22324 10492
rect 23937 10489 23949 10492
rect 23983 10489 23995 10523
rect 23937 10483 23995 10489
rect 20119 10424 20392 10452
rect 20119 10421 20131 10424
rect 20073 10415 20131 10421
rect 20806 10412 20812 10464
rect 20864 10452 20870 10464
rect 21821 10455 21879 10461
rect 21821 10452 21833 10455
rect 20864 10424 21833 10452
rect 20864 10412 20870 10424
rect 21821 10421 21833 10424
rect 21867 10421 21879 10455
rect 21821 10415 21879 10421
rect 22278 10412 22284 10464
rect 22336 10412 22342 10464
rect 22649 10455 22707 10461
rect 22649 10421 22661 10455
rect 22695 10452 22707 10455
rect 22830 10452 22836 10464
rect 22695 10424 22836 10452
rect 22695 10421 22707 10424
rect 22649 10415 22707 10421
rect 22830 10412 22836 10424
rect 22888 10412 22894 10464
rect 1104 10362 26220 10384
rect 1104 10310 5136 10362
rect 5188 10310 5200 10362
rect 5252 10310 5264 10362
rect 5316 10310 5328 10362
rect 5380 10310 5392 10362
rect 5444 10310 13508 10362
rect 13560 10310 13572 10362
rect 13624 10310 13636 10362
rect 13688 10310 13700 10362
rect 13752 10310 13764 10362
rect 13816 10310 21880 10362
rect 21932 10310 21944 10362
rect 21996 10310 22008 10362
rect 22060 10310 22072 10362
rect 22124 10310 22136 10362
rect 22188 10310 26220 10362
rect 1104 10288 26220 10310
rect 2866 10248 2872 10260
rect 2827 10220 2872 10248
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 5592 10220 7205 10248
rect 5592 10208 5598 10220
rect 7193 10217 7205 10220
rect 7239 10248 7251 10251
rect 8294 10248 8300 10260
rect 7239 10220 8300 10248
rect 7239 10217 7251 10220
rect 7193 10211 7251 10217
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 10226 10248 10232 10260
rect 9048 10220 10232 10248
rect 3326 10140 3332 10192
rect 3384 10180 3390 10192
rect 3602 10180 3608 10192
rect 3384 10152 3608 10180
rect 3384 10140 3390 10152
rect 3602 10140 3608 10152
rect 3660 10180 3666 10192
rect 3973 10183 4031 10189
rect 3973 10180 3985 10183
rect 3660 10152 3985 10180
rect 3660 10140 3666 10152
rect 3973 10149 3985 10152
rect 4019 10149 4031 10183
rect 3973 10143 4031 10149
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 9048 10189 9076 10220
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 11606 10208 11612 10260
rect 11664 10248 11670 10260
rect 12253 10251 12311 10257
rect 12253 10248 12265 10251
rect 11664 10220 12265 10248
rect 11664 10208 11670 10220
rect 12253 10217 12265 10220
rect 12299 10248 12311 10251
rect 12621 10251 12679 10257
rect 12299 10220 12434 10248
rect 12299 10217 12311 10220
rect 12253 10211 12311 10217
rect 9033 10183 9091 10189
rect 9033 10180 9045 10183
rect 8444 10152 9045 10180
rect 8444 10140 8450 10152
rect 9033 10149 9045 10152
rect 9079 10149 9091 10183
rect 12406 10180 12434 10220
rect 12621 10217 12633 10251
rect 12667 10248 12679 10251
rect 12710 10248 12716 10260
rect 12667 10220 12716 10248
rect 12667 10217 12679 10220
rect 12621 10211 12679 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 17034 10248 17040 10260
rect 16995 10220 17040 10248
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 18782 10208 18788 10260
rect 18840 10248 18846 10260
rect 19337 10251 19395 10257
rect 19337 10248 19349 10251
rect 18840 10220 19349 10248
rect 18840 10208 18846 10220
rect 19337 10217 19349 10220
rect 19383 10217 19395 10251
rect 19337 10211 19395 10217
rect 19610 10208 19616 10260
rect 19668 10248 19674 10260
rect 19668 10220 23612 10248
rect 19668 10208 19674 10220
rect 17586 10180 17592 10192
rect 12406 10152 17592 10180
rect 9033 10143 9091 10149
rect 17586 10140 17592 10152
rect 17644 10140 17650 10192
rect 21545 10183 21603 10189
rect 21545 10180 21557 10183
rect 20180 10152 21557 10180
rect 1486 10112 1492 10124
rect 1447 10084 1492 10112
rect 1486 10072 1492 10084
rect 1544 10072 1550 10124
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 3513 10115 3571 10121
rect 3513 10112 3525 10115
rect 3200 10084 3525 10112
rect 3200 10072 3206 10084
rect 3513 10081 3525 10084
rect 3559 10112 3571 10115
rect 4062 10112 4068 10124
rect 3559 10084 4068 10112
rect 3559 10081 3571 10084
rect 3513 10075 3571 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 9398 10112 9404 10124
rect 8527 10084 9404 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 14090 10072 14096 10124
rect 14148 10112 14154 10124
rect 14645 10115 14703 10121
rect 14645 10112 14657 10115
rect 14148 10084 14657 10112
rect 14148 10072 14154 10084
rect 14645 10081 14657 10084
rect 14691 10112 14703 10115
rect 15286 10112 15292 10124
rect 14691 10084 15292 10112
rect 14691 10081 14703 10084
rect 14645 10075 14703 10081
rect 15286 10072 15292 10084
rect 15344 10112 15350 10124
rect 15473 10115 15531 10121
rect 15473 10112 15485 10115
rect 15344 10084 15485 10112
rect 15344 10072 15350 10084
rect 15473 10081 15485 10084
rect 15519 10081 15531 10115
rect 15654 10112 15660 10124
rect 15615 10084 15660 10112
rect 15473 10075 15531 10081
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 16298 10112 16304 10124
rect 16259 10084 16304 10112
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 17126 10072 17132 10124
rect 17184 10112 17190 10124
rect 17497 10115 17555 10121
rect 17497 10112 17509 10115
rect 17184 10084 17509 10112
rect 17184 10072 17190 10084
rect 17497 10081 17509 10084
rect 17543 10081 17555 10115
rect 17681 10115 17739 10121
rect 17681 10112 17693 10115
rect 17497 10075 17555 10081
rect 17604 10084 17693 10112
rect 17604 10056 17632 10084
rect 17681 10081 17693 10084
rect 17727 10112 17739 10115
rect 17770 10112 17776 10124
rect 17727 10084 17776 10112
rect 17727 10081 17739 10084
rect 17681 10075 17739 10081
rect 17770 10072 17776 10084
rect 17828 10112 17834 10124
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 17828 10084 18429 10112
rect 17828 10072 17834 10084
rect 18417 10081 18429 10084
rect 18463 10112 18475 10115
rect 18969 10115 19027 10121
rect 18969 10112 18981 10115
rect 18463 10084 18981 10112
rect 18463 10081 18475 10084
rect 18417 10075 18475 10081
rect 18969 10081 18981 10084
rect 19015 10112 19027 10115
rect 19978 10112 19984 10124
rect 19015 10084 19984 10112
rect 19015 10081 19027 10084
rect 18969 10075 19027 10081
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 20180 10121 20208 10152
rect 21545 10149 21557 10152
rect 21591 10149 21603 10183
rect 21545 10143 21603 10149
rect 20165 10115 20223 10121
rect 20165 10081 20177 10115
rect 20211 10081 20223 10115
rect 20165 10075 20223 10081
rect 20622 10072 20628 10124
rect 20680 10112 20686 10124
rect 21177 10115 21235 10121
rect 21177 10112 21189 10115
rect 20680 10084 21189 10112
rect 20680 10072 20686 10084
rect 21177 10081 21189 10084
rect 21223 10081 21235 10115
rect 21177 10075 21235 10081
rect 21269 10115 21327 10121
rect 21269 10081 21281 10115
rect 21315 10112 21327 10115
rect 22005 10115 22063 10121
rect 22005 10112 22017 10115
rect 21315 10084 22017 10112
rect 21315 10081 21327 10084
rect 21269 10075 21327 10081
rect 22005 10081 22017 10084
rect 22051 10081 22063 10115
rect 22005 10075 22063 10081
rect 22189 10115 22247 10121
rect 22189 10081 22201 10115
rect 22235 10112 22247 10115
rect 22738 10112 22744 10124
rect 22235 10084 22744 10112
rect 22235 10081 22247 10084
rect 22189 10075 22247 10081
rect 3326 10044 3332 10056
rect 3287 10016 3332 10044
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 3418 10004 3424 10056
rect 3476 10044 3482 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3476 10016 3801 10044
rect 3476 10004 3482 10016
rect 3789 10013 3801 10016
rect 3835 10044 3847 10047
rect 4982 10044 4988 10056
rect 3835 10016 4988 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 5718 10044 5724 10056
rect 5679 10016 5724 10044
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 6914 10044 6920 10056
rect 5859 10016 6920 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10044 8263 10047
rect 8294 10044 8300 10056
rect 8251 10016 8300 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8574 10047 8632 10053
rect 8574 10013 8586 10047
rect 8620 10044 8632 10047
rect 8662 10044 8668 10056
rect 8620 10016 8668 10044
rect 8620 10013 8632 10016
rect 8574 10007 8632 10013
rect 1756 9979 1814 9985
rect 1756 9945 1768 9979
rect 1802 9976 1814 9979
rect 2498 9976 2504 9988
rect 1802 9948 2504 9976
rect 1802 9945 1814 9948
rect 1756 9939 1814 9945
rect 2498 9936 2504 9948
rect 2556 9936 2562 9988
rect 6086 9985 6092 9988
rect 6080 9976 6092 9985
rect 6047 9948 6092 9976
rect 6080 9939 6092 9948
rect 6086 9936 6092 9939
rect 6144 9936 6150 9988
rect 8404 9976 8432 10007
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 8754 10004 8760 10056
rect 8812 10044 8818 10056
rect 8812 10016 8857 10044
rect 8812 10004 8818 10016
rect 10134 10004 10140 10056
rect 10192 10053 10198 10056
rect 10192 10044 10204 10053
rect 10410 10044 10416 10056
rect 10192 10016 10237 10044
rect 10323 10016 10416 10044
rect 10192 10007 10204 10016
rect 10192 10004 10198 10007
rect 10410 10004 10416 10016
rect 10468 10044 10474 10056
rect 10873 10047 10931 10053
rect 10873 10044 10885 10047
rect 10468 10016 10885 10044
rect 10468 10004 10474 10016
rect 10873 10013 10885 10016
rect 10919 10013 10931 10047
rect 10873 10007 10931 10013
rect 10962 10004 10968 10056
rect 11020 10044 11026 10056
rect 11129 10047 11187 10053
rect 11129 10044 11141 10047
rect 11020 10016 11141 10044
rect 11020 10004 11026 10016
rect 11129 10013 11141 10016
rect 11175 10013 11187 10047
rect 11129 10007 11187 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 12526 10044 12532 10056
rect 12483 10016 12532 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 13538 10044 13544 10056
rect 13499 10016 13544 10044
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10044 13691 10047
rect 14182 10044 14188 10056
rect 13679 10016 14188 10044
rect 13679 10013 13691 10016
rect 13633 10007 13691 10013
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10044 14335 10047
rect 16022 10044 16028 10056
rect 14323 10016 16028 10044
rect 14323 10013 14335 10016
rect 14277 10007 14335 10013
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 16485 10047 16543 10053
rect 16485 10013 16497 10047
rect 16531 10044 16543 10047
rect 16666 10044 16672 10056
rect 16531 10016 16672 10044
rect 16531 10013 16543 10016
rect 16485 10007 16543 10013
rect 16666 10004 16672 10016
rect 16724 10044 16730 10056
rect 17402 10044 17408 10056
rect 16724 10016 16988 10044
rect 17363 10016 17408 10044
rect 16724 10004 16730 10016
rect 9122 9976 9128 9988
rect 8404 9948 9128 9976
rect 9122 9936 9128 9948
rect 9180 9976 9186 9988
rect 9582 9976 9588 9988
rect 9180 9948 9588 9976
rect 9180 9936 9186 9948
rect 9582 9936 9588 9948
rect 9640 9936 9646 9988
rect 14090 9976 14096 9988
rect 13280 9948 14096 9976
rect 13280 9920 13308 9948
rect 14090 9936 14096 9948
rect 14148 9936 14154 9988
rect 14366 9936 14372 9988
rect 14424 9976 14430 9988
rect 14734 9976 14740 9988
rect 14424 9948 14740 9976
rect 14424 9936 14430 9948
rect 14734 9936 14740 9948
rect 14792 9976 14798 9988
rect 14921 9979 14979 9985
rect 14921 9976 14933 9979
rect 14792 9948 14933 9976
rect 14792 9936 14798 9948
rect 14921 9945 14933 9948
rect 14967 9945 14979 9979
rect 15746 9976 15752 9988
rect 15707 9948 15752 9976
rect 14921 9939 14979 9945
rect 15746 9936 15752 9948
rect 15804 9936 15810 9988
rect 16577 9979 16635 9985
rect 16577 9976 16589 9979
rect 16132 9948 16589 9976
rect 2958 9868 2964 9920
rect 3016 9908 3022 9920
rect 3145 9911 3203 9917
rect 3145 9908 3157 9911
rect 3016 9880 3157 9908
rect 3016 9868 3022 9880
rect 3145 9877 3157 9880
rect 3191 9877 3203 9911
rect 3145 9871 3203 9877
rect 5537 9911 5595 9917
rect 5537 9877 5549 9911
rect 5583 9908 5595 9911
rect 5626 9908 5632 9920
rect 5583 9880 5632 9908
rect 5583 9877 5595 9880
rect 5537 9871 5595 9877
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 8113 9911 8171 9917
rect 8113 9877 8125 9911
rect 8159 9908 8171 9911
rect 8938 9908 8944 9920
rect 8159 9880 8944 9908
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 13262 9908 13268 9920
rect 13223 9880 13268 9908
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 13814 9908 13820 9920
rect 13775 9880 13820 9908
rect 13814 9868 13820 9880
rect 13872 9868 13878 9920
rect 14461 9911 14519 9917
rect 14461 9877 14473 9911
rect 14507 9908 14519 9911
rect 14829 9911 14887 9917
rect 14829 9908 14841 9911
rect 14507 9880 14841 9908
rect 14507 9877 14519 9880
rect 14461 9871 14519 9877
rect 14829 9877 14841 9880
rect 14875 9877 14887 9911
rect 15286 9908 15292 9920
rect 15247 9880 15292 9908
rect 14829 9871 14887 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 16132 9917 16160 9948
rect 16577 9945 16589 9948
rect 16623 9945 16635 9979
rect 16960 9976 16988 10016
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 17586 10004 17592 10056
rect 17644 10004 17650 10056
rect 17862 10004 17868 10056
rect 17920 10044 17926 10056
rect 18877 10047 18935 10053
rect 18877 10044 18889 10047
rect 17920 10016 18889 10044
rect 17920 10004 17926 10016
rect 18877 10013 18889 10016
rect 18923 10013 18935 10047
rect 18877 10007 18935 10013
rect 19058 10004 19064 10056
rect 19116 10044 19122 10056
rect 19521 10047 19579 10053
rect 19521 10044 19533 10047
rect 19116 10016 19533 10044
rect 19116 10004 19122 10016
rect 19521 10013 19533 10016
rect 19567 10013 19579 10047
rect 19521 10007 19579 10013
rect 19610 10004 19616 10056
rect 19668 10044 19674 10056
rect 19668 10016 19713 10044
rect 19668 10004 19674 10016
rect 19886 10004 19892 10056
rect 19944 10044 19950 10056
rect 20257 10047 20315 10053
rect 20257 10044 20269 10047
rect 19944 10016 20269 10044
rect 19944 10004 19950 10016
rect 20257 10013 20269 10016
rect 20303 10013 20315 10047
rect 20257 10007 20315 10013
rect 20990 10004 20996 10056
rect 21048 10044 21054 10056
rect 21284 10044 21312 10075
rect 22738 10072 22744 10084
rect 22796 10072 22802 10124
rect 23290 10112 23296 10124
rect 23251 10084 23296 10112
rect 23290 10072 23296 10084
rect 23348 10072 23354 10124
rect 23584 10121 23612 10220
rect 23569 10115 23627 10121
rect 23569 10081 23581 10115
rect 23615 10081 23627 10115
rect 23569 10075 23627 10081
rect 21726 10044 21732 10056
rect 21048 10016 21312 10044
rect 21687 10016 21732 10044
rect 21048 10004 21054 10016
rect 21726 10004 21732 10016
rect 21784 10004 21790 10056
rect 22278 10044 22284 10056
rect 22239 10016 22284 10044
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 22756 10044 22784 10072
rect 23109 10047 23167 10053
rect 23109 10044 23121 10047
rect 22756 10016 23121 10044
rect 23109 10013 23121 10016
rect 23155 10044 23167 10047
rect 23753 10047 23811 10053
rect 23753 10044 23765 10047
rect 23155 10016 23765 10044
rect 23155 10013 23167 10016
rect 23109 10007 23167 10013
rect 23753 10013 23765 10016
rect 23799 10013 23811 10047
rect 23753 10007 23811 10013
rect 23937 10047 23995 10053
rect 23937 10013 23949 10047
rect 23983 10044 23995 10047
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 23983 10016 24593 10044
rect 23983 10013 23995 10016
rect 23937 10007 23995 10013
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 17678 9976 17684 9988
rect 16960 9948 17684 9976
rect 16577 9939 16635 9945
rect 17678 9936 17684 9948
rect 17736 9976 17742 9988
rect 18233 9979 18291 9985
rect 18233 9976 18245 9979
rect 17736 9948 18245 9976
rect 17736 9936 17742 9948
rect 18233 9945 18245 9948
rect 18279 9945 18291 9979
rect 21085 9979 21143 9985
rect 21085 9976 21097 9979
rect 18233 9939 18291 9945
rect 20640 9948 21097 9976
rect 16117 9911 16175 9917
rect 16117 9877 16129 9911
rect 16163 9877 16175 9911
rect 16942 9908 16948 9920
rect 16903 9880 16948 9908
rect 16117 9871 16175 9877
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 17586 9868 17592 9920
rect 17644 9908 17650 9920
rect 20640 9917 20668 9948
rect 21085 9945 21097 9948
rect 21131 9945 21143 9979
rect 21085 9939 21143 9945
rect 23201 9979 23259 9985
rect 23201 9945 23213 9979
rect 23247 9976 23259 9979
rect 23247 9948 24440 9976
rect 23247 9945 23259 9948
rect 23201 9939 23259 9945
rect 17865 9911 17923 9917
rect 17865 9908 17877 9911
rect 17644 9880 17877 9908
rect 17644 9868 17650 9880
rect 17865 9877 17877 9880
rect 17911 9877 17923 9911
rect 17865 9871 17923 9877
rect 18325 9911 18383 9917
rect 18325 9877 18337 9911
rect 18371 9908 18383 9911
rect 18693 9911 18751 9917
rect 18693 9908 18705 9911
rect 18371 9880 18705 9908
rect 18371 9877 18383 9880
rect 18325 9871 18383 9877
rect 18693 9877 18705 9880
rect 18739 9877 18751 9911
rect 18693 9871 18751 9877
rect 20625 9911 20683 9917
rect 20625 9877 20637 9911
rect 20671 9877 20683 9911
rect 20625 9871 20683 9877
rect 20714 9868 20720 9920
rect 20772 9908 20778 9920
rect 20772 9880 20817 9908
rect 20772 9868 20778 9880
rect 22370 9868 22376 9920
rect 22428 9908 22434 9920
rect 22649 9911 22707 9917
rect 22649 9908 22661 9911
rect 22428 9880 22661 9908
rect 22428 9868 22434 9880
rect 22649 9877 22661 9880
rect 22695 9877 22707 9911
rect 22649 9871 22707 9877
rect 22738 9868 22744 9920
rect 22796 9908 22802 9920
rect 22796 9880 22841 9908
rect 22796 9868 22802 9880
rect 23290 9868 23296 9920
rect 23348 9908 23354 9920
rect 24412 9917 24440 9948
rect 24121 9911 24179 9917
rect 24121 9908 24133 9911
rect 23348 9880 24133 9908
rect 23348 9868 23354 9880
rect 24121 9877 24133 9880
rect 24167 9877 24179 9911
rect 24121 9871 24179 9877
rect 24397 9911 24455 9917
rect 24397 9877 24409 9911
rect 24443 9877 24455 9911
rect 24397 9871 24455 9877
rect 1104 9818 26220 9840
rect 1104 9766 9322 9818
rect 9374 9766 9386 9818
rect 9438 9766 9450 9818
rect 9502 9766 9514 9818
rect 9566 9766 9578 9818
rect 9630 9766 17694 9818
rect 17746 9766 17758 9818
rect 17810 9766 17822 9818
rect 17874 9766 17886 9818
rect 17938 9766 17950 9818
rect 18002 9766 26220 9818
rect 1104 9744 26220 9766
rect 2498 9704 2504 9716
rect 2459 9676 2504 9704
rect 2498 9664 2504 9676
rect 2556 9664 2562 9716
rect 11333 9707 11391 9713
rect 11333 9673 11345 9707
rect 11379 9704 11391 9707
rect 15197 9707 15255 9713
rect 11379 9676 12572 9704
rect 11379 9673 11391 9676
rect 11333 9667 11391 9673
rect 2866 9636 2872 9648
rect 2700 9608 2872 9636
rect 2700 9577 2728 9608
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 3418 9596 3424 9648
rect 3476 9636 3482 9648
rect 7374 9636 7380 9648
rect 3476 9608 7380 9636
rect 3476 9596 3482 9608
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 12434 9636 12440 9648
rect 8536 9608 10180 9636
rect 8536 9596 8542 9608
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 3050 9568 3056 9580
rect 2832 9540 2877 9568
rect 3011 9540 3056 9568
rect 2832 9528 2838 9540
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 3326 9568 3332 9580
rect 3287 9540 3332 9568
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3602 9568 3608 9580
rect 3563 9540 3608 9568
rect 3602 9528 3608 9540
rect 3660 9568 3666 9580
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 3660 9540 4261 9568
rect 3660 9528 3666 9540
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9568 4491 9571
rect 4614 9568 4620 9580
rect 4479 9540 4620 9568
rect 4479 9537 4491 9540
rect 4433 9531 4491 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 8938 9528 8944 9580
rect 8996 9568 9002 9580
rect 10152 9577 10180 9608
rect 11532 9608 12440 9636
rect 9870 9571 9928 9577
rect 9870 9568 9882 9571
rect 8996 9540 9882 9568
rect 8996 9528 9002 9540
rect 9870 9537 9882 9540
rect 9916 9537 9928 9571
rect 9870 9531 9928 9537
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9568 10195 9571
rect 10410 9568 10416 9580
rect 10183 9540 10416 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10594 9568 10600 9580
rect 10555 9540 10600 9568
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9568 10839 9571
rect 11146 9568 11152 9580
rect 10827 9540 10916 9568
rect 11107 9540 11152 9568
rect 10827 9537 10839 9540
rect 10781 9531 10839 9537
rect 2958 9500 2964 9512
rect 2919 9472 2964 9500
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9500 3479 9503
rect 4154 9500 4160 9512
rect 3467 9472 4160 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 4154 9460 4160 9472
rect 4212 9500 4218 9512
rect 4798 9500 4804 9512
rect 4212 9472 4804 9500
rect 4212 9460 4218 9472
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 3234 9392 3240 9444
rect 3292 9432 3298 9444
rect 4065 9435 4123 9441
rect 4065 9432 4077 9435
rect 3292 9404 4077 9432
rect 3292 9392 3298 9404
rect 4065 9401 4077 9404
rect 4111 9401 4123 9435
rect 4065 9395 4123 9401
rect 6086 9392 6092 9444
rect 6144 9432 6150 9444
rect 10778 9432 10784 9444
rect 6144 9404 8892 9432
rect 10739 9404 10784 9432
rect 6144 9392 6150 9404
rect 3145 9367 3203 9373
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 3694 9364 3700 9376
rect 3191 9336 3700 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 3789 9367 3847 9373
rect 3789 9333 3801 9367
rect 3835 9364 3847 9367
rect 3878 9364 3884 9376
rect 3835 9336 3884 9364
rect 3835 9333 3847 9336
rect 3789 9327 3847 9333
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 8294 9364 8300 9376
rect 4028 9336 8300 9364
rect 4028 9324 4034 9336
rect 8294 9324 8300 9336
rect 8352 9364 8358 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8352 9336 8769 9364
rect 8352 9324 8358 9336
rect 8757 9333 8769 9336
rect 8803 9333 8815 9367
rect 8864 9364 8892 9404
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 8864 9336 10425 9364
rect 8757 9327 8815 9333
rect 10413 9333 10425 9336
rect 10459 9364 10471 9367
rect 10888 9364 10916 9540
rect 11146 9528 11152 9540
rect 11204 9528 11210 9580
rect 11532 9577 11560 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 12544 9636 12572 9676
rect 15197 9673 15209 9707
rect 15243 9704 15255 9707
rect 15286 9704 15292 9716
rect 15243 9676 15292 9704
rect 15243 9673 15255 9676
rect 15197 9667 15255 9673
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 16669 9707 16727 9713
rect 16669 9704 16681 9707
rect 16632 9676 16681 9704
rect 16632 9664 16638 9676
rect 16669 9673 16681 9676
rect 16715 9673 16727 9707
rect 16669 9667 16727 9673
rect 17313 9707 17371 9713
rect 17313 9673 17325 9707
rect 17359 9704 17371 9707
rect 17402 9704 17408 9716
rect 17359 9676 17408 9704
rect 17359 9673 17371 9676
rect 17313 9667 17371 9673
rect 12618 9636 12624 9648
rect 12544 9608 12624 9636
rect 12618 9596 12624 9608
rect 12676 9596 12682 9648
rect 13170 9596 13176 9648
rect 13228 9636 13234 9648
rect 13228 9608 13400 9636
rect 13228 9596 13234 9608
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 11784 9571 11842 9577
rect 11784 9537 11796 9571
rect 11830 9568 11842 9571
rect 12342 9568 12348 9580
rect 11830 9540 12348 9568
rect 11830 9537 11842 9540
rect 11784 9531 11842 9537
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 13372 9577 13400 9608
rect 14182 9596 14188 9648
rect 14240 9636 14246 9648
rect 14369 9639 14427 9645
rect 14369 9636 14381 9639
rect 14240 9608 14381 9636
rect 14240 9596 14246 9608
rect 14369 9605 14381 9608
rect 14415 9605 14427 9639
rect 14369 9599 14427 9605
rect 15105 9639 15163 9645
rect 15105 9605 15117 9639
rect 15151 9636 15163 9639
rect 15746 9636 15752 9648
rect 15151 9608 15752 9636
rect 15151 9605 15163 9608
rect 15105 9599 15163 9605
rect 15746 9596 15752 9608
rect 15804 9596 15810 9648
rect 16022 9636 16028 9648
rect 15983 9608 16028 9636
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 16684 9636 16712 9667
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 18230 9704 18236 9716
rect 17512 9676 18236 9704
rect 17512 9648 17540 9676
rect 18230 9664 18236 9676
rect 18288 9704 18294 9716
rect 18509 9707 18567 9713
rect 18509 9704 18521 9707
rect 18288 9676 18521 9704
rect 18288 9664 18294 9676
rect 18509 9673 18521 9676
rect 18555 9673 18567 9707
rect 18966 9704 18972 9716
rect 18927 9676 18972 9704
rect 18509 9667 18567 9673
rect 18966 9664 18972 9676
rect 19024 9664 19030 9716
rect 19426 9704 19432 9716
rect 19387 9676 19432 9704
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 20806 9704 20812 9716
rect 20767 9676 20812 9704
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 22281 9707 22339 9713
rect 22281 9673 22293 9707
rect 22327 9704 22339 9707
rect 22554 9704 22560 9716
rect 22327 9676 22560 9704
rect 22327 9673 22339 9676
rect 22281 9667 22339 9673
rect 22554 9664 22560 9676
rect 22612 9664 22618 9716
rect 22738 9664 22744 9716
rect 22796 9704 22802 9716
rect 23017 9707 23075 9713
rect 23017 9704 23029 9707
rect 22796 9676 23029 9704
rect 22796 9664 22802 9676
rect 23017 9673 23029 9676
rect 23063 9673 23075 9707
rect 23017 9667 23075 9673
rect 23106 9664 23112 9716
rect 23164 9704 23170 9716
rect 23164 9676 23209 9704
rect 23164 9664 23170 9676
rect 17494 9636 17500 9648
rect 16684 9608 17500 9636
rect 17494 9596 17500 9608
rect 17552 9596 17558 9648
rect 18049 9639 18107 9645
rect 18049 9605 18061 9639
rect 18095 9636 18107 9639
rect 18598 9636 18604 9648
rect 18095 9608 18604 9636
rect 18095 9605 18107 9608
rect 18049 9599 18107 9605
rect 18598 9596 18604 9608
rect 18656 9596 18662 9648
rect 19981 9639 20039 9645
rect 19981 9605 19993 9639
rect 20027 9636 20039 9639
rect 20070 9636 20076 9648
rect 20027 9608 20076 9636
rect 20027 9605 20039 9608
rect 19981 9599 20039 9605
rect 20070 9596 20076 9608
rect 20128 9636 20134 9648
rect 20254 9636 20260 9648
rect 20128 9608 20260 9636
rect 20128 9596 20134 9608
rect 20254 9596 20260 9608
rect 20312 9636 20318 9648
rect 20901 9639 20959 9645
rect 20901 9636 20913 9639
rect 20312 9608 20913 9636
rect 20312 9596 20318 9608
rect 20901 9605 20913 9608
rect 20947 9605 20959 9639
rect 20901 9599 20959 9605
rect 22189 9639 22247 9645
rect 22189 9605 22201 9639
rect 22235 9636 22247 9639
rect 22462 9636 22468 9648
rect 22235 9608 22468 9636
rect 22235 9605 22247 9608
rect 22189 9599 22247 9605
rect 22462 9596 22468 9608
rect 22520 9596 22526 9648
rect 23198 9596 23204 9648
rect 23256 9596 23262 9648
rect 13357 9571 13415 9577
rect 13357 9537 13369 9571
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 13725 9571 13783 9577
rect 13725 9537 13737 9571
rect 13771 9568 13783 9571
rect 13814 9568 13820 9580
rect 13771 9540 13820 9568
rect 13771 9537 13783 9540
rect 13725 9531 13783 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 15657 9571 15715 9577
rect 15657 9568 15669 9571
rect 13924 9540 15669 9568
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 13078 9500 13084 9512
rect 12768 9472 13084 9500
rect 12768 9460 12774 9472
rect 13078 9460 13084 9472
rect 13136 9500 13142 9512
rect 13173 9503 13231 9509
rect 13173 9500 13185 9503
rect 13136 9472 13185 9500
rect 13136 9460 13142 9472
rect 13173 9469 13185 9472
rect 13219 9500 13231 9503
rect 13538 9500 13544 9512
rect 13219 9472 13544 9500
rect 13219 9469 13231 9472
rect 13173 9463 13231 9469
rect 13538 9460 13544 9472
rect 13596 9500 13602 9512
rect 13924 9500 13952 9540
rect 15657 9537 15669 9540
rect 15703 9537 15715 9571
rect 15657 9531 15715 9537
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9537 15899 9571
rect 15841 9531 15899 9537
rect 17221 9571 17279 9577
rect 17221 9537 17233 9571
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 14090 9500 14096 9512
rect 13596 9472 13952 9500
rect 14051 9472 14096 9500
rect 13596 9460 13602 9472
rect 14090 9460 14096 9472
rect 14148 9460 14154 9512
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9469 14335 9503
rect 14277 9463 14335 9469
rect 12802 9392 12808 9444
rect 12860 9432 12866 9444
rect 12897 9435 12955 9441
rect 12897 9432 12909 9435
rect 12860 9404 12909 9432
rect 12860 9392 12866 9404
rect 12897 9401 12909 9404
rect 12943 9401 12955 9435
rect 12897 9395 12955 9401
rect 13909 9435 13967 9441
rect 13909 9401 13921 9435
rect 13955 9432 13967 9435
rect 14292 9432 14320 9463
rect 14734 9460 14740 9512
rect 14792 9460 14798 9512
rect 15010 9500 15016 9512
rect 14971 9472 15016 9500
rect 15010 9460 15016 9472
rect 15068 9500 15074 9512
rect 15746 9500 15752 9512
rect 15068 9472 15752 9500
rect 15068 9460 15074 9472
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 13955 9404 14320 9432
rect 14752 9432 14780 9460
rect 15856 9432 15884 9531
rect 14752 9404 15884 9432
rect 17236 9432 17264 9531
rect 17310 9528 17316 9580
rect 17368 9568 17374 9580
rect 19058 9568 19064 9580
rect 17368 9540 19064 9568
rect 17368 9528 17374 9540
rect 19058 9528 19064 9540
rect 19116 9528 19122 9580
rect 23216 9568 23244 9596
rect 23661 9571 23719 9577
rect 23661 9568 23673 9571
rect 21560 9540 22416 9568
rect 23216 9540 23673 9568
rect 17402 9500 17408 9512
rect 17363 9472 17408 9500
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 18138 9500 18144 9512
rect 18099 9472 18144 9500
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 18785 9503 18843 9509
rect 18785 9500 18797 9503
rect 18288 9472 18797 9500
rect 18288 9460 18294 9472
rect 18785 9469 18797 9472
rect 18831 9469 18843 9503
rect 20070 9500 20076 9512
rect 20031 9472 20076 9500
rect 18785 9463 18843 9469
rect 17681 9435 17739 9441
rect 17681 9432 17693 9435
rect 17236 9404 17693 9432
rect 13955 9401 13967 9404
rect 13909 9395 13967 9401
rect 17681 9401 17693 9404
rect 17727 9401 17739 9435
rect 18800 9432 18828 9463
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 20165 9503 20223 9509
rect 20165 9469 20177 9503
rect 20211 9469 20223 9503
rect 20990 9500 20996 9512
rect 20951 9472 20996 9500
rect 20165 9463 20223 9469
rect 20180 9432 20208 9463
rect 20990 9460 20996 9472
rect 21048 9500 21054 9512
rect 21560 9509 21588 9540
rect 22388 9509 22416 9540
rect 23661 9537 23673 9540
rect 23707 9537 23719 9571
rect 23661 9531 23719 9537
rect 21361 9503 21419 9509
rect 21361 9500 21373 9503
rect 21048 9472 21373 9500
rect 21048 9460 21054 9472
rect 21361 9469 21373 9472
rect 21407 9500 21419 9503
rect 21545 9503 21603 9509
rect 21545 9500 21557 9503
rect 21407 9472 21557 9500
rect 21407 9469 21419 9472
rect 21361 9463 21419 9469
rect 21545 9469 21557 9472
rect 21591 9469 21603 9503
rect 21545 9463 21603 9469
rect 22373 9503 22431 9509
rect 22373 9469 22385 9503
rect 22419 9500 22431 9503
rect 23201 9503 23259 9509
rect 23201 9500 23213 9503
rect 22419 9472 23213 9500
rect 22419 9469 22431 9472
rect 22373 9463 22431 9469
rect 23201 9469 23213 9472
rect 23247 9469 23259 9503
rect 23201 9463 23259 9469
rect 23477 9503 23535 9509
rect 23477 9469 23489 9503
rect 23523 9469 23535 9503
rect 23477 9463 23535 9469
rect 18800 9404 20208 9432
rect 17681 9395 17739 9401
rect 20346 9392 20352 9444
rect 20404 9432 20410 9444
rect 23492 9432 23520 9463
rect 20404 9404 23520 9432
rect 20404 9392 20410 9404
rect 13354 9364 13360 9376
rect 10459 9336 13360 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 13541 9367 13599 9373
rect 13541 9333 13553 9367
rect 13587 9364 13599 9367
rect 14366 9364 14372 9376
rect 13587 9336 14372 9364
rect 13587 9333 13599 9336
rect 13541 9327 13599 9333
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 14737 9367 14795 9373
rect 14737 9364 14749 9367
rect 14516 9336 14749 9364
rect 14516 9324 14522 9336
rect 14737 9333 14749 9336
rect 14783 9333 14795 9367
rect 15562 9364 15568 9376
rect 15523 9336 15568 9364
rect 14737 9327 14795 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 15746 9324 15752 9376
rect 15804 9364 15810 9376
rect 16298 9364 16304 9376
rect 15804 9336 16304 9364
rect 15804 9324 15810 9336
rect 16298 9324 16304 9336
rect 16356 9364 16362 9376
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 16356 9336 16405 9364
rect 16356 9324 16362 9336
rect 16393 9333 16405 9336
rect 16439 9333 16451 9367
rect 16850 9364 16856 9376
rect 16811 9336 16856 9364
rect 16393 9327 16451 9333
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 19610 9364 19616 9376
rect 19571 9336 19616 9364
rect 19610 9324 19616 9336
rect 19668 9324 19674 9376
rect 20438 9364 20444 9376
rect 20399 9336 20444 9364
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 21726 9324 21732 9376
rect 21784 9364 21790 9376
rect 21821 9367 21879 9373
rect 21821 9364 21833 9367
rect 21784 9336 21833 9364
rect 21784 9324 21790 9336
rect 21821 9333 21833 9336
rect 21867 9333 21879 9367
rect 22646 9364 22652 9376
rect 22607 9336 22652 9364
rect 21821 9327 21879 9333
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 23474 9324 23480 9376
rect 23532 9364 23538 9376
rect 23845 9367 23903 9373
rect 23845 9364 23857 9367
rect 23532 9336 23857 9364
rect 23532 9324 23538 9336
rect 23845 9333 23857 9336
rect 23891 9333 23903 9367
rect 23845 9327 23903 9333
rect 1104 9274 26220 9296
rect 1104 9222 5136 9274
rect 5188 9222 5200 9274
rect 5252 9222 5264 9274
rect 5316 9222 5328 9274
rect 5380 9222 5392 9274
rect 5444 9222 13508 9274
rect 13560 9222 13572 9274
rect 13624 9222 13636 9274
rect 13688 9222 13700 9274
rect 13752 9222 13764 9274
rect 13816 9222 21880 9274
rect 21932 9222 21944 9274
rect 21996 9222 22008 9274
rect 22060 9222 22072 9274
rect 22124 9222 22136 9274
rect 22188 9222 26220 9274
rect 1104 9200 26220 9222
rect 2593 9163 2651 9169
rect 2593 9129 2605 9163
rect 2639 9160 2651 9163
rect 3050 9160 3056 9172
rect 2639 9132 3056 9160
rect 2639 9129 2651 9132
rect 2593 9123 2651 9129
rect 3050 9120 3056 9132
rect 3108 9120 3114 9172
rect 3234 9160 3240 9172
rect 3195 9132 3240 9160
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3878 9160 3884 9172
rect 3839 9132 3884 9160
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 5997 9163 6055 9169
rect 5997 9160 6009 9163
rect 5592 9132 6009 9160
rect 5592 9120 5598 9132
rect 5997 9129 6009 9132
rect 6043 9160 6055 9163
rect 6086 9160 6092 9172
rect 6043 9132 6092 9160
rect 6043 9129 6055 9132
rect 5997 9123 6055 9129
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 7834 9160 7840 9172
rect 7795 9132 7840 9160
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 12069 9163 12127 9169
rect 12069 9129 12081 9163
rect 12115 9160 12127 9163
rect 12526 9160 12532 9172
rect 12115 9132 12532 9160
rect 12115 9129 12127 9132
rect 12069 9123 12127 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 13354 9120 13360 9172
rect 13412 9160 13418 9172
rect 15194 9160 15200 9172
rect 13412 9132 15200 9160
rect 13412 9120 13418 9132
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 16298 9120 16304 9172
rect 16356 9160 16362 9172
rect 17221 9163 17279 9169
rect 17221 9160 17233 9163
rect 16356 9132 17233 9160
rect 16356 9120 16362 9132
rect 17221 9129 17233 9132
rect 17267 9160 17279 9163
rect 17313 9163 17371 9169
rect 17313 9160 17325 9163
rect 17267 9132 17325 9160
rect 17267 9129 17279 9132
rect 17221 9123 17279 9129
rect 17313 9129 17325 9132
rect 17359 9160 17371 9163
rect 17402 9160 17408 9172
rect 17359 9132 17408 9160
rect 17359 9129 17371 9132
rect 17313 9123 17371 9129
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 18877 9163 18935 9169
rect 18877 9160 18889 9163
rect 18196 9132 18889 9160
rect 18196 9120 18202 9132
rect 18877 9129 18889 9132
rect 18923 9129 18935 9163
rect 18877 9123 18935 9129
rect 20070 9120 20076 9172
rect 20128 9160 20134 9172
rect 20625 9163 20683 9169
rect 20625 9160 20637 9163
rect 20128 9132 20637 9160
rect 20128 9120 20134 9132
rect 20625 9129 20637 9132
rect 20671 9129 20683 9163
rect 20625 9123 20683 9129
rect 22922 9120 22928 9172
rect 22980 9160 22986 9172
rect 23293 9163 23351 9169
rect 23293 9160 23305 9163
rect 22980 9132 23305 9160
rect 22980 9120 22986 9132
rect 23293 9129 23305 9132
rect 23339 9129 23351 9163
rect 23293 9123 23351 9129
rect 4062 9092 4068 9104
rect 3068 9064 4068 9092
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3068 9024 3096 9064
rect 4062 9052 4068 9064
rect 4120 9052 4126 9104
rect 4525 9095 4583 9101
rect 4525 9061 4537 9095
rect 4571 9061 4583 9095
rect 12342 9092 12348 9104
rect 12303 9064 12348 9092
rect 4525 9055 4583 9061
rect 2832 8996 3096 9024
rect 2832 8984 2838 8996
rect 2409 8959 2467 8965
rect 2409 8925 2421 8959
rect 2455 8925 2467 8959
rect 2958 8956 2964 8968
rect 2919 8928 2964 8956
rect 2409 8919 2467 8925
rect 2424 8888 2452 8919
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 3068 8965 3096 8996
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 9024 3387 9027
rect 3789 9027 3847 9033
rect 3789 9024 3801 9027
rect 3375 8996 3801 9024
rect 3375 8993 3387 8996
rect 3329 8987 3387 8993
rect 3789 8993 3801 8996
rect 3835 9024 3847 9027
rect 4338 9024 4344 9036
rect 3835 8996 4344 9024
rect 3835 8993 3847 8996
rect 3789 8987 3847 8993
rect 4338 8984 4344 8996
rect 4396 9024 4402 9036
rect 4540 9024 4568 9055
rect 12342 9052 12348 9064
rect 12400 9052 12406 9104
rect 12710 9092 12716 9104
rect 12671 9064 12716 9092
rect 12710 9052 12716 9064
rect 12768 9052 12774 9104
rect 12802 9052 12808 9104
rect 12860 9052 12866 9104
rect 13556 9064 20116 9092
rect 4396 8996 4568 9024
rect 11793 9027 11851 9033
rect 4396 8984 4402 8996
rect 11793 8993 11805 9027
rect 11839 9024 11851 9027
rect 12820 9024 12848 9052
rect 11839 8996 12112 9024
rect 12820 8996 13400 9024
rect 11839 8993 11851 8996
rect 11793 8987 11851 8993
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8925 3663 8959
rect 4062 8956 4068 8968
rect 4023 8928 4068 8956
rect 3605 8919 3663 8925
rect 3620 8888 3648 8919
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4614 8956 4620 8968
rect 4203 8928 4620 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 4724 8888 4752 8919
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 5040 8928 5181 8956
rect 5040 8916 5046 8928
rect 5169 8925 5181 8928
rect 5215 8925 5227 8959
rect 6178 8956 6184 8968
rect 6139 8928 6184 8956
rect 5169 8919 5227 8925
rect 6178 8916 6184 8928
rect 6236 8916 6242 8968
rect 7466 8956 7472 8968
rect 7427 8928 7472 8956
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 7834 8956 7840 8968
rect 7699 8928 7840 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 12084 8956 12112 8996
rect 11204 8928 11928 8956
rect 12084 8928 12388 8956
rect 11204 8916 11210 8928
rect 5626 8888 5632 8900
rect 2424 8860 5632 8888
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 8386 8848 8392 8900
rect 8444 8888 8450 8900
rect 11900 8897 11928 8928
rect 11425 8891 11483 8897
rect 11425 8888 11437 8891
rect 8444 8860 11437 8888
rect 8444 8848 8450 8860
rect 11425 8857 11437 8860
rect 11471 8857 11483 8891
rect 11425 8851 11483 8857
rect 11885 8891 11943 8897
rect 11885 8857 11897 8891
rect 11931 8888 11943 8891
rect 12066 8888 12072 8900
rect 11931 8860 12072 8888
rect 11931 8857 11943 8860
rect 11885 8851 11943 8857
rect 12066 8848 12072 8860
rect 12124 8848 12130 8900
rect 12360 8888 12388 8928
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 12492 8928 12541 8956
rect 12492 8916 12498 8928
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 12618 8916 12624 8968
rect 12676 8956 12682 8968
rect 12676 8928 12721 8956
rect 12676 8916 12682 8928
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 13372 8965 13400 8996
rect 12989 8959 13047 8965
rect 12860 8928 12905 8956
rect 12860 8916 12866 8928
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13173 8959 13231 8965
rect 13173 8956 13185 8959
rect 13035 8928 13185 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 13173 8925 13185 8928
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 13556 8888 13584 9064
rect 14642 9024 14648 9036
rect 13648 8996 14648 9024
rect 13648 8965 13676 8996
rect 14642 8984 14648 8996
rect 14700 9024 14706 9036
rect 15010 9024 15016 9036
rect 14700 8996 15016 9024
rect 14700 8984 14706 8996
rect 15010 8984 15016 8996
rect 15068 9024 15074 9036
rect 18340 9033 18368 9064
rect 15197 9027 15255 9033
rect 15197 9024 15209 9027
rect 15068 8996 15209 9024
rect 15068 8984 15074 8996
rect 15197 8993 15209 8996
rect 15243 8993 15255 9027
rect 15197 8987 15255 8993
rect 17221 9027 17279 9033
rect 17221 8993 17233 9027
rect 17267 9024 17279 9027
rect 17589 9027 17647 9033
rect 17589 9024 17601 9027
rect 17267 8996 17601 9024
rect 17267 8993 17279 8996
rect 17221 8987 17279 8993
rect 17589 8993 17601 8996
rect 17635 8993 17647 9027
rect 17589 8987 17647 8993
rect 18325 9027 18383 9033
rect 18325 8993 18337 9027
rect 18371 8993 18383 9027
rect 19705 9027 19763 9033
rect 19705 9024 19717 9027
rect 18325 8987 18383 8993
rect 18616 8996 19717 9024
rect 18616 8968 18644 8996
rect 19705 8993 19717 8996
rect 19751 8993 19763 9027
rect 19886 9024 19892 9036
rect 19847 8996 19892 9024
rect 19705 8987 19763 8993
rect 19886 8984 19892 8996
rect 19944 8984 19950 9036
rect 20088 9033 20116 9064
rect 20073 9027 20131 9033
rect 20073 8993 20085 9027
rect 20119 9024 20131 9027
rect 20346 9024 20352 9036
rect 20119 8996 20352 9024
rect 20119 8993 20131 8996
rect 20073 8987 20131 8993
rect 20346 8984 20352 8996
rect 20404 8984 20410 9036
rect 23017 9027 23075 9033
rect 23017 9024 23029 9027
rect 22296 8996 23029 9024
rect 13633 8959 13691 8965
rect 13633 8925 13645 8959
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 13909 8959 13967 8965
rect 13909 8956 13921 8959
rect 13780 8928 13921 8956
rect 13780 8916 13786 8928
rect 13909 8925 13921 8928
rect 13955 8925 13967 8959
rect 14458 8956 14464 8968
rect 14419 8928 14464 8956
rect 13909 8919 13967 8925
rect 13924 8888 13952 8919
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8956 14611 8959
rect 14734 8956 14740 8968
rect 14599 8928 14740 8956
rect 14599 8925 14611 8928
rect 14553 8919 14611 8925
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 14921 8959 14979 8965
rect 14921 8925 14933 8959
rect 14967 8925 14979 8959
rect 14921 8919 14979 8925
rect 14936 8888 14964 8919
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17773 8959 17831 8965
rect 17773 8956 17785 8959
rect 17368 8928 17785 8956
rect 17368 8916 17374 8928
rect 17773 8925 17785 8928
rect 17819 8925 17831 8959
rect 17773 8919 17831 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8956 18567 8959
rect 18598 8956 18604 8968
rect 18555 8928 18604 8956
rect 18555 8925 18567 8928
rect 18509 8919 18567 8925
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8956 18751 8959
rect 19061 8959 19119 8965
rect 19061 8956 19073 8959
rect 18739 8928 19073 8956
rect 18739 8925 18751 8928
rect 18693 8919 18751 8925
rect 19061 8925 19073 8928
rect 19107 8925 19119 8959
rect 19610 8956 19616 8968
rect 19571 8928 19616 8956
rect 19061 8919 19119 8925
rect 19610 8916 19616 8928
rect 19668 8916 19674 8968
rect 20254 8956 20260 8968
rect 20215 8928 20260 8956
rect 20254 8916 20260 8928
rect 20312 8916 20318 8968
rect 20441 8959 20499 8965
rect 20441 8925 20453 8959
rect 20487 8956 20499 8959
rect 20809 8959 20867 8965
rect 20809 8956 20821 8959
rect 20487 8928 20821 8956
rect 20487 8925 20499 8928
rect 20441 8919 20499 8925
rect 20809 8925 20821 8928
rect 20855 8925 20867 8959
rect 20809 8919 20867 8925
rect 12360 8860 13768 8888
rect 13924 8860 14964 8888
rect 2682 8780 2688 8832
rect 2740 8820 2746 8832
rect 2777 8823 2835 8829
rect 2777 8820 2789 8823
rect 2740 8792 2789 8820
rect 2740 8780 2746 8792
rect 2777 8789 2789 8792
rect 2823 8789 2835 8823
rect 2777 8783 2835 8789
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 3326 8820 3332 8832
rect 2924 8792 3332 8820
rect 2924 8780 2930 8792
rect 3326 8780 3332 8792
rect 3384 8820 3390 8832
rect 3513 8823 3571 8829
rect 3513 8820 3525 8823
rect 3384 8792 3525 8820
rect 3384 8780 3390 8792
rect 3513 8789 3525 8792
rect 3559 8789 3571 8823
rect 3513 8783 3571 8789
rect 3602 8780 3608 8832
rect 3660 8820 3666 8832
rect 4341 8823 4399 8829
rect 4341 8820 4353 8823
rect 3660 8792 4353 8820
rect 3660 8780 3666 8792
rect 4341 8789 4353 8792
rect 4387 8789 4399 8823
rect 4341 8783 4399 8789
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 5353 8823 5411 8829
rect 5353 8820 5365 8823
rect 4948 8792 5365 8820
rect 4948 8780 4954 8792
rect 5353 8789 5365 8792
rect 5399 8789 5411 8823
rect 7374 8820 7380 8832
rect 7335 8792 7380 8820
rect 5353 8783 5411 8789
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 11698 8820 11704 8832
rect 11659 8792 11704 8820
rect 11698 8780 11704 8792
rect 11756 8820 11762 8832
rect 13262 8820 13268 8832
rect 11756 8792 13268 8820
rect 11756 8780 11762 8792
rect 13262 8780 13268 8792
rect 13320 8820 13326 8832
rect 13740 8829 13768 8860
rect 17586 8848 17592 8900
rect 17644 8888 17650 8900
rect 17865 8891 17923 8897
rect 17865 8888 17877 8891
rect 17644 8860 17877 8888
rect 17644 8848 17650 8860
rect 17865 8857 17877 8860
rect 17911 8857 17923 8891
rect 17865 8851 17923 8857
rect 19886 8848 19892 8900
rect 19944 8888 19950 8900
rect 20901 8891 20959 8897
rect 20901 8888 20913 8891
rect 19944 8860 20913 8888
rect 19944 8848 19950 8860
rect 20901 8857 20913 8860
rect 20947 8888 20959 8891
rect 20990 8888 20996 8900
rect 20947 8860 20996 8888
rect 20947 8857 20959 8860
rect 20901 8851 20959 8857
rect 20990 8848 20996 8860
rect 21048 8888 21054 8900
rect 22296 8897 22324 8996
rect 23017 8993 23029 8996
rect 23063 8993 23075 9027
rect 23017 8987 23075 8993
rect 22830 8956 22836 8968
rect 22791 8928 22836 8956
rect 22830 8916 22836 8928
rect 22888 8916 22894 8968
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8956 22983 8959
rect 23198 8956 23204 8968
rect 22971 8928 23204 8956
rect 22971 8925 22983 8928
rect 22925 8919 22983 8925
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 23474 8956 23480 8968
rect 23435 8928 23480 8956
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 21085 8891 21143 8897
rect 21085 8888 21097 8891
rect 21048 8860 21097 8888
rect 21048 8848 21054 8860
rect 21085 8857 21097 8860
rect 21131 8888 21143 8891
rect 21637 8891 21695 8897
rect 21637 8888 21649 8891
rect 21131 8860 21649 8888
rect 21131 8857 21143 8860
rect 21085 8851 21143 8857
rect 21637 8857 21649 8860
rect 21683 8888 21695 8891
rect 22281 8891 22339 8897
rect 22281 8888 22293 8891
rect 21683 8860 22293 8888
rect 21683 8857 21695 8860
rect 21637 8851 21695 8857
rect 22281 8857 22293 8860
rect 22327 8857 22339 8891
rect 22281 8851 22339 8857
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13320 8792 13553 8820
rect 13320 8780 13326 8792
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 13541 8783 13599 8789
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8789 13783 8823
rect 14090 8820 14096 8832
rect 14051 8792 14096 8820
rect 13725 8783 13783 8789
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 15105 8823 15163 8829
rect 15105 8789 15117 8823
rect 15151 8820 15163 8823
rect 16390 8820 16396 8832
rect 15151 8792 16396 8820
rect 15151 8789 15163 8792
rect 15105 8783 15163 8789
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 18046 8780 18052 8832
rect 18104 8820 18110 8832
rect 18233 8823 18291 8829
rect 18233 8820 18245 8823
rect 18104 8792 18245 8820
rect 18104 8780 18110 8792
rect 18233 8789 18245 8792
rect 18279 8789 18291 8823
rect 19242 8820 19248 8832
rect 19203 8792 19248 8820
rect 18233 8783 18291 8789
rect 19242 8780 19248 8792
rect 19300 8780 19306 8832
rect 22462 8820 22468 8832
rect 22423 8792 22468 8820
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 1104 8730 26220 8752
rect 1104 8678 9322 8730
rect 9374 8678 9386 8730
rect 9438 8678 9450 8730
rect 9502 8678 9514 8730
rect 9566 8678 9578 8730
rect 9630 8678 17694 8730
rect 17746 8678 17758 8730
rect 17810 8678 17822 8730
rect 17874 8678 17886 8730
rect 17938 8678 17950 8730
rect 18002 8678 26220 8730
rect 1104 8656 26220 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 2958 8616 2964 8628
rect 1627 8588 2964 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 4433 8619 4491 8625
rect 4433 8585 4445 8619
rect 4479 8616 4491 8619
rect 4614 8616 4620 8628
rect 4479 8588 4620 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 5994 8616 6000 8628
rect 5955 8588 6000 8616
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 9214 8616 9220 8628
rect 7616 8588 9220 8616
rect 7616 8576 7622 8588
rect 9214 8576 9220 8588
rect 9272 8616 9278 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 9272 8588 9321 8616
rect 9272 8576 9278 8588
rect 9309 8585 9321 8588
rect 9355 8585 9367 8619
rect 9309 8579 9367 8585
rect 10778 8576 10784 8628
rect 10836 8616 10842 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 10836 8588 11805 8616
rect 10836 8576 10842 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 11793 8579 11851 8585
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 12802 8616 12808 8628
rect 12492 8588 12537 8616
rect 12763 8588 12808 8616
rect 12492 8576 12498 8588
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 13078 8616 13084 8628
rect 13039 8588 13084 8616
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 13771 8588 14289 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 14277 8585 14289 8588
rect 14323 8585 14335 8619
rect 14277 8579 14335 8585
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15436 8588 15669 8616
rect 15436 8576 15442 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 19061 8619 19119 8625
rect 19061 8616 19073 8619
rect 17460 8588 19073 8616
rect 17460 8576 17466 8588
rect 19061 8585 19073 8588
rect 19107 8616 19119 8619
rect 19886 8616 19892 8628
rect 19107 8588 19892 8616
rect 19107 8585 19119 8588
rect 19061 8579 19119 8585
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 8478 8548 8484 8560
rect 3068 8520 3924 8548
rect 2682 8440 2688 8492
rect 2740 8489 2746 8492
rect 3068 8489 3096 8520
rect 3896 8492 3924 8520
rect 7116 8520 8484 8548
rect 2740 8480 2752 8489
rect 2961 8483 3019 8489
rect 2740 8452 2785 8480
rect 2740 8443 2752 8452
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 3053 8483 3111 8489
rect 3053 8480 3065 8483
rect 3007 8452 3065 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 3053 8449 3065 8452
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3320 8483 3378 8489
rect 3320 8449 3332 8483
rect 3366 8480 3378 8483
rect 3602 8480 3608 8492
rect 3366 8452 3608 8480
rect 3366 8449 3378 8452
rect 3320 8443 3378 8449
rect 2740 8440 2746 8443
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 3936 8452 4629 8480
rect 3936 8440 3942 8452
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 4873 8483 4931 8489
rect 4873 8480 4885 8483
rect 4764 8452 4885 8480
rect 4764 8440 4770 8452
rect 4873 8449 4885 8452
rect 4919 8449 4931 8483
rect 4873 8443 4931 8449
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 6730 8480 6736 8492
rect 5776 8452 6736 8480
rect 5776 8440 5782 8452
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7116 8489 7144 8520
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 9766 8548 9772 8560
rect 9048 8520 9772 8548
rect 7374 8489 7380 8492
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8449 7159 8483
rect 7368 8480 7380 8489
rect 7335 8452 7380 8480
rect 7101 8443 7159 8449
rect 7368 8443 7380 8452
rect 7374 8440 7380 8443
rect 7432 8440 7438 8492
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 9048 8489 9076 8520
rect 9766 8508 9772 8520
rect 9824 8548 9830 8560
rect 12621 8551 12679 8557
rect 12621 8548 12633 8551
rect 9824 8520 12633 8548
rect 9824 8508 9830 8520
rect 12621 8517 12633 8520
rect 12667 8517 12679 8551
rect 12621 8511 12679 8517
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8812 8452 8861 8480
rect 8812 8440 8818 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8449 9091 8483
rect 9214 8480 9220 8492
rect 9175 8452 9220 8480
rect 9033 8443 9091 8449
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11848 8452 11897 8480
rect 11848 8440 11854 8452
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 12250 8480 12256 8492
rect 11885 8443 11943 8449
rect 12084 8452 12256 8480
rect 6546 8412 6552 8424
rect 6507 8384 6552 8412
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 11333 8415 11391 8421
rect 11333 8381 11345 8415
rect 11379 8412 11391 8415
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 11379 8384 11713 8412
rect 11379 8381 11391 8384
rect 11333 8375 11391 8381
rect 11701 8381 11713 8384
rect 11747 8412 11759 8415
rect 11974 8412 11980 8424
rect 11747 8384 11980 8412
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 5684 8316 7052 8344
rect 5684 8304 5690 8316
rect 6914 8276 6920 8288
rect 6875 8248 6920 8276
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 7024 8276 7052 8316
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 8481 8347 8539 8353
rect 8481 8344 8493 8347
rect 8352 8316 8493 8344
rect 8352 8304 8358 8316
rect 8481 8313 8493 8316
rect 8527 8313 8539 8347
rect 8846 8344 8852 8356
rect 8807 8316 8852 8344
rect 8481 8307 8539 8313
rect 8846 8304 8852 8316
rect 8904 8304 8910 8356
rect 9030 8276 9036 8288
rect 7024 8248 9036 8276
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 11606 8236 11612 8288
rect 11664 8276 11670 8288
rect 12084 8276 12112 8452
rect 12250 8440 12256 8452
rect 12308 8480 12314 8492
rect 12820 8480 12848 8576
rect 13170 8508 13176 8560
rect 13228 8548 13234 8560
rect 13817 8551 13875 8557
rect 13817 8548 13829 8551
rect 13228 8520 13829 8548
rect 13228 8508 13234 8520
rect 13817 8517 13829 8520
rect 13863 8517 13875 8551
rect 13817 8511 13875 8517
rect 12308 8452 12848 8480
rect 13265 8483 13323 8489
rect 12308 8440 12314 8452
rect 13265 8449 13277 8483
rect 13311 8480 13323 8483
rect 13722 8480 13728 8492
rect 13311 8452 13728 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12216 8384 12909 8412
rect 12216 8372 12222 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 12621 8347 12679 8353
rect 12621 8313 12633 8347
rect 12667 8344 12679 8347
rect 13280 8344 13308 8443
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 14366 8440 14372 8492
rect 14424 8480 14430 8492
rect 14461 8483 14519 8489
rect 14461 8480 14473 8483
rect 14424 8452 14473 8480
rect 14424 8440 14430 8452
rect 14461 8449 14473 8452
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 12667 8316 13308 8344
rect 12667 8313 12679 8316
rect 12621 8307 12679 8313
rect 12250 8276 12256 8288
rect 11664 8248 12112 8276
rect 12211 8248 12256 8276
rect 11664 8236 11670 8248
rect 12250 8236 12256 8248
rect 12308 8236 12314 8288
rect 13078 8236 13084 8288
rect 13136 8276 13142 8288
rect 13354 8276 13360 8288
rect 13136 8248 13360 8276
rect 13136 8236 13142 8248
rect 13354 8236 13360 8248
rect 13412 8276 13418 8288
rect 13556 8276 13584 8375
rect 14829 8347 14887 8353
rect 14829 8313 14841 8347
rect 14875 8344 14887 8347
rect 14875 8316 16160 8344
rect 14875 8313 14887 8316
rect 14829 8307 14887 8313
rect 16132 8288 16160 8316
rect 14182 8276 14188 8288
rect 13412 8248 13584 8276
rect 14143 8248 14188 8276
rect 13412 8236 13418 8248
rect 14182 8236 14188 8248
rect 14240 8236 14246 8288
rect 14642 8276 14648 8288
rect 14603 8248 14648 8276
rect 14642 8236 14648 8248
rect 14700 8236 14706 8288
rect 16114 8276 16120 8288
rect 16075 8248 16120 8276
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 22097 8279 22155 8285
rect 22097 8245 22109 8279
rect 22143 8276 22155 8279
rect 22278 8276 22284 8288
rect 22143 8248 22284 8276
rect 22143 8245 22155 8248
rect 22097 8239 22155 8245
rect 22278 8236 22284 8248
rect 22336 8236 22342 8288
rect 1104 8186 26220 8208
rect 1104 8134 5136 8186
rect 5188 8134 5200 8186
rect 5252 8134 5264 8186
rect 5316 8134 5328 8186
rect 5380 8134 5392 8186
rect 5444 8134 13508 8186
rect 13560 8134 13572 8186
rect 13624 8134 13636 8186
rect 13688 8134 13700 8186
rect 13752 8134 13764 8186
rect 13816 8134 21880 8186
rect 21932 8134 21944 8186
rect 21996 8134 22008 8186
rect 22060 8134 22072 8186
rect 22124 8134 22136 8186
rect 22188 8134 26220 8186
rect 1104 8112 26220 8134
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4706 8072 4712 8084
rect 4571 8044 4712 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5353 8075 5411 8081
rect 5353 8072 5365 8075
rect 5040 8044 5365 8072
rect 5040 8032 5046 8044
rect 5353 8041 5365 8044
rect 5399 8041 5411 8075
rect 5353 8035 5411 8041
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 6546 8072 6552 8084
rect 6503 8044 6552 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 6972 8044 8125 8072
rect 6972 8032 6978 8044
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 8113 8035 8171 8041
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 8444 8044 8585 8072
rect 8444 8032 8450 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 8938 8032 8944 8084
rect 8996 8072 9002 8084
rect 9217 8075 9275 8081
rect 9217 8072 9229 8075
rect 8996 8044 9229 8072
rect 8996 8032 9002 8044
rect 9217 8041 9229 8044
rect 9263 8041 9275 8075
rect 9766 8072 9772 8084
rect 9217 8035 9275 8041
rect 9324 8044 9628 8072
rect 9727 8044 9772 8072
rect 4154 8004 4160 8016
rect 3252 7976 4160 8004
rect 2866 7868 2872 7880
rect 2827 7840 2872 7868
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 3252 7877 3280 7976
rect 4154 7964 4160 7976
rect 4212 7964 4218 8016
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 7377 8007 7435 8013
rect 7377 8004 7389 8007
rect 6788 7976 7389 8004
rect 6788 7964 6794 7976
rect 7377 7973 7389 7976
rect 7423 7973 7435 8007
rect 7377 7967 7435 7973
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7936 3571 7939
rect 4801 7939 4859 7945
rect 4801 7936 4813 7939
rect 3559 7908 4813 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 4801 7905 4813 7908
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 5994 7936 6000 7948
rect 5215 7908 6000 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 2774 7800 2780 7812
rect 2700 7772 2780 7800
rect 2700 7741 2728 7772
rect 2774 7760 2780 7772
rect 2832 7800 2838 7812
rect 3344 7800 3372 7831
rect 2832 7772 3372 7800
rect 3620 7800 3648 7831
rect 3694 7828 3700 7880
rect 3752 7868 3758 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3752 7840 3985 7868
rect 3752 7828 3758 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 4338 7868 4344 7880
rect 4396 7877 4402 7880
rect 3973 7831 4031 7837
rect 4080 7840 4344 7868
rect 4080 7800 4108 7840
rect 4338 7828 4344 7840
rect 4396 7868 4404 7877
rect 4982 7868 4988 7880
rect 4396 7840 4489 7868
rect 4943 7840 4988 7868
rect 4396 7831 4404 7840
rect 4396 7828 4402 7831
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 3620 7772 4108 7800
rect 4157 7803 4215 7809
rect 2832 7760 2838 7772
rect 4157 7769 4169 7803
rect 4203 7769 4215 7803
rect 4157 7763 4215 7769
rect 4249 7803 4307 7809
rect 4249 7769 4261 7803
rect 4295 7800 4307 7803
rect 5184 7800 5212 7899
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 7006 7896 7012 7948
rect 7064 7936 7070 7948
rect 7392 7936 7420 7967
rect 7466 7964 7472 8016
rect 7524 8004 7530 8016
rect 7653 8007 7711 8013
rect 7653 8004 7665 8007
rect 7524 7976 7665 8004
rect 7524 7964 7530 7976
rect 7653 7973 7665 7976
rect 7699 7973 7711 8007
rect 8754 8004 8760 8016
rect 7653 7967 7711 7973
rect 8128 7976 8760 8004
rect 8128 7936 8156 7976
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 9030 8004 9036 8016
rect 8991 7976 9036 8004
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 7064 7908 7109 7936
rect 7392 7908 8156 7936
rect 8205 7939 8263 7945
rect 7064 7896 7070 7908
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 8846 7936 8852 7948
rect 8251 7908 8852 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 9324 7945 9352 8044
rect 9600 8004 9628 8044
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 10229 8075 10287 8081
rect 10229 8041 10241 8075
rect 10275 8072 10287 8075
rect 11974 8072 11980 8084
rect 10275 8044 11980 8072
rect 10275 8041 10287 8044
rect 10229 8035 10287 8041
rect 9858 8004 9864 8016
rect 9600 7976 9864 8004
rect 9858 7964 9864 7976
rect 9916 8004 9922 8016
rect 10244 8004 10272 8035
rect 11974 8032 11980 8044
rect 12032 8072 12038 8084
rect 13078 8072 13084 8084
rect 12032 8044 13084 8072
rect 12032 8032 12038 8044
rect 13078 8032 13084 8044
rect 13136 8072 13142 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 13136 8044 13277 8072
rect 13136 8032 13142 8044
rect 13265 8041 13277 8044
rect 13311 8041 13323 8075
rect 13265 8035 13323 8041
rect 18141 8075 18199 8081
rect 18141 8041 18153 8075
rect 18187 8072 18199 8075
rect 18230 8072 18236 8084
rect 18187 8044 18236 8072
rect 18187 8041 18199 8044
rect 18141 8035 18199 8041
rect 18230 8032 18236 8044
rect 18288 8032 18294 8084
rect 9916 7976 10272 8004
rect 9916 7964 9922 7976
rect 10502 7964 10508 8016
rect 10560 8004 10566 8016
rect 12618 8004 12624 8016
rect 10560 7976 12624 8004
rect 10560 7964 10566 7976
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 13354 7964 13360 8016
rect 13412 8004 13418 8016
rect 14093 8007 14151 8013
rect 14093 8004 14105 8007
rect 13412 7976 14105 8004
rect 13412 7964 13418 7976
rect 14093 7973 14105 7976
rect 14139 7973 14151 8007
rect 22278 8004 22284 8016
rect 14093 7967 14151 7973
rect 21560 7976 22284 8004
rect 9309 7939 9367 7945
rect 9309 7905 9321 7939
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 9398 7896 9404 7948
rect 9456 7936 9462 7948
rect 12253 7939 12311 7945
rect 9456 7908 9904 7936
rect 9456 7896 9462 7908
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7868 5595 7871
rect 5718 7868 5724 7880
rect 5583 7840 5724 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7868 5871 7871
rect 5902 7868 5908 7880
rect 5859 7840 5908 7868
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6178 7868 6184 7880
rect 6139 7840 6184 7868
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 6362 7868 6368 7880
rect 6275 7840 6368 7868
rect 6362 7828 6368 7840
rect 6420 7868 6426 7880
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6420 7840 6837 7868
rect 6420 7828 6426 7840
rect 6825 7837 6837 7840
rect 6871 7837 6883 7871
rect 7466 7868 7472 7880
rect 7427 7840 7472 7868
rect 6825 7831 6883 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7800 7840 7849 7868
rect 7800 7828 7806 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8662 7868 8668 7880
rect 7975 7840 8524 7868
rect 8623 7840 8668 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 5994 7800 6000 7812
rect 4295 7772 5212 7800
rect 5955 7772 6000 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7701 2743 7735
rect 2685 7695 2743 7701
rect 3053 7735 3111 7741
rect 3053 7701 3065 7735
rect 3099 7732 3111 7735
rect 3234 7732 3240 7744
rect 3099 7704 3240 7732
rect 3099 7701 3111 7704
rect 3053 7695 3111 7701
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 4172 7732 4200 7763
rect 5994 7760 6000 7772
rect 6052 7760 6058 7812
rect 6730 7760 6736 7812
rect 6788 7800 6794 7812
rect 6917 7803 6975 7809
rect 6917 7800 6929 7803
rect 6788 7772 6929 7800
rect 6788 7760 6794 7772
rect 6917 7769 6929 7772
rect 6963 7769 6975 7803
rect 6917 7763 6975 7769
rect 5534 7732 5540 7744
rect 3927 7704 5540 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 5718 7732 5724 7744
rect 5679 7704 5724 7732
rect 5718 7692 5724 7704
rect 5776 7692 5782 7744
rect 5810 7692 5816 7744
rect 5868 7732 5874 7744
rect 8389 7735 8447 7741
rect 8389 7732 8401 7735
rect 5868 7704 8401 7732
rect 5868 7692 5874 7704
rect 8389 7701 8401 7704
rect 8435 7701 8447 7735
rect 8496 7732 8524 7840
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 8938 7868 8944 7880
rect 8803 7840 8944 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9217 7871 9275 7877
rect 9217 7868 9229 7871
rect 9088 7840 9229 7868
rect 9088 7828 9094 7840
rect 9217 7837 9229 7840
rect 9263 7868 9275 7871
rect 9582 7868 9588 7880
rect 9263 7840 9444 7868
rect 9543 7840 9588 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9416 7812 9444 7840
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 9876 7877 9904 7908
rect 12253 7905 12265 7939
rect 12299 7936 12311 7939
rect 12437 7939 12495 7945
rect 12299 7908 12333 7936
rect 12299 7905 12311 7908
rect 12253 7899 12311 7905
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 13170 7936 13176 7948
rect 12483 7908 13176 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7868 12127 7871
rect 12158 7868 12164 7880
rect 12115 7840 12164 7868
rect 12115 7837 12127 7840
rect 12069 7831 12127 7837
rect 12158 7828 12164 7840
rect 12216 7868 12222 7880
rect 12268 7868 12296 7899
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 14274 7896 14280 7948
rect 14332 7936 14338 7948
rect 14553 7939 14611 7945
rect 14553 7936 14565 7939
rect 14332 7908 14565 7936
rect 14332 7896 14338 7908
rect 14553 7905 14565 7908
rect 14599 7905 14611 7939
rect 14553 7899 14611 7905
rect 14642 7896 14648 7948
rect 14700 7936 14706 7948
rect 15565 7939 15623 7945
rect 14700 7908 14793 7936
rect 14700 7896 14706 7908
rect 15565 7905 15577 7939
rect 15611 7936 15623 7939
rect 16114 7936 16120 7948
rect 15611 7908 16120 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 16114 7896 16120 7908
rect 16172 7936 16178 7948
rect 16761 7939 16819 7945
rect 16761 7936 16773 7939
rect 16172 7908 16773 7936
rect 16172 7896 16178 7908
rect 16761 7905 16773 7908
rect 16807 7936 16819 7939
rect 18877 7939 18935 7945
rect 18877 7936 18889 7939
rect 16807 7908 18889 7936
rect 16807 7905 16819 7908
rect 16761 7899 16819 7905
rect 18877 7905 18889 7908
rect 18923 7936 18935 7939
rect 19705 7939 19763 7945
rect 19705 7936 19717 7939
rect 18923 7908 19717 7936
rect 18923 7905 18935 7908
rect 18877 7899 18935 7905
rect 19705 7905 19717 7908
rect 19751 7936 19763 7939
rect 20346 7936 20352 7948
rect 19751 7908 20352 7936
rect 19751 7905 19763 7908
rect 19705 7899 19763 7905
rect 20346 7896 20352 7908
rect 20404 7936 20410 7948
rect 21560 7945 21588 7976
rect 22278 7964 22284 7976
rect 22336 8004 22342 8016
rect 22336 7976 22784 8004
rect 22336 7964 22342 7976
rect 21269 7939 21327 7945
rect 21269 7936 21281 7939
rect 20404 7908 21281 7936
rect 20404 7896 20410 7908
rect 21269 7905 21281 7908
rect 21315 7936 21327 7939
rect 21545 7939 21603 7945
rect 21545 7936 21557 7939
rect 21315 7908 21557 7936
rect 21315 7905 21327 7908
rect 21269 7899 21327 7905
rect 21545 7905 21557 7908
rect 21591 7905 21603 7939
rect 21545 7899 21603 7905
rect 21634 7896 21640 7948
rect 21692 7936 21698 7948
rect 22756 7945 22784 7976
rect 22741 7939 22799 7945
rect 21692 7908 22692 7936
rect 21692 7896 21698 7908
rect 13817 7871 13875 7877
rect 13817 7868 13829 7871
rect 12216 7840 13829 7868
rect 12216 7828 12222 7840
rect 13817 7837 13829 7840
rect 13863 7837 13875 7871
rect 13817 7831 13875 7837
rect 9398 7760 9404 7812
rect 9456 7760 9462 7812
rect 9493 7803 9551 7809
rect 9493 7769 9505 7803
rect 9539 7800 9551 7803
rect 9674 7800 9680 7812
rect 9539 7772 9680 7800
rect 9539 7769 9551 7772
rect 9493 7763 9551 7769
rect 9674 7760 9680 7772
rect 9732 7760 9738 7812
rect 12250 7760 12256 7812
rect 12308 7800 12314 7812
rect 12529 7803 12587 7809
rect 12529 7800 12541 7803
rect 12308 7772 12541 7800
rect 12308 7760 12314 7772
rect 12529 7769 12541 7772
rect 12575 7769 12587 7803
rect 13832 7800 13860 7831
rect 14182 7828 14188 7880
rect 14240 7868 14246 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 14240 7840 14473 7868
rect 14240 7828 14246 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14660 7800 14688 7896
rect 15378 7828 15384 7880
rect 15436 7868 15442 7880
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 15436 7840 16037 7868
rect 15436 7828 15442 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 16850 7868 16856 7880
rect 16623 7840 16856 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 16850 7828 16856 7840
rect 16908 7828 16914 7880
rect 17218 7868 17224 7880
rect 17180 7840 17224 7868
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 17586 7868 17592 7880
rect 17547 7840 17592 7868
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7868 17739 7871
rect 18322 7868 18328 7880
rect 17727 7840 18328 7868
rect 17727 7837 17739 7840
rect 17681 7831 17739 7837
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7868 18475 7871
rect 18693 7871 18751 7877
rect 18693 7868 18705 7871
rect 18463 7840 18705 7868
rect 18463 7837 18475 7840
rect 18417 7831 18475 7837
rect 18693 7837 18705 7840
rect 18739 7837 18751 7871
rect 21726 7868 21732 7880
rect 21687 7840 21732 7868
rect 18693 7831 18751 7837
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 22462 7828 22468 7880
rect 22520 7868 22526 7880
rect 22557 7871 22615 7877
rect 22557 7868 22569 7871
rect 22520 7840 22569 7868
rect 22520 7828 22526 7840
rect 22557 7837 22569 7840
rect 22603 7837 22615 7871
rect 22664 7868 22692 7908
rect 22741 7905 22753 7939
rect 22787 7905 22799 7939
rect 22741 7899 22799 7905
rect 23017 7871 23075 7877
rect 23017 7868 23029 7871
rect 22664 7840 23029 7868
rect 22557 7831 22615 7837
rect 23017 7837 23029 7840
rect 23063 7837 23075 7871
rect 23017 7831 23075 7837
rect 13832 7772 14688 7800
rect 15289 7803 15347 7809
rect 12529 7763 12587 7769
rect 15289 7769 15301 7803
rect 15335 7800 15347 7803
rect 16482 7800 16488 7812
rect 15335 7772 16488 7800
rect 15335 7769 15347 7772
rect 15289 7763 15347 7769
rect 16482 7760 16488 7772
rect 16540 7760 16546 7812
rect 16669 7803 16727 7809
rect 16669 7769 16681 7803
rect 16715 7800 16727 7803
rect 17037 7803 17095 7809
rect 17037 7800 17049 7803
rect 16715 7772 17049 7800
rect 16715 7769 16727 7772
rect 16669 7763 16727 7769
rect 17037 7769 17049 7772
rect 17083 7769 17095 7803
rect 17037 7763 17095 7769
rect 17773 7803 17831 7809
rect 17773 7769 17785 7803
rect 17819 7769 17831 7803
rect 17773 7763 17831 7769
rect 18187 7803 18245 7809
rect 18187 7769 18199 7803
rect 18233 7800 18245 7803
rect 19426 7800 19432 7812
rect 18233 7772 19432 7800
rect 18233 7769 18245 7772
rect 18187 7763 18245 7769
rect 10045 7735 10103 7741
rect 10045 7732 10057 7735
rect 8496 7704 10057 7732
rect 8389 7695 8447 7701
rect 10045 7701 10057 7704
rect 10091 7732 10103 7735
rect 11698 7732 11704 7744
rect 10091 7704 11704 7732
rect 10091 7701 10103 7704
rect 10045 7695 10103 7701
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 12618 7692 12624 7744
rect 12676 7732 12682 7744
rect 12897 7735 12955 7741
rect 12897 7732 12909 7735
rect 12676 7704 12909 7732
rect 12676 7692 12682 7704
rect 12897 7701 12909 7704
rect 12943 7701 12955 7735
rect 14918 7732 14924 7744
rect 14879 7704 14924 7732
rect 12897 7695 12955 7701
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 15378 7692 15384 7744
rect 15436 7732 15442 7744
rect 15930 7732 15936 7744
rect 15436 7704 15481 7732
rect 15891 7704 15936 7732
rect 15436 7692 15442 7704
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 16206 7732 16212 7744
rect 16167 7704 16212 7732
rect 16206 7692 16212 7704
rect 16264 7692 16270 7744
rect 16390 7692 16396 7744
rect 16448 7732 16454 7744
rect 17788 7732 17816 7763
rect 19426 7760 19432 7772
rect 19484 7760 19490 7812
rect 21637 7803 21695 7809
rect 21637 7769 21649 7803
rect 21683 7800 21695 7803
rect 22278 7800 22284 7812
rect 21683 7772 22284 7800
rect 21683 7769 21695 7772
rect 21637 7763 21695 7769
rect 22278 7760 22284 7772
rect 22336 7760 22342 7812
rect 16448 7704 17816 7732
rect 16448 7692 16454 7704
rect 18414 7692 18420 7744
rect 18472 7732 18478 7744
rect 18509 7735 18567 7741
rect 18509 7732 18521 7735
rect 18472 7704 18521 7732
rect 18472 7692 18478 7704
rect 18509 7701 18521 7704
rect 18555 7701 18567 7735
rect 22094 7732 22100 7744
rect 22055 7704 22100 7732
rect 18509 7695 18567 7701
rect 22094 7692 22100 7704
rect 22152 7692 22158 7744
rect 22186 7692 22192 7744
rect 22244 7732 22250 7744
rect 22649 7735 22707 7741
rect 22244 7704 22289 7732
rect 22244 7692 22250 7704
rect 22649 7701 22661 7735
rect 22695 7732 22707 7735
rect 22922 7732 22928 7744
rect 22695 7704 22928 7732
rect 22695 7701 22707 7704
rect 22649 7695 22707 7701
rect 22922 7692 22928 7704
rect 22980 7692 22986 7744
rect 23198 7732 23204 7744
rect 23159 7704 23204 7732
rect 23198 7692 23204 7704
rect 23256 7692 23262 7744
rect 1104 7642 26220 7664
rect 1104 7590 9322 7642
rect 9374 7590 9386 7642
rect 9438 7590 9450 7642
rect 9502 7590 9514 7642
rect 9566 7590 9578 7642
rect 9630 7590 17694 7642
rect 17746 7590 17758 7642
rect 17810 7590 17822 7642
rect 17874 7590 17886 7642
rect 17938 7590 17950 7642
rect 18002 7590 26220 7642
rect 1104 7568 26220 7590
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4525 7531 4583 7537
rect 4525 7528 4537 7531
rect 4212 7500 4537 7528
rect 4212 7488 4218 7500
rect 4525 7497 4537 7500
rect 4571 7497 4583 7531
rect 4525 7491 4583 7497
rect 5718 7488 5724 7540
rect 5776 7528 5782 7540
rect 5776 7500 8340 7528
rect 5776 7488 5782 7500
rect 4985 7463 5043 7469
rect 3160 7432 3924 7460
rect 3160 7401 3188 7432
rect 3896 7404 3924 7432
rect 4985 7429 4997 7463
rect 5031 7460 5043 7463
rect 5736 7460 5764 7488
rect 5031 7432 5764 7460
rect 5031 7429 5043 7432
rect 4985 7423 5043 7429
rect 5902 7420 5908 7472
rect 5960 7460 5966 7472
rect 5997 7463 6055 7469
rect 5997 7460 6009 7463
rect 5960 7432 6009 7460
rect 5960 7420 5966 7432
rect 5997 7429 6009 7432
rect 6043 7429 6055 7463
rect 6362 7460 6368 7472
rect 6323 7432 6368 7460
rect 5997 7423 6055 7429
rect 6362 7420 6368 7432
rect 6420 7420 6426 7472
rect 7285 7463 7343 7469
rect 7285 7460 7297 7463
rect 6564 7432 7297 7460
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 3401 7395 3459 7401
rect 3401 7392 3413 7395
rect 3292 7364 3413 7392
rect 3292 7352 3298 7364
rect 3401 7361 3413 7364
rect 3447 7361 3459 7395
rect 3401 7355 3459 7361
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 6564 7401 6592 7432
rect 7285 7429 7297 7432
rect 7331 7429 7343 7463
rect 7285 7423 7343 7429
rect 7374 7420 7380 7472
rect 7432 7460 7438 7472
rect 7742 7460 7748 7472
rect 7432 7432 7604 7460
rect 7703 7432 7748 7460
rect 7432 7420 7438 7432
rect 4801 7395 4859 7401
rect 4801 7392 4813 7395
rect 3936 7364 4813 7392
rect 3936 7352 3942 7364
rect 4801 7361 4813 7364
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 7003 7395 7061 7401
rect 6779 7364 6960 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7293 6883 7327
rect 6932 7324 6960 7364
rect 7003 7361 7015 7395
rect 7049 7392 7061 7395
rect 7190 7392 7196 7404
rect 7049 7364 7196 7392
rect 7049 7361 7061 7364
rect 7003 7355 7061 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7466 7392 7472 7404
rect 7300 7364 7472 7392
rect 7300 7324 7328 7364
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 7576 7392 7604 7432
rect 7742 7420 7748 7432
rect 7800 7420 7806 7472
rect 8312 7469 8340 7500
rect 8386 7488 8392 7540
rect 8444 7528 8450 7540
rect 8444 7500 8984 7528
rect 8444 7488 8450 7500
rect 7929 7463 7987 7469
rect 7929 7429 7941 7463
rect 7975 7429 7987 7463
rect 7929 7423 7987 7429
rect 8297 7463 8355 7469
rect 8297 7429 8309 7463
rect 8343 7429 8355 7463
rect 8478 7460 8484 7472
rect 8439 7432 8484 7460
rect 8297 7423 8355 7429
rect 7944 7392 7972 7423
rect 8478 7420 8484 7432
rect 8536 7420 8542 7472
rect 8754 7392 8760 7404
rect 7576 7364 7972 7392
rect 8715 7364 8760 7392
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 8956 7392 8984 7500
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9309 7531 9367 7537
rect 9309 7528 9321 7531
rect 9272 7500 9321 7528
rect 9272 7488 9278 7500
rect 9309 7497 9321 7500
rect 9355 7497 9367 7531
rect 9309 7491 9367 7497
rect 11517 7531 11575 7537
rect 11517 7497 11529 7531
rect 11563 7528 11575 7531
rect 11882 7528 11888 7540
rect 11563 7500 11888 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 15102 7528 15108 7540
rect 12406 7500 15108 7528
rect 9033 7463 9091 7469
rect 9033 7429 9045 7463
rect 9079 7460 9091 7463
rect 12406 7460 12434 7500
rect 15102 7488 15108 7500
rect 15160 7488 15166 7540
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 15942 7531 16000 7537
rect 15942 7528 15954 7531
rect 15528 7500 15954 7528
rect 15528 7488 15534 7500
rect 15942 7497 15954 7500
rect 15988 7497 16000 7531
rect 15942 7491 16000 7497
rect 16485 7531 16543 7537
rect 16485 7497 16497 7531
rect 16531 7497 16543 7531
rect 18230 7528 18236 7540
rect 18191 7500 18236 7528
rect 16485 7491 16543 7497
rect 15010 7460 15016 7472
rect 9079 7432 9711 7460
rect 9079 7429 9091 7432
rect 9033 7423 9091 7429
rect 9683 7404 9711 7432
rect 10244 7432 12434 7460
rect 14016 7432 15016 7460
rect 9125 7395 9183 7401
rect 9125 7392 9137 7395
rect 8956 7364 9137 7392
rect 9048 7336 9076 7364
rect 9125 7361 9137 7364
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 9447 7364 9628 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 6932 7296 7328 7324
rect 7377 7327 7435 7333
rect 6825 7287 6883 7293
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 7742 7324 7748 7336
rect 7423 7296 7748 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 6840 7256 6868 7287
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 8018 7284 8024 7336
rect 8076 7324 8082 7336
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8076 7296 8585 7324
rect 8076 7284 8082 7296
rect 8573 7293 8585 7296
rect 8619 7324 8631 7327
rect 8662 7324 8668 7336
rect 8619 7296 8668 7324
rect 8619 7293 8631 7296
rect 8573 7287 8631 7293
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 9030 7284 9036 7336
rect 9088 7284 9094 7336
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 9493 7327 9551 7333
rect 9493 7324 9505 7327
rect 9272 7296 9505 7324
rect 9272 7284 9278 7296
rect 9493 7293 9505 7296
rect 9539 7293 9551 7327
rect 9600 7324 9628 7364
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10244 7401 10272 7432
rect 14016 7404 14044 7432
rect 15010 7420 15016 7432
rect 15068 7420 15074 7472
rect 16390 7460 16396 7472
rect 16132 7432 16396 7460
rect 10229 7395 10287 7401
rect 9732 7364 9825 7392
rect 9732 7352 9738 7364
rect 10229 7361 10241 7395
rect 10275 7361 10287 7395
rect 10410 7392 10416 7404
rect 10371 7364 10416 7392
rect 10229 7355 10287 7361
rect 10244 7324 10272 7355
rect 10410 7352 10416 7364
rect 10468 7392 10474 7404
rect 10689 7395 10747 7401
rect 10689 7392 10701 7395
rect 10468 7364 10701 7392
rect 10468 7352 10474 7364
rect 10689 7361 10701 7364
rect 10735 7361 10747 7395
rect 10870 7392 10876 7404
rect 10831 7364 10876 7392
rect 10689 7355 10747 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 11146 7392 11152 7404
rect 11107 7364 11152 7392
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11747 7364 11989 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 9600 7296 10272 7324
rect 10505 7327 10563 7333
rect 9493 7287 9551 7293
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 11716 7324 11744 7355
rect 10551 7296 11744 7324
rect 11992 7324 12020 7355
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 13725 7395 13783 7401
rect 12124 7364 12169 7392
rect 12124 7352 12130 7364
rect 13725 7361 13737 7395
rect 13771 7392 13783 7395
rect 13906 7392 13912 7404
rect 13771 7364 13912 7392
rect 13771 7361 13783 7364
rect 13725 7355 13783 7361
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 13998 7352 14004 7404
rect 14056 7392 14062 7404
rect 14274 7401 14280 7404
rect 14268 7392 14280 7401
rect 14056 7364 14149 7392
rect 14235 7364 14280 7392
rect 14056 7352 14062 7364
rect 14268 7355 14280 7364
rect 14274 7352 14280 7355
rect 14332 7352 14338 7404
rect 14826 7352 14832 7404
rect 14884 7392 14890 7404
rect 15565 7395 15623 7401
rect 15565 7392 15577 7395
rect 14884 7364 15577 7392
rect 14884 7352 14890 7364
rect 15565 7361 15577 7364
rect 15611 7392 15623 7395
rect 16132 7392 16160 7432
rect 16390 7420 16396 7432
rect 16448 7420 16454 7472
rect 16500 7460 16528 7491
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 18601 7531 18659 7537
rect 18601 7497 18613 7531
rect 18647 7528 18659 7531
rect 19242 7528 19248 7540
rect 18647 7500 19248 7528
rect 18647 7497 18659 7500
rect 18601 7491 18659 7497
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 19426 7488 19432 7540
rect 19484 7537 19490 7540
rect 19484 7528 19496 7537
rect 20165 7531 20223 7537
rect 19484 7500 20116 7528
rect 19484 7491 19496 7500
rect 19484 7488 19490 7491
rect 16914 7463 16972 7469
rect 16914 7460 16926 7463
rect 16500 7432 16926 7460
rect 16914 7429 16926 7432
rect 16960 7429 16972 7463
rect 20088 7460 20116 7500
rect 20165 7497 20177 7531
rect 20211 7528 20223 7531
rect 20438 7528 20444 7540
rect 20211 7500 20444 7528
rect 20211 7497 20223 7500
rect 20165 7491 20223 7497
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 20990 7488 20996 7540
rect 21048 7528 21054 7540
rect 21818 7528 21824 7540
rect 21048 7500 21824 7528
rect 21048 7488 21054 7500
rect 21818 7488 21824 7500
rect 21876 7488 21882 7540
rect 23198 7469 23204 7472
rect 21370 7463 21428 7469
rect 21370 7460 21382 7463
rect 20088 7432 21382 7460
rect 16914 7423 16972 7429
rect 21370 7429 21382 7432
rect 21416 7460 21428 7463
rect 22198 7463 22256 7469
rect 22198 7460 22210 7463
rect 21416 7432 22210 7460
rect 21416 7429 21428 7432
rect 21370 7423 21428 7429
rect 22198 7429 22210 7432
rect 22244 7429 22256 7463
rect 23192 7460 23204 7469
rect 23159 7432 23204 7460
rect 22198 7423 22256 7429
rect 23192 7423 23204 7432
rect 23198 7420 23204 7423
rect 23256 7420 23262 7472
rect 15611 7364 16160 7392
rect 16209 7395 16267 7401
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 16301 7395 16359 7401
rect 16301 7392 16313 7395
rect 16255 7364 16313 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 16301 7361 16313 7364
rect 16347 7361 16359 7395
rect 16408 7392 16436 7420
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 16408 7364 19073 7392
rect 16301 7355 16359 7361
rect 19061 7361 19073 7364
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20714 7392 20720 7404
rect 20303 7364 20720 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20714 7352 20720 7364
rect 20772 7352 20778 7404
rect 20990 7392 20996 7404
rect 20951 7364 20996 7392
rect 20990 7352 20996 7364
rect 21048 7352 21054 7404
rect 21634 7392 21640 7404
rect 21595 7364 21640 7392
rect 21634 7352 21640 7364
rect 21692 7352 21698 7404
rect 21818 7392 21824 7404
rect 21779 7364 21824 7392
rect 21818 7352 21824 7364
rect 21876 7352 21882 7404
rect 22465 7395 22523 7401
rect 22465 7361 22477 7395
rect 22511 7392 22523 7395
rect 22557 7395 22615 7401
rect 22557 7392 22569 7395
rect 22511 7364 22569 7392
rect 22511 7361 22523 7364
rect 22465 7355 22523 7361
rect 22557 7361 22569 7364
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 22925 7395 22983 7401
rect 22925 7361 22937 7395
rect 22971 7392 22983 7395
rect 23014 7392 23020 7404
rect 22971 7364 23020 7392
rect 22971 7361 22983 7364
rect 22925 7355 22983 7361
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 12250 7324 12256 7336
rect 11992 7296 12256 7324
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 16669 7327 16727 7333
rect 16669 7324 16681 7327
rect 15068 7296 16681 7324
rect 15068 7284 15074 7296
rect 16669 7293 16681 7296
rect 16715 7293 16727 7327
rect 16669 7287 16727 7293
rect 18506 7284 18512 7336
rect 18564 7324 18570 7336
rect 18693 7327 18751 7333
rect 18693 7324 18705 7327
rect 18564 7296 18705 7324
rect 18564 7284 18570 7296
rect 18693 7293 18705 7296
rect 18739 7293 18751 7327
rect 18693 7287 18751 7293
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 20346 7324 20352 7336
rect 18932 7296 20352 7324
rect 18932 7284 18938 7296
rect 20346 7284 20352 7296
rect 20404 7284 20410 7336
rect 22186 7324 22192 7336
rect 21376 7296 22192 7324
rect 8110 7256 8116 7268
rect 6840 7228 6960 7256
rect 8023 7228 8116 7256
rect 6932 7188 6960 7228
rect 8110 7216 8116 7228
rect 8168 7256 8174 7268
rect 9766 7256 9772 7268
rect 8168 7228 9772 7256
rect 8168 7216 8174 7228
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 9861 7259 9919 7265
rect 9861 7225 9873 7259
rect 9907 7256 9919 7259
rect 11238 7256 11244 7268
rect 9907 7228 11244 7256
rect 9907 7225 9919 7228
rect 9861 7219 9919 7225
rect 11238 7216 11244 7228
rect 11296 7216 11302 7268
rect 11606 7216 11612 7268
rect 11664 7256 11670 7268
rect 19797 7259 19855 7265
rect 19797 7256 19809 7259
rect 11664 7228 12296 7256
rect 11664 7216 11670 7228
rect 7006 7188 7012 7200
rect 6919 7160 7012 7188
rect 7006 7148 7012 7160
rect 7064 7188 7070 7200
rect 7745 7191 7803 7197
rect 7745 7188 7757 7191
rect 7064 7160 7757 7188
rect 7064 7148 7070 7160
rect 7745 7157 7757 7160
rect 7791 7157 7803 7191
rect 7745 7151 7803 7157
rect 8938 7148 8944 7200
rect 8996 7188 9002 7200
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 8996 7160 10057 7188
rect 8996 7148 9002 7160
rect 10045 7157 10057 7160
rect 10091 7157 10103 7191
rect 11054 7188 11060 7200
rect 11015 7160 11060 7188
rect 10045 7151 10103 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11330 7188 11336 7200
rect 11291 7160 11336 7188
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11790 7188 11796 7200
rect 11751 7160 11796 7188
rect 11790 7148 11796 7160
rect 11848 7188 11854 7200
rect 12066 7188 12072 7200
rect 11848 7160 12072 7188
rect 11848 7148 11854 7160
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 12268 7197 12296 7228
rect 19444 7228 19809 7256
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7157 12311 7191
rect 12253 7151 12311 7157
rect 13909 7191 13967 7197
rect 13909 7157 13921 7191
rect 13955 7188 13967 7191
rect 14274 7188 14280 7200
rect 13955 7160 14280 7188
rect 13955 7157 13967 7160
rect 13909 7151 13967 7157
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 15381 7191 15439 7197
rect 15381 7188 15393 7191
rect 15344 7160 15393 7188
rect 15344 7148 15350 7160
rect 15381 7157 15393 7160
rect 15427 7157 15439 7191
rect 15381 7151 15439 7157
rect 15933 7191 15991 7197
rect 15933 7157 15945 7191
rect 15979 7188 15991 7191
rect 16206 7188 16212 7200
rect 15979 7160 16212 7188
rect 15979 7157 15991 7160
rect 15933 7151 15991 7157
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 17034 7148 17040 7200
rect 17092 7188 17098 7200
rect 17586 7188 17592 7200
rect 17092 7160 17592 7188
rect 17092 7148 17098 7160
rect 17586 7148 17592 7160
rect 17644 7188 17650 7200
rect 19444 7197 19472 7228
rect 19797 7225 19809 7228
rect 19843 7225 19855 7259
rect 19797 7219 19855 7225
rect 18049 7191 18107 7197
rect 18049 7188 18061 7191
rect 17644 7160 18061 7188
rect 17644 7148 17650 7160
rect 18049 7157 18061 7160
rect 18095 7157 18107 7191
rect 18049 7151 18107 7157
rect 19429 7191 19487 7197
rect 19429 7157 19441 7191
rect 19475 7157 19487 7191
rect 19429 7151 19487 7157
rect 19518 7148 19524 7200
rect 19576 7188 19582 7200
rect 21376 7197 21404 7296
rect 22186 7284 22192 7296
rect 22244 7284 22250 7336
rect 22094 7216 22100 7268
rect 22152 7216 22158 7268
rect 19613 7191 19671 7197
rect 19613 7188 19625 7191
rect 19576 7160 19625 7188
rect 19576 7148 19582 7160
rect 19613 7157 19625 7160
rect 19659 7157 19671 7191
rect 19613 7151 19671 7157
rect 21361 7191 21419 7197
rect 21361 7157 21373 7191
rect 21407 7157 21419 7191
rect 22112 7188 22140 7216
rect 22189 7191 22247 7197
rect 22189 7188 22201 7191
rect 22112 7160 22201 7188
rect 21361 7151 21419 7157
rect 22189 7157 22201 7160
rect 22235 7157 22247 7191
rect 22738 7188 22744 7200
rect 22699 7160 22744 7188
rect 22189 7151 22247 7157
rect 22738 7148 22744 7160
rect 22796 7148 22802 7200
rect 23842 7148 23848 7200
rect 23900 7188 23906 7200
rect 24305 7191 24363 7197
rect 24305 7188 24317 7191
rect 23900 7160 24317 7188
rect 23900 7148 23906 7160
rect 24305 7157 24317 7160
rect 24351 7157 24363 7191
rect 24305 7151 24363 7157
rect 1104 7098 26220 7120
rect 1104 7046 5136 7098
rect 5188 7046 5200 7098
rect 5252 7046 5264 7098
rect 5316 7046 5328 7098
rect 5380 7046 5392 7098
rect 5444 7046 13508 7098
rect 13560 7046 13572 7098
rect 13624 7046 13636 7098
rect 13688 7046 13700 7098
rect 13752 7046 13764 7098
rect 13816 7046 21880 7098
rect 21932 7046 21944 7098
rect 21996 7046 22008 7098
rect 22060 7046 22072 7098
rect 22124 7046 22136 7098
rect 22188 7046 26220 7098
rect 1104 7024 26220 7046
rect 6730 6984 6736 6996
rect 6691 6956 6736 6984
rect 6730 6944 6736 6956
rect 6788 6944 6794 6996
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 8113 6987 8171 6993
rect 8113 6984 8125 6987
rect 7800 6956 8125 6984
rect 7800 6944 7806 6956
rect 8113 6953 8125 6956
rect 8159 6953 8171 6987
rect 8113 6947 8171 6953
rect 10321 6987 10379 6993
rect 10321 6953 10333 6987
rect 10367 6984 10379 6987
rect 11514 6984 11520 6996
rect 10367 6956 11520 6984
rect 10367 6953 10379 6956
rect 10321 6947 10379 6953
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 12437 6987 12495 6993
rect 12437 6953 12449 6987
rect 12483 6984 12495 6987
rect 12894 6984 12900 6996
rect 12483 6956 12900 6984
rect 12483 6953 12495 6956
rect 12437 6947 12495 6953
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 13906 6944 13912 6996
rect 13964 6984 13970 6996
rect 14185 6987 14243 6993
rect 14185 6984 14197 6987
rect 13964 6956 14197 6984
rect 13964 6944 13970 6956
rect 14185 6953 14197 6956
rect 14231 6953 14243 6987
rect 14185 6947 14243 6953
rect 14369 6987 14427 6993
rect 14369 6953 14381 6987
rect 14415 6984 14427 6987
rect 14918 6984 14924 6996
rect 14415 6956 14924 6984
rect 14415 6953 14427 6956
rect 14369 6947 14427 6953
rect 14918 6944 14924 6956
rect 14976 6944 14982 6996
rect 15102 6944 15108 6996
rect 15160 6984 15166 6996
rect 15565 6987 15623 6993
rect 15565 6984 15577 6987
rect 15160 6956 15577 6984
rect 15160 6944 15166 6956
rect 15565 6953 15577 6956
rect 15611 6953 15623 6987
rect 15565 6947 15623 6953
rect 17129 6987 17187 6993
rect 17129 6953 17141 6987
rect 17175 6984 17187 6987
rect 17310 6984 17316 6996
rect 17175 6956 17316 6984
rect 17175 6953 17187 6956
rect 17129 6947 17187 6953
rect 17310 6944 17316 6956
rect 17368 6944 17374 6996
rect 19426 6984 19432 6996
rect 19387 6956 19432 6984
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 22922 6944 22928 6996
rect 22980 6984 22986 6996
rect 23293 6987 23351 6993
rect 23293 6984 23305 6987
rect 22980 6956 23305 6984
rect 22980 6944 22986 6956
rect 23293 6953 23305 6956
rect 23339 6953 23351 6987
rect 23293 6947 23351 6953
rect 7834 6876 7840 6928
rect 7892 6916 7898 6928
rect 9125 6919 9183 6925
rect 9125 6916 9137 6919
rect 7892 6888 9137 6916
rect 7892 6876 7898 6888
rect 9125 6885 9137 6888
rect 9171 6885 9183 6919
rect 9125 6879 9183 6885
rect 14642 6876 14648 6928
rect 14700 6916 14706 6928
rect 15470 6916 15476 6928
rect 14700 6888 15476 6916
rect 14700 6876 14706 6888
rect 15470 6876 15476 6888
rect 15528 6876 15534 6928
rect 16758 6916 16764 6928
rect 16671 6888 16764 6916
rect 16758 6876 16764 6888
rect 16816 6916 16822 6928
rect 17218 6916 17224 6928
rect 16816 6888 17224 6916
rect 16816 6876 16822 6888
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 8110 6848 8116 6860
rect 6880 6820 8116 6848
rect 6880 6808 6886 6820
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 13998 6848 14004 6860
rect 12207 6820 14004 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 14921 6851 14979 6857
rect 14921 6817 14933 6851
rect 14967 6848 14979 6851
rect 15378 6848 15384 6860
rect 14967 6820 15384 6848
rect 14967 6817 14979 6820
rect 14921 6811 14979 6817
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 15988 6820 17356 6848
rect 15988 6808 15994 6820
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6549 6783 6607 6789
rect 6549 6780 6561 6783
rect 6052 6752 6561 6780
rect 6052 6740 6058 6752
rect 6549 6749 6561 6752
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 7285 6783 7343 6789
rect 7285 6749 7297 6783
rect 7331 6780 7343 6783
rect 7466 6780 7472 6792
rect 7331 6752 7472 6780
rect 7331 6749 7343 6752
rect 7285 6743 7343 6749
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 8481 6783 8539 6789
rect 8251 6752 8340 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 8312 6724 8340 6752
rect 8481 6749 8493 6783
rect 8527 6780 8539 6783
rect 8846 6780 8852 6792
rect 8527 6752 8852 6780
rect 8527 6749 8539 6752
rect 8481 6743 8539 6749
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 8938 6740 8944 6792
rect 8996 6780 9002 6792
rect 10597 6783 10655 6789
rect 8996 6752 9041 6780
rect 8996 6740 9002 6752
rect 10597 6749 10609 6783
rect 10643 6780 10655 6783
rect 11146 6780 11152 6792
rect 10643 6752 11152 6780
rect 10643 6749 10655 6752
rect 10597 6743 10655 6749
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11894 6783 11952 6789
rect 11894 6780 11906 6783
rect 11388 6752 11906 6780
rect 11388 6740 11394 6752
rect 11894 6749 11906 6752
rect 11940 6749 11952 6783
rect 12250 6780 12256 6792
rect 12211 6752 12256 6780
rect 11894 6743 11952 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 12526 6780 12532 6792
rect 12487 6752 12532 6780
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 13078 6780 13084 6792
rect 12943 6752 13084 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7248 6684 7696 6712
rect 7248 6672 7254 6684
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7101 6647 7159 6653
rect 7101 6644 7113 6647
rect 6972 6616 7113 6644
rect 6972 6604 6978 6616
rect 7101 6613 7113 6616
rect 7147 6644 7159 6647
rect 7558 6644 7564 6656
rect 7147 6616 7564 6644
rect 7147 6613 7159 6616
rect 7101 6607 7159 6613
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 7668 6644 7696 6684
rect 8294 6672 8300 6724
rect 8352 6672 8358 6724
rect 9953 6715 10011 6721
rect 9953 6681 9965 6715
rect 9999 6712 10011 6715
rect 10042 6712 10048 6724
rect 9999 6684 10048 6712
rect 9999 6681 10011 6684
rect 9953 6675 10011 6681
rect 10042 6672 10048 6684
rect 10100 6672 10106 6724
rect 10367 6715 10425 6721
rect 10367 6681 10379 6715
rect 10413 6712 10425 6715
rect 11790 6712 11796 6724
rect 10413 6684 11796 6712
rect 10413 6681 10425 6684
rect 10367 6675 10425 6681
rect 11790 6672 11796 6684
rect 11848 6672 11854 6724
rect 12820 6712 12848 6743
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 13262 6740 13268 6792
rect 13320 6780 13326 6792
rect 15105 6783 15163 6789
rect 15105 6780 15117 6783
rect 13320 6752 15117 6780
rect 13320 6740 13326 6752
rect 15105 6749 15117 6752
rect 15151 6749 15163 6783
rect 15286 6780 15292 6792
rect 15247 6752 15292 6780
rect 15105 6743 15163 6749
rect 15286 6740 15292 6752
rect 15344 6780 15350 6792
rect 15657 6783 15715 6789
rect 15657 6780 15669 6783
rect 15344 6752 15669 6780
rect 15344 6740 15350 6752
rect 15657 6749 15669 6752
rect 15703 6749 15715 6783
rect 15657 6743 15715 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6780 15899 6783
rect 16758 6780 16764 6792
rect 15887 6752 16764 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 12406 6684 12848 6712
rect 14360 6715 14418 6721
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 7668 6616 8401 6644
rect 8389 6613 8401 6616
rect 8435 6613 8447 6647
rect 8389 6607 8447 6613
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 10502 6644 10508 6656
rect 8812 6616 10508 6644
rect 8812 6604 8818 6616
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 10781 6647 10839 6653
rect 10781 6613 10793 6647
rect 10827 6644 10839 6647
rect 10962 6644 10968 6656
rect 10827 6616 10968 6644
rect 10827 6613 10839 6616
rect 10781 6607 10839 6613
rect 10962 6604 10968 6616
rect 11020 6644 11026 6656
rect 12406 6644 12434 6684
rect 14360 6681 14372 6715
rect 14406 6712 14418 6715
rect 14642 6712 14648 6724
rect 14406 6684 14648 6712
rect 14406 6681 14418 6684
rect 14360 6675 14418 6681
rect 14642 6672 14648 6684
rect 14700 6672 14706 6724
rect 14737 6715 14795 6721
rect 14737 6681 14749 6715
rect 14783 6712 14795 6715
rect 14826 6712 14832 6724
rect 14783 6684 14832 6712
rect 14783 6681 14795 6684
rect 14737 6675 14795 6681
rect 11020 6616 12434 6644
rect 12713 6647 12771 6653
rect 11020 6604 11026 6616
rect 12713 6613 12725 6647
rect 12759 6644 12771 6647
rect 14752 6644 14780 6675
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 15381 6715 15439 6721
rect 15381 6681 15393 6715
rect 15427 6712 15439 6715
rect 15856 6712 15884 6743
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 17034 6780 17040 6792
rect 16995 6752 17040 6780
rect 17034 6740 17040 6752
rect 17092 6740 17098 6792
rect 17126 6740 17132 6792
rect 17184 6780 17190 6792
rect 17328 6780 17356 6820
rect 18693 6783 18751 6789
rect 17184 6752 17229 6780
rect 17328 6752 18552 6780
rect 17184 6740 17190 6752
rect 18414 6712 18420 6724
rect 18472 6721 18478 6724
rect 15427 6684 15884 6712
rect 18384 6684 18420 6712
rect 15427 6681 15439 6684
rect 15381 6675 15439 6681
rect 18414 6672 18420 6684
rect 18472 6675 18484 6721
rect 18524 6712 18552 6752
rect 18693 6749 18705 6783
rect 18739 6780 18751 6783
rect 19242 6780 19248 6792
rect 18739 6752 19104 6780
rect 19203 6752 19248 6780
rect 18739 6749 18751 6752
rect 18693 6743 18751 6749
rect 19076 6721 19104 6752
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 19521 6783 19579 6789
rect 19521 6749 19533 6783
rect 19567 6780 19579 6783
rect 23014 6780 23020 6792
rect 19567 6752 23020 6780
rect 19567 6749 19579 6752
rect 19521 6743 19579 6749
rect 18877 6715 18935 6721
rect 18877 6712 18889 6715
rect 18524 6684 18889 6712
rect 18877 6681 18889 6684
rect 18923 6681 18935 6715
rect 18877 6675 18935 6681
rect 19061 6715 19119 6721
rect 19061 6681 19073 6715
rect 19107 6712 19119 6715
rect 19334 6712 19340 6724
rect 19107 6684 19340 6712
rect 19107 6681 19119 6684
rect 19061 6675 19119 6681
rect 18472 6672 18478 6675
rect 19334 6672 19340 6684
rect 19392 6712 19398 6724
rect 19536 6712 19564 6743
rect 23014 6740 23020 6752
rect 23072 6780 23078 6792
rect 23474 6789 23480 6792
rect 23109 6783 23167 6789
rect 23109 6780 23121 6783
rect 23072 6752 23121 6780
rect 23072 6740 23078 6752
rect 23109 6749 23121 6752
rect 23155 6749 23167 6783
rect 23109 6743 23167 6749
rect 23443 6783 23480 6789
rect 23443 6749 23455 6783
rect 23443 6743 23480 6749
rect 23474 6740 23480 6743
rect 23532 6740 23538 6792
rect 23750 6780 23756 6792
rect 23711 6752 23756 6780
rect 23750 6740 23756 6752
rect 23808 6740 23814 6792
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6749 23903 6783
rect 23845 6743 23903 6749
rect 19392 6684 19564 6712
rect 19392 6672 19398 6684
rect 19610 6672 19616 6724
rect 19668 6712 19674 6724
rect 19766 6715 19824 6721
rect 19766 6712 19778 6715
rect 19668 6684 19778 6712
rect 19668 6672 19674 6684
rect 19766 6681 19778 6684
rect 19812 6681 19824 6715
rect 19766 6675 19824 6681
rect 22738 6672 22744 6724
rect 22796 6712 22802 6724
rect 22842 6715 22900 6721
rect 22842 6712 22854 6715
rect 22796 6684 22854 6712
rect 22796 6672 22802 6684
rect 22842 6681 22854 6684
rect 22888 6681 22900 6715
rect 23860 6712 23888 6743
rect 22842 6675 22900 6681
rect 23400 6684 23888 6712
rect 23400 6656 23428 6684
rect 17310 6644 17316 6656
rect 12759 6616 14780 6644
rect 17271 6616 17316 6644
rect 12759 6613 12771 6616
rect 12713 6607 12771 6613
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 20901 6647 20959 6653
rect 20901 6613 20913 6647
rect 20947 6644 20959 6647
rect 21174 6644 21180 6656
rect 20947 6616 21180 6644
rect 20947 6613 20959 6616
rect 20901 6607 20959 6613
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 21726 6644 21732 6656
rect 21687 6616 21732 6644
rect 21726 6604 21732 6616
rect 21784 6604 21790 6656
rect 23382 6604 23388 6656
rect 23440 6604 23446 6656
rect 1104 6554 26220 6576
rect 1104 6502 9322 6554
rect 9374 6502 9386 6554
rect 9438 6502 9450 6554
rect 9502 6502 9514 6554
rect 9566 6502 9578 6554
rect 9630 6502 17694 6554
rect 17746 6502 17758 6554
rect 17810 6502 17822 6554
rect 17874 6502 17886 6554
rect 17938 6502 17950 6554
rect 18002 6502 26220 6554
rect 1104 6480 26220 6502
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5684 6412 6009 6440
rect 5684 6400 5690 6412
rect 5997 6409 6009 6412
rect 6043 6440 6055 6443
rect 6822 6440 6828 6452
rect 6043 6412 6828 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 7006 6440 7012 6452
rect 6967 6412 7012 6440
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 7469 6443 7527 6449
rect 7469 6409 7481 6443
rect 7515 6440 7527 6443
rect 8018 6440 8024 6452
rect 7515 6412 8024 6440
rect 7515 6409 7527 6412
rect 7469 6403 7527 6409
rect 8018 6400 8024 6412
rect 8076 6440 8082 6452
rect 9122 6440 9128 6452
rect 8076 6412 9128 6440
rect 8076 6400 8082 6412
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 10870 6400 10876 6452
rect 10928 6440 10934 6452
rect 10965 6443 11023 6449
rect 10965 6440 10977 6443
rect 10928 6412 10977 6440
rect 10928 6400 10934 6412
rect 10965 6409 10977 6412
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 11885 6443 11943 6449
rect 11885 6440 11897 6443
rect 11112 6412 11897 6440
rect 11112 6400 11118 6412
rect 11885 6409 11897 6412
rect 11931 6409 11943 6443
rect 11885 6403 11943 6409
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6440 12035 6443
rect 13078 6440 13084 6452
rect 12023 6412 13084 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 14737 6443 14795 6449
rect 14737 6409 14749 6443
rect 14783 6440 14795 6443
rect 15010 6440 15016 6452
rect 14783 6412 15016 6440
rect 14783 6409 14795 6412
rect 14737 6403 14795 6409
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 19429 6443 19487 6449
rect 17236 6412 18644 6440
rect 6178 6332 6184 6384
rect 6236 6372 6242 6384
rect 6549 6375 6607 6381
rect 6549 6372 6561 6375
rect 6236 6344 6561 6372
rect 6236 6332 6242 6344
rect 6549 6341 6561 6344
rect 6595 6341 6607 6375
rect 7926 6372 7932 6384
rect 6549 6335 6607 6341
rect 7300 6344 7932 6372
rect 6730 6304 6736 6316
rect 6691 6276 6736 6304
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 7300 6313 7328 6344
rect 7926 6332 7932 6344
rect 7984 6332 7990 6384
rect 8202 6372 8208 6384
rect 8163 6344 8208 6372
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 8938 6332 8944 6384
rect 8996 6372 9002 6384
rect 9214 6372 9220 6384
rect 8996 6344 9220 6372
rect 8996 6332 9002 6344
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 10134 6332 10140 6384
rect 10192 6372 10198 6384
rect 14829 6375 14887 6381
rect 10192 6344 12434 6372
rect 10192 6332 10198 6344
rect 7009 6307 7067 6313
rect 7009 6304 7021 6307
rect 6880 6276 7021 6304
rect 6880 6264 6886 6276
rect 7009 6273 7021 6276
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6304 7435 6307
rect 7466 6304 7472 6316
rect 7423 6276 7472 6304
rect 7423 6273 7435 6276
rect 7377 6267 7435 6273
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 7616 6276 7757 6304
rect 7616 6264 7622 6276
rect 7745 6273 7757 6276
rect 7791 6304 7803 6307
rect 8110 6304 8116 6316
rect 7791 6276 8116 6304
rect 7791 6273 7803 6276
rect 7745 6267 7803 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 10502 6264 10508 6316
rect 10560 6304 10566 6316
rect 10597 6307 10655 6313
rect 10597 6304 10609 6307
rect 10560 6276 10609 6304
rect 10560 6264 10566 6276
rect 10597 6273 10609 6276
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10744 6276 10793 6304
rect 10744 6264 10750 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 11238 6304 11244 6316
rect 11195 6276 11244 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 12406 6304 12434 6344
rect 14829 6341 14841 6375
rect 14875 6372 14887 6375
rect 15930 6372 15936 6384
rect 14875 6344 15936 6372
rect 14875 6341 14887 6344
rect 14829 6335 14887 6341
rect 15930 6332 15936 6344
rect 15988 6332 15994 6384
rect 17236 6304 17264 6412
rect 18506 6372 18512 6384
rect 18467 6344 18512 6372
rect 18506 6332 18512 6344
rect 18564 6332 18570 6384
rect 18616 6372 18644 6412
rect 19429 6409 19441 6443
rect 19475 6440 19487 6443
rect 19610 6440 19616 6452
rect 19475 6412 19616 6440
rect 19475 6409 19487 6412
rect 19429 6403 19487 6409
rect 19610 6400 19616 6412
rect 19668 6400 19674 6452
rect 20714 6440 20720 6452
rect 20675 6412 20720 6440
rect 20714 6400 20720 6412
rect 20772 6400 20778 6452
rect 21726 6400 21732 6452
rect 21784 6440 21790 6452
rect 21784 6412 22232 6440
rect 21784 6400 21790 6412
rect 22094 6372 22100 6384
rect 18616 6344 22100 6372
rect 22094 6332 22100 6344
rect 22152 6332 22158 6384
rect 22204 6372 22232 6412
rect 23474 6372 23480 6384
rect 22204 6344 22784 6372
rect 12406 6276 17264 6304
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 18322 6304 18328 6316
rect 17368 6276 18000 6304
rect 18283 6276 18328 6304
rect 17368 6264 17374 6276
rect 6365 6239 6423 6245
rect 6365 6205 6377 6239
rect 6411 6236 6423 6239
rect 9214 6236 9220 6248
rect 6411 6208 9220 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 12161 6239 12219 6245
rect 10704 6208 11652 6236
rect 5810 6128 5816 6180
rect 5868 6168 5874 6180
rect 6181 6171 6239 6177
rect 6181 6168 6193 6171
rect 5868 6140 6193 6168
rect 5868 6128 5874 6140
rect 6181 6137 6193 6140
rect 6227 6168 6239 6171
rect 8754 6168 8760 6180
rect 6227 6140 8760 6168
rect 6227 6137 6239 6140
rect 6181 6131 6239 6137
rect 8754 6128 8760 6140
rect 8812 6168 8818 6180
rect 10704 6168 10732 6208
rect 11514 6168 11520 6180
rect 8812 6140 10732 6168
rect 11475 6140 11520 6168
rect 8812 6128 8818 6140
rect 11514 6128 11520 6140
rect 11572 6128 11578 6180
rect 11624 6168 11652 6208
rect 12161 6205 12173 6239
rect 12207 6236 12219 6239
rect 12342 6236 12348 6248
rect 12207 6208 12348 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 17126 6196 17132 6248
rect 17184 6236 17190 6248
rect 17972 6245 18000 6276
rect 18322 6264 18328 6276
rect 18380 6304 18386 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 18380 6276 18613 6304
rect 18380 6264 18386 6276
rect 18601 6273 18613 6276
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 18969 6307 19027 6313
rect 18969 6273 18981 6307
rect 19015 6273 19027 6307
rect 18969 6267 19027 6273
rect 19245 6307 19303 6313
rect 19245 6273 19257 6307
rect 19291 6304 19303 6307
rect 19518 6304 19524 6316
rect 19291 6276 19524 6304
rect 19291 6273 19303 6276
rect 19245 6267 19303 6273
rect 17865 6239 17923 6245
rect 17865 6236 17877 6239
rect 17184 6208 17877 6236
rect 17184 6196 17190 6208
rect 17865 6205 17877 6208
rect 17911 6205 17923 6239
rect 17865 6199 17923 6205
rect 17957 6239 18015 6245
rect 17957 6205 17969 6239
rect 18003 6236 18015 6239
rect 18800 6236 18828 6267
rect 18003 6208 18828 6236
rect 18984 6236 19012 6267
rect 19518 6264 19524 6276
rect 19576 6264 19582 6316
rect 19610 6264 19616 6316
rect 19668 6304 19674 6316
rect 20898 6313 20904 6316
rect 19981 6307 20039 6313
rect 19981 6304 19993 6307
rect 19668 6276 19993 6304
rect 19668 6264 19674 6276
rect 19981 6273 19993 6276
rect 20027 6273 20039 6307
rect 20867 6307 20904 6313
rect 20867 6304 20879 6307
rect 19981 6267 20039 6273
rect 20088 6276 20879 6304
rect 20088 6236 20116 6276
rect 20867 6273 20879 6276
rect 20867 6267 20904 6273
rect 20898 6264 20904 6267
rect 20956 6264 20962 6316
rect 22756 6313 22784 6344
rect 22848 6344 23480 6372
rect 22848 6313 22876 6344
rect 23474 6332 23480 6344
rect 23532 6332 23538 6384
rect 23845 6375 23903 6381
rect 23845 6372 23857 6375
rect 23584 6344 23857 6372
rect 21269 6307 21327 6313
rect 21269 6273 21281 6307
rect 21315 6304 21327 6307
rect 22374 6307 22432 6313
rect 22374 6304 22386 6307
rect 21315 6276 22386 6304
rect 21315 6273 21327 6276
rect 21269 6267 21327 6273
rect 22374 6273 22386 6276
rect 22420 6304 22432 6307
rect 22741 6307 22799 6313
rect 22420 6276 22508 6304
rect 22420 6273 22432 6276
rect 22374 6267 22432 6273
rect 21174 6236 21180 6248
rect 18984 6208 20116 6236
rect 21135 6208 21180 6236
rect 18003 6205 18015 6208
rect 17957 6199 18015 6205
rect 16666 6168 16672 6180
rect 11624 6140 16672 6168
rect 16666 6128 16672 6140
rect 16724 6128 16730 6180
rect 17880 6168 17908 6199
rect 18984 6168 19012 6208
rect 21174 6196 21180 6208
rect 21232 6196 21238 6248
rect 22189 6239 22247 6245
rect 22189 6205 22201 6239
rect 22235 6236 22247 6239
rect 22278 6236 22284 6248
rect 22235 6208 22284 6236
rect 22235 6205 22247 6208
rect 22189 6199 22247 6205
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 17880 6140 19012 6168
rect 22480 6168 22508 6276
rect 22741 6273 22753 6307
rect 22787 6273 22799 6307
rect 22741 6267 22799 6273
rect 22833 6307 22891 6313
rect 22833 6273 22845 6307
rect 22879 6273 22891 6307
rect 23382 6304 23388 6316
rect 23343 6276 23388 6304
rect 22833 6267 22891 6273
rect 22756 6236 22784 6267
rect 23382 6264 23388 6276
rect 23440 6304 23446 6316
rect 23584 6304 23612 6344
rect 23845 6341 23857 6344
rect 23891 6341 23903 6375
rect 23845 6335 23903 6341
rect 23440 6276 23612 6304
rect 23661 6307 23719 6313
rect 23440 6264 23446 6276
rect 23661 6273 23673 6307
rect 23707 6304 23719 6307
rect 23750 6304 23756 6316
rect 23707 6276 23756 6304
rect 23707 6273 23719 6276
rect 23661 6267 23719 6273
rect 23293 6239 23351 6245
rect 23293 6236 23305 6239
rect 22756 6208 23305 6236
rect 23293 6205 23305 6208
rect 23339 6205 23351 6239
rect 23676 6236 23704 6267
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 23293 6199 23351 6205
rect 23492 6208 23704 6236
rect 23017 6171 23075 6177
rect 23017 6168 23029 6171
rect 22480 6140 23029 6168
rect 23017 6137 23029 6140
rect 23063 6137 23075 6171
rect 23017 6131 23075 6137
rect 23492 6112 23520 6208
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 7466 6100 7472 6112
rect 6696 6072 7472 6100
rect 6696 6060 6702 6072
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 7834 6100 7840 6112
rect 7795 6072 7840 6100
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8110 6100 8116 6112
rect 8071 6072 8116 6100
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 10100 6072 11345 6100
rect 10100 6060 10106 6072
rect 11333 6069 11345 6072
rect 11379 6100 11391 6103
rect 12526 6100 12532 6112
rect 11379 6072 12532 6100
rect 11379 6069 11391 6072
rect 11333 6063 11391 6069
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 20165 6103 20223 6109
rect 20165 6069 20177 6103
rect 20211 6100 20223 6103
rect 20714 6100 20720 6112
rect 20211 6072 20720 6100
rect 20211 6069 20223 6072
rect 20165 6063 20223 6069
rect 20714 6060 20720 6072
rect 20772 6100 20778 6112
rect 20990 6100 20996 6112
rect 20772 6072 20996 6100
rect 20772 6060 20778 6072
rect 20990 6060 20996 6072
rect 21048 6060 21054 6112
rect 23385 6103 23443 6109
rect 23385 6069 23397 6103
rect 23431 6100 23443 6103
rect 23474 6100 23480 6112
rect 23431 6072 23480 6100
rect 23431 6069 23443 6072
rect 23385 6063 23443 6069
rect 23474 6060 23480 6072
rect 23532 6060 23538 6112
rect 1104 6010 26220 6032
rect 1104 5958 5136 6010
rect 5188 5958 5200 6010
rect 5252 5958 5264 6010
rect 5316 5958 5328 6010
rect 5380 5958 5392 6010
rect 5444 5958 13508 6010
rect 13560 5958 13572 6010
rect 13624 5958 13636 6010
rect 13688 5958 13700 6010
rect 13752 5958 13764 6010
rect 13816 5958 21880 6010
rect 21932 5958 21944 6010
rect 21996 5958 22008 6010
rect 22060 5958 22072 6010
rect 22124 5958 22136 6010
rect 22188 5958 26220 6010
rect 1104 5936 26220 5958
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 5169 5899 5227 5905
rect 5169 5896 5181 5899
rect 4856 5868 5181 5896
rect 4856 5856 4862 5868
rect 5169 5865 5181 5868
rect 5215 5896 5227 5899
rect 5537 5899 5595 5905
rect 5215 5868 5304 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5276 5840 5304 5868
rect 5537 5865 5549 5899
rect 5583 5896 5595 5899
rect 5718 5896 5724 5908
rect 5583 5868 5724 5896
rect 5583 5865 5595 5868
rect 5537 5859 5595 5865
rect 5718 5856 5724 5868
rect 5776 5896 5782 5908
rect 6178 5896 6184 5908
rect 5776 5868 6184 5896
rect 5776 5856 5782 5868
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 8662 5896 8668 5908
rect 6748 5868 8668 5896
rect 5258 5788 5264 5840
rect 5316 5788 5322 5840
rect 5629 5831 5687 5837
rect 5629 5797 5641 5831
rect 5675 5828 5687 5831
rect 6748 5828 6776 5868
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 10137 5899 10195 5905
rect 10137 5896 10149 5899
rect 8864 5868 10149 5896
rect 7377 5831 7435 5837
rect 7377 5828 7389 5831
rect 5675 5800 6776 5828
rect 6840 5800 7389 5828
rect 5675 5797 5687 5800
rect 5629 5791 5687 5797
rect 6638 5760 6644 5772
rect 5368 5732 6644 5760
rect 5368 5704 5396 5732
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 6840 5769 6868 5800
rect 7377 5797 7389 5800
rect 7423 5797 7435 5831
rect 7377 5791 7435 5797
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 8202 5828 8208 5840
rect 7524 5800 7880 5828
rect 7524 5788 7530 5800
rect 6825 5763 6883 5769
rect 6825 5729 6837 5763
rect 6871 5729 6883 5763
rect 6825 5723 6883 5729
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7101 5763 7159 5769
rect 6972 5732 7017 5760
rect 6972 5720 6978 5732
rect 7101 5729 7113 5763
rect 7147 5760 7159 5763
rect 7190 5760 7196 5772
rect 7147 5732 7196 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7300 5711 7411 5726
rect 7281 5705 7411 5711
rect 5350 5692 5356 5704
rect 5311 5664 5356 5692
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5810 5692 5816 5704
rect 5771 5664 5816 5692
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 6086 5692 6092 5704
rect 6047 5664 6092 5692
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6270 5692 6276 5704
rect 6231 5664 6276 5692
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 7009 5695 7067 5701
rect 7009 5661 7021 5695
rect 7055 5692 7067 5695
rect 7055 5664 7236 5692
rect 7281 5671 7293 5705
rect 7327 5698 7411 5705
rect 7327 5671 7339 5698
rect 7281 5665 7339 5671
rect 7383 5692 7411 5698
rect 7558 5692 7564 5704
rect 7383 5664 7564 5692
rect 7055 5661 7067 5664
rect 7009 5655 7067 5661
rect 5997 5627 6055 5633
rect 5997 5593 6009 5627
rect 6043 5624 6055 5627
rect 6362 5624 6368 5636
rect 6043 5596 6368 5624
rect 6043 5593 6055 5596
rect 5997 5587 6055 5593
rect 6362 5584 6368 5596
rect 6420 5584 6426 5636
rect 6457 5627 6515 5633
rect 6457 5593 6469 5627
rect 6503 5624 6515 5627
rect 6546 5624 6552 5636
rect 6503 5596 6552 5624
rect 6503 5593 6515 5596
rect 6457 5587 6515 5593
rect 6546 5584 6552 5596
rect 6604 5584 6610 5636
rect 7208 5624 7236 5664
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7852 5692 7880 5800
rect 8036 5800 8208 5828
rect 8036 5769 8064 5800
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 8389 5831 8447 5837
rect 8389 5797 8401 5831
rect 8435 5828 8447 5831
rect 8754 5828 8760 5840
rect 8435 5800 8760 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 8754 5788 8760 5800
rect 8812 5788 8818 5840
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5729 8079 5763
rect 8021 5723 8079 5729
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 8864 5760 8892 5868
rect 10137 5865 10149 5868
rect 10183 5896 10195 5899
rect 21637 5899 21695 5905
rect 10183 5868 10916 5896
rect 10183 5865 10195 5868
rect 10137 5859 10195 5865
rect 9953 5831 10011 5837
rect 9953 5797 9965 5831
rect 9999 5828 10011 5831
rect 9999 5800 10640 5828
rect 9999 5797 10011 5800
rect 9953 5791 10011 5797
rect 8168 5732 8892 5760
rect 8168 5720 8174 5732
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 7852 5664 8217 5692
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8352 5664 8493 5692
rect 8352 5652 8358 5664
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8754 5692 8760 5704
rect 8715 5664 8760 5692
rect 8481 5655 8539 5661
rect 8754 5652 8760 5664
rect 8812 5692 8818 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8812 5664 8953 5692
rect 8812 5652 8818 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 9122 5692 9128 5704
rect 9083 5664 9128 5692
rect 8941 5655 8999 5661
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 10612 5701 10640 5800
rect 10888 5769 10916 5868
rect 21637 5865 21649 5899
rect 21683 5896 21695 5899
rect 23474 5896 23480 5908
rect 21683 5868 23480 5896
rect 21683 5865 21695 5868
rect 21637 5859 21695 5865
rect 23474 5856 23480 5868
rect 23532 5856 23538 5908
rect 10873 5763 10931 5769
rect 10873 5729 10885 5763
rect 10919 5760 10931 5763
rect 12158 5760 12164 5772
rect 10919 5732 12164 5760
rect 10919 5729 10931 5732
rect 10873 5723 10931 5729
rect 12158 5720 12164 5732
rect 12216 5720 12222 5772
rect 21358 5720 21364 5772
rect 21416 5760 21422 5772
rect 21453 5763 21511 5769
rect 21453 5760 21465 5763
rect 21416 5732 21465 5760
rect 21416 5720 21422 5732
rect 21453 5729 21465 5732
rect 21499 5729 21511 5763
rect 21453 5723 21511 5729
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5692 9367 5695
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9355 5664 9781 5692
rect 9355 5661 9367 5664
rect 9309 5655 9367 5661
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 10686 5692 10692 5704
rect 10643 5664 10692 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 10686 5652 10692 5664
rect 10744 5652 10750 5704
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 18601 5695 18659 5701
rect 18601 5692 18613 5695
rect 12860 5664 18613 5692
rect 12860 5652 12866 5664
rect 18601 5661 18613 5664
rect 18647 5692 18659 5695
rect 19242 5692 19248 5704
rect 18647 5664 19248 5692
rect 18647 5661 18659 5664
rect 18601 5655 18659 5661
rect 19242 5652 19248 5664
rect 19300 5652 19306 5704
rect 21637 5695 21695 5701
rect 21637 5661 21649 5695
rect 21683 5692 21695 5695
rect 21726 5692 21732 5704
rect 21683 5664 21732 5692
rect 21683 5661 21695 5664
rect 21637 5655 21695 5661
rect 21726 5652 21732 5664
rect 21784 5652 21790 5704
rect 8846 5624 8852 5636
rect 7208 5596 8852 5624
rect 8846 5584 8852 5596
rect 8904 5584 8910 5636
rect 11698 5624 11704 5636
rect 10704 5596 11704 5624
rect 6638 5556 6644 5568
rect 6599 5528 6644 5556
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 6880 5528 7757 5556
rect 6880 5516 6886 5528
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 7745 5519 7803 5525
rect 7837 5559 7895 5565
rect 7837 5525 7849 5559
rect 7883 5556 7895 5559
rect 8294 5556 8300 5568
rect 7883 5528 8300 5556
rect 7883 5525 7895 5528
rect 7837 5519 7895 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8481 5559 8539 5565
rect 8481 5525 8493 5559
rect 8527 5556 8539 5559
rect 8665 5559 8723 5565
rect 8665 5556 8677 5559
rect 8527 5528 8677 5556
rect 8527 5525 8539 5528
rect 8481 5519 8539 5525
rect 8665 5525 8677 5528
rect 8711 5525 8723 5559
rect 8665 5519 8723 5525
rect 10229 5559 10287 5565
rect 10229 5525 10241 5559
rect 10275 5556 10287 5559
rect 10410 5556 10416 5568
rect 10275 5528 10416 5556
rect 10275 5525 10287 5528
rect 10229 5519 10287 5525
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 10704 5565 10732 5596
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 20898 5584 20904 5636
rect 20956 5624 20962 5636
rect 21361 5627 21419 5633
rect 21361 5624 21373 5627
rect 20956 5596 21373 5624
rect 20956 5584 20962 5596
rect 21361 5593 21373 5596
rect 21407 5593 21419 5627
rect 21361 5587 21419 5593
rect 10689 5559 10747 5565
rect 10689 5525 10701 5559
rect 10735 5525 10747 5559
rect 10689 5519 10747 5525
rect 11425 5559 11483 5565
rect 11425 5525 11437 5559
rect 11471 5556 11483 5559
rect 12342 5556 12348 5568
rect 11471 5528 12348 5556
rect 11471 5525 11483 5528
rect 11425 5519 11483 5525
rect 12342 5516 12348 5528
rect 12400 5556 12406 5568
rect 13081 5559 13139 5565
rect 13081 5556 13093 5559
rect 12400 5528 13093 5556
rect 12400 5516 12406 5528
rect 13081 5525 13093 5528
rect 13127 5556 13139 5559
rect 13814 5556 13820 5568
rect 13127 5528 13820 5556
rect 13127 5525 13139 5528
rect 13081 5519 13139 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 18782 5556 18788 5568
rect 18743 5528 18788 5556
rect 18782 5516 18788 5528
rect 18840 5516 18846 5568
rect 21450 5516 21456 5568
rect 21508 5556 21514 5568
rect 21821 5559 21879 5565
rect 21821 5556 21833 5559
rect 21508 5528 21833 5556
rect 21508 5516 21514 5528
rect 21821 5525 21833 5528
rect 21867 5525 21879 5559
rect 21821 5519 21879 5525
rect 1104 5466 26220 5488
rect 1104 5414 9322 5466
rect 9374 5414 9386 5466
rect 9438 5414 9450 5466
rect 9502 5414 9514 5466
rect 9566 5414 9578 5466
rect 9630 5414 17694 5466
rect 17746 5414 17758 5466
rect 17810 5414 17822 5466
rect 17874 5414 17886 5466
rect 17938 5414 17950 5466
rect 18002 5414 26220 5466
rect 1104 5392 26220 5414
rect 4801 5355 4859 5361
rect 4801 5321 4813 5355
rect 4847 5352 4859 5355
rect 5350 5352 5356 5364
rect 4847 5324 5356 5352
rect 4847 5321 4859 5324
rect 4801 5315 4859 5321
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 6270 5352 6276 5364
rect 6227 5324 6276 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 6420 5324 6561 5352
rect 6420 5312 6426 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 6549 5315 6607 5321
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 8757 5355 8815 5361
rect 7616 5324 8340 5352
rect 7616 5312 7622 5324
rect 3878 5284 3884 5296
rect 3436 5256 3884 5284
rect 3436 5225 3464 5256
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 6638 5284 6644 5296
rect 5184 5256 6644 5284
rect 3694 5225 3700 5228
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 3688 5179 3700 5225
rect 3752 5216 3758 5228
rect 5184 5225 5212 5256
rect 6638 5244 6644 5256
rect 6696 5244 6702 5296
rect 6914 5244 6920 5296
rect 6972 5284 6978 5296
rect 6972 5256 7052 5284
rect 6972 5244 6978 5256
rect 5169 5219 5227 5225
rect 3752 5188 3788 5216
rect 3694 5176 3700 5179
rect 3752 5176 3758 5188
rect 5169 5185 5181 5219
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 5813 5219 5871 5225
rect 5316 5188 5361 5216
rect 5316 5176 5322 5188
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 5902 5216 5908 5228
rect 5859 5188 5908 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6328 5188 6377 5216
rect 6328 5176 6334 5188
rect 6365 5185 6377 5188
rect 6411 5216 6423 5219
rect 6822 5216 6828 5228
rect 6411 5188 6828 5216
rect 6411 5185 6423 5188
rect 6365 5179 6423 5185
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 7024 5225 7052 5256
rect 7190 5244 7196 5296
rect 7248 5284 7254 5296
rect 8312 5293 8340 5324
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 9030 5352 9036 5364
rect 8803 5324 9036 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 11609 5355 11667 5361
rect 11609 5352 11621 5355
rect 10520 5324 11621 5352
rect 8297 5287 8355 5293
rect 7248 5256 7880 5284
rect 7248 5244 7254 5256
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7374 5216 7380 5228
rect 7335 5188 7380 5216
rect 7009 5179 7067 5185
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 7650 5225 7656 5228
rect 7617 5219 7656 5225
rect 7524 5188 7569 5216
rect 7524 5176 7530 5188
rect 7617 5185 7629 5219
rect 7617 5179 7656 5185
rect 7650 5176 7656 5179
rect 7708 5176 7714 5228
rect 7742 5219 7800 5225
rect 7742 5185 7754 5219
rect 7788 5185 7800 5219
rect 7742 5179 7800 5185
rect 4982 5108 4988 5160
rect 5040 5148 5046 5160
rect 5276 5148 5304 5176
rect 5626 5148 5632 5160
rect 5040 5120 5304 5148
rect 5587 5120 5632 5148
rect 5040 5108 5046 5120
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 6638 5148 6644 5160
rect 5767 5120 6644 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 6914 5148 6920 5160
rect 6875 5120 6920 5148
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5148 7251 5151
rect 7282 5148 7288 5160
rect 7239 5120 7288 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 4430 5040 4436 5092
rect 4488 5080 4494 5092
rect 5077 5083 5135 5089
rect 5077 5080 5089 5083
rect 4488 5052 5089 5080
rect 4488 5040 4494 5052
rect 5077 5049 5089 5052
rect 5123 5049 5135 5083
rect 7116 5080 7144 5111
rect 7282 5108 7288 5120
rect 7340 5148 7346 5160
rect 7760 5148 7788 5179
rect 7852 5157 7880 5256
rect 8297 5253 8309 5287
rect 8343 5253 8355 5287
rect 8297 5247 8355 5253
rect 10134 5244 10140 5296
rect 10192 5284 10198 5296
rect 10422 5287 10480 5293
rect 10422 5284 10434 5287
rect 10192 5256 10434 5284
rect 10192 5244 10198 5256
rect 10422 5253 10434 5256
rect 10468 5284 10480 5287
rect 10520 5284 10548 5324
rect 11609 5321 11621 5324
rect 11655 5321 11667 5355
rect 11609 5315 11667 5321
rect 13354 5312 13360 5364
rect 13412 5352 13418 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 13412 5324 13553 5352
rect 13412 5312 13418 5324
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 13541 5315 13599 5321
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 14369 5355 14427 5361
rect 14369 5352 14381 5355
rect 14148 5324 14381 5352
rect 14148 5312 14154 5324
rect 14369 5321 14381 5324
rect 14415 5321 14427 5355
rect 14369 5315 14427 5321
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15562 5352 15568 5364
rect 15427 5324 15568 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 17957 5355 18015 5361
rect 17957 5321 17969 5355
rect 18003 5352 18015 5355
rect 18046 5352 18052 5364
rect 18003 5324 18052 5352
rect 18003 5321 18015 5324
rect 17957 5315 18015 5321
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 18874 5352 18880 5364
rect 18835 5324 18880 5352
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 19429 5355 19487 5361
rect 19429 5321 19441 5355
rect 19475 5352 19487 5355
rect 19794 5352 19800 5364
rect 19475 5324 19800 5352
rect 19475 5321 19487 5324
rect 19429 5315 19487 5321
rect 19794 5312 19800 5324
rect 19852 5312 19858 5364
rect 20990 5352 20996 5364
rect 20951 5324 20996 5352
rect 20990 5312 20996 5324
rect 21048 5312 21054 5364
rect 22646 5312 22652 5364
rect 22704 5352 22710 5364
rect 22741 5355 22799 5361
rect 22741 5352 22753 5355
rect 22704 5324 22753 5352
rect 22704 5312 22710 5324
rect 22741 5321 22753 5324
rect 22787 5321 22799 5355
rect 22741 5315 22799 5321
rect 11146 5284 11152 5296
rect 10468 5256 10548 5284
rect 10612 5256 11152 5284
rect 10468 5253 10480 5256
rect 10422 5247 10480 5253
rect 8018 5216 8024 5228
rect 7979 5188 8024 5216
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 8573 5219 8631 5225
rect 8573 5216 8585 5219
rect 8260 5188 8585 5216
rect 8260 5176 8266 5188
rect 8573 5185 8585 5188
rect 8619 5185 8631 5219
rect 9122 5216 9128 5228
rect 9083 5188 9128 5216
rect 8573 5179 8631 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 9272 5188 9413 5216
rect 9272 5176 9278 5188
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 10042 5216 10048 5228
rect 10003 5188 10048 5216
rect 9401 5179 9459 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 7340 5120 7788 5148
rect 7837 5151 7895 5157
rect 7340 5108 7346 5120
rect 7837 5117 7849 5151
rect 7883 5117 7895 5151
rect 8386 5148 8392 5160
rect 8347 5120 8392 5148
rect 7837 5111 7895 5117
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 7742 5080 7748 5092
rect 7116 5052 7748 5080
rect 5077 5043 5135 5049
rect 7742 5040 7748 5052
rect 7800 5040 7806 5092
rect 7926 5040 7932 5092
rect 7984 5080 7990 5092
rect 7984 5052 8248 5080
rect 7984 5040 7990 5052
rect 6638 4972 6644 5024
rect 6696 5012 6702 5024
rect 6733 5015 6791 5021
rect 6733 5012 6745 5015
rect 6696 4984 6745 5012
rect 6696 4972 6702 4984
rect 6733 4981 6745 4984
rect 6779 4981 6791 5015
rect 8110 5012 8116 5024
rect 8071 4984 8116 5012
rect 6733 4975 6791 4981
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 8220 5012 8248 5052
rect 8846 5040 8852 5092
rect 8904 5080 8910 5092
rect 10612 5089 10640 5256
rect 11146 5244 11152 5256
rect 11204 5244 11210 5296
rect 18693 5287 18751 5293
rect 12406 5256 12940 5284
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 10744 5188 10793 5216
rect 10744 5176 10750 5188
rect 10781 5185 10793 5188
rect 10827 5185 10839 5219
rect 11241 5219 11299 5225
rect 11241 5216 11253 5219
rect 10781 5179 10839 5185
rect 10980 5188 11253 5216
rect 10980 5089 11008 5188
rect 11241 5185 11253 5188
rect 11287 5185 11299 5219
rect 11241 5179 11299 5185
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 11882 5216 11888 5228
rect 11839 5188 11888 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 11882 5176 11888 5188
rect 11940 5216 11946 5228
rect 12406 5216 12434 5256
rect 12912 5225 12940 5256
rect 13556 5256 18644 5284
rect 11940 5188 12434 5216
rect 12805 5219 12863 5225
rect 11940 5176 11946 5188
rect 12805 5185 12817 5219
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 12820 5148 12848 5179
rect 13556 5148 13584 5256
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 14090 5216 14096 5228
rect 13679 5188 14096 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 14090 5176 14096 5188
rect 14148 5176 14154 5228
rect 18616 5225 18644 5256
rect 18693 5253 18705 5287
rect 18739 5284 18751 5287
rect 18892 5284 18920 5312
rect 21821 5287 21879 5293
rect 21821 5284 21833 5287
rect 18739 5256 21833 5284
rect 18739 5253 18751 5256
rect 18693 5247 18751 5253
rect 15473 5219 15531 5225
rect 14200 5188 14688 5216
rect 13814 5148 13820 5160
rect 11388 5120 13584 5148
rect 13727 5120 13820 5148
rect 11388 5108 11394 5120
rect 13814 5108 13820 5120
rect 13872 5148 13878 5160
rect 14200 5148 14228 5188
rect 14660 5157 14688 5188
rect 15473 5185 15485 5219
rect 15519 5216 15531 5219
rect 16669 5219 16727 5225
rect 16669 5216 16681 5219
rect 15519 5188 16681 5216
rect 15519 5185 15531 5188
rect 15473 5179 15531 5185
rect 16669 5185 16681 5188
rect 16715 5185 16727 5219
rect 16854 5219 16912 5225
rect 16854 5216 16866 5219
rect 16669 5179 16727 5185
rect 16776 5188 16866 5216
rect 13872 5120 14228 5148
rect 14461 5151 14519 5157
rect 13872 5108 13878 5120
rect 14461 5117 14473 5151
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 14645 5151 14703 5157
rect 14645 5117 14657 5151
rect 14691 5148 14703 5151
rect 14921 5151 14979 5157
rect 14921 5148 14933 5151
rect 14691 5120 14933 5148
rect 14691 5117 14703 5120
rect 14645 5111 14703 5117
rect 14921 5117 14933 5120
rect 14967 5148 14979 5151
rect 15657 5151 15715 5157
rect 15657 5148 15669 5151
rect 14967 5120 15669 5148
rect 14967 5117 14979 5120
rect 14921 5111 14979 5117
rect 15657 5117 15669 5120
rect 15703 5117 15715 5151
rect 15657 5111 15715 5117
rect 8941 5083 8999 5089
rect 8941 5080 8953 5083
rect 8904 5052 8953 5080
rect 8904 5040 8910 5052
rect 8941 5049 8953 5052
rect 8987 5049 8999 5083
rect 8941 5043 8999 5049
rect 10597 5083 10655 5089
rect 10597 5049 10609 5083
rect 10643 5049 10655 5083
rect 10597 5043 10655 5049
rect 10965 5083 11023 5089
rect 10965 5049 10977 5083
rect 11011 5049 11023 5083
rect 10965 5043 11023 5049
rect 12802 5040 12808 5092
rect 12860 5080 12866 5092
rect 13173 5083 13231 5089
rect 13173 5080 13185 5083
rect 12860 5052 13185 5080
rect 12860 5040 12866 5052
rect 13173 5049 13185 5052
rect 13219 5049 13231 5083
rect 14476 5080 14504 5111
rect 15470 5080 15476 5092
rect 14476 5052 15476 5080
rect 13173 5043 13231 5049
rect 15470 5040 15476 5052
rect 15528 5040 15534 5092
rect 15672 5080 15700 5111
rect 16206 5108 16212 5160
rect 16264 5148 16270 5160
rect 16776 5148 16804 5188
rect 16854 5185 16866 5188
rect 16900 5185 16912 5219
rect 16854 5179 16912 5185
rect 17497 5219 17555 5225
rect 17497 5185 17509 5219
rect 17543 5216 17555 5219
rect 18601 5219 18659 5225
rect 17543 5188 18276 5216
rect 17543 5185 17555 5188
rect 17497 5179 17555 5185
rect 17218 5148 17224 5160
rect 16264 5120 16804 5148
rect 17179 5120 17224 5148
rect 16264 5108 16270 5120
rect 17218 5108 17224 5120
rect 17276 5108 17282 5160
rect 17313 5151 17371 5157
rect 17313 5117 17325 5151
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 15672 5052 16252 5080
rect 8297 5015 8355 5021
rect 8297 5012 8309 5015
rect 8220 4984 8309 5012
rect 8297 4981 8309 4984
rect 8343 4981 8355 5015
rect 9214 5012 9220 5024
rect 9175 4984 9220 5012
rect 8297 4975 8355 4981
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 10226 4972 10232 5024
rect 10284 5012 10290 5024
rect 10413 5015 10471 5021
rect 10413 5012 10425 5015
rect 10284 4984 10425 5012
rect 10284 4972 10290 4984
rect 10413 4981 10425 4984
rect 10459 4981 10471 5015
rect 10413 4975 10471 4981
rect 10870 4972 10876 5024
rect 10928 5012 10934 5024
rect 11057 5015 11115 5021
rect 11057 5012 11069 5015
rect 10928 4984 11069 5012
rect 10928 4972 10934 4984
rect 11057 4981 11069 4984
rect 11103 4981 11115 5015
rect 11057 4975 11115 4981
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12621 5015 12679 5021
rect 12621 5012 12633 5015
rect 12492 4984 12633 5012
rect 12492 4972 12498 4984
rect 12621 4981 12633 4984
rect 12667 4981 12679 5015
rect 13078 5012 13084 5024
rect 13039 4984 13084 5012
rect 12621 4975 12679 4981
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 13998 5012 14004 5024
rect 13959 4984 14004 5012
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 15010 5012 15016 5024
rect 14971 4984 15016 5012
rect 15010 4972 15016 4984
rect 15068 4972 15074 5024
rect 16224 5021 16252 5052
rect 16482 5040 16488 5092
rect 16540 5080 16546 5092
rect 17328 5080 17356 5111
rect 17512 5080 17540 5179
rect 18248 5157 18276 5188
rect 18601 5185 18613 5219
rect 18647 5216 18659 5219
rect 19426 5216 19432 5228
rect 18647 5188 19432 5216
rect 18647 5185 18659 5188
rect 18601 5179 18659 5185
rect 19426 5176 19432 5188
rect 19484 5176 19490 5228
rect 19628 5160 19656 5256
rect 21821 5253 21833 5256
rect 21867 5284 21879 5287
rect 22189 5287 22247 5293
rect 22189 5284 22201 5287
rect 21867 5256 22201 5284
rect 21867 5253 21879 5256
rect 21821 5247 21879 5253
rect 22189 5253 22201 5256
rect 22235 5253 22247 5287
rect 24305 5287 24363 5293
rect 24305 5284 24317 5287
rect 22189 5247 22247 5253
rect 23768 5256 24317 5284
rect 20131 5219 20189 5225
rect 20131 5185 20143 5219
rect 20177 5216 20189 5219
rect 20622 5216 20628 5228
rect 20177 5188 20628 5216
rect 20177 5185 20189 5188
rect 20131 5179 20189 5185
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 21361 5219 21419 5225
rect 21361 5185 21373 5219
rect 21407 5185 21419 5219
rect 21361 5179 21419 5185
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 18233 5151 18291 5157
rect 18233 5117 18245 5151
rect 18279 5148 18291 5151
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18279 5120 18705 5148
rect 18279 5117 18291 5120
rect 18233 5111 18291 5117
rect 18693 5117 18705 5120
rect 18739 5117 18751 5151
rect 19518 5148 19524 5160
rect 19479 5120 19524 5148
rect 18693 5111 18751 5117
rect 16540 5052 17356 5080
rect 17420 5052 17540 5080
rect 18064 5080 18092 5111
rect 19518 5108 19524 5120
rect 19576 5108 19582 5160
rect 19610 5108 19616 5160
rect 19668 5148 19674 5160
rect 19668 5120 19761 5148
rect 19668 5108 19674 5120
rect 19794 5108 19800 5160
rect 19852 5148 19858 5160
rect 20441 5151 20499 5157
rect 20441 5148 20453 5151
rect 19852 5120 20453 5148
rect 19852 5108 19858 5120
rect 20441 5117 20453 5120
rect 20487 5117 20499 5151
rect 20441 5111 20499 5117
rect 20533 5151 20591 5157
rect 20533 5117 20545 5151
rect 20579 5117 20591 5151
rect 21266 5148 21272 5160
rect 21227 5120 21272 5148
rect 20533 5111 20591 5117
rect 19889 5083 19947 5089
rect 19889 5080 19901 5083
rect 18064 5052 19901 5080
rect 16540 5040 16546 5052
rect 16209 5015 16267 5021
rect 16209 4981 16221 5015
rect 16255 5012 16267 5015
rect 16390 5012 16396 5024
rect 16255 4984 16396 5012
rect 16255 4981 16267 4984
rect 16209 4975 16267 4981
rect 16390 4972 16396 4984
rect 16448 5012 16454 5024
rect 17420 5012 17448 5052
rect 19889 5049 19901 5052
rect 19935 5049 19947 5083
rect 19889 5043 19947 5049
rect 20346 5040 20352 5092
rect 20404 5080 20410 5092
rect 20548 5080 20576 5111
rect 21266 5108 21272 5120
rect 21324 5108 21330 5160
rect 21376 5080 21404 5179
rect 22204 5148 22232 5247
rect 22833 5219 22891 5225
rect 22833 5185 22845 5219
rect 22879 5216 22891 5219
rect 23201 5219 23259 5225
rect 23201 5216 23213 5219
rect 22879 5188 23213 5216
rect 22879 5185 22891 5188
rect 22833 5179 22891 5185
rect 23201 5185 23213 5188
rect 23247 5185 23259 5219
rect 23382 5216 23388 5228
rect 23353 5188 23388 5216
rect 23201 5179 23259 5185
rect 23382 5176 23388 5188
rect 23440 5225 23446 5228
rect 23440 5219 23501 5225
rect 23440 5185 23455 5219
rect 23489 5216 23501 5219
rect 23768 5216 23796 5256
rect 24305 5253 24317 5256
rect 24351 5253 24363 5287
rect 24305 5247 24363 5253
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 23489 5188 23796 5216
rect 23860 5188 23949 5216
rect 23489 5185 23501 5188
rect 23440 5179 23501 5185
rect 23440 5176 23446 5179
rect 23860 5160 23888 5188
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 24121 5219 24179 5225
rect 24121 5185 24133 5219
rect 24167 5185 24179 5219
rect 24121 5179 24179 5185
rect 22462 5148 22468 5160
rect 22204 5120 22468 5148
rect 22462 5108 22468 5120
rect 22520 5148 22526 5160
rect 22925 5151 22983 5157
rect 22925 5148 22937 5151
rect 22520 5120 22937 5148
rect 22520 5108 22526 5120
rect 22925 5117 22937 5120
rect 22971 5117 22983 5151
rect 22925 5111 22983 5117
rect 23753 5151 23811 5157
rect 23753 5117 23765 5151
rect 23799 5117 23811 5151
rect 23753 5111 23811 5117
rect 20404 5052 21404 5080
rect 20404 5040 20410 5052
rect 21726 5040 21732 5092
rect 21784 5080 21790 5092
rect 23768 5080 23796 5111
rect 23842 5108 23848 5160
rect 23900 5148 23906 5160
rect 23900 5120 23945 5148
rect 23900 5108 23906 5120
rect 24136 5092 24164 5179
rect 24118 5080 24124 5092
rect 21784 5052 24124 5080
rect 21784 5040 21790 5052
rect 24118 5040 24124 5052
rect 24176 5040 24182 5092
rect 16448 4984 17448 5012
rect 16448 4972 16454 4984
rect 17494 4972 17500 5024
rect 17552 5012 17558 5024
rect 17589 5015 17647 5021
rect 17589 5012 17601 5015
rect 17552 4984 17601 5012
rect 17552 4972 17558 4984
rect 17589 4981 17601 4984
rect 17635 4981 17647 5015
rect 18414 5012 18420 5024
rect 18375 4984 18420 5012
rect 17589 4975 17647 4981
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 19058 5012 19064 5024
rect 19019 4984 19064 5012
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 21361 5015 21419 5021
rect 21361 4981 21373 5015
rect 21407 5012 21419 5015
rect 21450 5012 21456 5024
rect 21407 4984 21456 5012
rect 21407 4981 21419 4984
rect 21361 4975 21419 4981
rect 21450 4972 21456 4984
rect 21508 4972 21514 5024
rect 22278 4972 22284 5024
rect 22336 5012 22342 5024
rect 22373 5015 22431 5021
rect 22373 5012 22385 5015
rect 22336 4984 22385 5012
rect 22336 4972 22342 4984
rect 22373 4981 22385 4984
rect 22419 4981 22431 5015
rect 22373 4975 22431 4981
rect 1104 4922 26220 4944
rect 1104 4870 5136 4922
rect 5188 4870 5200 4922
rect 5252 4870 5264 4922
rect 5316 4870 5328 4922
rect 5380 4870 5392 4922
rect 5444 4870 13508 4922
rect 13560 4870 13572 4922
rect 13624 4870 13636 4922
rect 13688 4870 13700 4922
rect 13752 4870 13764 4922
rect 13816 4870 21880 4922
rect 21932 4870 21944 4922
rect 21996 4870 22008 4922
rect 22060 4870 22072 4922
rect 22124 4870 22136 4922
rect 22188 4870 26220 4922
rect 1104 4848 26220 4870
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 3694 4808 3700 4820
rect 3651 4780 3700 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3694 4768 3700 4780
rect 3752 4768 3758 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 6270 4808 6276 4820
rect 5307 4780 6276 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 6730 4808 6736 4820
rect 6691 4780 6736 4808
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 7006 4808 7012 4820
rect 6880 4780 7012 4808
rect 6880 4768 6886 4780
rect 7006 4768 7012 4780
rect 7064 4808 7070 4820
rect 7190 4808 7196 4820
rect 7064 4780 7196 4808
rect 7064 4768 7070 4780
rect 7190 4768 7196 4780
rect 7248 4768 7254 4820
rect 7558 4808 7564 4820
rect 7519 4780 7564 4808
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 8076 4780 8677 4808
rect 8076 4768 8082 4780
rect 8665 4777 8677 4780
rect 8711 4808 8723 4811
rect 10226 4808 10232 4820
rect 8711 4780 9996 4808
rect 10187 4780 10232 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 5537 4743 5595 4749
rect 5537 4709 5549 4743
rect 5583 4740 5595 4743
rect 8205 4743 8263 4749
rect 5583 4712 7604 4740
rect 5583 4709 5595 4712
rect 5537 4703 5595 4709
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 6362 4672 6368 4684
rect 6043 4644 6368 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 6362 4632 6368 4644
rect 6420 4672 6426 4684
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6420 4644 7021 4672
rect 6420 4632 6426 4644
rect 7009 4641 7021 4644
rect 7055 4672 7067 4675
rect 7576 4672 7604 4712
rect 8205 4709 8217 4743
rect 8251 4740 8263 4743
rect 8754 4740 8760 4752
rect 8251 4712 8760 4740
rect 8251 4709 8263 4712
rect 8205 4703 8263 4709
rect 8754 4700 8760 4712
rect 8812 4700 8818 4752
rect 9030 4740 9036 4752
rect 8991 4712 9036 4740
rect 9030 4700 9036 4712
rect 9088 4700 9094 4752
rect 9968 4749 9996 4780
rect 10226 4768 10232 4780
rect 10284 4768 10290 4820
rect 12069 4811 12127 4817
rect 12069 4777 12081 4811
rect 12115 4808 12127 4811
rect 12342 4808 12348 4820
rect 12115 4780 12348 4808
rect 12115 4777 12127 4780
rect 12069 4771 12127 4777
rect 9953 4743 10011 4749
rect 9953 4709 9965 4743
rect 9999 4740 10011 4743
rect 10137 4743 10195 4749
rect 10137 4740 10149 4743
rect 9999 4712 10149 4740
rect 9999 4709 10011 4712
rect 9953 4703 10011 4709
rect 10137 4709 10149 4712
rect 10183 4740 10195 4743
rect 11054 4740 11060 4752
rect 10183 4712 11060 4740
rect 10183 4709 10195 4712
rect 10137 4703 10195 4709
rect 9122 4672 9128 4684
rect 7055 4644 7512 4672
rect 7576 4644 9128 4672
rect 7055 4641 7067 4644
rect 7009 4635 7067 4641
rect 3418 4604 3424 4616
rect 3379 4576 3424 4604
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3878 4604 3884 4616
rect 3839 4576 3884 4604
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 4148 4607 4206 4613
rect 4148 4573 4160 4607
rect 4194 4604 4206 4607
rect 4430 4604 4436 4616
rect 4194 4576 4436 4604
rect 4194 4573 4206 4576
rect 4148 4567 4206 4573
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 5718 4604 5724 4616
rect 5679 4576 5724 4604
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 5902 4604 5908 4616
rect 5863 4576 5908 4604
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4604 6607 4607
rect 6822 4604 6828 4616
rect 6595 4576 6828 4604
rect 6595 4573 6607 4576
rect 6549 4567 6607 4573
rect 5920 4468 5948 4564
rect 6196 4536 6224 4567
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 6932 4536 6960 4567
rect 7006 4536 7012 4548
rect 6196 4508 7012 4536
rect 7006 4496 7012 4508
rect 7064 4496 7070 4548
rect 6181 4471 6239 4477
rect 6181 4468 6193 4471
rect 5920 4440 6193 4468
rect 6181 4437 6193 4440
rect 6227 4437 6239 4471
rect 7116 4468 7144 4567
rect 7190 4564 7196 4616
rect 7248 4604 7254 4616
rect 7374 4604 7380 4616
rect 7248 4576 7293 4604
rect 7335 4576 7380 4604
rect 7248 4564 7254 4576
rect 7374 4564 7380 4576
rect 7432 4564 7438 4616
rect 7484 4613 7512 4644
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 10796 4681 10824 4712
rect 11054 4700 11060 4712
rect 11112 4740 11118 4752
rect 12084 4740 12112 4771
rect 12342 4768 12348 4780
rect 12400 4808 12406 4820
rect 13541 4811 13599 4817
rect 12400 4768 12434 4808
rect 13541 4777 13553 4811
rect 13587 4808 13599 4811
rect 13998 4808 14004 4820
rect 13587 4780 14004 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14645 4811 14703 4817
rect 14645 4777 14657 4811
rect 14691 4808 14703 4811
rect 15010 4808 15016 4820
rect 14691 4780 15016 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 15010 4768 15016 4780
rect 15068 4768 15074 4820
rect 15470 4768 15476 4820
rect 15528 4808 15534 4820
rect 15565 4811 15623 4817
rect 15565 4808 15577 4811
rect 15528 4780 15577 4808
rect 15528 4768 15534 4780
rect 15565 4777 15577 4780
rect 15611 4777 15623 4811
rect 17494 4808 17500 4820
rect 17455 4780 17500 4808
rect 15565 4771 15623 4777
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 18785 4811 18843 4817
rect 18785 4777 18797 4811
rect 18831 4808 18843 4811
rect 19058 4808 19064 4820
rect 18831 4780 19064 4808
rect 18831 4777 18843 4780
rect 18785 4771 18843 4777
rect 19058 4768 19064 4780
rect 19116 4768 19122 4820
rect 19518 4768 19524 4820
rect 19576 4808 19582 4820
rect 20533 4811 20591 4817
rect 20533 4808 20545 4811
rect 19576 4780 20545 4808
rect 19576 4768 19582 4780
rect 20533 4777 20545 4780
rect 20579 4777 20591 4811
rect 21266 4808 21272 4820
rect 21227 4780 21272 4808
rect 20533 4771 20591 4777
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 21726 4808 21732 4820
rect 21687 4780 21732 4808
rect 21726 4768 21732 4780
rect 21784 4768 21790 4820
rect 23014 4808 23020 4820
rect 22756 4780 23020 4808
rect 11112 4712 12112 4740
rect 11112 4700 11118 4712
rect 10781 4675 10839 4681
rect 10781 4641 10793 4675
rect 10827 4641 10839 4675
rect 10781 4635 10839 4641
rect 10962 4632 10968 4684
rect 11020 4672 11026 4684
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11020 4644 11713 4672
rect 11020 4632 11026 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 12406 4672 12434 4768
rect 14918 4700 14924 4752
rect 14976 4740 14982 4752
rect 16206 4740 16212 4752
rect 14976 4712 15056 4740
rect 16167 4712 16212 4740
rect 14976 4700 14982 4712
rect 12713 4675 12771 4681
rect 12713 4672 12725 4675
rect 12406 4644 12725 4672
rect 11701 4635 11759 4641
rect 12713 4641 12725 4644
rect 12759 4641 12771 4675
rect 12713 4635 12771 4641
rect 13078 4632 13084 4684
rect 13136 4672 13142 4684
rect 15028 4681 15056 4712
rect 16206 4700 16212 4712
rect 16264 4700 16270 4752
rect 19429 4743 19487 4749
rect 19429 4709 19441 4743
rect 19475 4740 19487 4743
rect 19610 4740 19616 4752
rect 19475 4712 19616 4740
rect 19475 4709 19487 4712
rect 19429 4703 19487 4709
rect 19610 4700 19616 4712
rect 19668 4700 19674 4752
rect 19794 4700 19800 4752
rect 19852 4740 19858 4752
rect 19852 4712 21588 4740
rect 19852 4700 19858 4712
rect 15013 4675 15071 4681
rect 13136 4644 14412 4672
rect 13136 4632 13142 4644
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7892 4576 7941 4604
rect 7892 4564 7898 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8202 4604 8208 4616
rect 8159 4576 8208 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8128 4468 8156 4567
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4604 8355 4607
rect 8386 4604 8392 4616
rect 8343 4576 8392 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 8662 4604 8668 4616
rect 8619 4576 8668 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4604 10655 4607
rect 10870 4604 10876 4616
rect 10643 4576 10876 4604
rect 10643 4573 10655 4576
rect 10597 4567 10655 4573
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 11330 4613 11336 4616
rect 11299 4607 11336 4613
rect 11299 4573 11311 4607
rect 11299 4567 11336 4573
rect 11330 4564 11336 4567
rect 11388 4564 11394 4616
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 12618 4604 12624 4616
rect 12575 4576 12624 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4604 13047 4607
rect 13265 4607 13323 4613
rect 13265 4604 13277 4607
rect 13035 4576 13277 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 13265 4573 13277 4576
rect 13311 4573 13323 4607
rect 13909 4607 13967 4613
rect 13909 4604 13921 4607
rect 13265 4567 13323 4573
rect 13372 4576 13921 4604
rect 10689 4539 10747 4545
rect 10689 4505 10701 4539
rect 10735 4536 10747 4539
rect 11057 4539 11115 4545
rect 11057 4536 11069 4539
rect 10735 4508 11069 4536
rect 10735 4505 10747 4508
rect 10689 4499 10747 4505
rect 11057 4505 11069 4508
rect 11103 4505 11115 4539
rect 11057 4499 11115 4505
rect 12434 4496 12440 4548
rect 12492 4536 12498 4548
rect 13372 4536 13400 4576
rect 13909 4573 13921 4576
rect 13955 4604 13967 4607
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13955 4576 14289 4604
rect 13955 4573 13967 4576
rect 13909 4567 13967 4573
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 12492 4508 13400 4536
rect 13532 4539 13590 4545
rect 12492 4496 12498 4508
rect 13532 4505 13544 4539
rect 13578 4536 13590 4539
rect 14384 4536 14412 4644
rect 15013 4641 15025 4675
rect 15059 4641 15071 4675
rect 16390 4672 16396 4684
rect 16351 4644 16396 4672
rect 15013 4635 15071 4641
rect 16390 4632 16396 4644
rect 16448 4632 16454 4684
rect 19628 4672 19656 4700
rect 20165 4675 20223 4681
rect 20165 4672 20177 4675
rect 19628 4644 20177 4672
rect 20165 4641 20177 4644
rect 20211 4641 20223 4675
rect 20165 4635 20223 4641
rect 20622 4632 20628 4684
rect 20680 4672 20686 4684
rect 20680 4644 21036 4672
rect 20680 4632 20686 4644
rect 14921 4607 14979 4613
rect 14921 4573 14933 4607
rect 14967 4573 14979 4607
rect 14921 4567 14979 4573
rect 14654 4539 14712 4545
rect 14654 4536 14666 4539
rect 13578 4508 14666 4536
rect 13578 4505 13590 4508
rect 13532 4499 13590 4505
rect 14654 4505 14666 4508
rect 14700 4536 14712 4539
rect 14826 4536 14832 4548
rect 14700 4508 14832 4536
rect 14700 4505 14712 4508
rect 14654 4499 14712 4505
rect 14826 4496 14832 4508
rect 14884 4496 14890 4548
rect 14936 4536 14964 4567
rect 15102 4564 15108 4616
rect 15160 4604 15166 4616
rect 15160 4576 15205 4604
rect 15160 4564 15166 4576
rect 15378 4564 15384 4616
rect 15436 4613 15442 4616
rect 15436 4607 15473 4613
rect 15461 4604 15473 4607
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15461 4576 15853 4604
rect 15461 4573 15473 4576
rect 15436 4567 15473 4573
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 16669 4607 16727 4613
rect 16669 4573 16681 4607
rect 16715 4604 16727 4607
rect 16942 4604 16948 4616
rect 16715 4576 16948 4604
rect 16715 4573 16727 4576
rect 16669 4567 16727 4573
rect 15436 4564 15442 4567
rect 16942 4564 16948 4576
rect 17000 4564 17006 4616
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4604 17187 4607
rect 17773 4607 17831 4613
rect 17175 4576 17724 4604
rect 17175 4573 17187 4576
rect 17129 4567 17187 4573
rect 15286 4536 15292 4548
rect 14936 4508 15292 4536
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 16025 4539 16083 4545
rect 16025 4505 16037 4539
rect 16071 4536 16083 4539
rect 17218 4536 17224 4548
rect 16071 4508 17224 4536
rect 16071 4505 16083 4508
rect 16025 4499 16083 4505
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 17696 4536 17724 4576
rect 17773 4573 17785 4607
rect 17819 4604 17831 4607
rect 17865 4607 17923 4613
rect 17865 4604 17877 4607
rect 17819 4576 17877 4604
rect 17819 4573 17831 4576
rect 17773 4567 17831 4573
rect 17865 4573 17877 4576
rect 17911 4573 17923 4607
rect 17865 4567 17923 4573
rect 19061 4607 19119 4613
rect 19061 4573 19073 4607
rect 19107 4604 19119 4607
rect 19518 4604 19524 4616
rect 19107 4576 19524 4604
rect 19107 4573 19119 4576
rect 19061 4567 19119 4573
rect 19518 4564 19524 4576
rect 19576 4564 19582 4616
rect 20438 4564 20444 4616
rect 20496 4604 20502 4616
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 20496 4576 20729 4604
rect 20496 4564 20502 4576
rect 20717 4573 20729 4576
rect 20763 4573 20775 4607
rect 20898 4604 20904 4616
rect 20859 4576 20904 4604
rect 20717 4567 20775 4573
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 21008 4613 21036 4644
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 18414 4536 18420 4548
rect 17696 4508 18420 4536
rect 18414 4496 18420 4508
rect 18472 4496 18478 4548
rect 18782 4496 18788 4548
rect 18840 4545 18846 4548
rect 18840 4536 18852 4545
rect 19981 4539 20039 4545
rect 18840 4508 18885 4536
rect 18840 4499 18852 4508
rect 19981 4505 19993 4539
rect 20027 4536 20039 4539
rect 20806 4536 20812 4548
rect 20027 4508 20812 4536
rect 20027 4505 20039 4508
rect 19981 4499 20039 4505
rect 18840 4496 18846 4499
rect 20806 4496 20812 4508
rect 20864 4496 20870 4548
rect 21008 4536 21036 4567
rect 21174 4564 21180 4616
rect 21232 4604 21238 4616
rect 21453 4607 21511 4613
rect 21453 4604 21465 4607
rect 21232 4576 21465 4604
rect 21232 4564 21238 4576
rect 21453 4573 21465 4576
rect 21499 4573 21511 4607
rect 21560 4604 21588 4712
rect 22756 4684 22784 4780
rect 23014 4768 23020 4780
rect 23072 4768 23078 4820
rect 24118 4808 24124 4820
rect 24079 4780 24124 4808
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 21637 4675 21695 4681
rect 21637 4641 21649 4675
rect 21683 4672 21695 4675
rect 22186 4672 22192 4684
rect 21683 4644 22192 4672
rect 21683 4641 21695 4644
rect 21637 4635 21695 4641
rect 22186 4632 22192 4644
rect 22244 4632 22250 4684
rect 22462 4672 22468 4684
rect 22423 4644 22468 4672
rect 22462 4632 22468 4644
rect 22520 4632 22526 4684
rect 22738 4672 22744 4684
rect 22651 4644 22744 4672
rect 22738 4632 22744 4644
rect 22796 4632 22802 4684
rect 21729 4607 21787 4613
rect 21729 4604 21741 4607
rect 21560 4576 21741 4604
rect 21453 4567 21511 4573
rect 21729 4573 21741 4576
rect 21775 4573 21787 4607
rect 21729 4567 21787 4573
rect 22281 4607 22339 4613
rect 22281 4573 22293 4607
rect 22327 4604 22339 4607
rect 22370 4604 22376 4616
rect 22327 4576 22376 4604
rect 22327 4573 22339 4576
rect 22281 4567 22339 4573
rect 22370 4564 22376 4576
rect 22428 4564 22434 4616
rect 24578 4604 24584 4616
rect 24539 4576 24584 4604
rect 24578 4564 24584 4576
rect 24636 4564 24642 4616
rect 21634 4536 21640 4548
rect 21008 4508 21640 4536
rect 21634 4496 21640 4508
rect 21692 4496 21698 4548
rect 23008 4539 23066 4545
rect 23008 4505 23020 4539
rect 23054 4536 23066 4539
rect 23054 4508 24440 4536
rect 23054 4505 23066 4508
rect 23008 4499 23066 4505
rect 7116 4440 8156 4468
rect 6181 4431 6239 4437
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 8389 4471 8447 4477
rect 8389 4468 8401 4471
rect 8352 4440 8401 4468
rect 8352 4428 8358 4440
rect 8389 4437 8401 4440
rect 8435 4437 8447 4471
rect 12158 4468 12164 4480
rect 12119 4440 12164 4468
rect 8389 4431 8447 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 12621 4471 12679 4477
rect 12621 4437 12633 4471
rect 12667 4468 12679 4471
rect 13078 4468 13084 4480
rect 12667 4440 13084 4468
rect 12667 4437 12679 4440
rect 12621 4431 12679 4437
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 13173 4471 13231 4477
rect 13173 4437 13185 4471
rect 13219 4468 13231 4471
rect 13998 4468 14004 4480
rect 13219 4440 14004 4468
rect 13219 4437 13231 4440
rect 13173 4431 13231 4437
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 16574 4468 16580 4480
rect 16535 4440 16580 4468
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 16942 4428 16948 4480
rect 17000 4468 17006 4480
rect 17037 4471 17095 4477
rect 17037 4468 17049 4471
rect 17000 4440 17049 4468
rect 17000 4428 17006 4440
rect 17037 4437 17049 4440
rect 17083 4437 17095 4471
rect 17037 4431 17095 4437
rect 17126 4428 17132 4480
rect 17184 4468 17190 4480
rect 17506 4471 17564 4477
rect 17506 4468 17518 4471
rect 17184 4440 17518 4468
rect 17184 4428 17190 4440
rect 17506 4437 17518 4440
rect 17552 4437 17564 4471
rect 18046 4468 18052 4480
rect 18007 4440 18052 4468
rect 17506 4431 17564 4437
rect 18046 4428 18052 4440
rect 18104 4428 18110 4480
rect 19610 4468 19616 4480
rect 19571 4440 19616 4468
rect 19610 4428 19616 4440
rect 19668 4428 19674 4480
rect 20070 4428 20076 4480
rect 20128 4468 20134 4480
rect 20128 4440 20173 4468
rect 20128 4428 20134 4440
rect 21358 4428 21364 4480
rect 21416 4468 21422 4480
rect 21913 4471 21971 4477
rect 21913 4468 21925 4471
rect 21416 4440 21925 4468
rect 21416 4428 21422 4440
rect 21913 4437 21925 4440
rect 21959 4437 21971 4471
rect 21913 4431 21971 4437
rect 22373 4471 22431 4477
rect 22373 4437 22385 4471
rect 22419 4468 22431 4471
rect 22646 4468 22652 4480
rect 22419 4440 22652 4468
rect 22419 4437 22431 4440
rect 22373 4431 22431 4437
rect 22646 4428 22652 4440
rect 22704 4428 22710 4480
rect 24412 4477 24440 4508
rect 24397 4471 24455 4477
rect 24397 4437 24409 4471
rect 24443 4437 24455 4471
rect 24397 4431 24455 4437
rect 1104 4378 26220 4400
rect 1104 4326 9322 4378
rect 9374 4326 9386 4378
rect 9438 4326 9450 4378
rect 9502 4326 9514 4378
rect 9566 4326 9578 4378
rect 9630 4326 17694 4378
rect 17746 4326 17758 4378
rect 17810 4326 17822 4378
rect 17874 4326 17886 4378
rect 17938 4326 17950 4378
rect 18002 4326 26220 4378
rect 1104 4304 26220 4326
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 6825 4267 6883 4273
rect 6825 4264 6837 4267
rect 6788 4236 6837 4264
rect 6788 4224 6794 4236
rect 6825 4233 6837 4236
rect 6871 4233 6883 4267
rect 6825 4227 6883 4233
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 7193 4267 7251 4273
rect 7193 4264 7205 4267
rect 6972 4236 7205 4264
rect 6972 4224 6978 4236
rect 7193 4233 7205 4236
rect 7239 4233 7251 4267
rect 7193 4227 7251 4233
rect 7374 4224 7380 4276
rect 7432 4264 7438 4276
rect 7745 4267 7803 4273
rect 7745 4264 7757 4267
rect 7432 4236 7757 4264
rect 7432 4224 7438 4236
rect 7745 4233 7757 4236
rect 7791 4233 7803 4267
rect 7745 4227 7803 4233
rect 9686 4267 9744 4273
rect 9686 4233 9698 4267
rect 9732 4264 9744 4267
rect 10134 4264 10140 4276
rect 9732 4236 10140 4264
rect 9732 4233 9744 4236
rect 9686 4227 9744 4233
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 10410 4264 10416 4276
rect 10371 4236 10416 4264
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 11968 4267 12026 4273
rect 11968 4264 11980 4267
rect 11164 4236 11980 4264
rect 3418 4156 3424 4208
rect 3476 4196 3482 4208
rect 3513 4199 3571 4205
rect 3513 4196 3525 4199
rect 3476 4168 3525 4196
rect 3476 4156 3482 4168
rect 3513 4165 3525 4168
rect 3559 4165 3571 4199
rect 7926 4196 7932 4208
rect 3513 4159 3571 4165
rect 7576 4168 7932 4196
rect 7576 4140 7604 4168
rect 7926 4156 7932 4168
rect 7984 4156 7990 4208
rect 9309 4199 9367 4205
rect 9309 4165 9321 4199
rect 9355 4196 9367 4199
rect 10042 4196 10048 4208
rect 9355 4168 10048 4196
rect 9355 4165 9367 4168
rect 9309 4159 9367 4165
rect 10042 4156 10048 4168
rect 10100 4156 10106 4208
rect 10152 4196 10180 4224
rect 11164 4196 11192 4236
rect 11968 4233 11980 4236
rect 12014 4264 12026 4267
rect 12814 4267 12872 4273
rect 12814 4264 12826 4267
rect 12014 4236 12826 4264
rect 12014 4233 12026 4236
rect 11968 4227 12026 4233
rect 12814 4233 12826 4236
rect 12860 4233 12872 4267
rect 12814 4227 12872 4233
rect 13078 4224 13084 4276
rect 13136 4264 13142 4276
rect 13725 4267 13783 4273
rect 13725 4264 13737 4267
rect 13136 4236 13737 4264
rect 13136 4224 13142 4236
rect 13725 4233 13737 4236
rect 13771 4233 13783 4267
rect 13725 4227 13783 4233
rect 14826 4224 14832 4276
rect 14884 4264 14890 4276
rect 16936 4267 16994 4273
rect 16936 4264 16948 4267
rect 14884 4236 16948 4264
rect 14884 4224 14890 4236
rect 16936 4233 16948 4236
rect 16982 4264 16994 4267
rect 17126 4264 17132 4276
rect 16982 4236 17132 4264
rect 16982 4233 16994 4236
rect 16936 4227 16994 4233
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 17328 4236 18460 4264
rect 11330 4196 11336 4208
rect 10152 4168 11192 4196
rect 11291 4168 11336 4196
rect 11330 4156 11336 4168
rect 11388 4156 11394 4208
rect 12345 4199 12403 4205
rect 12345 4165 12357 4199
rect 12391 4196 12403 4199
rect 12434 4196 12440 4208
rect 12391 4168 12440 4196
rect 12391 4165 12403 4168
rect 12345 4159 12403 4165
rect 12434 4156 12440 4168
rect 12492 4196 12498 4208
rect 12492 4168 12537 4196
rect 12492 4156 12498 4168
rect 15378 4156 15384 4208
rect 15436 4196 15442 4208
rect 16482 4196 16488 4208
rect 15436 4168 16488 4196
rect 15436 4156 15442 4168
rect 16482 4156 16488 4168
rect 16540 4196 16546 4208
rect 17328 4205 17356 4236
rect 18432 4208 18460 4236
rect 18782 4224 18788 4276
rect 18840 4264 18846 4276
rect 19990 4267 20048 4273
rect 19990 4264 20002 4267
rect 18840 4236 20002 4264
rect 18840 4224 18846 4236
rect 19990 4233 20002 4236
rect 20036 4264 20048 4267
rect 21370 4267 21428 4273
rect 21370 4264 21382 4267
rect 20036 4236 21382 4264
rect 20036 4233 20048 4236
rect 19990 4227 20048 4233
rect 21370 4233 21382 4236
rect 21416 4264 21428 4267
rect 22290 4267 22348 4273
rect 22290 4264 22302 4267
rect 21416 4236 22302 4264
rect 21416 4233 21428 4236
rect 21370 4227 21428 4233
rect 22290 4233 22302 4236
rect 22336 4233 22348 4267
rect 22290 4227 22348 4233
rect 17313 4199 17371 4205
rect 16540 4168 17172 4196
rect 16540 4156 16546 4168
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3145 4131 3203 4137
rect 3145 4128 3157 4131
rect 3016 4100 3157 4128
rect 3016 4088 3022 4100
rect 3145 4097 3157 4100
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 3375 4100 3709 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 3697 4097 3709 4100
rect 3743 4128 3755 4131
rect 4982 4128 4988 4140
rect 3743 4100 4988 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 4982 4088 4988 4100
rect 5040 4128 5046 4140
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5040 4100 5825 4128
rect 5040 4088 5046 4100
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4128 6147 4131
rect 6638 4128 6644 4140
rect 6135 4100 6644 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 7558 4128 7564 4140
rect 7519 4100 7564 4128
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 7837 4131 7895 4137
rect 7837 4128 7849 4131
rect 7800 4100 7849 4128
rect 7800 4088 7806 4100
rect 7837 4097 7849 4100
rect 7883 4128 7895 4131
rect 8202 4128 8208 4140
rect 7883 4100 8208 4128
rect 7883 4097 7895 4100
rect 7837 4091 7895 4097
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 10962 4128 10968 4140
rect 10923 4100 10968 4128
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11238 4128 11244 4140
rect 11195 4100 11244 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 11238 4088 11244 4100
rect 11296 4128 11302 4140
rect 11606 4128 11612 4140
rect 11296 4100 11612 4128
rect 11296 4088 11302 4100
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 13354 4088 13360 4140
rect 13412 4128 13418 4140
rect 13575 4131 13633 4137
rect 13575 4128 13587 4131
rect 13412 4100 13587 4128
rect 13412 4088 13418 4100
rect 13575 4097 13587 4100
rect 13621 4097 13633 4131
rect 13906 4128 13912 4140
rect 13867 4100 13912 4128
rect 13575 4091 13633 4097
rect 13906 4088 13912 4100
rect 13964 4088 13970 4140
rect 13998 4088 14004 4140
rect 14056 4128 14062 4140
rect 14165 4131 14223 4137
rect 14165 4128 14177 4131
rect 14056 4100 14177 4128
rect 14056 4088 14062 4100
rect 14165 4097 14177 4100
rect 14211 4097 14223 4131
rect 14165 4091 14223 4097
rect 15286 4088 15292 4140
rect 15344 4128 15350 4140
rect 15473 4131 15531 4137
rect 15473 4128 15485 4131
rect 15344 4100 15485 4128
rect 15344 4088 15350 4100
rect 15473 4097 15485 4100
rect 15519 4097 15531 4131
rect 15473 4091 15531 4097
rect 16083 4131 16141 4137
rect 16083 4097 16095 4131
rect 16129 4128 16141 4131
rect 16393 4131 16451 4137
rect 16129 4097 16160 4128
rect 16083 4091 16160 4097
rect 16393 4097 16405 4131
rect 16439 4128 16451 4131
rect 17144 4128 17172 4168
rect 17313 4165 17325 4199
rect 17359 4165 17371 4199
rect 17313 4159 17371 4165
rect 18046 4156 18052 4208
rect 18104 4196 18110 4208
rect 18294 4199 18352 4205
rect 18294 4196 18306 4199
rect 18104 4168 18306 4196
rect 18104 4156 18110 4168
rect 18294 4165 18306 4168
rect 18340 4165 18352 4199
rect 18294 4159 18352 4165
rect 18414 4156 18420 4208
rect 18472 4196 18478 4208
rect 19613 4199 19671 4205
rect 19613 4196 19625 4199
rect 18472 4168 19625 4196
rect 18472 4156 18478 4168
rect 19613 4165 19625 4168
rect 19659 4165 19671 4199
rect 19613 4159 19671 4165
rect 20714 4156 20720 4208
rect 20772 4196 20778 4208
rect 20993 4199 21051 4205
rect 20993 4196 21005 4199
rect 20772 4168 21005 4196
rect 20772 4156 20778 4168
rect 20993 4165 21005 4168
rect 21039 4196 21051 4199
rect 21913 4199 21971 4205
rect 21913 4196 21925 4199
rect 21039 4168 21925 4196
rect 21039 4165 21051 4168
rect 20993 4159 21051 4165
rect 21913 4165 21925 4168
rect 21959 4165 21971 4199
rect 22646 4196 22652 4208
rect 22607 4168 22652 4196
rect 21913 4159 21971 4165
rect 22646 4156 22652 4168
rect 22704 4156 22710 4208
rect 23753 4199 23811 4205
rect 23753 4196 23765 4199
rect 23308 4168 23765 4196
rect 17405 4131 17463 4137
rect 17405 4128 17417 4131
rect 16439 4100 17080 4128
rect 17144 4100 17417 4128
rect 16439 4097 16451 4100
rect 16393 4091 16451 4097
rect 6178 4060 6184 4072
rect 6139 4032 6184 4060
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 6549 4063 6607 4069
rect 6549 4029 6561 4063
rect 6595 4029 6607 4063
rect 6549 4023 6607 4029
rect 6733 4063 6791 4069
rect 6733 4029 6745 4063
rect 6779 4060 6791 4063
rect 9214 4060 9220 4072
rect 6779 4032 9220 4060
rect 6779 4029 6791 4032
rect 6733 4023 6791 4029
rect 4522 3952 4528 4004
rect 4580 3992 4586 4004
rect 6454 3992 6460 4004
rect 4580 3964 6460 3992
rect 4580 3952 4586 3964
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 2958 3924 2964 3936
rect 2919 3896 2964 3924
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 6564 3924 6592 4023
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4060 10747 4063
rect 11054 4060 11060 4072
rect 10735 4032 11060 4060
rect 10735 4029 10747 4032
rect 10689 4023 10747 4029
rect 7006 3952 7012 4004
rect 7064 3992 7070 4004
rect 7377 3995 7435 4001
rect 7377 3992 7389 3995
rect 7064 3964 7389 3992
rect 7064 3952 7070 3964
rect 7377 3961 7389 3964
rect 7423 3992 7435 3995
rect 7834 3992 7840 4004
rect 7423 3964 7840 3992
rect 7423 3961 7435 3964
rect 7377 3955 7435 3961
rect 7834 3952 7840 3964
rect 7892 3952 7898 4004
rect 10045 3995 10103 4001
rect 10045 3992 10057 3995
rect 9692 3964 10057 3992
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 5684 3896 7941 3924
rect 5684 3884 5690 3896
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 7929 3887 7987 3893
rect 8849 3927 8907 3933
rect 8849 3893 8861 3927
rect 8895 3924 8907 3927
rect 8938 3924 8944 3936
rect 8895 3896 8944 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9692 3933 9720 3964
rect 10045 3961 10057 3964
rect 10091 3961 10103 3995
rect 10520 3992 10548 4023
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 13170 4060 13176 4072
rect 13131 4032 13176 4060
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 13262 4020 13268 4072
rect 13320 4060 13326 4072
rect 13320 4032 13365 4060
rect 13320 4020 13326 4032
rect 11882 3992 11888 4004
rect 10520 3964 11888 3992
rect 10045 3955 10103 3961
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 16132 3992 16160 4091
rect 17052 4072 17080 4100
rect 17405 4097 17417 4100
rect 17451 4097 17463 4131
rect 20346 4128 20352 4140
rect 17405 4091 17463 4097
rect 17788 4100 20352 4128
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 16485 4063 16543 4069
rect 16485 4060 16497 4063
rect 16264 4032 16497 4060
rect 16264 4020 16270 4032
rect 16485 4029 16497 4032
rect 16531 4029 16543 4063
rect 16485 4023 16543 4029
rect 17034 4020 17040 4072
rect 17092 4060 17098 4072
rect 17497 4063 17555 4069
rect 17497 4060 17509 4063
rect 17092 4032 17509 4060
rect 17092 4020 17098 4032
rect 17497 4029 17509 4032
rect 17543 4029 17555 4063
rect 17497 4023 17555 4029
rect 17788 4001 17816 4100
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 20438 4088 20444 4140
rect 20496 4128 20502 4140
rect 20533 4131 20591 4137
rect 20533 4128 20545 4131
rect 20496 4100 20545 4128
rect 20496 4088 20502 4100
rect 20533 4097 20545 4100
rect 20579 4097 20591 4131
rect 20898 4128 20904 4140
rect 20859 4100 20904 4128
rect 20533 4091 20591 4097
rect 20898 4088 20904 4100
rect 20956 4088 20962 4140
rect 22891 4131 22949 4137
rect 22891 4097 22903 4131
rect 22937 4128 22949 4131
rect 23308 4128 23336 4168
rect 23753 4165 23765 4168
rect 23799 4196 23811 4199
rect 23842 4196 23848 4208
rect 23799 4168 23848 4196
rect 23799 4165 23811 4168
rect 23753 4159 23811 4165
rect 23842 4156 23848 4168
rect 23900 4156 23906 4208
rect 22937 4100 23336 4128
rect 23385 4131 23443 4137
rect 22937 4097 22949 4100
rect 22891 4091 22949 4097
rect 23385 4097 23397 4131
rect 23431 4097 23443 4131
rect 23385 4091 23443 4097
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 20717 4063 20775 4069
rect 20717 4029 20729 4063
rect 20763 4060 20775 4063
rect 21450 4060 21456 4072
rect 20763 4032 21456 4060
rect 20763 4029 20775 4032
rect 20717 4023 20775 4029
rect 17773 3995 17831 4001
rect 17773 3992 17785 3995
rect 16132 3964 17785 3992
rect 17773 3961 17785 3964
rect 17819 3961 17831 3995
rect 17773 3955 17831 3961
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3893 9735 3927
rect 9858 3924 9864 3936
rect 9819 3896 9864 3924
rect 9677 3887 9735 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 11790 3924 11796 3936
rect 11751 3896 11796 3924
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 11977 3927 12035 3933
rect 11977 3893 11989 3927
rect 12023 3924 12035 3927
rect 12158 3924 12164 3936
rect 12023 3896 12164 3924
rect 12023 3893 12035 3896
rect 11977 3887 12035 3893
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 12802 3924 12808 3936
rect 12763 3896 12808 3924
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 12986 3924 12992 3936
rect 12947 3896 12992 3924
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 15068 3896 15301 3924
rect 15068 3884 15074 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 15654 3924 15660 3936
rect 15615 3896 15660 3924
rect 15289 3887 15347 3893
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 15933 3927 15991 3933
rect 15933 3893 15945 3927
rect 15979 3924 15991 3927
rect 16574 3924 16580 3936
rect 15979 3896 16580 3924
rect 15979 3893 15991 3896
rect 15933 3887 15991 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 16761 3927 16819 3933
rect 16761 3924 16773 3927
rect 16724 3896 16773 3924
rect 16724 3884 16730 3896
rect 16761 3893 16773 3896
rect 16807 3893 16819 3927
rect 16942 3924 16948 3936
rect 16903 3896 16948 3924
rect 16761 3887 16819 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17218 3884 17224 3936
rect 17276 3924 17282 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 17276 3896 17417 3924
rect 17276 3884 17282 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 18064 3924 18092 4023
rect 21450 4020 21456 4032
rect 21508 4020 21514 4072
rect 22186 4020 22192 4072
rect 22244 4060 22250 4072
rect 23198 4060 23204 4072
rect 22244 4032 23204 4060
rect 22244 4020 22250 4032
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 23290 4020 23296 4072
rect 23348 4060 23354 4072
rect 23400 4060 23428 4091
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 23569 4131 23627 4137
rect 23569 4128 23581 4131
rect 23532 4100 23581 4128
rect 23532 4088 23538 4100
rect 23569 4097 23581 4100
rect 23615 4097 23627 4131
rect 23569 4091 23627 4097
rect 23348 4032 23428 4060
rect 23348 4020 23354 4032
rect 19429 3995 19487 4001
rect 19429 3961 19441 3995
rect 19475 3992 19487 3995
rect 19794 3992 19800 4004
rect 19475 3964 19800 3992
rect 19475 3961 19487 3964
rect 19429 3955 19487 3961
rect 19794 3952 19800 3964
rect 19852 3952 19858 4004
rect 20070 3952 20076 4004
rect 20128 3992 20134 4004
rect 20533 3995 20591 4001
rect 20533 3992 20545 3995
rect 20128 3964 20545 3992
rect 20128 3952 20134 3964
rect 20533 3961 20545 3964
rect 20579 3961 20591 3995
rect 20533 3955 20591 3961
rect 22465 3995 22523 4001
rect 22465 3961 22477 3995
rect 22511 3992 22523 3995
rect 24578 3992 24584 4004
rect 22511 3964 24584 3992
rect 22511 3961 22523 3964
rect 22465 3955 22523 3961
rect 24578 3952 24584 3964
rect 24636 3952 24642 4004
rect 19334 3924 19340 3936
rect 18064 3896 19340 3924
rect 17405 3887 17463 3893
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 19610 3884 19616 3936
rect 19668 3924 19674 3936
rect 19981 3927 20039 3933
rect 19981 3924 19993 3927
rect 19668 3896 19993 3924
rect 19668 3884 19674 3896
rect 19981 3893 19993 3896
rect 20027 3893 20039 3927
rect 20162 3924 20168 3936
rect 20123 3896 20168 3924
rect 19981 3887 20039 3893
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 21358 3924 21364 3936
rect 21319 3896 21364 3924
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 21542 3924 21548 3936
rect 21503 3896 21548 3924
rect 21542 3884 21548 3896
rect 21600 3884 21606 3936
rect 22278 3924 22284 3936
rect 22239 3896 22284 3924
rect 22278 3884 22284 3896
rect 22336 3884 22342 3936
rect 1104 3834 26220 3856
rect 1104 3782 5136 3834
rect 5188 3782 5200 3834
rect 5252 3782 5264 3834
rect 5316 3782 5328 3834
rect 5380 3782 5392 3834
rect 5444 3782 13508 3834
rect 13560 3782 13572 3834
rect 13624 3782 13636 3834
rect 13688 3782 13700 3834
rect 13752 3782 13764 3834
rect 13816 3782 21880 3834
rect 21932 3782 21944 3834
rect 21996 3782 22008 3834
rect 22060 3782 22072 3834
rect 22124 3782 22136 3834
rect 22188 3782 26220 3834
rect 1104 3760 26220 3782
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 6273 3723 6331 3729
rect 6273 3720 6285 3723
rect 5040 3692 6285 3720
rect 5040 3680 5046 3692
rect 6273 3689 6285 3692
rect 6319 3689 6331 3723
rect 6273 3683 6331 3689
rect 6825 3723 6883 3729
rect 6825 3689 6837 3723
rect 6871 3720 6883 3723
rect 7558 3720 7564 3732
rect 6871 3692 7564 3720
rect 6871 3689 6883 3692
rect 6825 3683 6883 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8389 3723 8447 3729
rect 8389 3689 8401 3723
rect 8435 3720 8447 3723
rect 8570 3720 8576 3732
rect 8435 3692 8576 3720
rect 8435 3689 8447 3692
rect 8389 3683 8447 3689
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 8754 3720 8760 3732
rect 8715 3692 8760 3720
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 11238 3720 11244 3732
rect 11199 3692 11244 3720
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 11977 3723 12035 3729
rect 11977 3720 11989 3723
rect 11940 3692 11989 3720
rect 11940 3680 11946 3692
rect 11977 3689 11989 3692
rect 12023 3689 12035 3723
rect 11977 3683 12035 3689
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 14829 3723 14887 3729
rect 14829 3720 14841 3723
rect 14700 3692 14841 3720
rect 14700 3680 14706 3692
rect 14829 3689 14841 3692
rect 14875 3689 14887 3723
rect 14829 3683 14887 3689
rect 15197 3723 15255 3729
rect 15197 3689 15209 3723
rect 15243 3720 15255 3723
rect 15378 3720 15384 3732
rect 15243 3692 15384 3720
rect 15243 3689 15255 3692
rect 15197 3683 15255 3689
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 17034 3720 17040 3732
rect 16995 3692 17040 3720
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 20898 3680 20904 3732
rect 20956 3720 20962 3732
rect 20993 3723 21051 3729
rect 20993 3720 21005 3723
rect 20956 3692 21005 3720
rect 20956 3680 20962 3692
rect 20993 3689 21005 3692
rect 21039 3689 21051 3723
rect 20993 3683 21051 3689
rect 13906 3612 13912 3664
rect 13964 3612 13970 3664
rect 14090 3652 14096 3664
rect 14051 3624 14096 3652
rect 14090 3612 14096 3624
rect 14148 3612 14154 3664
rect 16761 3655 16819 3661
rect 16761 3621 16773 3655
rect 16807 3652 16819 3655
rect 17218 3652 17224 3664
rect 16807 3624 17224 3652
rect 16807 3621 16819 3624
rect 16761 3615 16819 3621
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 21008 3652 21036 3683
rect 21082 3680 21088 3732
rect 21140 3720 21146 3732
rect 21177 3723 21235 3729
rect 21177 3720 21189 3723
rect 21140 3692 21189 3720
rect 21140 3680 21146 3692
rect 21177 3689 21189 3692
rect 21223 3689 21235 3723
rect 21177 3683 21235 3689
rect 21634 3680 21640 3732
rect 21692 3720 21698 3732
rect 21729 3723 21787 3729
rect 21729 3720 21741 3723
rect 21692 3692 21741 3720
rect 21692 3680 21698 3692
rect 21729 3689 21741 3692
rect 21775 3689 21787 3723
rect 23290 3720 23296 3732
rect 21729 3683 21787 3689
rect 22204 3692 23296 3720
rect 22204 3652 22232 3692
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 23382 3680 23388 3732
rect 23440 3720 23446 3732
rect 23569 3723 23627 3729
rect 23569 3720 23581 3723
rect 23440 3692 23581 3720
rect 23440 3680 23446 3692
rect 23569 3689 23581 3692
rect 23615 3689 23627 3723
rect 23569 3683 23627 3689
rect 21008 3624 22232 3652
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 8478 3584 8484 3596
rect 8251 3556 8484 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 8478 3544 8484 3556
rect 8536 3584 8542 3596
rect 9030 3584 9036 3596
rect 8536 3556 9036 3584
rect 8536 3544 8542 3556
rect 9030 3544 9036 3556
rect 9088 3584 9094 3596
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9088 3556 9873 3584
rect 9088 3544 9094 3556
rect 9861 3553 9873 3556
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 11425 3587 11483 3593
rect 11425 3584 11437 3587
rect 11388 3556 11437 3584
rect 11388 3544 11394 3556
rect 11425 3553 11437 3556
rect 11471 3553 11483 3587
rect 13924 3584 13952 3612
rect 15381 3587 15439 3593
rect 15381 3584 15393 3587
rect 11425 3547 11483 3553
rect 13832 3556 15393 3584
rect 7949 3519 8007 3525
rect 7949 3485 7961 3519
rect 7995 3516 8007 3519
rect 8110 3516 8116 3528
rect 7995 3488 8116 3516
rect 7995 3485 8007 3488
rect 7949 3479 8007 3485
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8570 3516 8576 3528
rect 8531 3488 8576 3516
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3516 8815 3519
rect 8846 3516 8852 3528
rect 8803 3488 8852 3516
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 5810 3408 5816 3460
rect 5868 3448 5874 3460
rect 8938 3448 8944 3460
rect 5868 3420 8944 3448
rect 5868 3408 5874 3420
rect 8938 3408 8944 3420
rect 8996 3448 9002 3460
rect 9140 3448 9168 3479
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9585 3519 9643 3525
rect 9272 3488 9317 3516
rect 9272 3476 9278 3488
rect 9585 3485 9597 3519
rect 9631 3516 9643 3519
rect 11514 3516 11520 3528
rect 9631 3488 9812 3516
rect 11475 3488 11520 3516
rect 9631 3485 9643 3488
rect 9585 3479 9643 3485
rect 8996 3420 9168 3448
rect 8996 3408 9002 3420
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 9033 3383 9091 3389
rect 9033 3380 9045 3383
rect 8720 3352 9045 3380
rect 8720 3340 8726 3352
rect 9033 3349 9045 3352
rect 9079 3349 9091 3383
rect 9033 3343 9091 3349
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 9784 3389 9812 3488
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 11884 3519 11942 3525
rect 11884 3485 11896 3519
rect 11930 3516 11942 3519
rect 12161 3519 12219 3525
rect 11930 3488 12112 3516
rect 11930 3485 11942 3488
rect 11884 3479 11942 3485
rect 10128 3451 10186 3457
rect 10128 3417 10140 3451
rect 10174 3448 10186 3451
rect 10962 3448 10968 3460
rect 10174 3420 10968 3448
rect 10174 3417 10186 3420
rect 10128 3411 10186 3417
rect 10962 3408 10968 3420
rect 11020 3408 11026 3460
rect 9769 3383 9827 3389
rect 9769 3380 9781 3383
rect 9180 3352 9781 3380
rect 9180 3340 9186 3352
rect 9769 3349 9781 3352
rect 9815 3380 9827 3383
rect 11606 3380 11612 3392
rect 9815 3352 11612 3380
rect 9815 3349 9827 3352
rect 9769 3343 9827 3349
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 12084 3380 12112 3488
rect 12161 3485 12173 3519
rect 12207 3516 12219 3519
rect 13832 3516 13860 3556
rect 15381 3553 15393 3556
rect 15427 3553 15439 3587
rect 15381 3547 15439 3553
rect 18417 3587 18475 3593
rect 18417 3553 18429 3587
rect 18463 3584 18475 3587
rect 19334 3584 19340 3596
rect 18463 3556 19340 3584
rect 18463 3553 18475 3556
rect 18417 3547 18475 3553
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 21634 3584 21640 3596
rect 21385 3556 21640 3584
rect 12207 3488 13860 3516
rect 13909 3519 13967 3525
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 13909 3485 13921 3519
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 14335 3519 14393 3525
rect 14335 3485 14347 3519
rect 14381 3516 14393 3519
rect 14642 3516 14648 3528
rect 14381 3488 14504 3516
rect 14603 3488 14648 3516
rect 14381 3485 14393 3488
rect 14335 3479 14393 3485
rect 12434 3457 12440 3460
rect 12428 3411 12440 3457
rect 12492 3448 12498 3460
rect 12492 3420 12528 3448
rect 12434 3408 12440 3411
rect 12492 3408 12498 3420
rect 12986 3408 12992 3460
rect 13044 3448 13050 3460
rect 13924 3448 13952 3479
rect 13044 3420 13952 3448
rect 14476 3448 14504 3488
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 14829 3519 14887 3525
rect 14829 3516 14841 3519
rect 14792 3488 14841 3516
rect 14792 3476 14798 3488
rect 14829 3485 14841 3488
rect 14875 3485 14887 3519
rect 15010 3516 15016 3528
rect 14971 3488 15016 3516
rect 14829 3479 14887 3485
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 15654 3525 15660 3528
rect 15648 3516 15660 3525
rect 15615 3488 15660 3516
rect 15648 3479 15660 3488
rect 15654 3476 15660 3479
rect 15712 3476 15718 3528
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3516 18935 3519
rect 20162 3516 20168 3528
rect 18923 3488 20168 3516
rect 18923 3485 18935 3488
rect 18877 3479 18935 3485
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 20346 3476 20352 3528
rect 20404 3516 20410 3528
rect 21385 3525 21413 3556
rect 21634 3544 21640 3556
rect 21692 3544 21698 3596
rect 21361 3519 21419 3525
rect 20404 3488 21312 3516
rect 20404 3476 20410 3488
rect 14918 3448 14924 3460
rect 14476 3420 14924 3448
rect 13044 3408 13050 3420
rect 14918 3408 14924 3420
rect 14976 3408 14982 3460
rect 16850 3408 16856 3460
rect 16908 3448 16914 3460
rect 19610 3457 19616 3460
rect 18150 3451 18208 3457
rect 18150 3448 18162 3451
rect 16908 3420 18162 3448
rect 16908 3408 16914 3420
rect 18150 3417 18162 3420
rect 18196 3417 18208 3451
rect 18150 3411 18208 3417
rect 19604 3411 19616 3457
rect 19668 3448 19674 3460
rect 19668 3420 19704 3448
rect 19610 3408 19616 3411
rect 19668 3408 19674 3420
rect 19794 3408 19800 3460
rect 19852 3448 19858 3460
rect 21284 3448 21312 3488
rect 21361 3485 21373 3519
rect 21407 3485 21419 3519
rect 21361 3479 21419 3485
rect 21542 3476 21548 3528
rect 21600 3516 21606 3528
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21600 3488 21925 3516
rect 21600 3476 21606 3488
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 22189 3519 22247 3525
rect 22189 3485 22201 3519
rect 22235 3516 22247 3519
rect 22738 3516 22744 3528
rect 22235 3488 22744 3516
rect 22235 3485 22247 3488
rect 22189 3479 22247 3485
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 24029 3519 24087 3525
rect 24029 3485 24041 3519
rect 24075 3516 24087 3519
rect 24118 3516 24124 3528
rect 24075 3488 24124 3516
rect 24075 3485 24087 3488
rect 24029 3479 24087 3485
rect 24118 3476 24124 3488
rect 24176 3476 24182 3528
rect 25133 3519 25191 3525
rect 25133 3485 25145 3519
rect 25179 3516 25191 3519
rect 26694 3516 26700 3528
rect 25179 3488 26700 3516
rect 25179 3485 25191 3488
rect 25133 3479 25191 3485
rect 26694 3476 26700 3488
rect 26752 3476 26758 3528
rect 21453 3451 21511 3457
rect 21453 3448 21465 3451
rect 19852 3420 21220 3448
rect 21284 3420 21465 3448
rect 19852 3408 19858 3420
rect 12526 3380 12532 3392
rect 12084 3352 12532 3380
rect 12526 3340 12532 3352
rect 12584 3380 12590 3392
rect 13170 3380 13176 3392
rect 12584 3352 13176 3380
rect 12584 3340 12590 3352
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 13262 3340 13268 3392
rect 13320 3380 13326 3392
rect 13541 3383 13599 3389
rect 13541 3380 13553 3383
rect 13320 3352 13553 3380
rect 13320 3340 13326 3352
rect 13541 3349 13553 3352
rect 13587 3349 13599 3383
rect 13722 3380 13728 3392
rect 13683 3352 13728 3380
rect 13541 3343 13599 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 19058 3380 19064 3392
rect 19019 3352 19064 3380
rect 19058 3340 19064 3352
rect 19116 3340 19122 3392
rect 20717 3383 20775 3389
rect 20717 3349 20729 3383
rect 20763 3380 20775 3383
rect 20898 3380 20904 3392
rect 20763 3352 20904 3380
rect 20763 3349 20775 3352
rect 20717 3343 20775 3349
rect 20898 3340 20904 3352
rect 20956 3380 20962 3392
rect 21082 3380 21088 3392
rect 20956 3352 21088 3380
rect 20956 3340 20962 3352
rect 21082 3340 21088 3352
rect 21140 3340 21146 3392
rect 21192 3380 21220 3420
rect 21453 3417 21465 3420
rect 21499 3417 21511 3451
rect 21453 3411 21511 3417
rect 21637 3451 21695 3457
rect 21637 3417 21649 3451
rect 21683 3417 21695 3451
rect 22434 3451 22492 3457
rect 22434 3448 22446 3451
rect 21637 3411 21695 3417
rect 22112 3420 22446 3448
rect 21652 3380 21680 3411
rect 22112 3389 22140 3420
rect 22434 3417 22446 3420
rect 22480 3417 22492 3451
rect 22434 3411 22492 3417
rect 21192 3352 21680 3380
rect 22097 3383 22155 3389
rect 22097 3349 22109 3383
rect 22143 3349 22155 3383
rect 22097 3343 22155 3349
rect 1104 3290 26220 3312
rect 1104 3238 9322 3290
rect 9374 3238 9386 3290
rect 9438 3238 9450 3290
rect 9502 3238 9514 3290
rect 9566 3238 9578 3290
rect 9630 3238 17694 3290
rect 17746 3238 17758 3290
rect 17810 3238 17822 3290
rect 17874 3238 17886 3290
rect 17938 3238 17950 3290
rect 18002 3238 26220 3290
rect 1104 3216 26220 3238
rect 7742 3176 7748 3188
rect 7703 3148 7748 3176
rect 7742 3136 7748 3148
rect 7800 3136 7806 3188
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 8849 3179 8907 3185
rect 8849 3176 8861 3179
rect 8812 3148 8861 3176
rect 8812 3136 8818 3148
rect 8849 3145 8861 3148
rect 8895 3176 8907 3179
rect 9214 3176 9220 3188
rect 8895 3148 9220 3176
rect 8895 3145 8907 3148
rect 8849 3139 8907 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 10962 3176 10968 3188
rect 10923 3148 10968 3176
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 12492 3148 12537 3176
rect 12492 3136 12498 3148
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 14461 3179 14519 3185
rect 13412 3148 14320 3176
rect 13412 3136 13418 3148
rect 6178 3068 6184 3120
rect 6236 3108 6242 3120
rect 6610 3111 6668 3117
rect 6610 3108 6622 3111
rect 6236 3080 6622 3108
rect 6236 3068 6242 3080
rect 6610 3077 6622 3080
rect 6656 3077 6668 3111
rect 6610 3071 6668 3077
rect 8570 3068 8576 3120
rect 8628 3108 8634 3120
rect 9122 3108 9128 3120
rect 8628 3080 9128 3108
rect 8628 3068 8634 3080
rect 9122 3068 9128 3080
rect 9180 3068 9186 3120
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 11517 3111 11575 3117
rect 11517 3108 11529 3111
rect 11388 3080 11529 3108
rect 11388 3068 11394 3080
rect 11517 3077 11529 3080
rect 11563 3077 11575 3111
rect 11517 3071 11575 3077
rect 11606 3068 11612 3120
rect 11664 3108 11670 3120
rect 13906 3108 13912 3120
rect 11664 3080 13032 3108
rect 11664 3068 11670 3080
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 3936 3012 6377 3040
rect 3936 3000 3942 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 6365 3003 6423 3009
rect 8404 3012 8769 3040
rect 8404 2913 8432 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 9674 3049 9680 3052
rect 9401 3043 9459 3049
rect 9401 3040 9413 3043
rect 9088 3012 9413 3040
rect 9088 3000 9094 3012
rect 9401 3009 9413 3012
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 9668 3003 9680 3049
rect 9732 3040 9738 3052
rect 11146 3040 11152 3052
rect 9732 3012 9768 3040
rect 11107 3012 11152 3040
rect 9674 3000 9680 3003
rect 9732 3000 9738 3012
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 8665 2975 8723 2981
rect 8665 2941 8677 2975
rect 8711 2972 8723 2975
rect 8846 2972 8852 2984
rect 8711 2944 8852 2972
rect 8711 2941 8723 2944
rect 8665 2935 8723 2941
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 11514 2972 11520 2984
rect 10796 2944 11520 2972
rect 10796 2913 10824 2944
rect 11514 2932 11520 2944
rect 11572 2972 11578 2984
rect 11716 2972 11744 3003
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 11848 3012 12633 3040
rect 11848 3000 11854 3012
rect 12621 3009 12633 3012
rect 12667 3009 12679 3043
rect 12621 3003 12679 3009
rect 11572 2944 11744 2972
rect 11885 2975 11943 2981
rect 11572 2932 11578 2944
rect 11885 2941 11897 2975
rect 11931 2972 11943 2975
rect 12526 2972 12532 2984
rect 11931 2944 12532 2972
rect 11931 2941 11943 2944
rect 11885 2935 11943 2941
rect 12526 2932 12532 2944
rect 12584 2932 12590 2984
rect 8389 2907 8447 2913
rect 8389 2904 8401 2907
rect 7668 2876 8401 2904
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 7668 2836 7696 2876
rect 8389 2873 8401 2876
rect 8435 2904 8447 2907
rect 10781 2907 10839 2913
rect 8435 2876 9167 2904
rect 8435 2873 8447 2876
rect 8389 2867 8447 2873
rect 2004 2808 7696 2836
rect 9139 2836 9167 2876
rect 10781 2873 10793 2907
rect 10827 2873 10839 2907
rect 10781 2867 10839 2873
rect 12894 2836 12900 2848
rect 9139 2808 12900 2836
rect 2004 2796 2010 2808
rect 12894 2796 12900 2808
rect 12952 2796 12958 2848
rect 13004 2836 13032 3080
rect 13096 3080 13912 3108
rect 13096 3049 13124 3080
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3009 13139 3043
rect 13081 3003 13139 3009
rect 13348 3043 13406 3049
rect 13348 3009 13360 3043
rect 13394 3040 13406 3043
rect 13722 3040 13728 3052
rect 13394 3012 13728 3040
rect 13394 3009 13406 3012
rect 13348 3003 13406 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14292 3040 14320 3148
rect 14461 3145 14473 3179
rect 14507 3176 14519 3179
rect 14642 3176 14648 3188
rect 14507 3148 14648 3176
rect 14507 3145 14519 3148
rect 14461 3139 14519 3145
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 16850 3176 16856 3188
rect 16811 3148 16856 3176
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 19521 3179 19579 3185
rect 19521 3145 19533 3179
rect 19567 3176 19579 3179
rect 19610 3176 19616 3188
rect 19567 3148 19616 3176
rect 19567 3145 19579 3148
rect 19521 3139 19579 3145
rect 19610 3136 19616 3148
rect 19668 3136 19674 3188
rect 21177 3179 21235 3185
rect 21177 3145 21189 3179
rect 21223 3176 21235 3179
rect 21266 3176 21272 3188
rect 21223 3148 21272 3176
rect 21223 3145 21235 3148
rect 21177 3139 21235 3145
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 21450 3176 21456 3188
rect 21411 3148 21456 3176
rect 21450 3136 21456 3148
rect 21508 3136 21514 3188
rect 14660 3108 14688 3136
rect 14829 3111 14887 3117
rect 14829 3108 14841 3111
rect 14660 3080 14841 3108
rect 14829 3077 14841 3080
rect 14875 3077 14887 3111
rect 14829 3071 14887 3077
rect 14918 3068 14924 3120
rect 14976 3108 14982 3120
rect 15013 3111 15071 3117
rect 15013 3108 15025 3111
rect 14976 3080 15025 3108
rect 14976 3068 14982 3080
rect 15013 3077 15025 3080
rect 15059 3077 15071 3111
rect 15013 3071 15071 3077
rect 19058 3068 19064 3120
rect 19116 3108 19122 3120
rect 20042 3111 20100 3117
rect 20042 3108 20054 3111
rect 19116 3080 20054 3108
rect 19116 3068 19122 3080
rect 20042 3077 20054 3080
rect 20088 3077 20100 3111
rect 20042 3071 20100 3077
rect 14645 3043 14703 3049
rect 14645 3040 14657 3043
rect 14292 3012 14657 3040
rect 14645 3009 14657 3012
rect 14691 3040 14703 3043
rect 14734 3040 14740 3052
rect 14691 3012 14740 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 19337 3043 19395 3049
rect 19337 3009 19349 3043
rect 19383 3009 19395 3043
rect 19337 3003 19395 3009
rect 19352 2972 19380 3003
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 19484 3012 19809 3040
rect 19484 3000 19490 3012
rect 19797 3009 19809 3012
rect 19843 3009 19855 3043
rect 21284 3040 21312 3136
rect 21361 3043 21419 3049
rect 21361 3040 21373 3043
rect 21284 3012 21373 3040
rect 19797 3003 19855 3009
rect 21361 3009 21373 3012
rect 21407 3009 21419 3043
rect 21361 3003 21419 3009
rect 19518 2972 19524 2984
rect 19352 2944 19524 2972
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 22094 2904 22100 2916
rect 20732 2876 22100 2904
rect 20732 2836 20760 2876
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 13004 2808 20760 2836
rect 21542 2796 21548 2848
rect 21600 2836 21606 2848
rect 21821 2839 21879 2845
rect 21821 2836 21833 2839
rect 21600 2808 21833 2836
rect 21600 2796 21606 2808
rect 21821 2805 21833 2808
rect 21867 2805 21879 2839
rect 21821 2799 21879 2805
rect 22741 2839 22799 2845
rect 22741 2805 22753 2839
rect 22787 2836 22799 2839
rect 22830 2836 22836 2848
rect 22787 2808 22836 2836
rect 22787 2805 22799 2808
rect 22741 2799 22799 2805
rect 22830 2796 22836 2808
rect 22888 2796 22894 2848
rect 1104 2746 26220 2768
rect 1104 2694 5136 2746
rect 5188 2694 5200 2746
rect 5252 2694 5264 2746
rect 5316 2694 5328 2746
rect 5380 2694 5392 2746
rect 5444 2694 13508 2746
rect 13560 2694 13572 2746
rect 13624 2694 13636 2746
rect 13688 2694 13700 2746
rect 13752 2694 13764 2746
rect 13816 2694 21880 2746
rect 21932 2694 21944 2746
rect 21996 2694 22008 2746
rect 22060 2694 22072 2746
rect 22124 2694 22136 2746
rect 22188 2694 26220 2746
rect 1104 2672 26220 2694
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 9861 2635 9919 2641
rect 9861 2632 9873 2635
rect 9732 2604 9873 2632
rect 9732 2592 9738 2604
rect 9861 2601 9873 2604
rect 9907 2601 9919 2635
rect 9861 2595 9919 2601
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13449 2635 13507 2641
rect 13449 2632 13461 2635
rect 13412 2604 13461 2632
rect 13412 2592 13418 2604
rect 13449 2601 13461 2604
rect 13495 2601 13507 2635
rect 13449 2595 13507 2601
rect 20438 2564 20444 2576
rect 20399 2536 20444 2564
rect 20438 2524 20444 2536
rect 20496 2524 20502 2576
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 10045 2431 10103 2437
rect 10045 2428 10057 2431
rect 9916 2400 10057 2428
rect 9916 2388 9922 2400
rect 10045 2397 10057 2400
rect 10091 2397 10103 2431
rect 13170 2428 13176 2440
rect 13131 2400 13176 2428
rect 10045 2391 10103 2397
rect 13170 2388 13176 2400
rect 13228 2388 13234 2440
rect 13262 2388 13268 2440
rect 13320 2428 13326 2440
rect 13357 2431 13415 2437
rect 13357 2428 13369 2431
rect 13320 2400 13369 2428
rect 13320 2388 13326 2400
rect 13357 2397 13369 2400
rect 13403 2397 13415 2431
rect 20162 2428 20168 2440
rect 20123 2400 20168 2428
rect 13357 2391 13415 2397
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 20533 2431 20591 2437
rect 20533 2397 20545 2431
rect 20579 2428 20591 2431
rect 20622 2428 20628 2440
rect 20579 2400 20628 2428
rect 20579 2397 20591 2400
rect 20533 2391 20591 2397
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2428 20775 2431
rect 20898 2428 20904 2440
rect 20763 2400 20904 2428
rect 20763 2397 20775 2400
rect 20717 2391 20775 2397
rect 20898 2388 20904 2400
rect 20956 2388 20962 2440
rect 1104 2202 26220 2224
rect 1104 2150 9322 2202
rect 9374 2150 9386 2202
rect 9438 2150 9450 2202
rect 9502 2150 9514 2202
rect 9566 2150 9578 2202
rect 9630 2150 17694 2202
rect 17746 2150 17758 2202
rect 17810 2150 17822 2202
rect 17874 2150 17886 2202
rect 17938 2150 17950 2202
rect 18002 2150 26220 2202
rect 1104 2128 26220 2150
rect 9214 1300 9220 1352
rect 9272 1340 9278 1352
rect 22094 1340 22100 1352
rect 9272 1312 22100 1340
rect 9272 1300 9278 1312
rect 22094 1300 22100 1312
rect 22152 1300 22158 1352
<< via1 >>
rect 26332 28747 26384 28756
rect 26332 28713 26341 28747
rect 26341 28713 26375 28747
rect 26375 28713 26384 28747
rect 26332 28704 26384 28713
rect 9322 27174 9374 27226
rect 9386 27174 9438 27226
rect 9450 27174 9502 27226
rect 9514 27174 9566 27226
rect 9578 27174 9630 27226
rect 17694 27174 17746 27226
rect 17758 27174 17810 27226
rect 17822 27174 17874 27226
rect 17886 27174 17938 27226
rect 17950 27174 18002 27226
rect 9772 26979 9824 26988
rect 9772 26945 9781 26979
rect 9781 26945 9815 26979
rect 9815 26945 9824 26979
rect 9772 26936 9824 26945
rect 14096 26979 14148 26988
rect 14096 26945 14105 26979
rect 14105 26945 14139 26979
rect 14139 26945 14148 26979
rect 14096 26936 14148 26945
rect 9956 26775 10008 26784
rect 9956 26741 9965 26775
rect 9965 26741 9999 26775
rect 9999 26741 10008 26775
rect 9956 26732 10008 26741
rect 14648 26732 14700 26784
rect 5136 26630 5188 26682
rect 5200 26630 5252 26682
rect 5264 26630 5316 26682
rect 5328 26630 5380 26682
rect 5392 26630 5444 26682
rect 13508 26630 13560 26682
rect 13572 26630 13624 26682
rect 13636 26630 13688 26682
rect 13700 26630 13752 26682
rect 13764 26630 13816 26682
rect 21880 26630 21932 26682
rect 21944 26630 21996 26682
rect 22008 26630 22060 26682
rect 22072 26630 22124 26682
rect 22136 26630 22188 26682
rect 14096 26528 14148 26580
rect 7012 26460 7064 26512
rect 9220 26460 9272 26512
rect 10692 26460 10744 26512
rect 13912 26460 13964 26512
rect 11244 26392 11296 26444
rect 14740 26460 14792 26512
rect 7104 26324 7156 26376
rect 7288 26367 7340 26376
rect 7288 26333 7297 26367
rect 7297 26333 7331 26367
rect 7331 26333 7340 26367
rect 7288 26324 7340 26333
rect 9680 26324 9732 26376
rect 10968 26367 11020 26376
rect 9128 26256 9180 26308
rect 10968 26333 10977 26367
rect 10977 26333 11011 26367
rect 11011 26333 11020 26367
rect 10968 26324 11020 26333
rect 11888 26256 11940 26308
rect 12440 26256 12492 26308
rect 14096 26299 14148 26308
rect 14096 26265 14105 26299
rect 14105 26265 14139 26299
rect 14139 26265 14148 26299
rect 14096 26256 14148 26265
rect 15108 26324 15160 26376
rect 14924 26256 14976 26308
rect 7196 26231 7248 26240
rect 7196 26197 7205 26231
rect 7205 26197 7239 26231
rect 7239 26197 7248 26231
rect 7196 26188 7248 26197
rect 9864 26231 9916 26240
rect 9864 26197 9873 26231
rect 9873 26197 9907 26231
rect 9907 26197 9916 26231
rect 9864 26188 9916 26197
rect 14740 26188 14792 26240
rect 9322 26086 9374 26138
rect 9386 26086 9438 26138
rect 9450 26086 9502 26138
rect 9514 26086 9566 26138
rect 9578 26086 9630 26138
rect 17694 26086 17746 26138
rect 17758 26086 17810 26138
rect 17822 26086 17874 26138
rect 17886 26086 17938 26138
rect 17950 26086 18002 26138
rect 1400 25984 1452 26036
rect 7104 25984 7156 26036
rect 7840 25984 7892 26036
rect 9680 26027 9732 26036
rect 9680 25993 9689 26027
rect 9689 25993 9723 26027
rect 9723 25993 9732 26027
rect 11244 26027 11296 26036
rect 9680 25984 9732 25993
rect 11244 25993 11253 26027
rect 11253 25993 11287 26027
rect 11287 25993 11296 26027
rect 11244 25984 11296 25993
rect 480 25848 532 25900
rect 1584 25848 1636 25900
rect 3332 25848 3384 25900
rect 4252 25848 4304 25900
rect 5632 25848 5684 25900
rect 8024 25891 8076 25900
rect 8024 25857 8033 25891
rect 8033 25857 8067 25891
rect 8067 25857 8076 25891
rect 8024 25848 8076 25857
rect 5816 25780 5868 25832
rect 9956 25916 10008 25968
rect 10968 25916 11020 25968
rect 15016 25984 15068 26036
rect 21272 25984 21324 26036
rect 11888 25959 11940 25968
rect 11888 25925 11897 25959
rect 11897 25925 11931 25959
rect 11931 25925 11940 25959
rect 11888 25916 11940 25925
rect 14004 25916 14056 25968
rect 14648 25959 14700 25968
rect 13084 25891 13136 25900
rect 13084 25857 13118 25891
rect 13118 25857 13136 25891
rect 14648 25925 14682 25959
rect 14682 25925 14700 25959
rect 14648 25916 14700 25925
rect 16120 25916 16172 25968
rect 17224 25916 17276 25968
rect 13084 25848 13136 25857
rect 16764 25848 16816 25900
rect 23940 25891 23992 25900
rect 23940 25857 23949 25891
rect 23949 25857 23983 25891
rect 23983 25857 23992 25891
rect 23940 25848 23992 25857
rect 24952 25891 25004 25900
rect 24952 25857 24961 25891
rect 24961 25857 24995 25891
rect 24995 25857 25004 25891
rect 24952 25848 25004 25857
rect 9588 25780 9640 25832
rect 12440 25780 12492 25832
rect 16672 25823 16724 25832
rect 16672 25789 16681 25823
rect 16681 25789 16715 25823
rect 16715 25789 16724 25823
rect 16672 25780 16724 25789
rect 26884 25780 26936 25832
rect 12624 25687 12676 25696
rect 12624 25653 12633 25687
rect 12633 25653 12667 25687
rect 12667 25653 12676 25687
rect 12624 25644 12676 25653
rect 13176 25644 13228 25696
rect 14740 25644 14792 25696
rect 15752 25687 15804 25696
rect 15752 25653 15761 25687
rect 15761 25653 15795 25687
rect 15795 25653 15804 25687
rect 15752 25644 15804 25653
rect 18052 25687 18104 25696
rect 18052 25653 18061 25687
rect 18061 25653 18095 25687
rect 18095 25653 18104 25687
rect 18052 25644 18104 25653
rect 5136 25542 5188 25594
rect 5200 25542 5252 25594
rect 5264 25542 5316 25594
rect 5328 25542 5380 25594
rect 5392 25542 5444 25594
rect 13508 25542 13560 25594
rect 13572 25542 13624 25594
rect 13636 25542 13688 25594
rect 13700 25542 13752 25594
rect 13764 25542 13816 25594
rect 21880 25542 21932 25594
rect 21944 25542 21996 25594
rect 22008 25542 22060 25594
rect 22072 25542 22124 25594
rect 22136 25542 22188 25594
rect 7288 25440 7340 25492
rect 8024 25440 8076 25492
rect 9772 25440 9824 25492
rect 10692 25483 10744 25492
rect 10692 25449 10701 25483
rect 10701 25449 10735 25483
rect 10735 25449 10744 25483
rect 10692 25440 10744 25449
rect 11336 25483 11388 25492
rect 11336 25449 11345 25483
rect 11345 25449 11379 25483
rect 11379 25449 11388 25483
rect 11336 25440 11388 25449
rect 13084 25483 13136 25492
rect 13084 25449 13093 25483
rect 13093 25449 13127 25483
rect 13127 25449 13136 25483
rect 13084 25440 13136 25449
rect 13176 25483 13228 25492
rect 13176 25449 13185 25483
rect 13185 25449 13219 25483
rect 13219 25449 13228 25483
rect 13176 25440 13228 25449
rect 13912 25440 13964 25492
rect 16764 25440 16816 25492
rect 5632 25415 5684 25424
rect 5632 25381 5641 25415
rect 5641 25381 5675 25415
rect 5675 25381 5684 25415
rect 5632 25372 5684 25381
rect 8484 25415 8536 25424
rect 8484 25381 8493 25415
rect 8493 25381 8527 25415
rect 8527 25381 8536 25415
rect 8484 25372 8536 25381
rect 9220 25415 9272 25424
rect 9220 25381 9229 25415
rect 9229 25381 9263 25415
rect 9263 25381 9272 25415
rect 9220 25372 9272 25381
rect 5816 25347 5868 25356
rect 5816 25313 5825 25347
rect 5825 25313 5859 25347
rect 5859 25313 5868 25347
rect 5816 25304 5868 25313
rect 7196 25304 7248 25356
rect 9864 25304 9916 25356
rect 5540 25236 5592 25288
rect 6460 25168 6512 25220
rect 7012 25168 7064 25220
rect 7748 25279 7800 25288
rect 7748 25245 7757 25279
rect 7757 25245 7791 25279
rect 7791 25245 7800 25279
rect 7932 25279 7984 25288
rect 7748 25236 7800 25245
rect 7932 25245 7941 25279
rect 7941 25245 7975 25279
rect 7975 25245 7984 25279
rect 7932 25236 7984 25245
rect 8116 25279 8168 25288
rect 8116 25245 8125 25279
rect 8125 25245 8159 25279
rect 8159 25245 8168 25279
rect 8116 25236 8168 25245
rect 9772 25236 9824 25288
rect 11888 25304 11940 25356
rect 12164 25304 12216 25356
rect 14924 25347 14976 25356
rect 11428 25279 11480 25288
rect 11428 25245 11437 25279
rect 11437 25245 11471 25279
rect 11471 25245 11480 25279
rect 11428 25236 11480 25245
rect 12624 25236 12676 25288
rect 14096 25236 14148 25288
rect 14924 25313 14933 25347
rect 14933 25313 14967 25347
rect 14967 25313 14976 25347
rect 14924 25304 14976 25313
rect 15200 25304 15252 25356
rect 15752 25304 15804 25356
rect 15476 25236 15528 25288
rect 16488 25279 16540 25288
rect 16488 25245 16497 25279
rect 16497 25245 16531 25279
rect 16531 25245 16540 25279
rect 16488 25236 16540 25245
rect 16672 25304 16724 25356
rect 16856 25236 16908 25288
rect 18144 25372 18196 25424
rect 19340 25347 19392 25356
rect 19340 25313 19349 25347
rect 19349 25313 19383 25347
rect 19383 25313 19392 25347
rect 19340 25304 19392 25313
rect 9220 25168 9272 25220
rect 11520 25168 11572 25220
rect 14740 25168 14792 25220
rect 15016 25168 15068 25220
rect 16764 25211 16816 25220
rect 16764 25177 16773 25211
rect 16773 25177 16807 25211
rect 16807 25177 16816 25211
rect 16764 25168 16816 25177
rect 17500 25236 17552 25288
rect 17592 25236 17644 25288
rect 18052 25279 18104 25288
rect 18052 25245 18061 25279
rect 18061 25245 18095 25279
rect 18095 25245 18104 25279
rect 18052 25236 18104 25245
rect 18144 25279 18196 25288
rect 18144 25245 18153 25279
rect 18153 25245 18187 25279
rect 18187 25245 18196 25279
rect 18144 25236 18196 25245
rect 18604 25236 18656 25288
rect 19708 25168 19760 25220
rect 9956 25143 10008 25152
rect 9956 25109 9965 25143
rect 9965 25109 9999 25143
rect 9999 25109 10008 25143
rect 9956 25100 10008 25109
rect 10416 25143 10468 25152
rect 10416 25109 10425 25143
rect 10425 25109 10459 25143
rect 10459 25109 10468 25143
rect 10416 25100 10468 25109
rect 11704 25143 11756 25152
rect 11704 25109 11713 25143
rect 11713 25109 11747 25143
rect 11747 25109 11756 25143
rect 11704 25100 11756 25109
rect 13176 25100 13228 25152
rect 16580 25100 16632 25152
rect 17408 25100 17460 25152
rect 18144 25100 18196 25152
rect 20720 25143 20772 25152
rect 20720 25109 20729 25143
rect 20729 25109 20763 25143
rect 20763 25109 20772 25143
rect 20720 25100 20772 25109
rect 9322 24998 9374 25050
rect 9386 24998 9438 25050
rect 9450 24998 9502 25050
rect 9514 24998 9566 25050
rect 9578 24998 9630 25050
rect 17694 24998 17746 25050
rect 17758 24998 17810 25050
rect 17822 24998 17874 25050
rect 17886 24998 17938 25050
rect 17950 24998 18002 25050
rect 6460 24939 6512 24948
rect 6460 24905 6469 24939
rect 6469 24905 6503 24939
rect 6503 24905 6512 24939
rect 6460 24896 6512 24905
rect 7196 24871 7248 24880
rect 7196 24837 7205 24871
rect 7205 24837 7239 24871
rect 7239 24837 7248 24871
rect 7196 24828 7248 24837
rect 6920 24803 6972 24812
rect 6920 24769 6929 24803
rect 6929 24769 6963 24803
rect 6963 24769 6972 24803
rect 8116 24896 8168 24948
rect 8484 24896 8536 24948
rect 11336 24896 11388 24948
rect 9312 24871 9364 24880
rect 9312 24837 9321 24871
rect 9321 24837 9355 24871
rect 9355 24837 9364 24871
rect 9312 24828 9364 24837
rect 9956 24828 10008 24880
rect 10416 24828 10468 24880
rect 14280 24896 14332 24948
rect 14924 24896 14976 24948
rect 15476 24939 15528 24948
rect 15476 24905 15485 24939
rect 15485 24905 15519 24939
rect 15519 24905 15528 24939
rect 15476 24896 15528 24905
rect 16488 24896 16540 24948
rect 18144 24896 18196 24948
rect 19708 24939 19760 24948
rect 19708 24905 19717 24939
rect 19717 24905 19751 24939
rect 19751 24905 19760 24939
rect 19708 24896 19760 24905
rect 6920 24760 6972 24769
rect 7840 24803 7892 24812
rect 7012 24692 7064 24744
rect 7840 24769 7849 24803
rect 7849 24769 7883 24803
rect 7883 24769 7892 24803
rect 7840 24760 7892 24769
rect 7748 24692 7800 24744
rect 9128 24692 9180 24744
rect 10692 24760 10744 24812
rect 11520 24803 11572 24812
rect 11520 24769 11529 24803
rect 11529 24769 11563 24803
rect 11563 24769 11572 24803
rect 11520 24760 11572 24769
rect 9588 24692 9640 24744
rect 12164 24803 12216 24812
rect 12164 24769 12173 24803
rect 12173 24769 12207 24803
rect 12207 24769 12216 24803
rect 12164 24760 12216 24769
rect 13912 24760 13964 24812
rect 12348 24624 12400 24676
rect 5632 24556 5684 24608
rect 7104 24556 7156 24608
rect 7932 24556 7984 24608
rect 8024 24556 8076 24608
rect 11704 24556 11756 24608
rect 14096 24692 14148 24744
rect 16580 24828 16632 24880
rect 18604 24871 18656 24880
rect 15108 24803 15160 24812
rect 15108 24769 15117 24803
rect 15117 24769 15151 24803
rect 15151 24769 15160 24803
rect 15108 24760 15160 24769
rect 15200 24803 15252 24812
rect 15200 24769 15209 24803
rect 15209 24769 15243 24803
rect 15243 24769 15252 24803
rect 16672 24803 16724 24812
rect 15200 24760 15252 24769
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 17316 24760 17368 24812
rect 17500 24760 17552 24812
rect 18604 24837 18613 24871
rect 18613 24837 18647 24871
rect 18647 24837 18656 24871
rect 18604 24828 18656 24837
rect 14556 24735 14608 24744
rect 14556 24701 14565 24735
rect 14565 24701 14599 24735
rect 14599 24701 14608 24735
rect 14556 24692 14608 24701
rect 14648 24692 14700 24744
rect 16580 24692 16632 24744
rect 18512 24692 18564 24744
rect 16212 24667 16264 24676
rect 14372 24599 14424 24608
rect 14372 24565 14381 24599
rect 14381 24565 14415 24599
rect 14415 24565 14424 24599
rect 14372 24556 14424 24565
rect 14832 24556 14884 24608
rect 15016 24556 15068 24608
rect 15200 24599 15252 24608
rect 15200 24565 15209 24599
rect 15209 24565 15243 24599
rect 15243 24565 15252 24599
rect 16212 24633 16221 24667
rect 16221 24633 16255 24667
rect 16255 24633 16264 24667
rect 16212 24624 16264 24633
rect 19248 24667 19300 24676
rect 19248 24633 19257 24667
rect 19257 24633 19291 24667
rect 19291 24633 19300 24667
rect 19248 24624 19300 24633
rect 20720 24871 20772 24880
rect 20720 24837 20729 24871
rect 20729 24837 20763 24871
rect 20763 24837 20772 24871
rect 20720 24828 20772 24837
rect 21180 24760 21232 24812
rect 15200 24556 15252 24565
rect 17316 24556 17368 24608
rect 17592 24556 17644 24608
rect 19708 24556 19760 24608
rect 26332 24531 26384 24540
rect 5136 24454 5188 24506
rect 5200 24454 5252 24506
rect 5264 24454 5316 24506
rect 5328 24454 5380 24506
rect 5392 24454 5444 24506
rect 13508 24454 13560 24506
rect 13572 24454 13624 24506
rect 13636 24454 13688 24506
rect 13700 24454 13752 24506
rect 13764 24454 13816 24506
rect 21880 24454 21932 24506
rect 21944 24454 21996 24506
rect 22008 24454 22060 24506
rect 22072 24454 22124 24506
rect 22136 24454 22188 24506
rect 26332 24497 26341 24531
rect 26341 24497 26375 24531
rect 26375 24497 26384 24531
rect 26332 24488 26384 24497
rect 5540 24352 5592 24404
rect 7472 24395 7524 24404
rect 7012 24284 7064 24336
rect 7472 24361 7481 24395
rect 7481 24361 7515 24395
rect 7515 24361 7524 24395
rect 7472 24352 7524 24361
rect 7840 24352 7892 24404
rect 9220 24352 9272 24404
rect 9312 24284 9364 24336
rect 9772 24352 9824 24404
rect 11428 24352 11480 24404
rect 7104 24216 7156 24268
rect 7196 24216 7248 24268
rect 8024 24216 8076 24268
rect 9220 24216 9272 24268
rect 9588 24216 9640 24268
rect 14556 24352 14608 24404
rect 14832 24352 14884 24404
rect 15200 24352 15252 24404
rect 16212 24352 16264 24404
rect 12624 24327 12676 24336
rect 12624 24293 12633 24327
rect 12633 24293 12667 24327
rect 12667 24293 12676 24327
rect 12624 24284 12676 24293
rect 14372 24284 14424 24336
rect 15108 24284 15160 24336
rect 19432 24352 19484 24404
rect 12348 24259 12400 24268
rect 5724 24148 5776 24200
rect 6000 24191 6052 24200
rect 4068 24123 4120 24132
rect 4068 24089 4102 24123
rect 4102 24089 4120 24123
rect 6000 24157 6009 24191
rect 6009 24157 6043 24191
rect 6043 24157 6052 24191
rect 6000 24148 6052 24157
rect 7288 24191 7340 24200
rect 7288 24157 7297 24191
rect 7297 24157 7331 24191
rect 7331 24157 7340 24191
rect 7288 24148 7340 24157
rect 7380 24148 7432 24200
rect 7564 24191 7616 24200
rect 7564 24157 7573 24191
rect 7573 24157 7607 24191
rect 7607 24157 7616 24191
rect 7564 24148 7616 24157
rect 9772 24148 9824 24200
rect 11704 24148 11756 24200
rect 12348 24225 12357 24259
rect 12357 24225 12391 24259
rect 12391 24225 12400 24259
rect 12348 24216 12400 24225
rect 15476 24259 15528 24268
rect 14096 24191 14148 24200
rect 14096 24157 14105 24191
rect 14105 24157 14139 24191
rect 14139 24157 14148 24191
rect 14096 24148 14148 24157
rect 4068 24080 4120 24089
rect 7656 24080 7708 24132
rect 9680 24080 9732 24132
rect 4252 24012 4304 24064
rect 5264 24012 5316 24064
rect 7104 24055 7156 24064
rect 7104 24021 7113 24055
rect 7113 24021 7147 24055
rect 7147 24021 7156 24055
rect 7104 24012 7156 24021
rect 12992 24123 13044 24132
rect 12992 24089 13001 24123
rect 13001 24089 13035 24123
rect 13035 24089 13044 24123
rect 12992 24080 13044 24089
rect 13912 24123 13964 24132
rect 13912 24089 13921 24123
rect 13921 24089 13955 24123
rect 13955 24089 13964 24123
rect 14648 24148 14700 24200
rect 15016 24191 15068 24200
rect 15016 24157 15026 24191
rect 15026 24157 15060 24191
rect 15060 24157 15068 24191
rect 15476 24225 15485 24259
rect 15485 24225 15519 24259
rect 15519 24225 15528 24259
rect 15476 24216 15528 24225
rect 17592 24284 17644 24336
rect 18880 24327 18932 24336
rect 18880 24293 18889 24327
rect 18889 24293 18923 24327
rect 18923 24293 18932 24327
rect 18880 24284 18932 24293
rect 19340 24284 19392 24336
rect 16764 24216 16816 24268
rect 17408 24259 17460 24268
rect 17408 24225 17417 24259
rect 17417 24225 17451 24259
rect 17451 24225 17460 24259
rect 17408 24216 17460 24225
rect 17500 24259 17552 24268
rect 17500 24225 17509 24259
rect 17509 24225 17543 24259
rect 17543 24225 17552 24259
rect 17500 24216 17552 24225
rect 15384 24191 15436 24200
rect 15016 24148 15068 24157
rect 15384 24157 15393 24191
rect 15393 24157 15427 24191
rect 15427 24157 15436 24191
rect 15384 24148 15436 24157
rect 18696 24216 18748 24268
rect 21088 24284 21140 24336
rect 21180 24259 21232 24268
rect 18052 24148 18104 24200
rect 18604 24148 18656 24200
rect 14832 24123 14884 24132
rect 13912 24080 13964 24089
rect 14832 24089 14841 24123
rect 14841 24089 14875 24123
rect 14875 24089 14884 24123
rect 14832 24080 14884 24089
rect 16580 24080 16632 24132
rect 18512 24123 18564 24132
rect 18512 24089 18521 24123
rect 18521 24089 18555 24123
rect 18555 24089 18564 24123
rect 18512 24080 18564 24089
rect 11796 24055 11848 24064
rect 11796 24021 11805 24055
rect 11805 24021 11839 24055
rect 11839 24021 11848 24055
rect 11796 24012 11848 24021
rect 11888 24012 11940 24064
rect 14648 24055 14700 24064
rect 14648 24021 14657 24055
rect 14657 24021 14691 24055
rect 14691 24021 14700 24055
rect 14648 24012 14700 24021
rect 16488 24055 16540 24064
rect 16488 24021 16497 24055
rect 16497 24021 16531 24055
rect 16531 24021 16540 24055
rect 16856 24055 16908 24064
rect 16488 24012 16540 24021
rect 16856 24021 16865 24055
rect 16865 24021 16899 24055
rect 16899 24021 16908 24055
rect 16856 24012 16908 24021
rect 21180 24225 21189 24259
rect 21189 24225 21223 24259
rect 21223 24225 21232 24259
rect 21180 24216 21232 24225
rect 21916 24148 21968 24200
rect 23204 24191 23256 24200
rect 22100 24080 22152 24132
rect 22560 24080 22612 24132
rect 23204 24157 23213 24191
rect 23213 24157 23247 24191
rect 23247 24157 23256 24191
rect 23204 24148 23256 24157
rect 24032 24080 24084 24132
rect 20536 24012 20588 24064
rect 9322 23910 9374 23962
rect 9386 23910 9438 23962
rect 9450 23910 9502 23962
rect 9514 23910 9566 23962
rect 9578 23910 9630 23962
rect 17694 23910 17746 23962
rect 17758 23910 17810 23962
rect 17822 23910 17874 23962
rect 17886 23910 17938 23962
rect 17950 23910 18002 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 4252 23808 4304 23860
rect 4068 23740 4120 23792
rect 4160 23715 4212 23724
rect 4160 23681 4169 23715
rect 4169 23681 4203 23715
rect 4203 23681 4212 23715
rect 4160 23672 4212 23681
rect 4436 23715 4488 23724
rect 4436 23681 4445 23715
rect 4445 23681 4479 23715
rect 4479 23681 4488 23715
rect 4436 23672 4488 23681
rect 5816 23740 5868 23792
rect 5264 23672 5316 23724
rect 6000 23808 6052 23860
rect 6828 23715 6880 23724
rect 6828 23681 6837 23715
rect 6837 23681 6871 23715
rect 6871 23681 6880 23715
rect 6828 23672 6880 23681
rect 8116 23808 8168 23860
rect 9772 23851 9824 23860
rect 9772 23817 9781 23851
rect 9781 23817 9815 23851
rect 9815 23817 9824 23851
rect 9772 23808 9824 23817
rect 11796 23808 11848 23860
rect 12440 23808 12492 23860
rect 12992 23808 13044 23860
rect 13912 23808 13964 23860
rect 15384 23851 15436 23860
rect 15384 23817 15393 23851
rect 15393 23817 15427 23851
rect 15427 23817 15436 23851
rect 15384 23808 15436 23817
rect 16764 23851 16816 23860
rect 16764 23817 16773 23851
rect 16773 23817 16807 23851
rect 16807 23817 16816 23851
rect 16764 23808 16816 23817
rect 17500 23808 17552 23860
rect 19340 23808 19392 23860
rect 19708 23851 19760 23860
rect 19708 23817 19717 23851
rect 19717 23817 19751 23851
rect 19751 23817 19760 23851
rect 19708 23808 19760 23817
rect 20536 23851 20588 23860
rect 7288 23740 7340 23792
rect 10784 23783 10836 23792
rect 10784 23749 10793 23783
rect 10793 23749 10827 23783
rect 10827 23749 10836 23783
rect 10784 23740 10836 23749
rect 7196 23715 7248 23724
rect 7196 23681 7205 23715
rect 7205 23681 7239 23715
rect 7239 23681 7248 23715
rect 7196 23672 7248 23681
rect 7380 23604 7432 23656
rect 8576 23672 8628 23724
rect 10692 23672 10744 23724
rect 9772 23604 9824 23656
rect 10048 23604 10100 23656
rect 11888 23715 11940 23724
rect 11888 23681 11897 23715
rect 11897 23681 11931 23715
rect 11931 23681 11940 23715
rect 11888 23672 11940 23681
rect 12164 23715 12216 23724
rect 12164 23681 12173 23715
rect 12173 23681 12207 23715
rect 12207 23681 12216 23715
rect 12164 23672 12216 23681
rect 16580 23740 16632 23792
rect 18880 23740 18932 23792
rect 20536 23817 20545 23851
rect 20545 23817 20579 23851
rect 20579 23817 20588 23851
rect 20536 23808 20588 23817
rect 21180 23808 21232 23860
rect 21088 23783 21140 23792
rect 21088 23749 21097 23783
rect 21097 23749 21131 23783
rect 21131 23749 21140 23783
rect 21088 23740 21140 23749
rect 21916 23740 21968 23792
rect 23204 23808 23256 23860
rect 24032 23783 24084 23792
rect 24032 23749 24041 23783
rect 24041 23749 24075 23783
rect 24075 23749 24084 23783
rect 24032 23740 24084 23749
rect 14004 23715 14056 23724
rect 14004 23681 14013 23715
rect 14013 23681 14047 23715
rect 14047 23681 14056 23715
rect 14004 23672 14056 23681
rect 14096 23672 14148 23724
rect 18328 23715 18380 23724
rect 18328 23681 18337 23715
rect 18337 23681 18371 23715
rect 18371 23681 18380 23715
rect 18328 23672 18380 23681
rect 19984 23672 20036 23724
rect 20812 23672 20864 23724
rect 21732 23672 21784 23724
rect 8208 23536 8260 23588
rect 16856 23579 16908 23588
rect 16856 23545 16865 23579
rect 16865 23545 16899 23579
rect 16899 23545 16908 23579
rect 16856 23536 16908 23545
rect 6736 23468 6788 23520
rect 7472 23511 7524 23520
rect 7472 23477 7481 23511
rect 7481 23477 7515 23511
rect 7515 23477 7524 23511
rect 7472 23468 7524 23477
rect 7748 23468 7800 23520
rect 8116 23511 8168 23520
rect 8116 23477 8125 23511
rect 8125 23477 8159 23511
rect 8159 23477 8168 23511
rect 8116 23468 8168 23477
rect 12164 23468 12216 23520
rect 19708 23604 19760 23656
rect 18512 23536 18564 23588
rect 19248 23579 19300 23588
rect 19248 23545 19257 23579
rect 19257 23545 19291 23579
rect 19291 23545 19300 23579
rect 19248 23536 19300 23545
rect 19432 23468 19484 23520
rect 20536 23604 20588 23656
rect 22100 23647 22152 23656
rect 22100 23613 22109 23647
rect 22109 23613 22143 23647
rect 22143 23613 22152 23647
rect 22100 23604 22152 23613
rect 22744 23468 22796 23520
rect 5136 23366 5188 23418
rect 5200 23366 5252 23418
rect 5264 23366 5316 23418
rect 5328 23366 5380 23418
rect 5392 23366 5444 23418
rect 13508 23366 13560 23418
rect 13572 23366 13624 23418
rect 13636 23366 13688 23418
rect 13700 23366 13752 23418
rect 13764 23366 13816 23418
rect 21880 23366 21932 23418
rect 21944 23366 21996 23418
rect 22008 23366 22060 23418
rect 22072 23366 22124 23418
rect 22136 23366 22188 23418
rect 4160 23239 4212 23248
rect 4160 23205 4169 23239
rect 4169 23205 4203 23239
rect 4203 23205 4212 23239
rect 4160 23196 4212 23205
rect 4436 23128 4488 23180
rect 7104 23264 7156 23316
rect 7196 23264 7248 23316
rect 7012 23196 7064 23248
rect 9772 23307 9824 23316
rect 9772 23273 9781 23307
rect 9781 23273 9815 23307
rect 9815 23273 9824 23307
rect 9772 23264 9824 23273
rect 12624 23307 12676 23316
rect 12624 23273 12633 23307
rect 12633 23273 12667 23307
rect 12667 23273 12676 23307
rect 12624 23264 12676 23273
rect 14096 23264 14148 23316
rect 5540 23128 5592 23180
rect 5816 23128 5868 23180
rect 8208 23171 8260 23180
rect 8208 23137 8217 23171
rect 8217 23137 8251 23171
rect 8251 23137 8260 23171
rect 8208 23128 8260 23137
rect 10784 23128 10836 23180
rect 15108 23264 15160 23316
rect 21732 23264 21784 23316
rect 20628 23196 20680 23248
rect 21456 23171 21508 23180
rect 21456 23137 21465 23171
rect 21465 23137 21499 23171
rect 21499 23137 21508 23171
rect 21456 23128 21508 23137
rect 22560 23171 22612 23180
rect 22560 23137 22569 23171
rect 22569 23137 22603 23171
rect 22603 23137 22612 23171
rect 22560 23128 22612 23137
rect 4712 23103 4764 23112
rect 4712 23069 4721 23103
rect 4721 23069 4755 23103
rect 4755 23069 4764 23103
rect 4712 23060 4764 23069
rect 5632 23103 5684 23112
rect 5632 23069 5641 23103
rect 5641 23069 5675 23103
rect 5675 23069 5684 23103
rect 5632 23060 5684 23069
rect 7840 23103 7892 23112
rect 7840 23069 7849 23103
rect 7849 23069 7883 23103
rect 7883 23069 7892 23103
rect 7840 23060 7892 23069
rect 7932 23103 7984 23112
rect 7932 23069 7941 23103
rect 7941 23069 7975 23103
rect 7975 23069 7984 23103
rect 7932 23060 7984 23069
rect 9956 23103 10008 23112
rect 9956 23069 9965 23103
rect 9965 23069 9999 23103
rect 9999 23069 10008 23103
rect 9956 23060 10008 23069
rect 12164 23060 12216 23112
rect 13820 23060 13872 23112
rect 14556 23060 14608 23112
rect 19708 23060 19760 23112
rect 20536 23060 20588 23112
rect 24032 23128 24084 23180
rect 25136 23171 25188 23180
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 23572 23103 23624 23112
rect 6920 22992 6972 23044
rect 9220 23035 9272 23044
rect 9220 23001 9229 23035
rect 9229 23001 9263 23035
rect 9263 23001 9272 23035
rect 9220 22992 9272 23001
rect 14648 22992 14700 23044
rect 18052 22992 18104 23044
rect 23020 23035 23072 23044
rect 23020 23001 23029 23035
rect 23029 23001 23063 23035
rect 23063 23001 23072 23035
rect 23020 22992 23072 23001
rect 23572 23069 23581 23103
rect 23581 23069 23615 23103
rect 23615 23069 23624 23103
rect 23572 23060 23624 23069
rect 23480 22992 23532 23044
rect 9864 22924 9916 22976
rect 12808 22924 12860 22976
rect 14096 22967 14148 22976
rect 14096 22933 14105 22967
rect 14105 22933 14139 22967
rect 14139 22933 14148 22967
rect 14096 22924 14148 22933
rect 14832 22924 14884 22976
rect 16672 22967 16724 22976
rect 16672 22933 16681 22967
rect 16681 22933 16715 22967
rect 16715 22933 16724 22967
rect 16672 22924 16724 22933
rect 18328 22924 18380 22976
rect 22468 22967 22520 22976
rect 22468 22933 22477 22967
rect 22477 22933 22511 22967
rect 22511 22933 22520 22967
rect 22468 22924 22520 22933
rect 9322 22822 9374 22874
rect 9386 22822 9438 22874
rect 9450 22822 9502 22874
rect 9514 22822 9566 22874
rect 9578 22822 9630 22874
rect 17694 22822 17746 22874
rect 17758 22822 17810 22874
rect 17822 22822 17874 22874
rect 17886 22822 17938 22874
rect 17950 22822 18002 22874
rect 5540 22763 5592 22772
rect 5540 22729 5549 22763
rect 5549 22729 5583 22763
rect 5583 22729 5592 22763
rect 5540 22720 5592 22729
rect 5816 22720 5868 22772
rect 6920 22652 6972 22704
rect 7840 22720 7892 22772
rect 8300 22720 8352 22772
rect 8852 22720 8904 22772
rect 8944 22720 8996 22772
rect 7196 22652 7248 22704
rect 3332 22627 3384 22636
rect 3332 22593 3341 22627
rect 3341 22593 3375 22627
rect 3375 22593 3384 22627
rect 3332 22584 3384 22593
rect 4344 22584 4396 22636
rect 7104 22584 7156 22636
rect 7656 22652 7708 22704
rect 9128 22652 9180 22704
rect 9956 22720 10008 22772
rect 13820 22763 13872 22772
rect 13820 22729 13829 22763
rect 13829 22729 13863 22763
rect 13863 22729 13872 22763
rect 13820 22720 13872 22729
rect 12992 22652 13044 22704
rect 14004 22652 14056 22704
rect 16672 22652 16724 22704
rect 17132 22695 17184 22704
rect 17132 22661 17141 22695
rect 17141 22661 17175 22695
rect 17175 22661 17184 22695
rect 17132 22652 17184 22661
rect 8300 22627 8352 22636
rect 8300 22593 8309 22627
rect 8309 22593 8343 22627
rect 8343 22593 8352 22627
rect 8300 22584 8352 22593
rect 8668 22627 8720 22636
rect 8668 22593 8677 22627
rect 8677 22593 8711 22627
rect 8711 22593 8720 22627
rect 8668 22584 8720 22593
rect 10048 22627 10100 22636
rect 8392 22559 8444 22568
rect 7564 22448 7616 22500
rect 8392 22525 8401 22559
rect 8401 22525 8435 22559
rect 8435 22525 8444 22559
rect 8392 22516 8444 22525
rect 8576 22448 8628 22500
rect 8668 22448 8720 22500
rect 10048 22593 10057 22627
rect 10057 22593 10091 22627
rect 10091 22593 10100 22627
rect 10048 22584 10100 22593
rect 10324 22627 10376 22636
rect 10324 22593 10333 22627
rect 10333 22593 10367 22627
rect 10367 22593 10376 22627
rect 10324 22584 10376 22593
rect 11888 22584 11940 22636
rect 19156 22652 19208 22704
rect 21456 22652 21508 22704
rect 18512 22627 18564 22636
rect 18512 22593 18521 22627
rect 18521 22593 18555 22627
rect 18555 22593 18564 22627
rect 18512 22584 18564 22593
rect 23572 22720 23624 22772
rect 22744 22627 22796 22636
rect 22744 22593 22753 22627
rect 22753 22593 22787 22627
rect 22787 22593 22796 22627
rect 22744 22584 22796 22593
rect 10416 22516 10468 22568
rect 15292 22516 15344 22568
rect 16212 22559 16264 22568
rect 16212 22525 16221 22559
rect 16221 22525 16255 22559
rect 16255 22525 16264 22559
rect 16212 22516 16264 22525
rect 14096 22448 14148 22500
rect 16672 22448 16724 22500
rect 17316 22491 17368 22500
rect 17316 22457 17325 22491
rect 17325 22457 17359 22491
rect 17359 22457 17368 22491
rect 17316 22448 17368 22457
rect 22284 22448 22336 22500
rect 4712 22423 4764 22432
rect 4712 22389 4721 22423
rect 4721 22389 4755 22423
rect 4755 22389 4764 22423
rect 4712 22380 4764 22389
rect 5632 22380 5684 22432
rect 6092 22423 6144 22432
rect 6092 22389 6101 22423
rect 6101 22389 6135 22423
rect 6135 22389 6144 22423
rect 6092 22380 6144 22389
rect 7012 22380 7064 22432
rect 8116 22380 8168 22432
rect 8944 22380 8996 22432
rect 15476 22380 15528 22432
rect 16764 22423 16816 22432
rect 16764 22389 16773 22423
rect 16773 22389 16807 22423
rect 16807 22389 16816 22423
rect 16764 22380 16816 22389
rect 18328 22423 18380 22432
rect 18328 22389 18337 22423
rect 18337 22389 18371 22423
rect 18371 22389 18380 22423
rect 18328 22380 18380 22389
rect 5136 22278 5188 22330
rect 5200 22278 5252 22330
rect 5264 22278 5316 22330
rect 5328 22278 5380 22330
rect 5392 22278 5444 22330
rect 13508 22278 13560 22330
rect 13572 22278 13624 22330
rect 13636 22278 13688 22330
rect 13700 22278 13752 22330
rect 13764 22278 13816 22330
rect 21880 22278 21932 22330
rect 21944 22278 21996 22330
rect 22008 22278 22060 22330
rect 22072 22278 22124 22330
rect 22136 22278 22188 22330
rect 4344 22219 4396 22228
rect 4344 22185 4353 22219
rect 4353 22185 4387 22219
rect 4387 22185 4396 22219
rect 4344 22176 4396 22185
rect 7104 22176 7156 22228
rect 9772 22176 9824 22228
rect 17132 22219 17184 22228
rect 6092 22108 6144 22160
rect 7748 22108 7800 22160
rect 3976 22040 4028 22092
rect 6920 22083 6972 22092
rect 6920 22049 6929 22083
rect 6929 22049 6963 22083
rect 6963 22049 6972 22083
rect 6920 22040 6972 22049
rect 9312 22040 9364 22092
rect 17132 22185 17141 22219
rect 17141 22185 17175 22219
rect 17175 22185 17184 22219
rect 17132 22176 17184 22185
rect 22284 22219 22336 22228
rect 22284 22185 22293 22219
rect 22293 22185 22327 22219
rect 22327 22185 22336 22219
rect 22284 22176 22336 22185
rect 23480 22219 23532 22228
rect 23480 22185 23489 22219
rect 23489 22185 23523 22219
rect 23523 22185 23532 22219
rect 23480 22176 23532 22185
rect 12348 22083 12400 22092
rect 1492 21972 1544 22024
rect 3332 21972 3384 22024
rect 3424 21972 3476 22024
rect 8852 21972 8904 22024
rect 9128 21972 9180 22024
rect 2688 21904 2740 21956
rect 3700 21904 3752 21956
rect 4712 21904 4764 21956
rect 7656 21904 7708 21956
rect 8300 21904 8352 21956
rect 10048 21972 10100 22024
rect 10324 21972 10376 22024
rect 11152 21972 11204 22024
rect 11888 21972 11940 22024
rect 12348 22049 12357 22083
rect 12357 22049 12391 22083
rect 12391 22049 12400 22083
rect 12348 22040 12400 22049
rect 12440 22040 12492 22092
rect 14004 22040 14056 22092
rect 15016 22040 15068 22092
rect 22836 22083 22888 22092
rect 22836 22049 22845 22083
rect 22845 22049 22879 22083
rect 22879 22049 22888 22083
rect 22836 22040 22888 22049
rect 3332 21879 3384 21888
rect 3332 21845 3341 21879
rect 3341 21845 3375 21879
rect 3375 21845 3384 21879
rect 3332 21836 3384 21845
rect 8392 21836 8444 21888
rect 9128 21836 9180 21888
rect 9680 21836 9732 21888
rect 15292 21972 15344 22024
rect 15476 22015 15528 22024
rect 15476 21981 15485 22015
rect 15485 21981 15519 22015
rect 15519 21981 15528 22015
rect 15476 21972 15528 21981
rect 17316 22015 17368 22024
rect 17316 21981 17325 22015
rect 17325 21981 17359 22015
rect 17359 21981 17368 22015
rect 17316 21972 17368 21981
rect 19248 22015 19300 22024
rect 19248 21981 19257 22015
rect 19257 21981 19291 22015
rect 19291 21981 19300 22015
rect 19248 21972 19300 21981
rect 23020 21972 23072 22024
rect 23572 22015 23624 22024
rect 23572 21981 23581 22015
rect 23581 21981 23615 22015
rect 23615 21981 23624 22015
rect 23572 21972 23624 21981
rect 24032 21972 24084 22024
rect 11980 21836 12032 21888
rect 12716 21879 12768 21888
rect 12716 21845 12725 21879
rect 12725 21845 12759 21879
rect 12759 21845 12768 21879
rect 12716 21836 12768 21845
rect 18328 21904 18380 21956
rect 19064 21904 19116 21956
rect 17500 21879 17552 21888
rect 17500 21845 17509 21879
rect 17509 21845 17543 21879
rect 17543 21845 17552 21879
rect 17500 21836 17552 21845
rect 19248 21836 19300 21888
rect 19340 21836 19392 21888
rect 20076 21836 20128 21888
rect 22652 21879 22704 21888
rect 22652 21845 22661 21879
rect 22661 21845 22695 21879
rect 22695 21845 22704 21879
rect 22652 21836 22704 21845
rect 9322 21734 9374 21786
rect 9386 21734 9438 21786
rect 9450 21734 9502 21786
rect 9514 21734 9566 21786
rect 9578 21734 9630 21786
rect 17694 21734 17746 21786
rect 17758 21734 17810 21786
rect 17822 21734 17874 21786
rect 17886 21734 17938 21786
rect 17950 21734 18002 21786
rect 2688 21675 2740 21684
rect 2688 21641 2697 21675
rect 2697 21641 2731 21675
rect 2731 21641 2740 21675
rect 2688 21632 2740 21641
rect 3700 21675 3752 21684
rect 3700 21641 3709 21675
rect 3709 21641 3743 21675
rect 3743 21641 3752 21675
rect 3700 21632 3752 21641
rect 7932 21632 7984 21684
rect 2872 21539 2924 21548
rect 2872 21505 2881 21539
rect 2881 21505 2915 21539
rect 2915 21505 2924 21539
rect 2872 21496 2924 21505
rect 2964 21539 3016 21548
rect 2964 21505 2973 21539
rect 2973 21505 3007 21539
rect 3007 21505 3016 21539
rect 3332 21564 3384 21616
rect 9680 21632 9732 21684
rect 10048 21632 10100 21684
rect 11152 21632 11204 21684
rect 12348 21632 12400 21684
rect 12440 21632 12492 21684
rect 14188 21632 14240 21684
rect 16672 21675 16724 21684
rect 16672 21641 16681 21675
rect 16681 21641 16715 21675
rect 16715 21641 16724 21675
rect 16672 21632 16724 21641
rect 16764 21632 16816 21684
rect 18512 21632 18564 21684
rect 2964 21496 3016 21505
rect 8668 21496 8720 21548
rect 8852 21539 8904 21548
rect 8852 21505 8861 21539
rect 8861 21505 8895 21539
rect 8895 21505 8904 21539
rect 8852 21496 8904 21505
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9864 21564 9916 21616
rect 9036 21496 9088 21505
rect 11888 21564 11940 21616
rect 12716 21607 12768 21616
rect 12716 21573 12734 21607
rect 12734 21573 12768 21607
rect 12716 21564 12768 21573
rect 16212 21564 16264 21616
rect 10232 21539 10284 21548
rect 10232 21505 10241 21539
rect 10241 21505 10275 21539
rect 10275 21505 10284 21539
rect 10232 21496 10284 21505
rect 11980 21496 12032 21548
rect 14004 21496 14056 21548
rect 16120 21496 16172 21548
rect 17132 21496 17184 21548
rect 18328 21496 18380 21548
rect 4160 21471 4212 21480
rect 4160 21437 4169 21471
rect 4169 21437 4203 21471
rect 4203 21437 4212 21471
rect 4160 21428 4212 21437
rect 15016 21471 15068 21480
rect 4436 21360 4488 21412
rect 9128 21360 9180 21412
rect 15016 21437 15025 21471
rect 15025 21437 15059 21471
rect 15059 21437 15068 21471
rect 15016 21428 15068 21437
rect 17500 21428 17552 21480
rect 18880 21428 18932 21480
rect 10048 21403 10100 21412
rect 10048 21369 10057 21403
rect 10057 21369 10091 21403
rect 10091 21369 10100 21403
rect 19156 21496 19208 21548
rect 19432 21539 19484 21548
rect 19432 21505 19441 21539
rect 19441 21505 19475 21539
rect 19475 21505 19484 21539
rect 19432 21496 19484 21505
rect 19708 21539 19760 21548
rect 19708 21505 19718 21539
rect 19718 21505 19752 21539
rect 19752 21505 19760 21539
rect 19708 21496 19760 21505
rect 21364 21496 21416 21548
rect 19248 21428 19300 21480
rect 20076 21471 20128 21480
rect 10048 21360 10100 21369
rect 20076 21437 20085 21471
rect 20085 21437 20119 21471
rect 20119 21437 20128 21471
rect 20076 21428 20128 21437
rect 20168 21471 20220 21480
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 21272 21471 21324 21480
rect 21272 21437 21281 21471
rect 21281 21437 21315 21471
rect 21315 21437 21324 21471
rect 21824 21564 21876 21616
rect 22284 21564 22336 21616
rect 22560 21539 22612 21548
rect 22560 21505 22569 21539
rect 22569 21505 22603 21539
rect 22603 21505 22612 21539
rect 22560 21496 22612 21505
rect 21272 21428 21324 21437
rect 23204 21496 23256 21548
rect 23480 21539 23532 21548
rect 23480 21505 23489 21539
rect 23489 21505 23523 21539
rect 23523 21505 23532 21539
rect 23480 21496 23532 21505
rect 23296 21428 23348 21480
rect 3148 21335 3200 21344
rect 3148 21301 3157 21335
rect 3157 21301 3191 21335
rect 3191 21301 3200 21335
rect 3148 21292 3200 21301
rect 3332 21335 3384 21344
rect 3332 21301 3341 21335
rect 3341 21301 3375 21335
rect 3375 21301 3384 21335
rect 3332 21292 3384 21301
rect 7656 21292 7708 21344
rect 8944 21335 8996 21344
rect 8944 21301 8953 21335
rect 8953 21301 8987 21335
rect 8987 21301 8996 21335
rect 8944 21292 8996 21301
rect 16028 21292 16080 21344
rect 19340 21335 19392 21344
rect 19340 21301 19349 21335
rect 19349 21301 19383 21335
rect 19383 21301 19392 21335
rect 19340 21292 19392 21301
rect 19616 21335 19668 21344
rect 19616 21301 19625 21335
rect 19625 21301 19659 21335
rect 19659 21301 19668 21335
rect 19616 21292 19668 21301
rect 21456 21360 21508 21412
rect 21640 21292 21692 21344
rect 22836 21292 22888 21344
rect 22928 21335 22980 21344
rect 22928 21301 22937 21335
rect 22937 21301 22971 21335
rect 22971 21301 22980 21335
rect 22928 21292 22980 21301
rect 5136 21190 5188 21242
rect 5200 21190 5252 21242
rect 5264 21190 5316 21242
rect 5328 21190 5380 21242
rect 5392 21190 5444 21242
rect 13508 21190 13560 21242
rect 13572 21190 13624 21242
rect 13636 21190 13688 21242
rect 13700 21190 13752 21242
rect 13764 21190 13816 21242
rect 21880 21190 21932 21242
rect 21944 21190 21996 21242
rect 22008 21190 22060 21242
rect 22072 21190 22124 21242
rect 22136 21190 22188 21242
rect 2872 21088 2924 21140
rect 4160 21088 4212 21140
rect 4804 21088 4856 21140
rect 9036 21088 9088 21140
rect 10048 21131 10100 21140
rect 10048 21097 10057 21131
rect 10057 21097 10091 21131
rect 10091 21097 10100 21131
rect 10048 21088 10100 21097
rect 1492 20995 1544 21004
rect 1492 20961 1501 20995
rect 1501 20961 1535 20995
rect 1535 20961 1544 20995
rect 1492 20952 1544 20961
rect 3148 20952 3200 21004
rect 4436 20995 4488 21004
rect 3424 20927 3476 20936
rect 3424 20893 3433 20927
rect 3433 20893 3467 20927
rect 3467 20893 3476 20927
rect 3424 20884 3476 20893
rect 4436 20961 4445 20995
rect 4445 20961 4479 20995
rect 4479 20961 4488 20995
rect 4436 20952 4488 20961
rect 9220 21020 9272 21072
rect 8300 20995 8352 21004
rect 8300 20961 8309 20995
rect 8309 20961 8343 20995
rect 8343 20961 8352 20995
rect 8300 20952 8352 20961
rect 8944 20952 8996 21004
rect 5540 20884 5592 20936
rect 6828 20884 6880 20936
rect 6920 20884 6972 20936
rect 7840 20884 7892 20936
rect 8852 20884 8904 20936
rect 10232 20884 10284 20936
rect 11428 20884 11480 20936
rect 12440 21088 12492 21140
rect 17500 21131 17552 21140
rect 17500 21097 17509 21131
rect 17509 21097 17543 21131
rect 17543 21097 17552 21131
rect 17500 21088 17552 21097
rect 11980 20995 12032 21004
rect 11980 20961 11989 20995
rect 11989 20961 12023 20995
rect 12023 20961 12032 20995
rect 11980 20952 12032 20961
rect 16212 20952 16264 21004
rect 12164 20927 12216 20936
rect 2504 20816 2556 20868
rect 3056 20816 3108 20868
rect 6000 20816 6052 20868
rect 6092 20859 6144 20868
rect 6092 20825 6110 20859
rect 6110 20825 6144 20859
rect 6092 20816 6144 20825
rect 6276 20816 6328 20868
rect 9864 20816 9916 20868
rect 10968 20816 11020 20868
rect 4436 20748 4488 20800
rect 9680 20791 9732 20800
rect 9680 20757 9689 20791
rect 9689 20757 9723 20791
rect 9723 20757 9732 20791
rect 9680 20748 9732 20757
rect 12164 20893 12173 20927
rect 12173 20893 12207 20927
rect 12207 20893 12216 20927
rect 12164 20884 12216 20893
rect 15016 20884 15068 20936
rect 15476 20884 15528 20936
rect 18880 21020 18932 21072
rect 19064 21063 19116 21072
rect 19064 21029 19073 21063
rect 19073 21029 19107 21063
rect 19107 21029 19116 21063
rect 19064 21020 19116 21029
rect 19616 20952 19668 21004
rect 20904 21020 20956 21072
rect 20536 20952 20588 21004
rect 12532 20816 12584 20868
rect 14372 20816 14424 20868
rect 15292 20816 15344 20868
rect 13636 20748 13688 20800
rect 14096 20748 14148 20800
rect 15200 20748 15252 20800
rect 20168 20816 20220 20868
rect 20628 20816 20680 20868
rect 21640 20884 21692 20936
rect 23296 21088 23348 21140
rect 22836 20927 22888 20936
rect 22836 20893 22870 20927
rect 22870 20893 22888 20927
rect 21732 20816 21784 20868
rect 22836 20884 22888 20893
rect 19616 20791 19668 20800
rect 19616 20757 19625 20791
rect 19625 20757 19659 20791
rect 19659 20757 19668 20791
rect 19616 20748 19668 20757
rect 21364 20748 21416 20800
rect 9322 20646 9374 20698
rect 9386 20646 9438 20698
rect 9450 20646 9502 20698
rect 9514 20646 9566 20698
rect 9578 20646 9630 20698
rect 17694 20646 17746 20698
rect 17758 20646 17810 20698
rect 17822 20646 17874 20698
rect 17886 20646 17938 20698
rect 17950 20646 18002 20698
rect 2504 20587 2556 20596
rect 2504 20553 2513 20587
rect 2513 20553 2547 20587
rect 2547 20553 2556 20587
rect 2504 20544 2556 20553
rect 4344 20587 4396 20596
rect 2964 20476 3016 20528
rect 4068 20476 4120 20528
rect 4344 20553 4353 20587
rect 4353 20553 4387 20587
rect 4387 20553 4396 20587
rect 4344 20544 4396 20553
rect 4528 20544 4580 20596
rect 6092 20544 6144 20596
rect 6368 20544 6420 20596
rect 8576 20544 8628 20596
rect 8852 20544 8904 20596
rect 9956 20544 10008 20596
rect 10416 20544 10468 20596
rect 10600 20587 10652 20596
rect 10600 20553 10609 20587
rect 10609 20553 10643 20587
rect 10643 20553 10652 20587
rect 10600 20544 10652 20553
rect 13268 20544 13320 20596
rect 13636 20587 13688 20596
rect 13636 20553 13645 20587
rect 13645 20553 13679 20587
rect 13679 20553 13688 20587
rect 13636 20544 13688 20553
rect 3056 20451 3108 20460
rect 3056 20417 3065 20451
rect 3065 20417 3099 20451
rect 3099 20417 3108 20451
rect 3056 20408 3108 20417
rect 3516 20451 3568 20460
rect 3516 20417 3525 20451
rect 3525 20417 3559 20451
rect 3559 20417 3568 20451
rect 3516 20408 3568 20417
rect 3976 20451 4028 20460
rect 3976 20417 3985 20451
rect 3985 20417 4019 20451
rect 4019 20417 4028 20451
rect 3976 20408 4028 20417
rect 4252 20408 4304 20460
rect 4804 20451 4856 20460
rect 3608 20383 3660 20392
rect 3608 20349 3617 20383
rect 3617 20349 3651 20383
rect 3651 20349 3660 20383
rect 3608 20340 3660 20349
rect 4344 20340 4396 20392
rect 4436 20340 4488 20392
rect 4804 20417 4813 20451
rect 4813 20417 4847 20451
rect 4847 20417 4856 20451
rect 4804 20408 4856 20417
rect 5264 20408 5316 20460
rect 5448 20451 5500 20460
rect 5448 20417 5457 20451
rect 5457 20417 5491 20451
rect 5491 20417 5500 20451
rect 5448 20408 5500 20417
rect 5632 20451 5684 20460
rect 5632 20417 5640 20451
rect 5640 20417 5674 20451
rect 5674 20417 5684 20451
rect 5632 20408 5684 20417
rect 6000 20451 6052 20460
rect 6000 20417 6009 20451
rect 6009 20417 6043 20451
rect 6043 20417 6052 20451
rect 6000 20408 6052 20417
rect 6276 20476 6328 20528
rect 6644 20476 6696 20528
rect 6552 20451 6604 20460
rect 6552 20417 6561 20451
rect 6561 20417 6595 20451
rect 6595 20417 6604 20451
rect 6552 20408 6604 20417
rect 7104 20451 7156 20460
rect 6736 20383 6788 20392
rect 6736 20349 6745 20383
rect 6745 20349 6779 20383
rect 6779 20349 6788 20383
rect 6736 20340 6788 20349
rect 7104 20417 7113 20451
rect 7113 20417 7147 20451
rect 7147 20417 7156 20451
rect 7104 20408 7156 20417
rect 9220 20476 9272 20528
rect 14372 20544 14424 20596
rect 15292 20587 15344 20596
rect 15292 20553 15301 20587
rect 15301 20553 15335 20587
rect 15335 20553 15344 20587
rect 15292 20544 15344 20553
rect 15384 20544 15436 20596
rect 16120 20587 16172 20596
rect 8392 20340 8444 20392
rect 5540 20204 5592 20256
rect 7104 20272 7156 20324
rect 7288 20272 7340 20324
rect 9680 20408 9732 20460
rect 9864 20408 9916 20460
rect 10508 20408 10560 20460
rect 9128 20340 9180 20392
rect 10232 20340 10284 20392
rect 11428 20340 11480 20392
rect 12532 20451 12584 20460
rect 12532 20417 12566 20451
rect 12566 20417 12584 20451
rect 12532 20408 12584 20417
rect 12900 20408 12952 20460
rect 14096 20451 14148 20460
rect 14096 20417 14105 20451
rect 14105 20417 14139 20451
rect 14139 20417 14148 20451
rect 14096 20408 14148 20417
rect 14188 20383 14240 20392
rect 14188 20349 14197 20383
rect 14197 20349 14231 20383
rect 14231 20349 14240 20383
rect 14188 20340 14240 20349
rect 9680 20272 9732 20324
rect 10600 20272 10652 20324
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 14832 20451 14884 20460
rect 14832 20417 14840 20451
rect 14840 20417 14874 20451
rect 14874 20417 14884 20451
rect 15200 20451 15252 20460
rect 14832 20408 14884 20417
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 16120 20553 16129 20587
rect 16129 20553 16163 20587
rect 16163 20553 16172 20587
rect 16120 20544 16172 20553
rect 18880 20544 18932 20596
rect 19708 20519 19760 20528
rect 19708 20485 19717 20519
rect 19717 20485 19751 20519
rect 19751 20485 19760 20519
rect 19708 20476 19760 20485
rect 20076 20544 20128 20596
rect 20536 20544 20588 20596
rect 20904 20587 20956 20596
rect 16028 20451 16080 20460
rect 15292 20340 15344 20392
rect 6552 20204 6604 20256
rect 9956 20204 10008 20256
rect 10324 20247 10376 20256
rect 10324 20213 10333 20247
rect 10333 20213 10367 20247
rect 10367 20213 10376 20247
rect 10324 20204 10376 20213
rect 11888 20204 11940 20256
rect 12164 20204 12216 20256
rect 15200 20272 15252 20324
rect 16028 20417 16037 20451
rect 16037 20417 16071 20451
rect 16071 20417 16080 20451
rect 16028 20408 16080 20417
rect 20260 20408 20312 20460
rect 15752 20383 15804 20392
rect 15752 20349 15761 20383
rect 15761 20349 15795 20383
rect 15795 20349 15804 20383
rect 15752 20340 15804 20349
rect 20904 20553 20913 20587
rect 20913 20553 20947 20587
rect 20947 20553 20956 20587
rect 20904 20544 20956 20553
rect 21456 20544 21508 20596
rect 22928 20544 22980 20596
rect 23204 20519 23256 20528
rect 23204 20485 23213 20519
rect 23213 20485 23247 20519
rect 23247 20485 23256 20519
rect 23204 20476 23256 20485
rect 23296 20476 23348 20528
rect 23480 20476 23532 20528
rect 21272 20451 21324 20460
rect 21272 20417 21281 20451
rect 21281 20417 21315 20451
rect 21315 20417 21324 20451
rect 21272 20408 21324 20417
rect 22376 20408 22428 20460
rect 22744 20383 22796 20392
rect 22744 20349 22753 20383
rect 22753 20349 22787 20383
rect 22787 20349 22796 20383
rect 22744 20340 22796 20349
rect 14924 20204 14976 20256
rect 17316 20272 17368 20324
rect 22284 20204 22336 20256
rect 5136 20102 5188 20154
rect 5200 20102 5252 20154
rect 5264 20102 5316 20154
rect 5328 20102 5380 20154
rect 5392 20102 5444 20154
rect 13508 20102 13560 20154
rect 13572 20102 13624 20154
rect 13636 20102 13688 20154
rect 13700 20102 13752 20154
rect 13764 20102 13816 20154
rect 21880 20102 21932 20154
rect 21944 20102 21996 20154
rect 22008 20102 22060 20154
rect 22072 20102 22124 20154
rect 22136 20102 22188 20154
rect 3608 20000 3660 20052
rect 6460 20000 6512 20052
rect 7104 20000 7156 20052
rect 3516 19932 3568 19984
rect 3976 19932 4028 19984
rect 4436 19864 4488 19916
rect 3424 19796 3476 19848
rect 3700 19796 3752 19848
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 4344 19796 4396 19848
rect 2136 19728 2188 19780
rect 6828 19907 6880 19916
rect 6828 19873 6837 19907
rect 6837 19873 6871 19907
rect 6871 19873 6880 19907
rect 6828 19864 6880 19873
rect 7840 19864 7892 19916
rect 6552 19839 6604 19848
rect 9128 20000 9180 20052
rect 9680 20043 9732 20052
rect 8944 19975 8996 19984
rect 8944 19941 8953 19975
rect 8953 19941 8987 19975
rect 8987 19941 8996 19975
rect 8944 19932 8996 19941
rect 9680 20009 9689 20043
rect 9689 20009 9723 20043
rect 9723 20009 9732 20043
rect 9680 20000 9732 20009
rect 10692 20043 10744 20052
rect 10692 20009 10701 20043
rect 10701 20009 10735 20043
rect 10735 20009 10744 20043
rect 10692 20000 10744 20009
rect 11704 20000 11756 20052
rect 14832 20000 14884 20052
rect 6552 19805 6570 19839
rect 6570 19805 6604 19839
rect 6552 19796 6604 19805
rect 3792 19660 3844 19712
rect 7288 19728 7340 19780
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 9036 19796 9088 19848
rect 9772 19839 9824 19848
rect 8852 19728 8904 19780
rect 9220 19728 9272 19780
rect 9772 19805 9781 19839
rect 9781 19805 9815 19839
rect 9815 19805 9824 19839
rect 9772 19796 9824 19805
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 11796 19839 11848 19848
rect 11796 19805 11805 19839
rect 11805 19805 11839 19839
rect 11839 19805 11848 19839
rect 11796 19796 11848 19805
rect 14096 19864 14148 19916
rect 15200 20000 15252 20052
rect 15752 20000 15804 20052
rect 22376 20043 22428 20052
rect 22376 20009 22385 20043
rect 22385 20009 22419 20043
rect 22419 20009 22428 20043
rect 22376 20000 22428 20009
rect 22284 19932 22336 19984
rect 12992 19796 13044 19848
rect 15292 19864 15344 19916
rect 15476 19907 15528 19916
rect 15476 19873 15485 19907
rect 15485 19873 15519 19907
rect 15519 19873 15528 19907
rect 15476 19864 15528 19873
rect 16672 19864 16724 19916
rect 20168 19864 20220 19916
rect 22376 19864 22428 19916
rect 15200 19839 15252 19848
rect 7472 19703 7524 19712
rect 7472 19669 7481 19703
rect 7481 19669 7515 19703
rect 7515 19669 7524 19703
rect 7472 19660 7524 19669
rect 8668 19660 8720 19712
rect 10324 19660 10376 19712
rect 12164 19728 12216 19780
rect 14004 19728 14056 19780
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 14924 19728 14976 19780
rect 16764 19728 16816 19780
rect 12624 19660 12676 19712
rect 13268 19660 13320 19712
rect 16672 19660 16724 19712
rect 16856 19703 16908 19712
rect 16856 19669 16865 19703
rect 16865 19669 16899 19703
rect 16899 19669 16908 19703
rect 16856 19660 16908 19669
rect 17040 19703 17092 19712
rect 17040 19669 17049 19703
rect 17049 19669 17083 19703
rect 17083 19669 17092 19703
rect 17040 19660 17092 19669
rect 17408 19703 17460 19712
rect 17408 19669 17417 19703
rect 17417 19669 17451 19703
rect 17451 19669 17460 19703
rect 17408 19660 17460 19669
rect 18052 19703 18104 19712
rect 18052 19669 18061 19703
rect 18061 19669 18095 19703
rect 18095 19669 18104 19703
rect 18052 19660 18104 19669
rect 18420 19703 18472 19712
rect 18420 19669 18429 19703
rect 18429 19669 18463 19703
rect 18463 19669 18472 19703
rect 18420 19660 18472 19669
rect 22468 19660 22520 19712
rect 22560 19660 22612 19712
rect 22836 19703 22888 19712
rect 22836 19669 22845 19703
rect 22845 19669 22879 19703
rect 22879 19669 22888 19703
rect 25044 19703 25096 19712
rect 22836 19660 22888 19669
rect 25044 19669 25053 19703
rect 25053 19669 25087 19703
rect 25087 19669 25096 19703
rect 25044 19660 25096 19669
rect 9322 19558 9374 19610
rect 9386 19558 9438 19610
rect 9450 19558 9502 19610
rect 9514 19558 9566 19610
rect 9578 19558 9630 19610
rect 17694 19558 17746 19610
rect 17758 19558 17810 19610
rect 17822 19558 17874 19610
rect 17886 19558 17938 19610
rect 17950 19558 18002 19610
rect 4344 19499 4396 19508
rect 4344 19465 4353 19499
rect 4353 19465 4387 19499
rect 4387 19465 4396 19499
rect 4344 19456 4396 19465
rect 4528 19499 4580 19508
rect 4528 19465 4537 19499
rect 4537 19465 4571 19499
rect 4571 19465 4580 19499
rect 4528 19456 4580 19465
rect 7104 19456 7156 19508
rect 12164 19499 12216 19508
rect 2964 19363 3016 19372
rect 2964 19329 2973 19363
rect 2973 19329 3007 19363
rect 3007 19329 3016 19363
rect 2964 19320 3016 19329
rect 3240 19320 3292 19372
rect 3976 19363 4028 19372
rect 3976 19329 3985 19363
rect 3985 19329 4019 19363
rect 4019 19329 4028 19363
rect 3976 19320 4028 19329
rect 6736 19363 6788 19372
rect 6736 19329 6745 19363
rect 6745 19329 6779 19363
rect 6779 19329 6788 19363
rect 6736 19320 6788 19329
rect 6920 19363 6972 19372
rect 6920 19329 6930 19363
rect 6930 19329 6964 19363
rect 6964 19329 6972 19363
rect 6920 19320 6972 19329
rect 7288 19320 7340 19372
rect 8392 19388 8444 19440
rect 8944 19388 8996 19440
rect 8668 19363 8720 19372
rect 4528 19252 4580 19304
rect 4712 19295 4764 19304
rect 4712 19261 4721 19295
rect 4721 19261 4755 19295
rect 4755 19261 4764 19295
rect 4712 19252 4764 19261
rect 6644 19252 6696 19304
rect 4068 19184 4120 19236
rect 7380 19252 7432 19304
rect 8668 19329 8677 19363
rect 8677 19329 8711 19363
rect 8711 19329 8720 19363
rect 8668 19320 8720 19329
rect 10232 19320 10284 19372
rect 12164 19465 12173 19499
rect 12173 19465 12207 19499
rect 12207 19465 12216 19499
rect 12164 19456 12216 19465
rect 12624 19499 12676 19508
rect 12624 19465 12633 19499
rect 12633 19465 12667 19499
rect 12667 19465 12676 19499
rect 12624 19456 12676 19465
rect 14648 19456 14700 19508
rect 15200 19456 15252 19508
rect 16856 19456 16908 19508
rect 18236 19456 18288 19508
rect 18604 19456 18656 19508
rect 19340 19456 19392 19508
rect 20352 19499 20404 19508
rect 20352 19465 20361 19499
rect 20361 19465 20395 19499
rect 20395 19465 20404 19499
rect 20352 19456 20404 19465
rect 22376 19456 22428 19508
rect 22560 19499 22612 19508
rect 22560 19465 22569 19499
rect 22569 19465 22603 19499
rect 22603 19465 22612 19499
rect 22560 19456 22612 19465
rect 11428 19320 11480 19372
rect 11704 19363 11756 19372
rect 11704 19329 11712 19363
rect 11712 19329 11746 19363
rect 11746 19329 11756 19363
rect 11704 19320 11756 19329
rect 12440 19388 12492 19440
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 8944 19252 8996 19304
rect 9128 19295 9180 19304
rect 9128 19261 9137 19295
rect 9137 19261 9171 19295
rect 9171 19261 9180 19295
rect 9128 19252 9180 19261
rect 11888 19295 11940 19304
rect 11888 19261 11897 19295
rect 11897 19261 11931 19295
rect 11931 19261 11940 19295
rect 11888 19252 11940 19261
rect 2780 19159 2832 19168
rect 2780 19125 2789 19159
rect 2789 19125 2823 19159
rect 2823 19125 2832 19159
rect 2780 19116 2832 19125
rect 7840 19116 7892 19168
rect 8668 19116 8720 19168
rect 8852 19116 8904 19168
rect 12164 19184 12216 19236
rect 12624 19320 12676 19372
rect 14004 19363 14056 19372
rect 14004 19329 14013 19363
rect 14013 19329 14047 19363
rect 14047 19329 14056 19363
rect 14004 19320 14056 19329
rect 15752 19388 15804 19440
rect 17960 19388 18012 19440
rect 23112 19388 23164 19440
rect 14188 19363 14240 19372
rect 14188 19329 14196 19363
rect 14196 19329 14230 19363
rect 14230 19329 14240 19363
rect 14188 19320 14240 19329
rect 14464 19320 14516 19372
rect 16672 19320 16724 19372
rect 18236 19320 18288 19372
rect 22468 19320 22520 19372
rect 22836 19320 22888 19372
rect 15292 19252 15344 19304
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 23296 19252 23348 19304
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 12440 19116 12492 19168
rect 12900 19116 12952 19168
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 14832 19116 14884 19168
rect 25044 19184 25096 19236
rect 22376 19116 22428 19168
rect 23204 19116 23256 19168
rect 5136 19014 5188 19066
rect 5200 19014 5252 19066
rect 5264 19014 5316 19066
rect 5328 19014 5380 19066
rect 5392 19014 5444 19066
rect 13508 19014 13560 19066
rect 13572 19014 13624 19066
rect 13636 19014 13688 19066
rect 13700 19014 13752 19066
rect 13764 19014 13816 19066
rect 21880 19014 21932 19066
rect 21944 19014 21996 19066
rect 22008 19014 22060 19066
rect 22072 19014 22124 19066
rect 22136 19014 22188 19066
rect 3976 18912 4028 18964
rect 6736 18912 6788 18964
rect 7748 18912 7800 18964
rect 8852 18912 8904 18964
rect 10232 18955 10284 18964
rect 10232 18921 10241 18955
rect 10241 18921 10275 18955
rect 10275 18921 10284 18955
rect 10232 18912 10284 18921
rect 12072 18912 12124 18964
rect 15292 18912 15344 18964
rect 15752 18912 15804 18964
rect 17132 18912 17184 18964
rect 17868 18912 17920 18964
rect 7196 18844 7248 18896
rect 8392 18844 8444 18896
rect 6920 18819 6972 18828
rect 6920 18785 6929 18819
rect 6929 18785 6963 18819
rect 6963 18785 6972 18819
rect 6920 18776 6972 18785
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 4712 18708 4764 18760
rect 6552 18708 6604 18760
rect 7012 18708 7064 18760
rect 7380 18708 7432 18760
rect 7656 18708 7708 18760
rect 8024 18708 8076 18760
rect 8392 18751 8444 18760
rect 8392 18717 8401 18751
rect 8401 18717 8435 18751
rect 8435 18717 8444 18751
rect 8392 18708 8444 18717
rect 8944 18751 8996 18760
rect 3424 18640 3476 18692
rect 2504 18572 2556 18624
rect 8668 18640 8720 18692
rect 8944 18717 8953 18751
rect 8953 18717 8987 18751
rect 8987 18717 8996 18751
rect 8944 18708 8996 18717
rect 9220 18751 9272 18760
rect 9220 18717 9229 18751
rect 9229 18717 9263 18751
rect 9263 18717 9272 18751
rect 9220 18708 9272 18717
rect 8852 18640 8904 18692
rect 9680 18844 9732 18896
rect 18512 18912 18564 18964
rect 10232 18776 10284 18828
rect 10784 18819 10836 18828
rect 10784 18785 10793 18819
rect 10793 18785 10827 18819
rect 10827 18785 10836 18819
rect 10784 18776 10836 18785
rect 11704 18776 11756 18828
rect 11888 18776 11940 18828
rect 14188 18776 14240 18828
rect 9772 18708 9824 18760
rect 10140 18708 10192 18760
rect 12532 18751 12584 18760
rect 7380 18615 7432 18624
rect 7380 18581 7389 18615
rect 7389 18581 7423 18615
rect 7423 18581 7432 18615
rect 7380 18572 7432 18581
rect 9956 18615 10008 18624
rect 9956 18581 9965 18615
rect 9965 18581 9999 18615
rect 9999 18581 10008 18615
rect 9956 18572 10008 18581
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 12900 18751 12952 18760
rect 12900 18717 12910 18751
rect 12910 18717 12944 18751
rect 12944 18717 12952 18751
rect 12900 18708 12952 18717
rect 13084 18751 13136 18760
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 13084 18708 13136 18717
rect 14096 18708 14148 18760
rect 15844 18751 15896 18760
rect 15844 18717 15853 18751
rect 15853 18717 15887 18751
rect 15887 18717 15896 18751
rect 15844 18708 15896 18717
rect 12348 18640 12400 18692
rect 11060 18572 11112 18624
rect 11612 18572 11664 18624
rect 12440 18615 12492 18624
rect 12440 18581 12449 18615
rect 12449 18581 12483 18615
rect 12483 18581 12492 18615
rect 12992 18640 13044 18692
rect 12440 18572 12492 18581
rect 14464 18572 14516 18624
rect 14648 18640 14700 18692
rect 15660 18640 15712 18692
rect 18144 18776 18196 18828
rect 17040 18708 17092 18760
rect 17316 18708 17368 18760
rect 17592 18751 17644 18760
rect 17592 18717 17600 18751
rect 17600 18717 17634 18751
rect 17634 18717 17644 18751
rect 17960 18751 18012 18760
rect 17592 18708 17644 18717
rect 17960 18717 17969 18751
rect 17969 18717 18003 18751
rect 18003 18717 18012 18751
rect 17960 18708 18012 18717
rect 18880 18844 18932 18896
rect 18144 18640 18196 18692
rect 18512 18751 18564 18760
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 21180 18912 21232 18964
rect 21732 18912 21784 18964
rect 22928 18912 22980 18964
rect 20720 18844 20772 18896
rect 21640 18844 21692 18896
rect 18512 18708 18564 18717
rect 18972 18708 19024 18760
rect 20720 18708 20772 18760
rect 17132 18572 17184 18624
rect 17408 18572 17460 18624
rect 17500 18572 17552 18624
rect 19892 18640 19944 18692
rect 21640 18708 21692 18760
rect 24216 18751 24268 18760
rect 24216 18717 24225 18751
rect 24225 18717 24259 18751
rect 24259 18717 24268 18751
rect 24216 18708 24268 18717
rect 22376 18683 22428 18692
rect 22376 18649 22394 18683
rect 22394 18649 22428 18683
rect 22376 18640 22428 18649
rect 23388 18640 23440 18692
rect 22560 18572 22612 18624
rect 22836 18615 22888 18624
rect 22836 18581 22845 18615
rect 22845 18581 22879 18615
rect 22879 18581 22888 18615
rect 22836 18572 22888 18581
rect 9322 18470 9374 18522
rect 9386 18470 9438 18522
rect 9450 18470 9502 18522
rect 9514 18470 9566 18522
rect 9578 18470 9630 18522
rect 17694 18470 17746 18522
rect 17758 18470 17810 18522
rect 17822 18470 17874 18522
rect 17886 18470 17938 18522
rect 17950 18470 18002 18522
rect 2964 18368 3016 18420
rect 3424 18368 3476 18420
rect 8668 18411 8720 18420
rect 8668 18377 8677 18411
rect 8677 18377 8711 18411
rect 8711 18377 8720 18411
rect 8668 18368 8720 18377
rect 9680 18368 9732 18420
rect 11888 18368 11940 18420
rect 14188 18368 14240 18420
rect 15568 18411 15620 18420
rect 15568 18377 15577 18411
rect 15577 18377 15611 18411
rect 15611 18377 15620 18411
rect 15568 18368 15620 18377
rect 17500 18368 17552 18420
rect 2780 18300 2832 18352
rect 4712 18300 4764 18352
rect 7380 18300 7432 18352
rect 12440 18343 12492 18352
rect 12440 18309 12474 18343
rect 12474 18309 12492 18343
rect 12440 18300 12492 18309
rect 16764 18300 16816 18352
rect 1952 18232 2004 18284
rect 3700 18275 3752 18284
rect 3700 18241 3709 18275
rect 3709 18241 3743 18275
rect 3743 18241 3752 18275
rect 3700 18232 3752 18241
rect 3792 18275 3844 18284
rect 3792 18241 3801 18275
rect 3801 18241 3835 18275
rect 3835 18241 3844 18275
rect 3792 18232 3844 18241
rect 3976 18232 4028 18284
rect 6552 18275 6604 18284
rect 6552 18241 6561 18275
rect 6561 18241 6595 18275
rect 6595 18241 6604 18275
rect 6552 18232 6604 18241
rect 7012 18275 7064 18284
rect 7012 18241 7021 18275
rect 7021 18241 7055 18275
rect 7055 18241 7064 18275
rect 7012 18232 7064 18241
rect 8668 18232 8720 18284
rect 9680 18275 9732 18284
rect 9680 18241 9689 18275
rect 9689 18241 9723 18275
rect 9723 18241 9732 18275
rect 9680 18232 9732 18241
rect 9772 18275 9824 18284
rect 9772 18241 9781 18275
rect 9781 18241 9815 18275
rect 9815 18241 9824 18275
rect 9772 18232 9824 18241
rect 10232 18275 10284 18284
rect 10232 18241 10241 18275
rect 10241 18241 10275 18275
rect 10275 18241 10284 18275
rect 10232 18232 10284 18241
rect 10508 18232 10560 18284
rect 12992 18232 13044 18284
rect 14280 18232 14332 18284
rect 17500 18275 17552 18284
rect 17500 18241 17509 18275
rect 17509 18241 17543 18275
rect 17543 18241 17552 18275
rect 17500 18232 17552 18241
rect 18512 18368 18564 18420
rect 19616 18368 19668 18420
rect 18604 18300 18656 18352
rect 20996 18368 21048 18420
rect 21364 18368 21416 18420
rect 3148 18164 3200 18216
rect 7656 18164 7708 18216
rect 9128 18096 9180 18148
rect 9404 18139 9456 18148
rect 9404 18105 9413 18139
rect 9413 18105 9447 18139
rect 9447 18105 9456 18139
rect 9404 18096 9456 18105
rect 10600 18096 10652 18148
rect 11796 18164 11848 18216
rect 14096 18164 14148 18216
rect 17868 18207 17920 18216
rect 17868 18173 17877 18207
rect 17877 18173 17911 18207
rect 17911 18173 17920 18207
rect 17868 18164 17920 18173
rect 18144 18164 18196 18216
rect 18788 18275 18840 18284
rect 18788 18241 18797 18275
rect 18797 18241 18831 18275
rect 18831 18241 18840 18275
rect 18788 18232 18840 18241
rect 19248 18232 19300 18284
rect 19892 18232 19944 18284
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20168 18232 20220 18241
rect 20352 18232 20404 18284
rect 21088 18232 21140 18284
rect 22284 18232 22336 18284
rect 22560 18368 22612 18420
rect 4436 18028 4488 18080
rect 5816 18028 5868 18080
rect 6736 18071 6788 18080
rect 6736 18037 6745 18071
rect 6745 18037 6779 18071
rect 6779 18037 6788 18071
rect 6736 18028 6788 18037
rect 6828 18071 6880 18080
rect 6828 18037 6837 18071
rect 6837 18037 6871 18071
rect 6871 18037 6880 18071
rect 7656 18071 7708 18080
rect 6828 18028 6880 18037
rect 7656 18037 7665 18071
rect 7665 18037 7699 18071
rect 7699 18037 7708 18071
rect 7656 18028 7708 18037
rect 9312 18028 9364 18080
rect 10324 18028 10376 18080
rect 11704 18028 11756 18080
rect 14004 18096 14056 18148
rect 18236 18139 18288 18148
rect 18236 18105 18245 18139
rect 18245 18105 18279 18139
rect 18279 18105 18288 18139
rect 18236 18096 18288 18105
rect 20904 18164 20956 18216
rect 20996 18164 21048 18216
rect 22744 18300 22796 18352
rect 23388 18300 23440 18352
rect 18604 18139 18656 18148
rect 18604 18105 18613 18139
rect 18613 18105 18647 18139
rect 18647 18105 18656 18139
rect 18604 18096 18656 18105
rect 18788 18096 18840 18148
rect 21732 18096 21784 18148
rect 22192 18096 22244 18148
rect 22836 18232 22888 18284
rect 22744 18207 22796 18216
rect 22744 18173 22753 18207
rect 22753 18173 22787 18207
rect 22787 18173 22796 18207
rect 22744 18164 22796 18173
rect 15108 18028 15160 18080
rect 22836 18096 22888 18148
rect 5136 17926 5188 17978
rect 5200 17926 5252 17978
rect 5264 17926 5316 17978
rect 5328 17926 5380 17978
rect 5392 17926 5444 17978
rect 13508 17926 13560 17978
rect 13572 17926 13624 17978
rect 13636 17926 13688 17978
rect 13700 17926 13752 17978
rect 13764 17926 13816 17978
rect 21880 17926 21932 17978
rect 21944 17926 21996 17978
rect 22008 17926 22060 17978
rect 22072 17926 22124 17978
rect 22136 17926 22188 17978
rect 4528 17824 4580 17876
rect 8392 17824 8444 17876
rect 9956 17867 10008 17876
rect 9956 17833 9965 17867
rect 9965 17833 9999 17867
rect 9999 17833 10008 17867
rect 9956 17824 10008 17833
rect 3332 17731 3384 17740
rect 3332 17697 3341 17731
rect 3341 17697 3375 17731
rect 3375 17697 3384 17731
rect 3332 17688 3384 17697
rect 4344 17688 4396 17740
rect 9404 17756 9456 17808
rect 11796 17824 11848 17876
rect 12256 17824 12308 17876
rect 12716 17824 12768 17876
rect 8300 17688 8352 17740
rect 3148 17663 3200 17672
rect 3148 17629 3157 17663
rect 3157 17629 3191 17663
rect 3191 17629 3200 17663
rect 3148 17620 3200 17629
rect 4160 17620 4212 17672
rect 6368 17620 6420 17672
rect 8760 17620 8812 17672
rect 9312 17663 9364 17672
rect 9312 17629 9321 17663
rect 9321 17629 9355 17663
rect 9355 17629 9364 17663
rect 17592 17824 17644 17876
rect 17868 17824 17920 17876
rect 18144 17824 18196 17876
rect 18420 17824 18472 17876
rect 19248 17824 19300 17876
rect 20168 17867 20220 17876
rect 20168 17833 20177 17867
rect 20177 17833 20211 17867
rect 20211 17833 20220 17867
rect 20168 17824 20220 17833
rect 20260 17824 20312 17876
rect 15384 17756 15436 17808
rect 17408 17756 17460 17808
rect 22376 17824 22428 17876
rect 14096 17731 14148 17740
rect 9312 17620 9364 17629
rect 10600 17663 10652 17672
rect 7932 17595 7984 17604
rect 2872 17527 2924 17536
rect 2872 17493 2881 17527
rect 2881 17493 2915 17527
rect 2915 17493 2924 17527
rect 2872 17484 2924 17493
rect 2964 17484 3016 17536
rect 6092 17484 6144 17536
rect 7932 17561 7950 17595
rect 7950 17561 7984 17595
rect 7932 17552 7984 17561
rect 9036 17552 9088 17604
rect 8116 17484 8168 17536
rect 8944 17484 8996 17536
rect 9680 17552 9732 17604
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 12256 17620 12308 17672
rect 13084 17620 13136 17672
rect 14096 17697 14105 17731
rect 14105 17697 14139 17731
rect 14139 17697 14148 17731
rect 14096 17688 14148 17697
rect 20904 17688 20956 17740
rect 21640 17731 21692 17740
rect 21640 17697 21649 17731
rect 21649 17697 21683 17731
rect 21683 17697 21692 17731
rect 21640 17688 21692 17697
rect 22376 17688 22428 17740
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 16672 17620 16724 17672
rect 9956 17484 10008 17536
rect 11244 17552 11296 17604
rect 12164 17552 12216 17604
rect 13544 17552 13596 17604
rect 18420 17620 18472 17672
rect 19064 17663 19116 17672
rect 19064 17629 19073 17663
rect 19073 17629 19107 17663
rect 19107 17629 19116 17663
rect 19064 17620 19116 17629
rect 21088 17663 21140 17672
rect 18604 17552 18656 17604
rect 11060 17484 11112 17536
rect 12256 17484 12308 17536
rect 12716 17484 12768 17536
rect 21088 17629 21097 17663
rect 21097 17629 21131 17663
rect 21131 17629 21140 17663
rect 21088 17620 21140 17629
rect 21364 17663 21416 17672
rect 21364 17629 21373 17663
rect 21373 17629 21407 17663
rect 21407 17629 21416 17663
rect 21364 17620 21416 17629
rect 21916 17663 21968 17672
rect 21916 17629 21925 17663
rect 21925 17629 21959 17663
rect 21959 17629 21968 17663
rect 21916 17620 21968 17629
rect 22284 17620 22336 17672
rect 23020 17756 23072 17808
rect 24216 17688 24268 17740
rect 22744 17663 22796 17672
rect 22744 17629 22753 17663
rect 22753 17629 22787 17663
rect 22787 17629 22796 17663
rect 22744 17620 22796 17629
rect 22836 17663 22888 17672
rect 22836 17629 22845 17663
rect 22845 17629 22879 17663
rect 22879 17629 22888 17663
rect 22836 17620 22888 17629
rect 20720 17552 20772 17604
rect 20536 17527 20588 17536
rect 20536 17493 20545 17527
rect 20545 17493 20579 17527
rect 20579 17493 20588 17527
rect 20536 17484 20588 17493
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 21180 17484 21232 17536
rect 21916 17484 21968 17536
rect 22284 17484 22336 17536
rect 22376 17527 22428 17536
rect 22376 17493 22385 17527
rect 22385 17493 22419 17527
rect 22419 17493 22428 17527
rect 22376 17484 22428 17493
rect 22836 17484 22888 17536
rect 25780 17527 25832 17536
rect 25780 17493 25789 17527
rect 25789 17493 25823 17527
rect 25823 17493 25832 17527
rect 25780 17484 25832 17493
rect 9322 17382 9374 17434
rect 9386 17382 9438 17434
rect 9450 17382 9502 17434
rect 9514 17382 9566 17434
rect 9578 17382 9630 17434
rect 17694 17382 17746 17434
rect 17758 17382 17810 17434
rect 17822 17382 17874 17434
rect 17886 17382 17938 17434
rect 17950 17382 18002 17434
rect 3700 17280 3752 17332
rect 2872 17212 2924 17264
rect 3148 17212 3200 17264
rect 1952 17144 2004 17196
rect 3516 17144 3568 17196
rect 4344 17119 4396 17128
rect 4344 17085 4353 17119
rect 4353 17085 4387 17119
rect 4387 17085 4396 17119
rect 4344 17076 4396 17085
rect 4436 17076 4488 17128
rect 6184 17280 6236 17332
rect 7932 17255 7984 17264
rect 7932 17221 7941 17255
rect 7941 17221 7975 17255
rect 7975 17221 7984 17255
rect 7932 17212 7984 17221
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 5816 17187 5868 17196
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 6092 17144 6144 17196
rect 6184 17187 6236 17196
rect 6184 17153 6193 17187
rect 6193 17153 6227 17187
rect 6227 17153 6236 17187
rect 6184 17144 6236 17153
rect 6368 17144 6420 17196
rect 6736 17144 6788 17196
rect 4068 17008 4120 17060
rect 6828 17076 6880 17128
rect 8300 17280 8352 17332
rect 8116 17187 8168 17196
rect 8116 17153 8125 17187
rect 8125 17153 8159 17187
rect 8159 17153 8168 17187
rect 8116 17144 8168 17153
rect 9128 17280 9180 17332
rect 11244 17323 11296 17332
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 8668 17144 8720 17153
rect 4160 16940 4212 16992
rect 4804 16940 4856 16992
rect 7932 17008 7984 17060
rect 8760 17076 8812 17128
rect 9496 17212 9548 17264
rect 9404 17187 9456 17196
rect 9404 17153 9413 17187
rect 9413 17153 9447 17187
rect 9447 17153 9456 17187
rect 9956 17212 10008 17264
rect 9404 17144 9456 17153
rect 9128 17119 9180 17128
rect 9128 17085 9137 17119
rect 9137 17085 9171 17119
rect 9171 17085 9180 17119
rect 9128 17076 9180 17085
rect 11244 17289 11253 17323
rect 11253 17289 11287 17323
rect 11287 17289 11296 17323
rect 11244 17280 11296 17289
rect 10508 17144 10560 17196
rect 11060 17187 11112 17196
rect 11060 17153 11069 17187
rect 11069 17153 11103 17187
rect 11103 17153 11112 17187
rect 11060 17144 11112 17153
rect 13084 17144 13136 17196
rect 10140 17076 10192 17128
rect 12716 17076 12768 17128
rect 13268 17076 13320 17128
rect 13544 17144 13596 17196
rect 15568 17280 15620 17332
rect 17224 17280 17276 17332
rect 17592 17280 17644 17332
rect 14280 17212 14332 17264
rect 16948 17212 17000 17264
rect 18604 17280 18656 17332
rect 20720 17280 20772 17332
rect 21180 17323 21232 17332
rect 21180 17289 21189 17323
rect 21189 17289 21223 17323
rect 21223 17289 21232 17323
rect 21180 17280 21232 17289
rect 21272 17280 21324 17332
rect 22652 17323 22704 17332
rect 22652 17289 22661 17323
rect 22661 17289 22695 17323
rect 22695 17289 22704 17323
rect 22652 17280 22704 17289
rect 13912 17144 13964 17196
rect 9680 17008 9732 17060
rect 12348 17008 12400 17060
rect 14096 17076 14148 17128
rect 17500 17076 17552 17128
rect 17776 17144 17828 17196
rect 18144 17144 18196 17196
rect 17960 17119 18012 17128
rect 17960 17085 17969 17119
rect 17969 17085 18003 17119
rect 18003 17085 18012 17119
rect 17960 17076 18012 17085
rect 14372 17008 14424 17060
rect 17408 17008 17460 17060
rect 18512 17144 18564 17196
rect 20996 17212 21048 17264
rect 22284 17212 22336 17264
rect 23204 17212 23256 17264
rect 20720 17187 20772 17196
rect 20720 17153 20729 17187
rect 20729 17153 20763 17187
rect 20763 17153 20772 17187
rect 20720 17144 20772 17153
rect 23020 17187 23072 17196
rect 23020 17153 23029 17187
rect 23029 17153 23063 17187
rect 23063 17153 23072 17187
rect 23020 17144 23072 17153
rect 18880 17076 18932 17128
rect 20260 17076 20312 17128
rect 21548 17076 21600 17128
rect 22376 17076 22428 17128
rect 23112 17076 23164 17128
rect 20996 17008 21048 17060
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 10324 16940 10376 16949
rect 12992 16983 13044 16992
rect 12992 16949 13001 16983
rect 13001 16949 13035 16983
rect 13035 16949 13044 16983
rect 12992 16940 13044 16949
rect 13912 16940 13964 16992
rect 17224 16940 17276 16992
rect 17776 16940 17828 16992
rect 18880 16940 18932 16992
rect 5136 16838 5188 16890
rect 5200 16838 5252 16890
rect 5264 16838 5316 16890
rect 5328 16838 5380 16890
rect 5392 16838 5444 16890
rect 13508 16838 13560 16890
rect 13572 16838 13624 16890
rect 13636 16838 13688 16890
rect 13700 16838 13752 16890
rect 13764 16838 13816 16890
rect 21880 16838 21932 16890
rect 21944 16838 21996 16890
rect 22008 16838 22060 16890
rect 22072 16838 22124 16890
rect 22136 16838 22188 16890
rect 3516 16779 3568 16788
rect 3516 16745 3525 16779
rect 3525 16745 3559 16779
rect 3559 16745 3568 16779
rect 3516 16736 3568 16745
rect 2136 16643 2188 16652
rect 2136 16609 2145 16643
rect 2145 16609 2179 16643
rect 2179 16609 2188 16643
rect 2136 16600 2188 16609
rect 6552 16736 6604 16788
rect 6828 16736 6880 16788
rect 7932 16736 7984 16788
rect 8668 16736 8720 16788
rect 8760 16779 8812 16788
rect 8760 16745 8769 16779
rect 8769 16745 8803 16779
rect 8803 16745 8812 16779
rect 8760 16736 8812 16745
rect 9312 16736 9364 16788
rect 11520 16736 11572 16788
rect 11888 16736 11940 16788
rect 12900 16736 12952 16788
rect 13268 16736 13320 16788
rect 16212 16736 16264 16788
rect 17040 16736 17092 16788
rect 20904 16779 20956 16788
rect 4344 16668 4396 16720
rect 4712 16600 4764 16652
rect 8300 16600 8352 16652
rect 15568 16668 15620 16720
rect 16580 16711 16632 16720
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 8024 16532 8076 16584
rect 8208 16575 8260 16584
rect 8208 16541 8217 16575
rect 8217 16541 8251 16575
rect 8251 16541 8260 16575
rect 8208 16532 8260 16541
rect 15476 16600 15528 16652
rect 16580 16677 16589 16711
rect 16589 16677 16623 16711
rect 16623 16677 16632 16711
rect 16580 16668 16632 16677
rect 20904 16745 20913 16779
rect 20913 16745 20947 16779
rect 20947 16745 20956 16779
rect 20904 16736 20956 16745
rect 22376 16736 22428 16788
rect 18512 16668 18564 16720
rect 19064 16668 19116 16720
rect 23112 16736 23164 16788
rect 23296 16736 23348 16788
rect 4804 16464 4856 16516
rect 6276 16464 6328 16516
rect 7288 16464 7340 16516
rect 3792 16439 3844 16448
rect 3792 16405 3801 16439
rect 3801 16405 3835 16439
rect 3835 16405 3844 16439
rect 3792 16396 3844 16405
rect 6368 16396 6420 16448
rect 9220 16396 9272 16448
rect 9496 16464 9548 16516
rect 9772 16464 9824 16516
rect 10600 16532 10652 16584
rect 12256 16464 12308 16516
rect 15752 16532 15804 16584
rect 16212 16575 16264 16584
rect 15292 16464 15344 16516
rect 16212 16541 16221 16575
rect 16221 16541 16255 16575
rect 16255 16541 16264 16575
rect 16212 16532 16264 16541
rect 16396 16575 16448 16584
rect 16396 16541 16405 16575
rect 16405 16541 16439 16575
rect 16439 16541 16448 16575
rect 16396 16532 16448 16541
rect 16856 16575 16908 16584
rect 16856 16541 16864 16575
rect 16864 16541 16898 16575
rect 16898 16541 16908 16575
rect 16856 16532 16908 16541
rect 17040 16575 17092 16584
rect 17040 16541 17049 16575
rect 17049 16541 17083 16575
rect 17083 16541 17092 16575
rect 17040 16532 17092 16541
rect 17224 16575 17276 16584
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 17592 16532 17644 16584
rect 22836 16668 22888 16720
rect 22744 16600 22796 16652
rect 19892 16532 19944 16584
rect 20628 16532 20680 16584
rect 21364 16532 21416 16584
rect 22836 16575 22888 16584
rect 22836 16541 22845 16575
rect 22845 16541 22879 16575
rect 22879 16541 22888 16575
rect 22836 16532 22888 16541
rect 23388 16575 23440 16584
rect 10600 16396 10652 16448
rect 11704 16396 11756 16448
rect 12808 16396 12860 16448
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 13268 16396 13320 16448
rect 15476 16439 15528 16448
rect 15476 16405 15485 16439
rect 15485 16405 15519 16439
rect 15519 16405 15528 16439
rect 15476 16396 15528 16405
rect 15936 16396 15988 16448
rect 16764 16396 16816 16448
rect 17224 16396 17276 16448
rect 18328 16439 18380 16448
rect 18328 16405 18337 16439
rect 18337 16405 18371 16439
rect 18371 16405 18380 16439
rect 18328 16396 18380 16405
rect 18420 16396 18472 16448
rect 18788 16439 18840 16448
rect 18788 16405 18797 16439
rect 18797 16405 18831 16439
rect 18831 16405 18840 16439
rect 20720 16464 20772 16516
rect 23388 16541 23397 16575
rect 23397 16541 23431 16575
rect 23431 16541 23440 16575
rect 23388 16532 23440 16541
rect 23296 16464 23348 16516
rect 24124 16464 24176 16516
rect 18788 16396 18840 16405
rect 21272 16439 21324 16448
rect 21272 16405 21281 16439
rect 21281 16405 21315 16439
rect 21315 16405 21324 16439
rect 21272 16396 21324 16405
rect 21548 16396 21600 16448
rect 22284 16396 22336 16448
rect 9322 16294 9374 16346
rect 9386 16294 9438 16346
rect 9450 16294 9502 16346
rect 9514 16294 9566 16346
rect 9578 16294 9630 16346
rect 17694 16294 17746 16346
rect 17758 16294 17810 16346
rect 17822 16294 17874 16346
rect 17886 16294 17938 16346
rect 17950 16294 18002 16346
rect 2136 16192 2188 16244
rect 3424 16192 3476 16244
rect 4988 16192 5040 16244
rect 6276 16192 6328 16244
rect 7288 16235 7340 16244
rect 7288 16201 7297 16235
rect 7297 16201 7331 16235
rect 7331 16201 7340 16235
rect 7288 16192 7340 16201
rect 7380 16192 7432 16244
rect 7748 16192 7800 16244
rect 6368 16124 6420 16176
rect 2872 16056 2924 16108
rect 4344 16099 4396 16108
rect 4344 16065 4353 16099
rect 4353 16065 4387 16099
rect 4387 16065 4396 16099
rect 4344 16056 4396 16065
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 6828 16099 6880 16108
rect 6828 16065 6837 16099
rect 6837 16065 6871 16099
rect 6871 16065 6880 16099
rect 6828 16056 6880 16065
rect 6920 16099 6972 16108
rect 6920 16065 6930 16099
rect 6930 16065 6964 16099
rect 6964 16065 6972 16099
rect 6920 16056 6972 16065
rect 7288 16056 7340 16108
rect 5816 15988 5868 16040
rect 8300 16099 8352 16108
rect 8300 16065 8309 16099
rect 8309 16065 8343 16099
rect 8343 16065 8352 16099
rect 8300 16056 8352 16065
rect 8668 16056 8720 16108
rect 9128 16099 9180 16108
rect 8576 15988 8628 16040
rect 9128 16065 9136 16099
rect 9136 16065 9170 16099
rect 9170 16065 9180 16099
rect 9128 16056 9180 16065
rect 10140 16192 10192 16244
rect 9588 16124 9640 16176
rect 9772 16099 9824 16108
rect 9220 16031 9272 16040
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 9772 16065 9781 16099
rect 9781 16065 9815 16099
rect 9815 16065 9824 16099
rect 9772 16056 9824 16065
rect 10324 16124 10376 16176
rect 12624 16192 12676 16244
rect 14372 16235 14424 16244
rect 14372 16201 14381 16235
rect 14381 16201 14415 16235
rect 14415 16201 14424 16235
rect 14372 16192 14424 16201
rect 16212 16192 16264 16244
rect 16396 16192 16448 16244
rect 18236 16192 18288 16244
rect 18420 16235 18472 16244
rect 18420 16201 18429 16235
rect 18429 16201 18463 16235
rect 18463 16201 18472 16235
rect 18420 16192 18472 16201
rect 18880 16235 18932 16244
rect 18880 16201 18889 16235
rect 18889 16201 18923 16235
rect 18923 16201 18932 16235
rect 18880 16192 18932 16201
rect 20260 16192 20312 16244
rect 10784 16056 10836 16108
rect 9588 15988 9640 16040
rect 8760 15920 8812 15972
rect 9496 15920 9548 15972
rect 6920 15852 6972 15904
rect 8024 15895 8076 15904
rect 8024 15861 8033 15895
rect 8033 15861 8067 15895
rect 8067 15861 8076 15895
rect 8024 15852 8076 15861
rect 8208 15852 8260 15904
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 12164 16056 12216 16108
rect 12808 16031 12860 16040
rect 12808 15997 12817 16031
rect 12817 15997 12851 16031
rect 12851 15997 12860 16031
rect 12808 15988 12860 15997
rect 14188 16056 14240 16108
rect 14280 16056 14332 16108
rect 13360 15988 13412 16040
rect 14372 15988 14424 16040
rect 15200 15988 15252 16040
rect 15568 16099 15620 16108
rect 15568 16065 15577 16099
rect 15577 16065 15611 16099
rect 15611 16065 15620 16099
rect 15568 16056 15620 16065
rect 15936 16056 15988 16108
rect 16580 16124 16632 16176
rect 19064 16124 19116 16176
rect 16672 16099 16724 16108
rect 16212 15988 16264 16040
rect 16672 16065 16681 16099
rect 16681 16065 16715 16099
rect 16715 16065 16724 16099
rect 16672 16056 16724 16065
rect 18604 16056 18656 16108
rect 18788 16099 18840 16108
rect 18788 16065 18797 16099
rect 18797 16065 18831 16099
rect 18831 16065 18840 16099
rect 18788 16056 18840 16065
rect 19340 16056 19392 16108
rect 19892 16099 19944 16108
rect 19892 16065 19901 16099
rect 19901 16065 19935 16099
rect 19935 16065 19944 16099
rect 19892 16056 19944 16065
rect 16580 15988 16632 16040
rect 13176 15920 13228 15972
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 12900 15852 12952 15904
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 15936 15895 15988 15904
rect 15936 15861 15945 15895
rect 15945 15861 15979 15895
rect 15979 15861 15988 15895
rect 15936 15852 15988 15861
rect 18788 15920 18840 15972
rect 18144 15852 18196 15904
rect 20628 16056 20680 16108
rect 20352 16031 20404 16040
rect 20352 15997 20361 16031
rect 20361 15997 20395 16031
rect 20395 15997 20404 16031
rect 20352 15988 20404 15997
rect 20076 15920 20128 15972
rect 20536 15920 20588 15972
rect 21732 16056 21784 16108
rect 21456 15988 21508 16040
rect 22376 16099 22428 16108
rect 22376 16065 22410 16099
rect 22410 16065 22428 16099
rect 24216 16192 24268 16244
rect 24124 16124 24176 16176
rect 22376 16056 22428 16065
rect 23388 15920 23440 15972
rect 21088 15852 21140 15904
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 23480 15895 23532 15904
rect 23480 15861 23489 15895
rect 23489 15861 23523 15895
rect 23523 15861 23532 15895
rect 23480 15852 23532 15861
rect 5136 15750 5188 15802
rect 5200 15750 5252 15802
rect 5264 15750 5316 15802
rect 5328 15750 5380 15802
rect 5392 15750 5444 15802
rect 13508 15750 13560 15802
rect 13572 15750 13624 15802
rect 13636 15750 13688 15802
rect 13700 15750 13752 15802
rect 13764 15750 13816 15802
rect 21880 15750 21932 15802
rect 21944 15750 21996 15802
rect 22008 15750 22060 15802
rect 22072 15750 22124 15802
rect 22136 15750 22188 15802
rect 2872 15691 2924 15700
rect 2872 15657 2881 15691
rect 2881 15657 2915 15691
rect 2915 15657 2924 15691
rect 2872 15648 2924 15657
rect 3332 15691 3384 15700
rect 3332 15657 3341 15691
rect 3341 15657 3375 15691
rect 3375 15657 3384 15691
rect 3332 15648 3384 15657
rect 7196 15648 7248 15700
rect 7748 15691 7800 15700
rect 7748 15657 7757 15691
rect 7757 15657 7791 15691
rect 7791 15657 7800 15691
rect 7748 15648 7800 15657
rect 9496 15648 9548 15700
rect 3792 15580 3844 15632
rect 3424 15555 3476 15564
rect 3424 15521 3433 15555
rect 3433 15521 3467 15555
rect 3467 15521 3476 15555
rect 3424 15512 3476 15521
rect 8576 15580 8628 15632
rect 12716 15580 12768 15632
rect 13084 15648 13136 15700
rect 15292 15648 15344 15700
rect 16764 15648 16816 15700
rect 17316 15648 17368 15700
rect 17500 15648 17552 15700
rect 18512 15691 18564 15700
rect 8024 15512 8076 15564
rect 9680 15512 9732 15564
rect 9772 15512 9824 15564
rect 13360 15580 13412 15632
rect 18512 15657 18521 15691
rect 18521 15657 18555 15691
rect 18555 15657 18564 15691
rect 18512 15648 18564 15657
rect 18880 15648 18932 15700
rect 20352 15648 20404 15700
rect 20536 15648 20588 15700
rect 21456 15648 21508 15700
rect 22376 15648 22428 15700
rect 23020 15648 23072 15700
rect 22284 15623 22336 15632
rect 14372 15512 14424 15564
rect 14832 15555 14884 15564
rect 14832 15521 14841 15555
rect 14841 15521 14875 15555
rect 14875 15521 14884 15555
rect 14832 15512 14884 15521
rect 18236 15512 18288 15564
rect 20628 15555 20680 15564
rect 3148 15487 3200 15496
rect 3148 15453 3157 15487
rect 3157 15453 3191 15487
rect 3191 15453 3200 15487
rect 3148 15444 3200 15453
rect 9588 15444 9640 15496
rect 12624 15487 12676 15496
rect 12624 15453 12633 15487
rect 12633 15453 12667 15487
rect 12667 15453 12676 15487
rect 12624 15444 12676 15453
rect 13912 15444 13964 15496
rect 14280 15444 14332 15496
rect 16672 15444 16724 15496
rect 17224 15444 17276 15496
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 18972 15444 19024 15496
rect 20628 15521 20637 15555
rect 20637 15521 20671 15555
rect 20671 15521 20680 15555
rect 20628 15512 20680 15521
rect 21088 15512 21140 15564
rect 20536 15487 20588 15496
rect 20536 15453 20545 15487
rect 20545 15453 20579 15487
rect 20579 15453 20588 15487
rect 20536 15444 20588 15453
rect 20720 15444 20772 15496
rect 22284 15589 22293 15623
rect 22293 15589 22327 15623
rect 22327 15589 22336 15623
rect 22284 15580 22336 15589
rect 23112 15580 23164 15632
rect 10692 15376 10744 15428
rect 11152 15376 11204 15428
rect 5540 15308 5592 15360
rect 9128 15308 9180 15360
rect 10048 15308 10100 15360
rect 12808 15308 12860 15360
rect 13268 15376 13320 15428
rect 15384 15376 15436 15428
rect 15936 15376 15988 15428
rect 18328 15376 18380 15428
rect 19064 15419 19116 15428
rect 19064 15385 19073 15419
rect 19073 15385 19107 15419
rect 19107 15385 19116 15419
rect 19064 15376 19116 15385
rect 21272 15376 21324 15428
rect 21456 15376 21508 15428
rect 21824 15444 21876 15496
rect 23480 15444 23532 15496
rect 13176 15308 13228 15360
rect 14188 15308 14240 15360
rect 18604 15308 18656 15360
rect 21364 15308 21416 15360
rect 23204 15351 23256 15360
rect 23204 15317 23213 15351
rect 23213 15317 23247 15351
rect 23247 15317 23256 15351
rect 23204 15308 23256 15317
rect 23296 15351 23348 15360
rect 23296 15317 23305 15351
rect 23305 15317 23339 15351
rect 23339 15317 23348 15351
rect 23296 15308 23348 15317
rect 9322 15206 9374 15258
rect 9386 15206 9438 15258
rect 9450 15206 9502 15258
rect 9514 15206 9566 15258
rect 9578 15206 9630 15258
rect 17694 15206 17746 15258
rect 17758 15206 17810 15258
rect 17822 15206 17874 15258
rect 17886 15206 17938 15258
rect 17950 15206 18002 15258
rect 26332 15215 26384 15224
rect 26332 15181 26341 15215
rect 26341 15181 26375 15215
rect 26375 15181 26384 15215
rect 26332 15172 26384 15181
rect 4896 15104 4948 15156
rect 5540 15036 5592 15088
rect 2872 14900 2924 14952
rect 4712 14968 4764 15020
rect 5632 14968 5684 15020
rect 9864 15104 9916 15156
rect 10600 15104 10652 15156
rect 12624 15104 12676 15156
rect 18880 15104 18932 15156
rect 19340 15104 19392 15156
rect 23296 15147 23348 15156
rect 23296 15113 23305 15147
rect 23305 15113 23339 15147
rect 23339 15113 23348 15147
rect 23296 15104 23348 15113
rect 23388 15104 23440 15156
rect 7748 15036 7800 15088
rect 7380 14968 7432 15020
rect 4344 14832 4396 14884
rect 5816 14900 5868 14952
rect 6552 14900 6604 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 7288 14900 7340 14952
rect 8668 15036 8720 15088
rect 8852 15036 8904 15088
rect 9496 15036 9548 15088
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 10140 14968 10192 15020
rect 10232 15011 10284 15020
rect 10232 14977 10241 15011
rect 10241 14977 10275 15011
rect 10275 14977 10284 15011
rect 10692 15011 10744 15020
rect 10232 14968 10284 14977
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 12348 14968 12400 15020
rect 12716 14968 12768 15020
rect 4804 14832 4856 14884
rect 9220 14900 9272 14952
rect 10600 14900 10652 14952
rect 12808 14900 12860 14952
rect 4068 14764 4120 14816
rect 4712 14764 4764 14816
rect 11428 14832 11480 14884
rect 18052 15036 18104 15088
rect 15108 15011 15160 15020
rect 15108 14977 15117 15011
rect 15117 14977 15151 15011
rect 15151 14977 15160 15011
rect 15108 14968 15160 14977
rect 16580 14968 16632 15020
rect 14004 14900 14056 14952
rect 14924 14900 14976 14952
rect 15200 14943 15252 14952
rect 15200 14909 15209 14943
rect 15209 14909 15243 14943
rect 15243 14909 15252 14943
rect 15200 14900 15252 14909
rect 9496 14807 9548 14816
rect 9496 14773 9505 14807
rect 9505 14773 9539 14807
rect 9539 14773 9548 14807
rect 9496 14764 9548 14773
rect 10324 14807 10376 14816
rect 10324 14773 10333 14807
rect 10333 14773 10367 14807
rect 10367 14773 10376 14807
rect 10324 14764 10376 14773
rect 10600 14764 10652 14816
rect 12072 14807 12124 14816
rect 12072 14773 12081 14807
rect 12081 14773 12115 14807
rect 12115 14773 12124 14807
rect 12072 14764 12124 14773
rect 14464 14764 14516 14816
rect 14832 14764 14884 14816
rect 15752 14900 15804 14952
rect 18328 15011 18380 15020
rect 18328 14977 18337 15011
rect 18337 14977 18380 15011
rect 18328 14968 18380 14977
rect 18512 14968 18564 15020
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 17500 14900 17552 14952
rect 19064 14900 19116 14952
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 21272 15036 21324 15088
rect 17408 14764 17460 14816
rect 19156 14764 19208 14816
rect 21272 14943 21324 14952
rect 21272 14909 21281 14943
rect 21281 14909 21315 14943
rect 21315 14909 21324 14943
rect 21272 14900 21324 14909
rect 21732 14968 21784 15020
rect 23388 14764 23440 14816
rect 5136 14662 5188 14714
rect 5200 14662 5252 14714
rect 5264 14662 5316 14714
rect 5328 14662 5380 14714
rect 5392 14662 5444 14714
rect 13508 14662 13560 14714
rect 13572 14662 13624 14714
rect 13636 14662 13688 14714
rect 13700 14662 13752 14714
rect 13764 14662 13816 14714
rect 21880 14662 21932 14714
rect 21944 14662 21996 14714
rect 22008 14662 22060 14714
rect 22072 14662 22124 14714
rect 22136 14662 22188 14714
rect 5540 14560 5592 14612
rect 8484 14560 8536 14612
rect 9680 14560 9732 14612
rect 12716 14560 12768 14612
rect 13084 14603 13136 14612
rect 4896 14492 4948 14544
rect 10324 14424 10376 14476
rect 13084 14569 13093 14603
rect 13093 14569 13127 14603
rect 13127 14569 13136 14603
rect 13084 14560 13136 14569
rect 13912 14535 13964 14544
rect 13912 14501 13921 14535
rect 13921 14501 13955 14535
rect 13955 14501 13964 14535
rect 13912 14492 13964 14501
rect 3424 14356 3476 14408
rect 4068 14399 4120 14408
rect 4068 14365 4102 14399
rect 4102 14365 4120 14399
rect 4068 14356 4120 14365
rect 6552 14399 6604 14408
rect 6552 14365 6570 14399
rect 6570 14365 6604 14399
rect 6552 14356 6604 14365
rect 7932 14356 7984 14408
rect 9220 14356 9272 14408
rect 13820 14424 13872 14476
rect 14372 14560 14424 14612
rect 14740 14560 14792 14612
rect 17500 14560 17552 14612
rect 21272 14560 21324 14612
rect 21732 14560 21784 14612
rect 14648 14492 14700 14544
rect 19340 14492 19392 14544
rect 22376 14492 22428 14544
rect 22836 14492 22888 14544
rect 12164 14399 12216 14408
rect 12164 14365 12173 14399
rect 12173 14365 12207 14399
rect 12207 14365 12216 14399
rect 12164 14356 12216 14365
rect 12532 14356 12584 14408
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 12808 14356 12860 14365
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 13452 14356 13504 14408
rect 14004 14356 14056 14408
rect 15108 14424 15160 14476
rect 14464 14399 14516 14408
rect 14464 14365 14473 14399
rect 14473 14365 14507 14399
rect 14507 14365 14516 14399
rect 14464 14356 14516 14365
rect 14832 14356 14884 14408
rect 18144 14356 18196 14408
rect 21088 14356 21140 14408
rect 21916 14356 21968 14408
rect 23112 14424 23164 14476
rect 23480 14399 23532 14408
rect 23480 14365 23489 14399
rect 23489 14365 23523 14399
rect 23523 14365 23532 14399
rect 23480 14356 23532 14365
rect 7288 14288 7340 14340
rect 8208 14288 8260 14340
rect 8300 14288 8352 14340
rect 10232 14220 10284 14272
rect 12072 14220 12124 14272
rect 12348 14288 12400 14340
rect 15108 14288 15160 14340
rect 22468 14288 22520 14340
rect 14464 14220 14516 14272
rect 14832 14220 14884 14272
rect 15200 14220 15252 14272
rect 20168 14220 20220 14272
rect 22008 14220 22060 14272
rect 23296 14288 23348 14340
rect 9322 14118 9374 14170
rect 9386 14118 9438 14170
rect 9450 14118 9502 14170
rect 9514 14118 9566 14170
rect 9578 14118 9630 14170
rect 17694 14118 17746 14170
rect 17758 14118 17810 14170
rect 17822 14118 17874 14170
rect 17886 14118 17938 14170
rect 17950 14118 18002 14170
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 4804 14059 4856 14068
rect 4804 14025 4813 14059
rect 4813 14025 4847 14059
rect 4847 14025 4856 14059
rect 4804 14016 4856 14025
rect 6828 13948 6880 14000
rect 2320 13880 2372 13932
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 4436 13880 4488 13932
rect 6920 13923 6972 13932
rect 6920 13889 6929 13923
rect 6929 13889 6963 13923
rect 6963 13889 6972 13923
rect 6920 13880 6972 13889
rect 8668 14016 8720 14068
rect 8300 13991 8352 14000
rect 8300 13957 8309 13991
rect 8309 13957 8343 13991
rect 8343 13957 8352 13991
rect 8300 13948 8352 13957
rect 8484 13948 8536 14000
rect 8760 13991 8812 14000
rect 8760 13957 8769 13991
rect 8769 13957 8803 13991
rect 8803 13957 8812 13991
rect 8760 13948 8812 13957
rect 7196 13923 7248 13932
rect 7196 13889 7205 13923
rect 7205 13889 7239 13923
rect 7239 13889 7248 13923
rect 7196 13880 7248 13889
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 7012 13812 7064 13864
rect 7380 13676 7432 13728
rect 7748 13923 7800 13932
rect 7748 13889 7756 13923
rect 7756 13889 7790 13923
rect 7790 13889 7800 13923
rect 7748 13880 7800 13889
rect 8024 13880 8076 13932
rect 9312 13948 9364 14000
rect 14280 14016 14332 14068
rect 14372 14016 14424 14068
rect 16856 14016 16908 14068
rect 18144 14016 18196 14068
rect 19248 14016 19300 14068
rect 19616 14059 19668 14068
rect 19616 14025 19625 14059
rect 19625 14025 19659 14059
rect 19659 14025 19668 14059
rect 19616 14016 19668 14025
rect 19984 14059 20036 14068
rect 19984 14025 19993 14059
rect 19993 14025 20027 14059
rect 20027 14025 20036 14059
rect 19984 14016 20036 14025
rect 20812 14059 20864 14068
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 21916 14016 21968 14068
rect 13452 13991 13504 14000
rect 9036 13880 9088 13932
rect 12256 13880 12308 13932
rect 12624 13880 12676 13932
rect 13452 13957 13461 13991
rect 13461 13957 13495 13991
rect 13495 13957 13504 13991
rect 13452 13948 13504 13957
rect 8208 13812 8260 13864
rect 8484 13812 8536 13864
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 13544 13880 13596 13932
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 14464 13923 14516 13932
rect 8944 13812 8996 13821
rect 8300 13744 8352 13796
rect 13268 13744 13320 13796
rect 13728 13812 13780 13864
rect 14464 13889 14473 13923
rect 14473 13889 14507 13923
rect 14507 13889 14516 13923
rect 14464 13880 14516 13889
rect 14832 13991 14884 14000
rect 14832 13957 14841 13991
rect 14841 13957 14875 13991
rect 14875 13957 14884 13991
rect 14832 13948 14884 13957
rect 18512 13948 18564 14000
rect 20444 13923 20496 13932
rect 14740 13812 14792 13864
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 20812 13880 20864 13932
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 22284 13880 22336 13932
rect 22836 13880 22888 13932
rect 19892 13812 19944 13864
rect 20168 13855 20220 13864
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 20352 13855 20404 13864
rect 20352 13821 20361 13855
rect 20361 13821 20395 13855
rect 20395 13821 20404 13855
rect 20352 13812 20404 13821
rect 22560 13855 22612 13864
rect 22560 13821 22569 13855
rect 22569 13821 22603 13855
rect 22603 13821 22612 13855
rect 22560 13812 22612 13821
rect 14464 13744 14516 13796
rect 14648 13744 14700 13796
rect 17224 13744 17276 13796
rect 8208 13676 8260 13728
rect 11520 13719 11572 13728
rect 11520 13685 11529 13719
rect 11529 13685 11563 13719
rect 11563 13685 11572 13719
rect 11520 13676 11572 13685
rect 11980 13676 12032 13728
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 17500 13676 17552 13728
rect 20904 13676 20956 13728
rect 20996 13676 21048 13728
rect 23020 13744 23072 13796
rect 21640 13676 21692 13728
rect 22652 13719 22704 13728
rect 22652 13685 22661 13719
rect 22661 13685 22695 13719
rect 22695 13685 22704 13719
rect 22652 13676 22704 13685
rect 5136 13574 5188 13626
rect 5200 13574 5252 13626
rect 5264 13574 5316 13626
rect 5328 13574 5380 13626
rect 5392 13574 5444 13626
rect 13508 13574 13560 13626
rect 13572 13574 13624 13626
rect 13636 13574 13688 13626
rect 13700 13574 13752 13626
rect 13764 13574 13816 13626
rect 21880 13574 21932 13626
rect 21944 13574 21996 13626
rect 22008 13574 22060 13626
rect 22072 13574 22124 13626
rect 22136 13574 22188 13626
rect 3332 13472 3384 13524
rect 8484 13472 8536 13524
rect 8668 13472 8720 13524
rect 8944 13472 8996 13524
rect 2504 13404 2556 13456
rect 8116 13404 8168 13456
rect 3424 13336 3476 13388
rect 7932 13379 7984 13388
rect 7932 13345 7941 13379
rect 7941 13345 7975 13379
rect 7975 13345 7984 13379
rect 7932 13336 7984 13345
rect 8300 13336 8352 13388
rect 1492 13311 1544 13320
rect 1492 13277 1501 13311
rect 1501 13277 1535 13311
rect 1535 13277 1544 13311
rect 1492 13268 1544 13277
rect 3240 13268 3292 13320
rect 4988 13268 5040 13320
rect 6460 13268 6512 13320
rect 2136 13200 2188 13252
rect 3424 13200 3476 13252
rect 7012 13200 7064 13252
rect 8024 13200 8076 13252
rect 8576 13311 8628 13320
rect 8576 13277 8586 13311
rect 8586 13277 8620 13311
rect 8620 13277 8628 13311
rect 10416 13472 10468 13524
rect 12164 13472 12216 13524
rect 14004 13472 14056 13524
rect 14372 13472 14424 13524
rect 14556 13515 14608 13524
rect 14556 13481 14565 13515
rect 14565 13481 14599 13515
rect 14599 13481 14608 13515
rect 14556 13472 14608 13481
rect 16488 13472 16540 13524
rect 9220 13336 9272 13388
rect 8576 13268 8628 13277
rect 9036 13268 9088 13320
rect 12900 13404 12952 13456
rect 13084 13404 13136 13456
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 12072 13379 12124 13388
rect 12072 13345 12081 13379
rect 12081 13345 12115 13379
rect 12115 13345 12124 13379
rect 12072 13336 12124 13345
rect 11888 13311 11940 13320
rect 11888 13277 11896 13311
rect 11896 13277 11930 13311
rect 11930 13277 11940 13311
rect 11888 13268 11940 13277
rect 9680 13243 9732 13252
rect 9680 13209 9714 13243
rect 9714 13209 9732 13243
rect 9680 13200 9732 13209
rect 11244 13200 11296 13252
rect 12256 13311 12308 13320
rect 12256 13277 12265 13311
rect 12265 13277 12299 13311
rect 12299 13277 12308 13311
rect 12256 13268 12308 13277
rect 3148 13175 3200 13184
rect 3148 13141 3157 13175
rect 3157 13141 3191 13175
rect 3191 13141 3200 13175
rect 3148 13132 3200 13141
rect 6920 13132 6972 13184
rect 7196 13132 7248 13184
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 8944 13132 8996 13184
rect 9864 13132 9916 13184
rect 10692 13132 10744 13184
rect 11428 13175 11480 13184
rect 11428 13141 11437 13175
rect 11437 13141 11471 13175
rect 11471 13141 11480 13175
rect 11428 13132 11480 13141
rect 11888 13132 11940 13184
rect 14372 13336 14424 13388
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 14004 13268 14056 13320
rect 14280 13268 14332 13320
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 15844 13336 15896 13388
rect 16856 13379 16908 13388
rect 16856 13345 16865 13379
rect 16865 13345 16899 13379
rect 16899 13345 16908 13379
rect 16856 13336 16908 13345
rect 13268 13200 13320 13252
rect 15108 13200 15160 13252
rect 16580 13200 16632 13252
rect 17500 13472 17552 13524
rect 17592 13472 17644 13524
rect 18696 13472 18748 13524
rect 19616 13472 19668 13524
rect 20444 13472 20496 13524
rect 20996 13515 21048 13524
rect 17408 13379 17460 13388
rect 17408 13345 17417 13379
rect 17417 13345 17451 13379
rect 17451 13345 17460 13379
rect 17408 13336 17460 13345
rect 17592 13336 17644 13388
rect 18512 13379 18564 13388
rect 18512 13345 18521 13379
rect 18521 13345 18555 13379
rect 18555 13345 18564 13379
rect 18512 13336 18564 13345
rect 17224 13268 17276 13320
rect 19524 13404 19576 13456
rect 19248 13336 19300 13388
rect 20996 13481 21005 13515
rect 21005 13481 21039 13515
rect 21039 13481 21048 13515
rect 20996 13472 21048 13481
rect 22284 13472 22336 13524
rect 18236 13200 18288 13252
rect 19892 13200 19944 13252
rect 20352 13268 20404 13320
rect 20628 13268 20680 13320
rect 21272 13404 21324 13456
rect 21640 13404 21692 13456
rect 20904 13268 20956 13320
rect 21456 13277 21462 13296
rect 21462 13277 21496 13296
rect 21496 13277 21508 13296
rect 21456 13244 21508 13277
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 22008 13311 22060 13320
rect 22008 13277 22017 13311
rect 22017 13277 22051 13311
rect 22051 13277 22060 13311
rect 22008 13268 22060 13277
rect 22560 13268 22612 13320
rect 23388 13268 23440 13320
rect 23480 13268 23532 13320
rect 23664 13268 23716 13320
rect 14832 13132 14884 13184
rect 15292 13132 15344 13184
rect 16028 13175 16080 13184
rect 16028 13141 16037 13175
rect 16037 13141 16071 13175
rect 16071 13141 16080 13175
rect 16028 13132 16080 13141
rect 16948 13132 17000 13184
rect 18052 13132 18104 13184
rect 19800 13175 19852 13184
rect 19800 13141 19809 13175
rect 19809 13141 19843 13175
rect 19843 13141 19852 13175
rect 19800 13132 19852 13141
rect 21824 13200 21876 13252
rect 21640 13132 21692 13184
rect 23112 13132 23164 13184
rect 23296 13132 23348 13184
rect 9322 13030 9374 13082
rect 9386 13030 9438 13082
rect 9450 13030 9502 13082
rect 9514 13030 9566 13082
rect 9578 13030 9630 13082
rect 17694 13030 17746 13082
rect 17758 13030 17810 13082
rect 17822 13030 17874 13082
rect 17886 13030 17938 13082
rect 17950 13030 18002 13082
rect 2136 12971 2188 12980
rect 2136 12937 2145 12971
rect 2145 12937 2179 12971
rect 2179 12937 2188 12971
rect 2136 12928 2188 12937
rect 2504 12860 2556 12912
rect 2596 12792 2648 12844
rect 2964 12928 3016 12980
rect 3424 12971 3476 12980
rect 3424 12937 3433 12971
rect 3433 12937 3467 12971
rect 3467 12937 3476 12971
rect 3424 12928 3476 12937
rect 2872 12724 2924 12776
rect 3332 12835 3384 12844
rect 3332 12801 3341 12835
rect 3341 12801 3375 12835
rect 3375 12801 3384 12835
rect 3332 12792 3384 12801
rect 3516 12792 3568 12844
rect 3792 12835 3844 12844
rect 3792 12801 3800 12835
rect 3800 12801 3834 12835
rect 3834 12801 3844 12835
rect 3792 12792 3844 12801
rect 3976 12928 4028 12980
rect 4896 12928 4948 12980
rect 6460 12971 6512 12980
rect 6460 12937 6469 12971
rect 6469 12937 6503 12971
rect 6503 12937 6512 12971
rect 6460 12928 6512 12937
rect 7748 12928 7800 12980
rect 8392 12928 8444 12980
rect 9680 12928 9732 12980
rect 9772 12928 9824 12980
rect 10508 12928 10560 12980
rect 11152 12928 11204 12980
rect 11704 12928 11756 12980
rect 12256 12928 12308 12980
rect 4436 12903 4488 12912
rect 4436 12869 4445 12903
rect 4445 12869 4479 12903
rect 4479 12869 4488 12903
rect 4436 12860 4488 12869
rect 4528 12792 4580 12844
rect 4804 12860 4856 12912
rect 8116 12860 8168 12912
rect 4988 12835 5040 12844
rect 4988 12801 4998 12835
rect 4998 12801 5032 12835
rect 5032 12801 5040 12835
rect 4988 12792 5040 12801
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5724 12792 5776 12844
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 7932 12792 7984 12844
rect 8760 12792 8812 12844
rect 9404 12792 9456 12844
rect 2964 12656 3016 12708
rect 4344 12724 4396 12776
rect 4804 12767 4856 12776
rect 4804 12733 4813 12767
rect 4813 12733 4847 12767
rect 4847 12733 4856 12767
rect 4804 12724 4856 12733
rect 4896 12767 4948 12776
rect 4896 12733 4905 12767
rect 4905 12733 4939 12767
rect 4939 12733 4948 12767
rect 4896 12724 4948 12733
rect 4712 12656 4764 12708
rect 3332 12588 3384 12640
rect 4160 12588 4212 12640
rect 4528 12588 4580 12640
rect 4988 12588 5040 12640
rect 8484 12724 8536 12776
rect 8668 12724 8720 12776
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 9036 12656 9088 12708
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 9956 12835 10008 12844
rect 9956 12801 9964 12835
rect 9964 12801 9998 12835
rect 9998 12801 10008 12835
rect 9956 12792 10008 12801
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 10508 12792 10560 12844
rect 10692 12792 10744 12844
rect 11520 12860 11572 12912
rect 11336 12792 11388 12844
rect 13268 12860 13320 12912
rect 14556 12928 14608 12980
rect 15108 12971 15160 12980
rect 15108 12937 15117 12971
rect 15117 12937 15151 12971
rect 15151 12937 15160 12971
rect 15108 12928 15160 12937
rect 16396 12928 16448 12980
rect 17500 12928 17552 12980
rect 18052 12971 18104 12980
rect 18052 12937 18061 12971
rect 18061 12937 18095 12971
rect 18095 12937 18104 12971
rect 18052 12928 18104 12937
rect 21272 12928 21324 12980
rect 11244 12724 11296 12776
rect 12440 12792 12492 12844
rect 16028 12860 16080 12912
rect 17592 12860 17644 12912
rect 10232 12656 10284 12708
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 16764 12767 16816 12776
rect 16764 12733 16773 12767
rect 16773 12733 16807 12767
rect 16807 12733 16816 12767
rect 16764 12724 16816 12733
rect 18052 12792 18104 12844
rect 22008 12860 22060 12912
rect 18236 12792 18288 12844
rect 19984 12835 20036 12844
rect 19984 12801 19993 12835
rect 19993 12801 20036 12835
rect 19984 12792 20036 12801
rect 20812 12835 20864 12844
rect 17500 12724 17552 12776
rect 19708 12699 19760 12708
rect 10416 12588 10468 12640
rect 12256 12588 12308 12640
rect 12348 12588 12400 12640
rect 15384 12588 15436 12640
rect 16856 12588 16908 12640
rect 19708 12665 19717 12699
rect 19717 12665 19751 12699
rect 19751 12665 19760 12699
rect 19708 12656 19760 12665
rect 20352 12767 20404 12776
rect 20352 12733 20361 12767
rect 20361 12733 20395 12767
rect 20395 12733 20404 12767
rect 20352 12724 20404 12733
rect 20812 12801 20821 12835
rect 20821 12801 20855 12835
rect 20855 12801 20864 12835
rect 20812 12792 20864 12801
rect 20996 12792 21048 12844
rect 21640 12835 21692 12844
rect 21640 12801 21649 12835
rect 21649 12801 21683 12835
rect 21683 12801 21692 12835
rect 21640 12792 21692 12801
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 22376 12792 22428 12844
rect 21456 12767 21508 12776
rect 21456 12733 21465 12767
rect 21465 12733 21499 12767
rect 21499 12733 21508 12767
rect 21456 12724 21508 12733
rect 21732 12724 21784 12776
rect 22744 12792 22796 12844
rect 22928 12724 22980 12776
rect 23296 12792 23348 12844
rect 23480 12835 23532 12844
rect 23480 12801 23489 12835
rect 23489 12801 23523 12835
rect 23523 12801 23532 12835
rect 23480 12792 23532 12801
rect 23664 12835 23716 12844
rect 23664 12801 23673 12835
rect 23673 12801 23707 12835
rect 23707 12801 23716 12835
rect 23664 12792 23716 12801
rect 19800 12588 19852 12640
rect 22744 12656 22796 12708
rect 23020 12656 23072 12708
rect 25136 12631 25188 12640
rect 25136 12597 25145 12631
rect 25145 12597 25179 12631
rect 25179 12597 25188 12631
rect 25136 12588 25188 12597
rect 5136 12486 5188 12538
rect 5200 12486 5252 12538
rect 5264 12486 5316 12538
rect 5328 12486 5380 12538
rect 5392 12486 5444 12538
rect 13508 12486 13560 12538
rect 13572 12486 13624 12538
rect 13636 12486 13688 12538
rect 13700 12486 13752 12538
rect 13764 12486 13816 12538
rect 21880 12486 21932 12538
rect 21944 12486 21996 12538
rect 22008 12486 22060 12538
rect 22072 12486 22124 12538
rect 22136 12486 22188 12538
rect 2320 12427 2372 12436
rect 2320 12393 2329 12427
rect 2329 12393 2363 12427
rect 2363 12393 2372 12427
rect 2320 12384 2372 12393
rect 3148 12384 3200 12436
rect 3332 12427 3384 12436
rect 3332 12393 3341 12427
rect 3341 12393 3375 12427
rect 3375 12393 3384 12427
rect 3332 12384 3384 12393
rect 4804 12384 4856 12436
rect 4988 12384 5040 12436
rect 5540 12384 5592 12436
rect 5908 12384 5960 12436
rect 7656 12384 7708 12436
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 8024 12384 8076 12436
rect 8484 12427 8536 12436
rect 8484 12393 8493 12427
rect 8493 12393 8527 12427
rect 8527 12393 8536 12427
rect 8484 12384 8536 12393
rect 9404 12384 9456 12436
rect 10324 12384 10376 12436
rect 12348 12384 12400 12436
rect 14832 12384 14884 12436
rect 16948 12427 17000 12436
rect 16948 12393 16957 12427
rect 16957 12393 16991 12427
rect 16991 12393 17000 12427
rect 16948 12384 17000 12393
rect 2872 12316 2924 12368
rect 2688 12248 2740 12300
rect 6276 12316 6328 12368
rect 10968 12316 11020 12368
rect 14740 12316 14792 12368
rect 4896 12248 4948 12300
rect 7564 12248 7616 12300
rect 8484 12248 8536 12300
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 15016 12248 15068 12300
rect 3056 12180 3108 12232
rect 3240 12180 3292 12232
rect 3424 12180 3476 12232
rect 3884 12223 3936 12232
rect 3884 12189 3893 12223
rect 3893 12189 3927 12223
rect 3927 12189 3936 12223
rect 3884 12180 3936 12189
rect 4160 12223 4212 12232
rect 4160 12189 4194 12223
rect 4194 12189 4212 12223
rect 5632 12223 5684 12232
rect 4160 12180 4212 12189
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 5632 12180 5684 12189
rect 5724 12180 5776 12232
rect 2688 12112 2740 12164
rect 4712 12112 4764 12164
rect 5908 12155 5960 12164
rect 5908 12121 5917 12155
rect 5917 12121 5951 12155
rect 5951 12121 5960 12155
rect 5908 12112 5960 12121
rect 6184 12180 6236 12232
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 9128 12180 9180 12232
rect 10324 12180 10376 12232
rect 10508 12180 10560 12232
rect 10232 12112 10284 12164
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 6276 12044 6328 12096
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 9220 12087 9272 12096
rect 9220 12053 9229 12087
rect 9229 12053 9263 12087
rect 9263 12053 9272 12087
rect 9956 12087 10008 12096
rect 9220 12044 9272 12053
rect 9956 12053 9965 12087
rect 9965 12053 9999 12087
rect 9999 12053 10008 12087
rect 9956 12044 10008 12053
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 12440 12180 12492 12232
rect 15292 12223 15344 12232
rect 15292 12189 15301 12223
rect 15301 12189 15335 12223
rect 15335 12189 15344 12223
rect 15292 12180 15344 12189
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 16672 12316 16724 12368
rect 17500 12316 17552 12368
rect 17684 12316 17736 12368
rect 18236 12316 18288 12368
rect 16396 12291 16448 12300
rect 16396 12257 16405 12291
rect 16405 12257 16439 12291
rect 16439 12257 16448 12291
rect 16396 12248 16448 12257
rect 15384 12180 15436 12189
rect 16580 12180 16632 12232
rect 16764 12180 16816 12232
rect 18328 12248 18380 12300
rect 17224 12180 17276 12232
rect 17500 12180 17552 12232
rect 17040 12155 17092 12164
rect 17040 12121 17049 12155
rect 17049 12121 17083 12155
rect 17083 12121 17092 12155
rect 17040 12112 17092 12121
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 20352 12384 20404 12436
rect 21272 12427 21324 12436
rect 21272 12393 21281 12427
rect 21281 12393 21315 12427
rect 21315 12393 21324 12427
rect 21272 12384 21324 12393
rect 21640 12427 21692 12436
rect 21640 12393 21649 12427
rect 21649 12393 21683 12427
rect 21683 12393 21692 12427
rect 21640 12384 21692 12393
rect 19524 12316 19576 12368
rect 20168 12316 20220 12368
rect 19708 12180 19760 12232
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 20996 12291 21048 12300
rect 20996 12257 21005 12291
rect 21005 12257 21039 12291
rect 21039 12257 21048 12291
rect 20996 12248 21048 12257
rect 21456 12316 21508 12368
rect 22468 12359 22520 12368
rect 22468 12325 22477 12359
rect 22477 12325 22511 12359
rect 22511 12325 22520 12359
rect 22468 12316 22520 12325
rect 22836 12316 22888 12368
rect 21732 12180 21784 12232
rect 22652 12180 22704 12232
rect 12348 12044 12400 12096
rect 15936 12044 15988 12096
rect 16488 12044 16540 12096
rect 16764 12044 16816 12096
rect 18052 12044 18104 12096
rect 18236 12044 18288 12096
rect 19892 12044 19944 12096
rect 20352 12044 20404 12096
rect 9322 11942 9374 11994
rect 9386 11942 9438 11994
rect 9450 11942 9502 11994
rect 9514 11942 9566 11994
rect 9578 11942 9630 11994
rect 17694 11942 17746 11994
rect 17758 11942 17810 11994
rect 17822 11942 17874 11994
rect 17886 11942 17938 11994
rect 17950 11942 18002 11994
rect 2872 11883 2924 11892
rect 2872 11849 2881 11883
rect 2881 11849 2915 11883
rect 2915 11849 2924 11883
rect 2872 11840 2924 11849
rect 4436 11840 4488 11892
rect 5172 11883 5224 11892
rect 5172 11849 5181 11883
rect 5181 11849 5215 11883
rect 5215 11849 5224 11883
rect 5172 11840 5224 11849
rect 5264 11840 5316 11892
rect 7104 11840 7156 11892
rect 1492 11772 1544 11824
rect 2320 11704 2372 11756
rect 3884 11772 3936 11824
rect 9588 11772 9640 11824
rect 9956 11772 10008 11824
rect 11060 11840 11112 11892
rect 11336 11840 11388 11892
rect 16396 11883 16448 11892
rect 4528 11704 4580 11756
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 6184 11704 6236 11756
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 1492 11679 1544 11688
rect 1492 11645 1501 11679
rect 1501 11645 1535 11679
rect 1535 11645 1544 11679
rect 1492 11636 1544 11645
rect 4804 11636 4856 11688
rect 5264 11636 5316 11688
rect 5540 11636 5592 11688
rect 9496 11747 9548 11756
rect 9496 11713 9505 11747
rect 9505 11713 9539 11747
rect 9539 11713 9548 11747
rect 9496 11704 9548 11713
rect 9864 11704 9916 11756
rect 8024 11636 8076 11688
rect 9404 11636 9456 11688
rect 9772 11636 9824 11688
rect 11704 11772 11756 11824
rect 10784 11704 10836 11756
rect 11888 11704 11940 11756
rect 12440 11772 12492 11824
rect 12256 11747 12308 11756
rect 12256 11713 12290 11747
rect 12290 11713 12308 11747
rect 12256 11704 12308 11713
rect 13912 11704 13964 11756
rect 11612 11636 11664 11688
rect 16396 11849 16405 11883
rect 16405 11849 16439 11883
rect 16439 11849 16448 11883
rect 16396 11840 16448 11849
rect 16856 11840 16908 11892
rect 17592 11840 17644 11892
rect 19984 11840 20036 11892
rect 23112 11840 23164 11892
rect 23388 11840 23440 11892
rect 16672 11772 16724 11824
rect 15384 11704 15436 11756
rect 15936 11747 15988 11756
rect 15936 11713 15945 11747
rect 15945 11713 15979 11747
rect 15979 11713 15988 11747
rect 15936 11704 15988 11713
rect 17500 11772 17552 11824
rect 17040 11704 17092 11756
rect 17224 11747 17276 11756
rect 17224 11713 17233 11747
rect 17233 11713 17267 11747
rect 17267 11713 17276 11747
rect 17224 11704 17276 11713
rect 17592 11747 17644 11756
rect 17592 11713 17601 11747
rect 17601 11713 17635 11747
rect 17635 11713 17644 11747
rect 17592 11704 17644 11713
rect 18052 11747 18104 11756
rect 18052 11713 18061 11747
rect 18061 11713 18095 11747
rect 18095 11713 18104 11747
rect 18052 11704 18104 11713
rect 20352 11747 20404 11756
rect 20352 11713 20361 11747
rect 20361 11713 20395 11747
rect 20395 11713 20404 11747
rect 20352 11704 20404 11713
rect 20812 11704 20864 11756
rect 23020 11747 23072 11756
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 15844 11679 15896 11688
rect 4988 11568 5040 11620
rect 5632 11543 5684 11552
rect 5632 11509 5641 11543
rect 5641 11509 5675 11543
rect 5675 11509 5684 11543
rect 5632 11500 5684 11509
rect 8668 11500 8720 11552
rect 9404 11500 9456 11552
rect 9588 11500 9640 11552
rect 10232 11543 10284 11552
rect 10232 11509 10241 11543
rect 10241 11509 10275 11543
rect 10275 11509 10284 11543
rect 10232 11500 10284 11509
rect 15568 11568 15620 11620
rect 15844 11645 15853 11679
rect 15853 11645 15887 11679
rect 15887 11645 15896 11679
rect 15844 11636 15896 11645
rect 18328 11636 18380 11688
rect 16948 11611 17000 11620
rect 15476 11500 15528 11552
rect 16672 11500 16724 11552
rect 16948 11577 16957 11611
rect 16957 11577 16991 11611
rect 16991 11577 17000 11611
rect 16948 11568 17000 11577
rect 17316 11568 17368 11620
rect 17408 11500 17460 11552
rect 20628 11500 20680 11552
rect 5136 11398 5188 11450
rect 5200 11398 5252 11450
rect 5264 11398 5316 11450
rect 5328 11398 5380 11450
rect 5392 11398 5444 11450
rect 13508 11398 13560 11450
rect 13572 11398 13624 11450
rect 13636 11398 13688 11450
rect 13700 11398 13752 11450
rect 13764 11398 13816 11450
rect 21880 11398 21932 11450
rect 21944 11398 21996 11450
rect 22008 11398 22060 11450
rect 22072 11398 22124 11450
rect 22136 11398 22188 11450
rect 2320 11296 2372 11348
rect 2872 11296 2924 11348
rect 4528 11339 4580 11348
rect 4528 11305 4537 11339
rect 4537 11305 4571 11339
rect 4571 11305 4580 11339
rect 4528 11296 4580 11305
rect 7472 11339 7524 11348
rect 2872 11203 2924 11212
rect 2872 11169 2881 11203
rect 2881 11169 2915 11203
rect 2915 11169 2924 11203
rect 2872 11160 2924 11169
rect 3056 11160 3108 11212
rect 3516 11160 3568 11212
rect 2780 11092 2832 11144
rect 3700 11092 3752 11144
rect 3976 11160 4028 11212
rect 4620 11160 4672 11212
rect 5632 11203 5684 11212
rect 4068 11135 4120 11144
rect 4068 11101 4076 11135
rect 4076 11101 4110 11135
rect 4110 11101 4120 11135
rect 4068 11092 4120 11101
rect 4436 11135 4488 11144
rect 4436 11101 4445 11135
rect 4445 11101 4479 11135
rect 4479 11101 4488 11135
rect 4436 11092 4488 11101
rect 4896 11092 4948 11144
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 5540 11135 5592 11144
rect 5540 11101 5549 11135
rect 5549 11101 5583 11135
rect 5583 11101 5592 11135
rect 7472 11305 7481 11339
rect 7481 11305 7515 11339
rect 7515 11305 7524 11339
rect 7472 11296 7524 11305
rect 9312 11296 9364 11348
rect 7748 11228 7800 11280
rect 9864 11296 9916 11348
rect 13912 11296 13964 11348
rect 17592 11296 17644 11348
rect 21548 11296 21600 11348
rect 5540 11092 5592 11101
rect 6920 11092 6972 11144
rect 14924 11228 14976 11280
rect 8484 11160 8536 11212
rect 9036 11160 9088 11212
rect 9588 11160 9640 11212
rect 11336 11092 11388 11144
rect 15844 11228 15896 11280
rect 17132 11228 17184 11280
rect 17408 11228 17460 11280
rect 15292 11160 15344 11212
rect 15752 11160 15804 11212
rect 21180 11228 21232 11280
rect 22192 11228 22244 11280
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 15568 11135 15620 11144
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 5632 11024 5684 11076
rect 6184 11024 6236 11076
rect 7564 11024 7616 11076
rect 6460 10956 6512 11008
rect 7748 11024 7800 11076
rect 12348 11024 12400 11076
rect 16580 11092 16632 11144
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 19616 11092 19668 11144
rect 19892 11135 19944 11144
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 17132 11067 17184 11076
rect 17132 11033 17141 11067
rect 17141 11033 17175 11067
rect 17175 11033 17184 11067
rect 17132 11024 17184 11033
rect 8300 10956 8352 11008
rect 9680 10956 9732 11008
rect 10508 10956 10560 11008
rect 15200 10956 15252 11008
rect 20352 11092 20404 11144
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 23296 11203 23348 11212
rect 23296 11169 23305 11203
rect 23305 11169 23339 11203
rect 23339 11169 23348 11203
rect 23296 11160 23348 11169
rect 22560 11092 22612 11144
rect 23204 11092 23256 11144
rect 21732 11024 21784 11076
rect 20536 10999 20588 11008
rect 20536 10965 20545 10999
rect 20545 10965 20579 10999
rect 20579 10965 20588 10999
rect 20536 10956 20588 10965
rect 21456 10956 21508 11008
rect 22376 11024 22428 11076
rect 22928 11067 22980 11076
rect 22928 11033 22937 11067
rect 22937 11033 22971 11067
rect 22971 11033 22980 11067
rect 22928 11024 22980 11033
rect 22468 10999 22520 11008
rect 22468 10965 22477 10999
rect 22477 10965 22511 10999
rect 22511 10965 22520 10999
rect 22468 10956 22520 10965
rect 9322 10854 9374 10906
rect 9386 10854 9438 10906
rect 9450 10854 9502 10906
rect 9514 10854 9566 10906
rect 9578 10854 9630 10906
rect 17694 10854 17746 10906
rect 17758 10854 17810 10906
rect 17822 10854 17874 10906
rect 17886 10854 17938 10906
rect 17950 10854 18002 10906
rect 2872 10795 2924 10804
rect 2872 10761 2881 10795
rect 2881 10761 2915 10795
rect 2915 10761 2924 10795
rect 2872 10752 2924 10761
rect 4804 10752 4856 10804
rect 3332 10616 3384 10668
rect 4804 10659 4856 10668
rect 4804 10625 4812 10659
rect 4812 10625 4846 10659
rect 4846 10625 4856 10659
rect 4804 10616 4856 10625
rect 5540 10752 5592 10804
rect 5632 10752 5684 10804
rect 2872 10548 2924 10600
rect 3792 10548 3844 10600
rect 5264 10616 5316 10668
rect 7472 10752 7524 10804
rect 7748 10795 7800 10804
rect 7748 10761 7757 10795
rect 7757 10761 7791 10795
rect 7791 10761 7800 10795
rect 7748 10752 7800 10761
rect 9772 10752 9824 10804
rect 9864 10752 9916 10804
rect 14096 10752 14148 10804
rect 17040 10752 17092 10804
rect 19892 10752 19944 10804
rect 20536 10795 20588 10804
rect 20536 10761 20545 10795
rect 20545 10761 20579 10795
rect 20579 10761 20588 10795
rect 20536 10752 20588 10761
rect 21180 10752 21232 10804
rect 22192 10795 22244 10804
rect 22192 10761 22201 10795
rect 22201 10761 22235 10795
rect 22235 10761 22244 10795
rect 22192 10752 22244 10761
rect 22560 10752 22612 10804
rect 23020 10752 23072 10804
rect 6184 10727 6236 10736
rect 6184 10693 6193 10727
rect 6193 10693 6227 10727
rect 6227 10693 6236 10727
rect 6184 10684 6236 10693
rect 6920 10684 6972 10736
rect 5540 10480 5592 10532
rect 6460 10616 6512 10668
rect 7932 10659 7984 10668
rect 7932 10625 7941 10659
rect 7941 10625 7975 10659
rect 7975 10625 7984 10659
rect 7932 10616 7984 10625
rect 8024 10616 8076 10668
rect 8760 10616 8812 10668
rect 9680 10659 9732 10668
rect 9680 10625 9688 10659
rect 9688 10625 9722 10659
rect 9722 10625 9732 10659
rect 9680 10616 9732 10625
rect 10232 10616 10284 10668
rect 13084 10684 13136 10736
rect 16396 10684 16448 10736
rect 10508 10659 10560 10668
rect 10508 10625 10516 10659
rect 10516 10625 10550 10659
rect 10550 10625 10560 10659
rect 10508 10616 10560 10625
rect 5724 10591 5776 10600
rect 5724 10557 5733 10591
rect 5733 10557 5767 10591
rect 5767 10557 5776 10591
rect 5724 10548 5776 10557
rect 9404 10548 9456 10600
rect 6000 10480 6052 10532
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 11612 10616 11664 10668
rect 11888 10616 11940 10668
rect 12716 10659 12768 10668
rect 12716 10625 12750 10659
rect 12750 10625 12768 10659
rect 12716 10616 12768 10625
rect 15200 10616 15252 10668
rect 15568 10659 15620 10668
rect 15568 10625 15577 10659
rect 15577 10625 15611 10659
rect 15611 10625 15620 10659
rect 15568 10616 15620 10625
rect 16580 10616 16632 10668
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 17592 10684 17644 10736
rect 22652 10684 22704 10736
rect 17684 10659 17736 10668
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 6092 10412 6144 10464
rect 10140 10455 10192 10464
rect 10140 10421 10149 10455
rect 10149 10421 10183 10455
rect 10183 10421 10192 10455
rect 10140 10412 10192 10421
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 15476 10480 15528 10532
rect 15660 10480 15712 10532
rect 17684 10625 17693 10659
rect 17693 10625 17727 10659
rect 17727 10625 17736 10659
rect 17684 10616 17736 10625
rect 17776 10616 17828 10668
rect 18788 10659 18840 10668
rect 18788 10625 18797 10659
rect 18797 10625 18831 10659
rect 18831 10625 18840 10659
rect 18788 10616 18840 10625
rect 19432 10659 19484 10668
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 20628 10659 20680 10668
rect 20628 10625 20637 10659
rect 20637 10625 20671 10659
rect 20671 10625 20680 10659
rect 20628 10616 20680 10625
rect 21180 10659 21232 10668
rect 21180 10625 21189 10659
rect 21189 10625 21223 10659
rect 21223 10625 21232 10659
rect 21180 10616 21232 10625
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 23020 10659 23072 10668
rect 19616 10548 19668 10600
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 15292 10412 15344 10464
rect 16304 10455 16356 10464
rect 16304 10421 16313 10455
rect 16313 10421 16347 10455
rect 16347 10421 16356 10455
rect 16304 10412 16356 10421
rect 16488 10412 16540 10464
rect 17868 10455 17920 10464
rect 17868 10421 17877 10455
rect 17877 10421 17911 10455
rect 17911 10421 17920 10455
rect 17868 10412 17920 10421
rect 18972 10455 19024 10464
rect 18972 10421 18981 10455
rect 18981 10421 19015 10455
rect 19015 10421 19024 10455
rect 18972 10412 19024 10421
rect 19800 10455 19852 10464
rect 19800 10421 19809 10455
rect 19809 10421 19843 10455
rect 19843 10421 19852 10455
rect 19800 10412 19852 10421
rect 19984 10455 20036 10464
rect 19984 10421 19993 10455
rect 19993 10421 20027 10455
rect 20027 10421 20036 10455
rect 19984 10412 20036 10421
rect 21456 10548 21508 10600
rect 22376 10591 22428 10600
rect 22376 10557 22385 10591
rect 22385 10557 22419 10591
rect 22419 10557 22428 10591
rect 22376 10548 22428 10557
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 23296 10591 23348 10600
rect 23296 10557 23305 10591
rect 23305 10557 23339 10591
rect 23339 10557 23348 10591
rect 23296 10548 23348 10557
rect 20812 10412 20864 10464
rect 22284 10412 22336 10464
rect 22836 10412 22888 10464
rect 5136 10310 5188 10362
rect 5200 10310 5252 10362
rect 5264 10310 5316 10362
rect 5328 10310 5380 10362
rect 5392 10310 5444 10362
rect 13508 10310 13560 10362
rect 13572 10310 13624 10362
rect 13636 10310 13688 10362
rect 13700 10310 13752 10362
rect 13764 10310 13816 10362
rect 21880 10310 21932 10362
rect 21944 10310 21996 10362
rect 22008 10310 22060 10362
rect 22072 10310 22124 10362
rect 22136 10310 22188 10362
rect 2872 10251 2924 10260
rect 2872 10217 2881 10251
rect 2881 10217 2915 10251
rect 2915 10217 2924 10251
rect 2872 10208 2924 10217
rect 5540 10208 5592 10260
rect 8300 10208 8352 10260
rect 3332 10140 3384 10192
rect 3608 10140 3660 10192
rect 8392 10140 8444 10192
rect 10232 10208 10284 10260
rect 11612 10208 11664 10260
rect 12716 10208 12768 10260
rect 17040 10251 17092 10260
rect 17040 10217 17049 10251
rect 17049 10217 17083 10251
rect 17083 10217 17092 10251
rect 17040 10208 17092 10217
rect 18788 10208 18840 10260
rect 19616 10208 19668 10260
rect 17592 10140 17644 10192
rect 1492 10115 1544 10124
rect 1492 10081 1501 10115
rect 1501 10081 1535 10115
rect 1535 10081 1544 10115
rect 1492 10072 1544 10081
rect 3148 10072 3200 10124
rect 4068 10072 4120 10124
rect 9404 10072 9456 10124
rect 14096 10072 14148 10124
rect 15292 10072 15344 10124
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 17132 10072 17184 10124
rect 17776 10072 17828 10124
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 20628 10072 20680 10124
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 3424 10004 3476 10056
rect 4988 10004 5040 10056
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 6920 10004 6972 10056
rect 8300 10004 8352 10056
rect 2504 9936 2556 9988
rect 6092 9979 6144 9988
rect 6092 9945 6126 9979
rect 6126 9945 6144 9979
rect 6092 9936 6144 9945
rect 8668 10004 8720 10056
rect 8760 10047 8812 10056
rect 8760 10013 8769 10047
rect 8769 10013 8803 10047
rect 8803 10013 8812 10047
rect 8760 10004 8812 10013
rect 10140 10047 10192 10056
rect 10140 10013 10158 10047
rect 10158 10013 10192 10047
rect 10416 10047 10468 10056
rect 10140 10004 10192 10013
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 10968 10004 11020 10056
rect 12532 10004 12584 10056
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 14188 10004 14240 10056
rect 16028 10004 16080 10056
rect 16672 10004 16724 10056
rect 17408 10047 17460 10056
rect 9128 9936 9180 9988
rect 9588 9936 9640 9988
rect 14096 9979 14148 9988
rect 14096 9945 14105 9979
rect 14105 9945 14139 9979
rect 14139 9945 14148 9979
rect 14096 9936 14148 9945
rect 14372 9936 14424 9988
rect 14740 9936 14792 9988
rect 15752 9979 15804 9988
rect 15752 9945 15761 9979
rect 15761 9945 15795 9979
rect 15795 9945 15804 9979
rect 15752 9936 15804 9945
rect 2964 9868 3016 9920
rect 5632 9868 5684 9920
rect 8944 9868 8996 9920
rect 13268 9911 13320 9920
rect 13268 9877 13277 9911
rect 13277 9877 13311 9911
rect 13311 9877 13320 9911
rect 13268 9868 13320 9877
rect 13820 9911 13872 9920
rect 13820 9877 13829 9911
rect 13829 9877 13863 9911
rect 13863 9877 13872 9911
rect 13820 9868 13872 9877
rect 15292 9911 15344 9920
rect 15292 9877 15301 9911
rect 15301 9877 15335 9911
rect 15335 9877 15344 9911
rect 15292 9868 15344 9877
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 17592 10004 17644 10056
rect 17868 10004 17920 10056
rect 19064 10004 19116 10056
rect 19616 10047 19668 10056
rect 19616 10013 19625 10047
rect 19625 10013 19659 10047
rect 19659 10013 19668 10047
rect 19616 10004 19668 10013
rect 19892 10004 19944 10056
rect 20996 10004 21048 10056
rect 22744 10072 22796 10124
rect 23296 10115 23348 10124
rect 23296 10081 23305 10115
rect 23305 10081 23339 10115
rect 23339 10081 23348 10115
rect 23296 10072 23348 10081
rect 21732 10047 21784 10056
rect 21732 10013 21741 10047
rect 21741 10013 21775 10047
rect 21775 10013 21784 10047
rect 21732 10004 21784 10013
rect 22284 10047 22336 10056
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 17684 9936 17736 9988
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 17592 9868 17644 9920
rect 20720 9911 20772 9920
rect 20720 9877 20729 9911
rect 20729 9877 20763 9911
rect 20763 9877 20772 9911
rect 20720 9868 20772 9877
rect 22376 9868 22428 9920
rect 22744 9911 22796 9920
rect 22744 9877 22753 9911
rect 22753 9877 22787 9911
rect 22787 9877 22796 9911
rect 22744 9868 22796 9877
rect 23296 9868 23348 9920
rect 9322 9766 9374 9818
rect 9386 9766 9438 9818
rect 9450 9766 9502 9818
rect 9514 9766 9566 9818
rect 9578 9766 9630 9818
rect 17694 9766 17746 9818
rect 17758 9766 17810 9818
rect 17822 9766 17874 9818
rect 17886 9766 17938 9818
rect 17950 9766 18002 9818
rect 2504 9707 2556 9716
rect 2504 9673 2513 9707
rect 2513 9673 2547 9707
rect 2547 9673 2556 9707
rect 2504 9664 2556 9673
rect 2872 9596 2924 9648
rect 3424 9596 3476 9648
rect 7380 9596 7432 9648
rect 8484 9596 8536 9648
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 3056 9571 3108 9580
rect 2780 9528 2832 9537
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 4620 9528 4672 9580
rect 8944 9528 8996 9580
rect 10416 9528 10468 9580
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 11152 9571 11204 9580
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 4160 9460 4212 9512
rect 4804 9460 4856 9512
rect 3240 9392 3292 9444
rect 6092 9392 6144 9444
rect 10784 9435 10836 9444
rect 3700 9324 3752 9376
rect 3884 9324 3936 9376
rect 3976 9324 4028 9376
rect 8300 9324 8352 9376
rect 10784 9401 10793 9435
rect 10793 9401 10827 9435
rect 10827 9401 10836 9435
rect 10784 9392 10836 9401
rect 11152 9537 11161 9571
rect 11161 9537 11195 9571
rect 11195 9537 11204 9571
rect 11152 9528 11204 9537
rect 12440 9596 12492 9648
rect 15292 9664 15344 9716
rect 16580 9664 16632 9716
rect 12624 9596 12676 9648
rect 13176 9596 13228 9648
rect 12348 9528 12400 9580
rect 14188 9596 14240 9648
rect 15752 9596 15804 9648
rect 16028 9639 16080 9648
rect 16028 9605 16037 9639
rect 16037 9605 16071 9639
rect 16071 9605 16080 9639
rect 16028 9596 16080 9605
rect 17408 9664 17460 9716
rect 18236 9664 18288 9716
rect 18972 9707 19024 9716
rect 18972 9673 18981 9707
rect 18981 9673 19015 9707
rect 19015 9673 19024 9707
rect 18972 9664 19024 9673
rect 19432 9707 19484 9716
rect 19432 9673 19441 9707
rect 19441 9673 19475 9707
rect 19475 9673 19484 9707
rect 19432 9664 19484 9673
rect 20812 9707 20864 9716
rect 20812 9673 20821 9707
rect 20821 9673 20855 9707
rect 20855 9673 20864 9707
rect 20812 9664 20864 9673
rect 22560 9664 22612 9716
rect 22744 9664 22796 9716
rect 23112 9707 23164 9716
rect 23112 9673 23121 9707
rect 23121 9673 23155 9707
rect 23155 9673 23164 9707
rect 23112 9664 23164 9673
rect 17500 9596 17552 9648
rect 18604 9596 18656 9648
rect 20076 9596 20128 9648
rect 20260 9596 20312 9648
rect 22468 9596 22520 9648
rect 23204 9596 23256 9648
rect 13820 9528 13872 9580
rect 12716 9460 12768 9512
rect 13084 9460 13136 9512
rect 13544 9460 13596 9512
rect 14096 9503 14148 9512
rect 14096 9469 14105 9503
rect 14105 9469 14139 9503
rect 14139 9469 14148 9503
rect 14096 9460 14148 9469
rect 12808 9392 12860 9444
rect 14740 9460 14792 9512
rect 15016 9503 15068 9512
rect 15016 9469 15025 9503
rect 15025 9469 15059 9503
rect 15059 9469 15068 9503
rect 15016 9460 15068 9469
rect 15752 9460 15804 9512
rect 17316 9528 17368 9580
rect 19064 9571 19116 9580
rect 19064 9537 19073 9571
rect 19073 9537 19107 9571
rect 19107 9537 19116 9571
rect 19064 9528 19116 9537
rect 17408 9503 17460 9512
rect 17408 9469 17417 9503
rect 17417 9469 17451 9503
rect 17451 9469 17460 9503
rect 17408 9460 17460 9469
rect 18144 9503 18196 9512
rect 18144 9469 18153 9503
rect 18153 9469 18187 9503
rect 18187 9469 18196 9503
rect 18144 9460 18196 9469
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 20996 9503 21048 9512
rect 20996 9469 21005 9503
rect 21005 9469 21039 9503
rect 21039 9469 21048 9503
rect 20996 9460 21048 9469
rect 20352 9392 20404 9444
rect 13360 9324 13412 9376
rect 14372 9324 14424 9376
rect 14464 9324 14516 9376
rect 15568 9367 15620 9376
rect 15568 9333 15577 9367
rect 15577 9333 15611 9367
rect 15611 9333 15620 9367
rect 15568 9324 15620 9333
rect 15752 9324 15804 9376
rect 16304 9324 16356 9376
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 19616 9367 19668 9376
rect 19616 9333 19625 9367
rect 19625 9333 19659 9367
rect 19659 9333 19668 9367
rect 19616 9324 19668 9333
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 21732 9324 21784 9376
rect 22652 9367 22704 9376
rect 22652 9333 22661 9367
rect 22661 9333 22695 9367
rect 22695 9333 22704 9367
rect 22652 9324 22704 9333
rect 23480 9324 23532 9376
rect 5136 9222 5188 9274
rect 5200 9222 5252 9274
rect 5264 9222 5316 9274
rect 5328 9222 5380 9274
rect 5392 9222 5444 9274
rect 13508 9222 13560 9274
rect 13572 9222 13624 9274
rect 13636 9222 13688 9274
rect 13700 9222 13752 9274
rect 13764 9222 13816 9274
rect 21880 9222 21932 9274
rect 21944 9222 21996 9274
rect 22008 9222 22060 9274
rect 22072 9222 22124 9274
rect 22136 9222 22188 9274
rect 3056 9120 3108 9172
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 3884 9163 3936 9172
rect 3884 9129 3893 9163
rect 3893 9129 3927 9163
rect 3927 9129 3936 9163
rect 3884 9120 3936 9129
rect 5540 9120 5592 9172
rect 6092 9120 6144 9172
rect 7840 9163 7892 9172
rect 7840 9129 7849 9163
rect 7849 9129 7883 9163
rect 7883 9129 7892 9163
rect 7840 9120 7892 9129
rect 12532 9120 12584 9172
rect 13360 9120 13412 9172
rect 15200 9120 15252 9172
rect 16304 9120 16356 9172
rect 17408 9120 17460 9172
rect 18144 9120 18196 9172
rect 20076 9120 20128 9172
rect 22928 9120 22980 9172
rect 2780 8984 2832 9036
rect 4068 9052 4120 9104
rect 12348 9095 12400 9104
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 4344 8984 4396 9036
rect 12348 9061 12357 9095
rect 12357 9061 12391 9095
rect 12391 9061 12400 9095
rect 12348 9052 12400 9061
rect 12716 9095 12768 9104
rect 12716 9061 12725 9095
rect 12725 9061 12759 9095
rect 12759 9061 12768 9095
rect 12716 9052 12768 9061
rect 12808 9052 12860 9104
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 4620 8916 4672 8968
rect 4988 8916 5040 8968
rect 6184 8959 6236 8968
rect 6184 8925 6193 8959
rect 6193 8925 6227 8959
rect 6227 8925 6236 8959
rect 6184 8916 6236 8925
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 7840 8916 7892 8968
rect 11152 8916 11204 8968
rect 5632 8848 5684 8900
rect 8392 8848 8444 8900
rect 12072 8848 12124 8900
rect 12440 8916 12492 8968
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 12808 8959 12860 8968
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 14648 9027 14700 9036
rect 14648 8993 14657 9027
rect 14657 8993 14691 9027
rect 14691 8993 14700 9027
rect 14648 8984 14700 8993
rect 15016 8984 15068 9036
rect 19892 9027 19944 9036
rect 19892 8993 19901 9027
rect 19901 8993 19935 9027
rect 19935 8993 19944 9027
rect 19892 8984 19944 8993
rect 20352 8984 20404 9036
rect 13728 8916 13780 8968
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 14740 8916 14792 8968
rect 17316 8916 17368 8968
rect 18604 8916 18656 8968
rect 19616 8959 19668 8968
rect 19616 8925 19625 8959
rect 19625 8925 19659 8959
rect 19659 8925 19668 8959
rect 19616 8916 19668 8925
rect 20260 8959 20312 8968
rect 20260 8925 20269 8959
rect 20269 8925 20303 8959
rect 20303 8925 20312 8959
rect 20260 8916 20312 8925
rect 2688 8780 2740 8832
rect 2872 8780 2924 8832
rect 3332 8780 3384 8832
rect 3608 8780 3660 8832
rect 4896 8780 4948 8832
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 11704 8823 11756 8832
rect 11704 8789 11713 8823
rect 11713 8789 11747 8823
rect 11747 8789 11756 8823
rect 11704 8780 11756 8789
rect 13268 8780 13320 8832
rect 17592 8848 17644 8900
rect 19892 8848 19944 8900
rect 20996 8848 21048 8900
rect 22836 8959 22888 8968
rect 22836 8925 22845 8959
rect 22845 8925 22879 8959
rect 22879 8925 22888 8959
rect 22836 8916 22888 8925
rect 23204 8916 23256 8968
rect 23480 8959 23532 8968
rect 23480 8925 23489 8959
rect 23489 8925 23523 8959
rect 23523 8925 23532 8959
rect 23480 8916 23532 8925
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 16396 8780 16448 8832
rect 18052 8780 18104 8832
rect 19248 8823 19300 8832
rect 19248 8789 19257 8823
rect 19257 8789 19291 8823
rect 19291 8789 19300 8823
rect 19248 8780 19300 8789
rect 22468 8823 22520 8832
rect 22468 8789 22477 8823
rect 22477 8789 22511 8823
rect 22511 8789 22520 8823
rect 22468 8780 22520 8789
rect 9322 8678 9374 8730
rect 9386 8678 9438 8730
rect 9450 8678 9502 8730
rect 9514 8678 9566 8730
rect 9578 8678 9630 8730
rect 17694 8678 17746 8730
rect 17758 8678 17810 8730
rect 17822 8678 17874 8730
rect 17886 8678 17938 8730
rect 17950 8678 18002 8730
rect 2964 8576 3016 8628
rect 4620 8576 4672 8628
rect 6000 8619 6052 8628
rect 6000 8585 6009 8619
rect 6009 8585 6043 8619
rect 6043 8585 6052 8619
rect 6000 8576 6052 8585
rect 7564 8576 7616 8628
rect 9220 8576 9272 8628
rect 10784 8576 10836 8628
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12808 8619 12860 8628
rect 12440 8576 12492 8585
rect 12808 8585 12817 8619
rect 12817 8585 12851 8619
rect 12851 8585 12860 8619
rect 12808 8576 12860 8585
rect 13084 8619 13136 8628
rect 13084 8585 13093 8619
rect 13093 8585 13127 8619
rect 13127 8585 13136 8619
rect 13084 8576 13136 8585
rect 15384 8576 15436 8628
rect 17408 8576 17460 8628
rect 19892 8576 19944 8628
rect 2688 8483 2740 8492
rect 2688 8449 2706 8483
rect 2706 8449 2740 8483
rect 2688 8440 2740 8449
rect 3608 8440 3660 8492
rect 3884 8440 3936 8492
rect 4712 8440 4764 8492
rect 5724 8440 5776 8492
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 8484 8508 8536 8560
rect 7380 8483 7432 8492
rect 7380 8449 7414 8483
rect 7414 8449 7432 8483
rect 7380 8440 7432 8449
rect 8760 8440 8812 8492
rect 9772 8508 9824 8560
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 11796 8440 11848 8492
rect 6552 8415 6604 8424
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 11980 8372 12032 8424
rect 5632 8304 5684 8356
rect 6920 8279 6972 8288
rect 6920 8245 6929 8279
rect 6929 8245 6963 8279
rect 6963 8245 6972 8279
rect 6920 8236 6972 8245
rect 8300 8304 8352 8356
rect 8852 8347 8904 8356
rect 8852 8313 8861 8347
rect 8861 8313 8895 8347
rect 8895 8313 8904 8347
rect 8852 8304 8904 8313
rect 9036 8236 9088 8288
rect 11612 8236 11664 8288
rect 12256 8440 12308 8492
rect 13176 8508 13228 8560
rect 12164 8372 12216 8424
rect 13728 8440 13780 8492
rect 14372 8440 14424 8492
rect 12256 8279 12308 8288
rect 12256 8245 12265 8279
rect 12265 8245 12299 8279
rect 12299 8245 12308 8279
rect 12256 8236 12308 8245
rect 13084 8236 13136 8288
rect 13360 8236 13412 8288
rect 14188 8279 14240 8288
rect 14188 8245 14197 8279
rect 14197 8245 14231 8279
rect 14231 8245 14240 8279
rect 14188 8236 14240 8245
rect 14648 8279 14700 8288
rect 14648 8245 14657 8279
rect 14657 8245 14691 8279
rect 14691 8245 14700 8279
rect 14648 8236 14700 8245
rect 16120 8279 16172 8288
rect 16120 8245 16129 8279
rect 16129 8245 16163 8279
rect 16163 8245 16172 8279
rect 16120 8236 16172 8245
rect 22284 8236 22336 8288
rect 5136 8134 5188 8186
rect 5200 8134 5252 8186
rect 5264 8134 5316 8186
rect 5328 8134 5380 8186
rect 5392 8134 5444 8186
rect 13508 8134 13560 8186
rect 13572 8134 13624 8186
rect 13636 8134 13688 8186
rect 13700 8134 13752 8186
rect 13764 8134 13816 8186
rect 21880 8134 21932 8186
rect 21944 8134 21996 8186
rect 22008 8134 22060 8186
rect 22072 8134 22124 8186
rect 22136 8134 22188 8186
rect 4712 8032 4764 8084
rect 4988 8032 5040 8084
rect 6552 8032 6604 8084
rect 6920 8032 6972 8084
rect 8392 8032 8444 8084
rect 8944 8032 8996 8084
rect 9772 8075 9824 8084
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 4160 7964 4212 8016
rect 6736 7964 6788 8016
rect 2780 7760 2832 7812
rect 3700 7828 3752 7880
rect 4344 7871 4396 7880
rect 4344 7837 4358 7871
rect 4358 7837 4392 7871
rect 4392 7837 4396 7871
rect 4988 7871 5040 7880
rect 4344 7828 4396 7837
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 6000 7896 6052 7948
rect 7012 7939 7064 7948
rect 7012 7905 7021 7939
rect 7021 7905 7055 7939
rect 7055 7905 7064 7939
rect 7472 7964 7524 8016
rect 8760 7964 8812 8016
rect 9036 8007 9088 8016
rect 9036 7973 9045 8007
rect 9045 7973 9079 8007
rect 9079 7973 9088 8007
rect 9036 7964 9088 7973
rect 7012 7896 7064 7905
rect 8852 7896 8904 7948
rect 9772 8041 9781 8075
rect 9781 8041 9815 8075
rect 9815 8041 9824 8075
rect 9772 8032 9824 8041
rect 9864 7964 9916 8016
rect 11980 8032 12032 8084
rect 13084 8032 13136 8084
rect 18236 8032 18288 8084
rect 10508 7964 10560 8016
rect 12624 7964 12676 8016
rect 13360 7964 13412 8016
rect 9404 7896 9456 7948
rect 5724 7828 5776 7880
rect 5908 7828 5960 7880
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 7748 7828 7800 7880
rect 8668 7871 8720 7880
rect 6000 7803 6052 7812
rect 3240 7692 3292 7744
rect 6000 7769 6009 7803
rect 6009 7769 6043 7803
rect 6043 7769 6052 7803
rect 6000 7760 6052 7769
rect 6736 7760 6788 7812
rect 5540 7692 5592 7744
rect 5724 7735 5776 7744
rect 5724 7701 5733 7735
rect 5733 7701 5767 7735
rect 5767 7701 5776 7735
rect 5724 7692 5776 7701
rect 5816 7692 5868 7744
rect 8668 7837 8677 7871
rect 8677 7837 8711 7871
rect 8711 7837 8720 7871
rect 8668 7828 8720 7837
rect 8944 7828 8996 7880
rect 9036 7828 9088 7880
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 12164 7828 12216 7880
rect 13176 7896 13228 7948
rect 14280 7896 14332 7948
rect 14648 7939 14700 7948
rect 14648 7905 14657 7939
rect 14657 7905 14691 7939
rect 14691 7905 14700 7939
rect 14648 7896 14700 7905
rect 16120 7896 16172 7948
rect 20352 7896 20404 7948
rect 22284 7964 22336 8016
rect 21640 7896 21692 7948
rect 9404 7760 9456 7812
rect 9680 7760 9732 7812
rect 12256 7760 12308 7812
rect 14188 7828 14240 7880
rect 15384 7828 15436 7880
rect 16856 7828 16908 7880
rect 17224 7871 17276 7880
rect 17224 7837 17234 7871
rect 17234 7837 17268 7871
rect 17268 7837 17276 7871
rect 17224 7828 17276 7837
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 18328 7828 18380 7880
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 22468 7828 22520 7880
rect 16488 7760 16540 7812
rect 11704 7692 11756 7744
rect 12624 7692 12676 7744
rect 14924 7735 14976 7744
rect 14924 7701 14933 7735
rect 14933 7701 14967 7735
rect 14967 7701 14976 7735
rect 14924 7692 14976 7701
rect 15384 7735 15436 7744
rect 15384 7701 15393 7735
rect 15393 7701 15427 7735
rect 15427 7701 15436 7735
rect 15936 7735 15988 7744
rect 15384 7692 15436 7701
rect 15936 7701 15945 7735
rect 15945 7701 15979 7735
rect 15979 7701 15988 7735
rect 15936 7692 15988 7701
rect 16212 7735 16264 7744
rect 16212 7701 16221 7735
rect 16221 7701 16255 7735
rect 16255 7701 16264 7735
rect 16212 7692 16264 7701
rect 16396 7692 16448 7744
rect 19432 7760 19484 7812
rect 22284 7760 22336 7812
rect 18420 7692 18472 7744
rect 22100 7735 22152 7744
rect 22100 7701 22109 7735
rect 22109 7701 22143 7735
rect 22143 7701 22152 7735
rect 22100 7692 22152 7701
rect 22192 7735 22244 7744
rect 22192 7701 22201 7735
rect 22201 7701 22235 7735
rect 22235 7701 22244 7735
rect 22192 7692 22244 7701
rect 22928 7692 22980 7744
rect 23204 7735 23256 7744
rect 23204 7701 23213 7735
rect 23213 7701 23247 7735
rect 23247 7701 23256 7735
rect 23204 7692 23256 7701
rect 9322 7590 9374 7642
rect 9386 7590 9438 7642
rect 9450 7590 9502 7642
rect 9514 7590 9566 7642
rect 9578 7590 9630 7642
rect 17694 7590 17746 7642
rect 17758 7590 17810 7642
rect 17822 7590 17874 7642
rect 17886 7590 17938 7642
rect 17950 7590 18002 7642
rect 4160 7488 4212 7540
rect 5724 7488 5776 7540
rect 5908 7420 5960 7472
rect 6368 7463 6420 7472
rect 6368 7429 6377 7463
rect 6377 7429 6411 7463
rect 6411 7429 6420 7463
rect 6368 7420 6420 7429
rect 3240 7352 3292 7404
rect 3884 7352 3936 7404
rect 7380 7420 7432 7472
rect 7748 7463 7800 7472
rect 7196 7352 7248 7404
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 7748 7429 7757 7463
rect 7757 7429 7791 7463
rect 7791 7429 7800 7463
rect 7748 7420 7800 7429
rect 8392 7488 8444 7540
rect 8484 7463 8536 7472
rect 8484 7429 8493 7463
rect 8493 7429 8527 7463
rect 8527 7429 8536 7463
rect 8484 7420 8536 7429
rect 8760 7395 8812 7404
rect 8760 7361 8769 7395
rect 8769 7361 8803 7395
rect 8803 7361 8812 7395
rect 8760 7352 8812 7361
rect 9220 7488 9272 7540
rect 11888 7488 11940 7540
rect 15108 7488 15160 7540
rect 15476 7488 15528 7540
rect 18236 7531 18288 7540
rect 7748 7284 7800 7336
rect 8024 7284 8076 7336
rect 8668 7284 8720 7336
rect 9036 7284 9088 7336
rect 9220 7284 9272 7336
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 15016 7420 15068 7472
rect 9680 7352 9732 7361
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 12072 7395 12124 7404
rect 12072 7361 12081 7395
rect 12081 7361 12115 7395
rect 12115 7361 12124 7395
rect 12072 7352 12124 7361
rect 13912 7352 13964 7404
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14280 7395 14332 7404
rect 14004 7352 14056 7361
rect 14280 7361 14314 7395
rect 14314 7361 14332 7395
rect 14280 7352 14332 7361
rect 14832 7352 14884 7404
rect 16396 7420 16448 7472
rect 18236 7497 18245 7531
rect 18245 7497 18279 7531
rect 18279 7497 18288 7531
rect 18236 7488 18288 7497
rect 19248 7488 19300 7540
rect 19432 7531 19484 7540
rect 19432 7497 19450 7531
rect 19450 7497 19484 7531
rect 19432 7488 19484 7497
rect 20444 7488 20496 7540
rect 20996 7488 21048 7540
rect 21824 7488 21876 7540
rect 23204 7463 23256 7472
rect 23204 7429 23238 7463
rect 23238 7429 23256 7463
rect 23204 7420 23256 7429
rect 20720 7352 20772 7404
rect 20996 7395 21048 7404
rect 20996 7361 21005 7395
rect 21005 7361 21039 7395
rect 21039 7361 21048 7395
rect 20996 7352 21048 7361
rect 21640 7395 21692 7404
rect 21640 7361 21649 7395
rect 21649 7361 21683 7395
rect 21683 7361 21692 7395
rect 21640 7352 21692 7361
rect 21824 7395 21876 7404
rect 21824 7361 21833 7395
rect 21833 7361 21867 7395
rect 21867 7361 21876 7395
rect 21824 7352 21876 7361
rect 23020 7352 23072 7404
rect 12256 7284 12308 7336
rect 15016 7284 15068 7336
rect 18512 7284 18564 7336
rect 18880 7327 18932 7336
rect 18880 7293 18889 7327
rect 18889 7293 18923 7327
rect 18923 7293 18932 7327
rect 20352 7327 20404 7336
rect 18880 7284 18932 7293
rect 20352 7293 20361 7327
rect 20361 7293 20395 7327
rect 20395 7293 20404 7327
rect 20352 7284 20404 7293
rect 8116 7259 8168 7268
rect 8116 7225 8125 7259
rect 8125 7225 8159 7259
rect 8159 7225 8168 7259
rect 8116 7216 8168 7225
rect 9772 7216 9824 7268
rect 11244 7216 11296 7268
rect 11612 7216 11664 7268
rect 7012 7148 7064 7200
rect 8944 7148 8996 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 12072 7148 12124 7200
rect 14280 7148 14332 7200
rect 15292 7148 15344 7200
rect 16212 7148 16264 7200
rect 17040 7148 17092 7200
rect 17592 7148 17644 7200
rect 19524 7148 19576 7200
rect 22192 7284 22244 7336
rect 22100 7216 22152 7268
rect 22744 7191 22796 7200
rect 22744 7157 22753 7191
rect 22753 7157 22787 7191
rect 22787 7157 22796 7191
rect 22744 7148 22796 7157
rect 23848 7148 23900 7200
rect 5136 7046 5188 7098
rect 5200 7046 5252 7098
rect 5264 7046 5316 7098
rect 5328 7046 5380 7098
rect 5392 7046 5444 7098
rect 13508 7046 13560 7098
rect 13572 7046 13624 7098
rect 13636 7046 13688 7098
rect 13700 7046 13752 7098
rect 13764 7046 13816 7098
rect 21880 7046 21932 7098
rect 21944 7046 21996 7098
rect 22008 7046 22060 7098
rect 22072 7046 22124 7098
rect 22136 7046 22188 7098
rect 6736 6987 6788 6996
rect 6736 6953 6745 6987
rect 6745 6953 6779 6987
rect 6779 6953 6788 6987
rect 6736 6944 6788 6953
rect 7748 6944 7800 6996
rect 11520 6944 11572 6996
rect 12900 6944 12952 6996
rect 13912 6944 13964 6996
rect 14924 6944 14976 6996
rect 15108 6944 15160 6996
rect 17316 6944 17368 6996
rect 19432 6987 19484 6996
rect 19432 6953 19441 6987
rect 19441 6953 19475 6987
rect 19475 6953 19484 6987
rect 19432 6944 19484 6953
rect 22928 6944 22980 6996
rect 7840 6876 7892 6928
rect 14648 6876 14700 6928
rect 15476 6876 15528 6928
rect 16764 6919 16816 6928
rect 16764 6885 16773 6919
rect 16773 6885 16807 6919
rect 16807 6885 16816 6919
rect 16764 6876 16816 6885
rect 17224 6876 17276 6928
rect 6828 6808 6880 6860
rect 8116 6808 8168 6860
rect 14004 6808 14056 6860
rect 15384 6808 15436 6860
rect 15936 6808 15988 6860
rect 6000 6740 6052 6792
rect 7472 6740 7524 6792
rect 8852 6740 8904 6792
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 11152 6740 11204 6792
rect 11336 6740 11388 6792
rect 12256 6783 12308 6792
rect 12256 6749 12265 6783
rect 12265 6749 12299 6783
rect 12299 6749 12308 6783
rect 12256 6740 12308 6749
rect 12532 6783 12584 6792
rect 12532 6749 12541 6783
rect 12541 6749 12575 6783
rect 12575 6749 12584 6783
rect 12532 6740 12584 6749
rect 7196 6672 7248 6724
rect 6920 6604 6972 6656
rect 7564 6604 7616 6656
rect 8300 6672 8352 6724
rect 10048 6672 10100 6724
rect 11796 6672 11848 6724
rect 13084 6740 13136 6792
rect 13268 6740 13320 6792
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 8760 6604 8812 6656
rect 10508 6604 10560 6656
rect 10968 6604 11020 6656
rect 14648 6672 14700 6724
rect 14832 6672 14884 6724
rect 16764 6740 16816 6792
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 17132 6783 17184 6792
rect 17132 6749 17141 6783
rect 17141 6749 17175 6783
rect 17175 6749 17184 6783
rect 17132 6740 17184 6749
rect 18420 6715 18472 6724
rect 18420 6681 18438 6715
rect 18438 6681 18472 6715
rect 18420 6672 18472 6681
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 19340 6672 19392 6724
rect 23020 6740 23072 6792
rect 23480 6783 23532 6792
rect 23480 6749 23489 6783
rect 23489 6749 23532 6783
rect 23480 6740 23532 6749
rect 23756 6783 23808 6792
rect 23756 6749 23765 6783
rect 23765 6749 23799 6783
rect 23799 6749 23808 6783
rect 23756 6740 23808 6749
rect 19616 6672 19668 6724
rect 22744 6672 22796 6724
rect 17316 6647 17368 6656
rect 17316 6613 17325 6647
rect 17325 6613 17359 6647
rect 17359 6613 17368 6647
rect 17316 6604 17368 6613
rect 21180 6604 21232 6656
rect 21732 6647 21784 6656
rect 21732 6613 21741 6647
rect 21741 6613 21775 6647
rect 21775 6613 21784 6647
rect 21732 6604 21784 6613
rect 23388 6604 23440 6656
rect 9322 6502 9374 6554
rect 9386 6502 9438 6554
rect 9450 6502 9502 6554
rect 9514 6502 9566 6554
rect 9578 6502 9630 6554
rect 17694 6502 17746 6554
rect 17758 6502 17810 6554
rect 17822 6502 17874 6554
rect 17886 6502 17938 6554
rect 17950 6502 18002 6554
rect 5632 6400 5684 6452
rect 6828 6400 6880 6452
rect 7012 6443 7064 6452
rect 7012 6409 7021 6443
rect 7021 6409 7055 6443
rect 7055 6409 7064 6443
rect 7012 6400 7064 6409
rect 8024 6400 8076 6452
rect 9128 6400 9180 6452
rect 10876 6400 10928 6452
rect 11060 6400 11112 6452
rect 13084 6400 13136 6452
rect 15016 6400 15068 6452
rect 6184 6332 6236 6384
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 6828 6264 6880 6316
rect 7932 6332 7984 6384
rect 8208 6375 8260 6384
rect 8208 6341 8217 6375
rect 8217 6341 8251 6375
rect 8251 6341 8260 6375
rect 8208 6332 8260 6341
rect 8944 6332 8996 6384
rect 9220 6332 9272 6384
rect 10140 6332 10192 6384
rect 7472 6264 7524 6316
rect 7564 6264 7616 6316
rect 8116 6264 8168 6316
rect 10508 6264 10560 6316
rect 10692 6264 10744 6316
rect 11244 6264 11296 6316
rect 15936 6332 15988 6384
rect 18512 6375 18564 6384
rect 18512 6341 18521 6375
rect 18521 6341 18555 6375
rect 18555 6341 18564 6375
rect 18512 6332 18564 6341
rect 19616 6400 19668 6452
rect 20720 6443 20772 6452
rect 20720 6409 20729 6443
rect 20729 6409 20763 6443
rect 20763 6409 20772 6443
rect 20720 6400 20772 6409
rect 21732 6400 21784 6452
rect 22100 6332 22152 6384
rect 23480 6375 23532 6384
rect 17316 6264 17368 6316
rect 18328 6307 18380 6316
rect 9220 6196 9272 6248
rect 5816 6128 5868 6180
rect 8760 6128 8812 6180
rect 11520 6171 11572 6180
rect 11520 6137 11529 6171
rect 11529 6137 11563 6171
rect 11563 6137 11572 6171
rect 11520 6128 11572 6137
rect 12348 6196 12400 6248
rect 17132 6196 17184 6248
rect 18328 6273 18336 6307
rect 18336 6273 18370 6307
rect 18370 6273 18380 6307
rect 18328 6264 18380 6273
rect 19524 6264 19576 6316
rect 19616 6264 19668 6316
rect 20904 6307 20956 6316
rect 20904 6273 20913 6307
rect 20913 6273 20956 6307
rect 20904 6264 20956 6273
rect 23480 6341 23489 6375
rect 23489 6341 23523 6375
rect 23523 6341 23532 6375
rect 23480 6332 23532 6341
rect 21180 6239 21232 6248
rect 16672 6128 16724 6180
rect 21180 6205 21189 6239
rect 21189 6205 21223 6239
rect 21223 6205 21232 6239
rect 21180 6196 21232 6205
rect 22284 6196 22336 6248
rect 23388 6307 23440 6316
rect 23388 6273 23397 6307
rect 23397 6273 23431 6307
rect 23431 6273 23440 6307
rect 23388 6264 23440 6273
rect 23756 6264 23808 6316
rect 6644 6060 6696 6112
rect 7472 6060 7524 6112
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 8116 6103 8168 6112
rect 8116 6069 8125 6103
rect 8125 6069 8159 6103
rect 8159 6069 8168 6103
rect 8116 6060 8168 6069
rect 10048 6060 10100 6112
rect 12532 6060 12584 6112
rect 20720 6060 20772 6112
rect 20996 6060 21048 6112
rect 23480 6060 23532 6112
rect 5136 5958 5188 6010
rect 5200 5958 5252 6010
rect 5264 5958 5316 6010
rect 5328 5958 5380 6010
rect 5392 5958 5444 6010
rect 13508 5958 13560 6010
rect 13572 5958 13624 6010
rect 13636 5958 13688 6010
rect 13700 5958 13752 6010
rect 13764 5958 13816 6010
rect 21880 5958 21932 6010
rect 21944 5958 21996 6010
rect 22008 5958 22060 6010
rect 22072 5958 22124 6010
rect 22136 5958 22188 6010
rect 4804 5856 4856 5908
rect 5724 5856 5776 5908
rect 6184 5856 6236 5908
rect 5264 5788 5316 5840
rect 8668 5856 8720 5908
rect 6644 5720 6696 5772
rect 7472 5788 7524 5840
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 7196 5720 7248 5772
rect 5356 5695 5408 5704
rect 5356 5661 5365 5695
rect 5365 5661 5399 5695
rect 5399 5661 5408 5695
rect 5356 5652 5408 5661
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 6368 5584 6420 5636
rect 6552 5584 6604 5636
rect 7564 5652 7616 5704
rect 8208 5788 8260 5840
rect 8760 5788 8812 5840
rect 8116 5720 8168 5772
rect 8300 5652 8352 5704
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 23480 5856 23532 5908
rect 12164 5720 12216 5772
rect 21364 5720 21416 5772
rect 10692 5652 10744 5704
rect 12808 5652 12860 5704
rect 19248 5652 19300 5704
rect 21732 5652 21784 5704
rect 8852 5584 8904 5636
rect 6644 5559 6696 5568
rect 6644 5525 6653 5559
rect 6653 5525 6687 5559
rect 6687 5525 6696 5559
rect 6644 5516 6696 5525
rect 6828 5516 6880 5568
rect 8300 5516 8352 5568
rect 10416 5516 10468 5568
rect 11704 5584 11756 5636
rect 20904 5584 20956 5636
rect 12348 5516 12400 5568
rect 13820 5559 13872 5568
rect 13820 5525 13829 5559
rect 13829 5525 13863 5559
rect 13863 5525 13872 5559
rect 13820 5516 13872 5525
rect 18788 5559 18840 5568
rect 18788 5525 18797 5559
rect 18797 5525 18831 5559
rect 18831 5525 18840 5559
rect 18788 5516 18840 5525
rect 21456 5516 21508 5568
rect 9322 5414 9374 5466
rect 9386 5414 9438 5466
rect 9450 5414 9502 5466
rect 9514 5414 9566 5466
rect 9578 5414 9630 5466
rect 17694 5414 17746 5466
rect 17758 5414 17810 5466
rect 17822 5414 17874 5466
rect 17886 5414 17938 5466
rect 17950 5414 18002 5466
rect 5356 5312 5408 5364
rect 6276 5312 6328 5364
rect 6368 5312 6420 5364
rect 7564 5312 7616 5364
rect 3884 5244 3936 5296
rect 3700 5219 3752 5228
rect 3700 5185 3734 5219
rect 3734 5185 3752 5219
rect 6644 5244 6696 5296
rect 6920 5244 6972 5296
rect 3700 5176 3752 5185
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 5908 5176 5960 5228
rect 6276 5176 6328 5228
rect 6828 5176 6880 5228
rect 7196 5244 7248 5296
rect 9036 5312 9088 5364
rect 7380 5219 7432 5228
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7656 5219 7708 5228
rect 7472 5176 7524 5185
rect 7656 5185 7663 5219
rect 7663 5185 7708 5219
rect 7656 5176 7708 5185
rect 4988 5108 5040 5160
rect 5632 5151 5684 5160
rect 5632 5117 5641 5151
rect 5641 5117 5675 5151
rect 5675 5117 5684 5151
rect 5632 5108 5684 5117
rect 6644 5108 6696 5160
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 4436 5040 4488 5092
rect 7288 5108 7340 5160
rect 10140 5244 10192 5296
rect 13360 5312 13412 5364
rect 14096 5312 14148 5364
rect 15568 5312 15620 5364
rect 18052 5312 18104 5364
rect 18880 5355 18932 5364
rect 18880 5321 18889 5355
rect 18889 5321 18923 5355
rect 18923 5321 18932 5355
rect 18880 5312 18932 5321
rect 19800 5312 19852 5364
rect 20996 5355 21048 5364
rect 20996 5321 21005 5355
rect 21005 5321 21039 5355
rect 21039 5321 21048 5355
rect 20996 5312 21048 5321
rect 22652 5312 22704 5364
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 8208 5176 8260 5228
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 9220 5176 9272 5228
rect 10048 5219 10100 5228
rect 10048 5185 10057 5219
rect 10057 5185 10091 5219
rect 10091 5185 10100 5219
rect 10048 5176 10100 5185
rect 8392 5151 8444 5160
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 7748 5040 7800 5092
rect 7932 5040 7984 5092
rect 6644 4972 6696 5024
rect 8116 5015 8168 5024
rect 8116 4981 8125 5015
rect 8125 4981 8159 5015
rect 8159 4981 8168 5015
rect 8116 4972 8168 4981
rect 8852 5040 8904 5092
rect 11152 5244 11204 5296
rect 10692 5176 10744 5228
rect 11888 5176 11940 5228
rect 11336 5108 11388 5160
rect 14096 5176 14148 5228
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 12808 5040 12860 5092
rect 15476 5040 15528 5092
rect 16212 5108 16264 5160
rect 17224 5151 17276 5160
rect 17224 5117 17233 5151
rect 17233 5117 17267 5151
rect 17267 5117 17276 5151
rect 17224 5108 17276 5117
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 10232 4972 10284 5024
rect 10876 4972 10928 5024
rect 12440 4972 12492 5024
rect 13084 5015 13136 5024
rect 13084 4981 13093 5015
rect 13093 4981 13127 5015
rect 13127 4981 13136 5015
rect 13084 4972 13136 4981
rect 14004 5015 14056 5024
rect 14004 4981 14013 5015
rect 14013 4981 14047 5015
rect 14047 4981 14056 5015
rect 14004 4972 14056 4981
rect 15016 5015 15068 5024
rect 15016 4981 15025 5015
rect 15025 4981 15059 5015
rect 15059 4981 15068 5015
rect 15016 4972 15068 4981
rect 16488 5040 16540 5092
rect 19432 5176 19484 5228
rect 20628 5176 20680 5228
rect 19524 5151 19576 5160
rect 19524 5117 19533 5151
rect 19533 5117 19567 5151
rect 19567 5117 19576 5151
rect 19524 5108 19576 5117
rect 19616 5151 19668 5160
rect 19616 5117 19625 5151
rect 19625 5117 19659 5151
rect 19659 5117 19668 5151
rect 19616 5108 19668 5117
rect 19800 5108 19852 5160
rect 21272 5151 21324 5160
rect 16396 4972 16448 5024
rect 20352 5040 20404 5092
rect 21272 5117 21281 5151
rect 21281 5117 21315 5151
rect 21315 5117 21324 5151
rect 21272 5108 21324 5117
rect 23388 5176 23440 5228
rect 22468 5108 22520 5160
rect 21732 5040 21784 5092
rect 23848 5151 23900 5160
rect 23848 5117 23857 5151
rect 23857 5117 23891 5151
rect 23891 5117 23900 5151
rect 23848 5108 23900 5117
rect 24124 5040 24176 5092
rect 17500 4972 17552 5024
rect 18420 5015 18472 5024
rect 18420 4981 18429 5015
rect 18429 4981 18463 5015
rect 18463 4981 18472 5015
rect 18420 4972 18472 4981
rect 19064 5015 19116 5024
rect 19064 4981 19073 5015
rect 19073 4981 19107 5015
rect 19107 4981 19116 5015
rect 19064 4972 19116 4981
rect 21456 4972 21508 5024
rect 22284 4972 22336 5024
rect 5136 4870 5188 4922
rect 5200 4870 5252 4922
rect 5264 4870 5316 4922
rect 5328 4870 5380 4922
rect 5392 4870 5444 4922
rect 13508 4870 13560 4922
rect 13572 4870 13624 4922
rect 13636 4870 13688 4922
rect 13700 4870 13752 4922
rect 13764 4870 13816 4922
rect 21880 4870 21932 4922
rect 21944 4870 21996 4922
rect 22008 4870 22060 4922
rect 22072 4870 22124 4922
rect 22136 4870 22188 4922
rect 3700 4768 3752 4820
rect 6276 4768 6328 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 6828 4768 6880 4820
rect 7012 4768 7064 4820
rect 7196 4768 7248 4820
rect 7564 4811 7616 4820
rect 7564 4777 7573 4811
rect 7573 4777 7607 4811
rect 7607 4777 7616 4811
rect 7564 4768 7616 4777
rect 8024 4768 8076 4820
rect 10232 4811 10284 4820
rect 6368 4632 6420 4684
rect 8760 4700 8812 4752
rect 9036 4743 9088 4752
rect 9036 4709 9045 4743
rect 9045 4709 9079 4743
rect 9079 4709 9088 4743
rect 9036 4700 9088 4709
rect 10232 4777 10241 4811
rect 10241 4777 10275 4811
rect 10275 4777 10284 4811
rect 10232 4768 10284 4777
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 3884 4607 3936 4616
rect 3884 4573 3893 4607
rect 3893 4573 3927 4607
rect 3927 4573 3936 4607
rect 3884 4564 3936 4573
rect 4436 4564 4488 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6828 4564 6880 4616
rect 7012 4496 7064 4548
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7380 4607 7432 4616
rect 7196 4564 7248 4573
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 9128 4632 9180 4684
rect 11060 4700 11112 4752
rect 12348 4768 12400 4820
rect 14004 4768 14056 4820
rect 15016 4768 15068 4820
rect 15476 4768 15528 4820
rect 17500 4811 17552 4820
rect 17500 4777 17509 4811
rect 17509 4777 17543 4811
rect 17543 4777 17552 4811
rect 17500 4768 17552 4777
rect 19064 4768 19116 4820
rect 19524 4768 19576 4820
rect 21272 4811 21324 4820
rect 21272 4777 21281 4811
rect 21281 4777 21315 4811
rect 21315 4777 21324 4811
rect 21272 4768 21324 4777
rect 21732 4811 21784 4820
rect 21732 4777 21741 4811
rect 21741 4777 21775 4811
rect 21775 4777 21784 4811
rect 21732 4768 21784 4777
rect 10968 4632 11020 4684
rect 14924 4700 14976 4752
rect 16212 4743 16264 4752
rect 13084 4632 13136 4684
rect 16212 4709 16221 4743
rect 16221 4709 16255 4743
rect 16255 4709 16264 4743
rect 16212 4700 16264 4709
rect 19616 4700 19668 4752
rect 19800 4700 19852 4752
rect 7840 4564 7892 4616
rect 8208 4564 8260 4616
rect 8392 4564 8444 4616
rect 8668 4564 8720 4616
rect 10876 4564 10928 4616
rect 11336 4607 11388 4616
rect 11336 4573 11345 4607
rect 11345 4573 11388 4607
rect 11336 4564 11388 4573
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 12624 4564 12676 4616
rect 12440 4496 12492 4548
rect 16396 4675 16448 4684
rect 16396 4641 16405 4675
rect 16405 4641 16439 4675
rect 16439 4641 16448 4675
rect 16396 4632 16448 4641
rect 20628 4632 20680 4684
rect 14832 4496 14884 4548
rect 15108 4607 15160 4616
rect 15108 4573 15117 4607
rect 15117 4573 15151 4607
rect 15151 4573 15160 4607
rect 15108 4564 15160 4573
rect 15384 4607 15436 4616
rect 15384 4573 15427 4607
rect 15427 4573 15436 4607
rect 15384 4564 15436 4573
rect 16948 4564 17000 4616
rect 15292 4496 15344 4548
rect 17224 4496 17276 4548
rect 19524 4564 19576 4616
rect 20444 4564 20496 4616
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 18420 4539 18472 4548
rect 18420 4505 18429 4539
rect 18429 4505 18463 4539
rect 18463 4505 18472 4539
rect 18420 4496 18472 4505
rect 18788 4539 18840 4548
rect 18788 4505 18806 4539
rect 18806 4505 18840 4539
rect 18788 4496 18840 4505
rect 20812 4496 20864 4548
rect 21180 4564 21232 4616
rect 23020 4768 23072 4820
rect 24124 4811 24176 4820
rect 24124 4777 24133 4811
rect 24133 4777 24167 4811
rect 24167 4777 24176 4811
rect 24124 4768 24176 4777
rect 22192 4632 22244 4684
rect 22468 4675 22520 4684
rect 22468 4641 22477 4675
rect 22477 4641 22511 4675
rect 22511 4641 22520 4675
rect 22468 4632 22520 4641
rect 22744 4675 22796 4684
rect 22744 4641 22753 4675
rect 22753 4641 22787 4675
rect 22787 4641 22796 4675
rect 22744 4632 22796 4641
rect 22376 4564 22428 4616
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 21640 4496 21692 4548
rect 8300 4428 8352 4480
rect 12164 4471 12216 4480
rect 12164 4437 12173 4471
rect 12173 4437 12207 4471
rect 12207 4437 12216 4471
rect 12164 4428 12216 4437
rect 13084 4428 13136 4480
rect 14004 4428 14056 4480
rect 16580 4471 16632 4480
rect 16580 4437 16589 4471
rect 16589 4437 16623 4471
rect 16623 4437 16632 4471
rect 16580 4428 16632 4437
rect 16948 4428 17000 4480
rect 17132 4428 17184 4480
rect 18052 4471 18104 4480
rect 18052 4437 18061 4471
rect 18061 4437 18095 4471
rect 18095 4437 18104 4471
rect 18052 4428 18104 4437
rect 19616 4471 19668 4480
rect 19616 4437 19625 4471
rect 19625 4437 19659 4471
rect 19659 4437 19668 4471
rect 19616 4428 19668 4437
rect 20076 4471 20128 4480
rect 20076 4437 20085 4471
rect 20085 4437 20119 4471
rect 20119 4437 20128 4471
rect 20076 4428 20128 4437
rect 21364 4428 21416 4480
rect 22652 4428 22704 4480
rect 9322 4326 9374 4378
rect 9386 4326 9438 4378
rect 9450 4326 9502 4378
rect 9514 4326 9566 4378
rect 9578 4326 9630 4378
rect 17694 4326 17746 4378
rect 17758 4326 17810 4378
rect 17822 4326 17874 4378
rect 17886 4326 17938 4378
rect 17950 4326 18002 4378
rect 6736 4224 6788 4276
rect 6920 4224 6972 4276
rect 7380 4224 7432 4276
rect 10140 4224 10192 4276
rect 10416 4267 10468 4276
rect 10416 4233 10425 4267
rect 10425 4233 10459 4267
rect 10459 4233 10468 4267
rect 10416 4224 10468 4233
rect 3424 4156 3476 4208
rect 7932 4156 7984 4208
rect 10048 4156 10100 4208
rect 13084 4224 13136 4276
rect 14832 4224 14884 4276
rect 17132 4224 17184 4276
rect 11336 4199 11388 4208
rect 11336 4165 11345 4199
rect 11345 4165 11379 4199
rect 11379 4165 11388 4199
rect 11336 4156 11388 4165
rect 12440 4199 12492 4208
rect 12440 4165 12449 4199
rect 12449 4165 12483 4199
rect 12483 4165 12492 4199
rect 12440 4156 12492 4165
rect 15384 4156 15436 4208
rect 16488 4156 16540 4208
rect 18788 4224 18840 4276
rect 2964 4088 3016 4140
rect 4988 4088 5040 4140
rect 6644 4088 6696 4140
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 7748 4088 7800 4140
rect 8208 4088 8260 4140
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 11244 4088 11296 4140
rect 11612 4088 11664 4140
rect 13360 4088 13412 4140
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 14004 4088 14056 4140
rect 15292 4088 15344 4140
rect 18052 4156 18104 4208
rect 18420 4156 18472 4208
rect 20720 4156 20772 4208
rect 22652 4199 22704 4208
rect 22652 4165 22661 4199
rect 22661 4165 22695 4199
rect 22695 4165 22704 4199
rect 22652 4156 22704 4165
rect 6184 4063 6236 4072
rect 6184 4029 6193 4063
rect 6193 4029 6227 4063
rect 6227 4029 6236 4063
rect 6184 4020 6236 4029
rect 4528 3952 4580 4004
rect 6460 3952 6512 4004
rect 2964 3927 3016 3936
rect 2964 3893 2973 3927
rect 2973 3893 3007 3927
rect 3007 3893 3016 3927
rect 2964 3884 3016 3893
rect 5632 3884 5684 3936
rect 9220 4020 9272 4072
rect 7012 3952 7064 4004
rect 7840 3952 7892 4004
rect 8944 3884 8996 3936
rect 11060 4020 11112 4072
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 13176 4020 13228 4029
rect 13268 4063 13320 4072
rect 13268 4029 13277 4063
rect 13277 4029 13311 4063
rect 13311 4029 13320 4063
rect 13268 4020 13320 4029
rect 11888 3952 11940 4004
rect 16212 4020 16264 4072
rect 17040 4020 17092 4072
rect 20352 4088 20404 4140
rect 20444 4088 20496 4140
rect 20904 4131 20956 4140
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 23848 4156 23900 4208
rect 9864 3927 9916 3936
rect 9864 3893 9873 3927
rect 9873 3893 9907 3927
rect 9907 3893 9916 3927
rect 9864 3884 9916 3893
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 12164 3884 12216 3936
rect 12808 3927 12860 3936
rect 12808 3893 12817 3927
rect 12817 3893 12851 3927
rect 12851 3893 12860 3927
rect 12808 3884 12860 3893
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 15016 3884 15068 3936
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 16580 3884 16632 3936
rect 16672 3884 16724 3936
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 17224 3884 17276 3936
rect 21456 4020 21508 4072
rect 22192 4020 22244 4072
rect 23204 4063 23256 4072
rect 23204 4029 23213 4063
rect 23213 4029 23247 4063
rect 23247 4029 23256 4063
rect 23204 4020 23256 4029
rect 23296 4063 23348 4072
rect 23296 4029 23305 4063
rect 23305 4029 23339 4063
rect 23339 4029 23348 4063
rect 23480 4088 23532 4140
rect 23296 4020 23348 4029
rect 19800 3952 19852 4004
rect 20076 3952 20128 4004
rect 24584 3952 24636 4004
rect 19340 3884 19392 3936
rect 19616 3884 19668 3936
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 21364 3927 21416 3936
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 21548 3927 21600 3936
rect 21548 3893 21557 3927
rect 21557 3893 21591 3927
rect 21591 3893 21600 3927
rect 21548 3884 21600 3893
rect 22284 3927 22336 3936
rect 22284 3893 22293 3927
rect 22293 3893 22327 3927
rect 22327 3893 22336 3927
rect 22284 3884 22336 3893
rect 5136 3782 5188 3834
rect 5200 3782 5252 3834
rect 5264 3782 5316 3834
rect 5328 3782 5380 3834
rect 5392 3782 5444 3834
rect 13508 3782 13560 3834
rect 13572 3782 13624 3834
rect 13636 3782 13688 3834
rect 13700 3782 13752 3834
rect 13764 3782 13816 3834
rect 21880 3782 21932 3834
rect 21944 3782 21996 3834
rect 22008 3782 22060 3834
rect 22072 3782 22124 3834
rect 22136 3782 22188 3834
rect 4988 3680 5040 3732
rect 7564 3680 7616 3732
rect 8576 3680 8628 3732
rect 8760 3723 8812 3732
rect 8760 3689 8769 3723
rect 8769 3689 8803 3723
rect 8803 3689 8812 3723
rect 8760 3680 8812 3689
rect 11244 3723 11296 3732
rect 11244 3689 11253 3723
rect 11253 3689 11287 3723
rect 11287 3689 11296 3723
rect 11244 3680 11296 3689
rect 11888 3680 11940 3732
rect 14648 3680 14700 3732
rect 15384 3680 15436 3732
rect 17040 3723 17092 3732
rect 17040 3689 17049 3723
rect 17049 3689 17083 3723
rect 17083 3689 17092 3723
rect 17040 3680 17092 3689
rect 20904 3680 20956 3732
rect 13912 3612 13964 3664
rect 14096 3655 14148 3664
rect 14096 3621 14105 3655
rect 14105 3621 14139 3655
rect 14139 3621 14148 3655
rect 14096 3612 14148 3621
rect 17224 3612 17276 3664
rect 21088 3680 21140 3732
rect 21640 3680 21692 3732
rect 23296 3680 23348 3732
rect 23388 3680 23440 3732
rect 8484 3544 8536 3596
rect 9036 3544 9088 3596
rect 11336 3544 11388 3596
rect 8116 3476 8168 3528
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 8852 3476 8904 3528
rect 5816 3408 5868 3460
rect 8944 3408 8996 3460
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 11520 3519 11572 3528
rect 8668 3340 8720 3392
rect 9128 3340 9180 3392
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 10968 3408 11020 3460
rect 11612 3340 11664 3392
rect 19340 3587 19392 3596
rect 19340 3553 19349 3587
rect 19349 3553 19383 3587
rect 19383 3553 19392 3587
rect 19340 3544 19392 3553
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 14648 3519 14700 3528
rect 12440 3451 12492 3460
rect 12440 3417 12474 3451
rect 12474 3417 12492 3451
rect 12440 3408 12492 3417
rect 12992 3408 13044 3460
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 14740 3519 14792 3528
rect 14740 3485 14749 3519
rect 14749 3485 14783 3519
rect 14783 3485 14792 3519
rect 14740 3476 14792 3485
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 15660 3519 15712 3528
rect 15660 3485 15694 3519
rect 15694 3485 15712 3519
rect 15660 3476 15712 3485
rect 20168 3476 20220 3528
rect 20352 3476 20404 3528
rect 21640 3544 21692 3596
rect 14924 3408 14976 3460
rect 16856 3408 16908 3460
rect 19616 3451 19668 3460
rect 19616 3417 19650 3451
rect 19650 3417 19668 3451
rect 19616 3408 19668 3417
rect 19800 3408 19852 3460
rect 21548 3476 21600 3528
rect 22744 3476 22796 3528
rect 24124 3476 24176 3528
rect 26700 3476 26752 3528
rect 12532 3340 12584 3392
rect 13176 3340 13228 3392
rect 13268 3340 13320 3392
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 19064 3383 19116 3392
rect 19064 3349 19073 3383
rect 19073 3349 19107 3383
rect 19107 3349 19116 3383
rect 19064 3340 19116 3349
rect 20904 3340 20956 3392
rect 21088 3340 21140 3392
rect 9322 3238 9374 3290
rect 9386 3238 9438 3290
rect 9450 3238 9502 3290
rect 9514 3238 9566 3290
rect 9578 3238 9630 3290
rect 17694 3238 17746 3290
rect 17758 3238 17810 3290
rect 17822 3238 17874 3290
rect 17886 3238 17938 3290
rect 17950 3238 18002 3290
rect 7748 3179 7800 3188
rect 7748 3145 7757 3179
rect 7757 3145 7791 3179
rect 7791 3145 7800 3179
rect 7748 3136 7800 3145
rect 8760 3136 8812 3188
rect 9220 3179 9272 3188
rect 9220 3145 9229 3179
rect 9229 3145 9263 3179
rect 9263 3145 9272 3179
rect 9220 3136 9272 3145
rect 10968 3179 11020 3188
rect 10968 3145 10977 3179
rect 10977 3145 11011 3179
rect 11011 3145 11020 3179
rect 10968 3136 11020 3145
rect 12440 3179 12492 3188
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 12440 3136 12492 3145
rect 13360 3136 13412 3188
rect 6184 3068 6236 3120
rect 8576 3068 8628 3120
rect 9128 3111 9180 3120
rect 9128 3077 9137 3111
rect 9137 3077 9171 3111
rect 9171 3077 9180 3111
rect 9128 3068 9180 3077
rect 11336 3068 11388 3120
rect 11612 3068 11664 3120
rect 3884 3000 3936 3052
rect 9036 3000 9088 3052
rect 9680 3043 9732 3052
rect 9680 3009 9714 3043
rect 9714 3009 9732 3043
rect 11152 3043 11204 3052
rect 9680 3000 9732 3009
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 8852 2932 8904 2984
rect 11520 2932 11572 2984
rect 11796 3000 11848 3052
rect 12532 2932 12584 2984
rect 1952 2796 2004 2848
rect 12900 2796 12952 2848
rect 13912 3068 13964 3120
rect 13728 3000 13780 3052
rect 14648 3136 14700 3188
rect 16856 3179 16908 3188
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 19616 3136 19668 3188
rect 21272 3136 21324 3188
rect 21456 3179 21508 3188
rect 21456 3145 21465 3179
rect 21465 3145 21499 3179
rect 21499 3145 21508 3179
rect 21456 3136 21508 3145
rect 14924 3068 14976 3120
rect 19064 3068 19116 3120
rect 14740 3000 14792 3052
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 19432 3000 19484 3052
rect 19524 2932 19576 2984
rect 22100 2864 22152 2916
rect 21548 2796 21600 2848
rect 22836 2796 22888 2848
rect 5136 2694 5188 2746
rect 5200 2694 5252 2746
rect 5264 2694 5316 2746
rect 5328 2694 5380 2746
rect 5392 2694 5444 2746
rect 13508 2694 13560 2746
rect 13572 2694 13624 2746
rect 13636 2694 13688 2746
rect 13700 2694 13752 2746
rect 13764 2694 13816 2746
rect 21880 2694 21932 2746
rect 21944 2694 21996 2746
rect 22008 2694 22060 2746
rect 22072 2694 22124 2746
rect 22136 2694 22188 2746
rect 9680 2592 9732 2644
rect 13360 2592 13412 2644
rect 20444 2567 20496 2576
rect 20444 2533 20453 2567
rect 20453 2533 20487 2567
rect 20487 2533 20496 2567
rect 20444 2524 20496 2533
rect 9864 2388 9916 2440
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 13268 2388 13320 2440
rect 20168 2431 20220 2440
rect 20168 2397 20177 2431
rect 20177 2397 20211 2431
rect 20211 2397 20220 2431
rect 20168 2388 20220 2397
rect 20628 2388 20680 2440
rect 20904 2388 20956 2440
rect 9322 2150 9374 2202
rect 9386 2150 9438 2202
rect 9450 2150 9502 2202
rect 9514 2150 9566 2202
rect 9578 2150 9630 2202
rect 17694 2150 17746 2202
rect 17758 2150 17810 2202
rect 17822 2150 17874 2202
rect 17886 2150 17938 2202
rect 17950 2150 18002 2202
rect 9220 1300 9272 1352
rect 22100 1300 22152 1352
<< metal2 >>
rect 478 28739 534 29539
rect 1398 28739 1454 29539
rect 2410 28739 2466 29539
rect 3330 28739 3386 29539
rect 4342 28739 4398 29539
rect 4908 28750 5304 28778
rect 492 25906 520 28739
rect 1412 26042 1440 28739
rect 1400 26036 1452 26042
rect 1400 25978 1452 25984
rect 480 25900 532 25906
rect 480 25842 532 25848
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1596 23866 1624 25842
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1492 22024 1544 22030
rect 1492 21966 1544 21972
rect 1504 21010 1532 21966
rect 1492 21004 1544 21010
rect 1492 20946 1544 20952
rect 2424 20482 2452 28739
rect 3344 25906 3372 28739
rect 3332 25900 3384 25906
rect 3332 25842 3384 25848
rect 4252 25900 4304 25906
rect 4252 25842 4304 25848
rect 4068 24132 4120 24138
rect 4068 24074 4120 24080
rect 4080 23798 4108 24074
rect 4264 24070 4292 25842
rect 4252 24064 4304 24070
rect 4252 24006 4304 24012
rect 4264 23866 4292 24006
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 4172 23254 4200 23666
rect 4356 23474 4384 28739
rect 4436 23724 4488 23730
rect 4436 23666 4488 23672
rect 4264 23446 4384 23474
rect 4160 23248 4212 23254
rect 4160 23190 4212 23196
rect 3332 22636 3384 22642
rect 3332 22578 3384 22584
rect 3344 22030 3372 22578
rect 3976 22092 4028 22098
rect 3976 22034 4028 22040
rect 3332 22024 3384 22030
rect 3332 21966 3384 21972
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 2688 21956 2740 21962
rect 2688 21898 2740 21904
rect 2700 21690 2728 21898
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 3344 21622 3372 21830
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 2872 21548 2924 21554
rect 2872 21490 2924 21496
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 2884 21146 2912 21490
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 2504 20868 2556 20874
rect 2504 20810 2556 20816
rect 2516 20602 2544 20810
rect 2504 20596 2556 20602
rect 2504 20538 2556 20544
rect 2976 20534 3004 21490
rect 3436 21434 3464 21966
rect 3700 21956 3752 21962
rect 3700 21898 3752 21904
rect 3712 21690 3740 21898
rect 3700 21684 3752 21690
rect 3700 21626 3752 21632
rect 3344 21406 3464 21434
rect 3344 21350 3372 21406
rect 3148 21344 3200 21350
rect 3148 21286 3200 21292
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 3160 21010 3188 21286
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3056 20868 3108 20874
rect 3056 20810 3108 20816
rect 2964 20528 3016 20534
rect 2424 20454 2544 20482
rect 2964 20470 3016 20476
rect 3068 20466 3096 20810
rect 2136 19780 2188 19786
rect 2136 19722 2188 19728
rect 2148 18766 2176 19722
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 1952 18284 2004 18290
rect 2148 18272 2176 18702
rect 2516 18630 2544 20454
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 3240 19372 3292 19378
rect 3344 19360 3372 21286
rect 3424 20936 3476 20942
rect 3424 20878 3476 20884
rect 3436 19854 3464 20878
rect 3988 20466 4016 22034
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4172 21146 4200 21422
rect 4160 21140 4212 21146
rect 4160 21082 4212 21088
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3528 19990 3556 20402
rect 3608 20392 3660 20398
rect 3608 20334 3660 20340
rect 3620 20058 3648 20334
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3988 19990 4016 20402
rect 3516 19984 3568 19990
rect 3976 19984 4028 19990
rect 3516 19926 3568 19932
rect 3712 19932 3976 19938
rect 3712 19926 4028 19932
rect 3712 19910 4016 19926
rect 3712 19854 3740 19910
rect 4080 19854 4108 20470
rect 4264 20466 4292 23446
rect 4448 23186 4476 23666
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 4344 22636 4396 22642
rect 4344 22578 4396 22584
rect 4356 22234 4384 22578
rect 4724 22438 4752 23054
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4344 22228 4396 22234
rect 4344 22170 4396 22176
rect 4724 21962 4752 22374
rect 4712 21956 4764 21962
rect 4712 21898 4764 21904
rect 4436 21412 4488 21418
rect 4436 21354 4488 21360
rect 4448 21010 4476 21354
rect 4804 21140 4856 21146
rect 4804 21082 4856 21088
rect 4436 21004 4488 21010
rect 4356 20964 4436 20992
rect 4356 20602 4384 20964
rect 4436 20946 4488 20952
rect 4436 20800 4488 20806
rect 4436 20742 4488 20748
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4356 20398 4384 20538
rect 4448 20398 4476 20742
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 4436 20392 4488 20398
rect 4436 20334 4488 20340
rect 4448 19922 4476 20334
rect 4436 19916 4488 19922
rect 4436 19858 4488 19864
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3292 19332 3372 19360
rect 3240 19314 3292 19320
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2792 18358 2820 19110
rect 2976 18426 3004 19314
rect 2964 18420 3016 18426
rect 2964 18362 3016 18368
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2004 18244 2176 18272
rect 1952 18226 2004 18232
rect 2148 17218 2176 18244
rect 2976 17542 3004 18362
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 3160 17678 3188 18158
rect 3344 17746 3372 19332
rect 3424 18692 3476 18698
rect 3424 18634 3476 18640
rect 3436 18426 3464 18634
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3804 18290 3832 19654
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3988 18970 4016 19314
rect 4080 19242 4108 19790
rect 4356 19514 4384 19790
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3988 18290 4016 18906
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3792 18284 3844 18290
rect 3792 18226 3844 18232
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2884 17270 2912 17478
rect 3160 17270 3188 17614
rect 1964 17202 2176 17218
rect 2872 17264 2924 17270
rect 2872 17206 2924 17212
rect 3148 17264 3200 17270
rect 3148 17206 3200 17212
rect 1952 17196 2176 17202
rect 2004 17190 2176 17196
rect 1952 17138 2004 17144
rect 2148 16658 2176 17190
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 2148 16250 2176 16594
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2884 15706 2912 16050
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 3160 15502 3188 17206
rect 3344 15706 3372 17682
rect 3712 17338 3740 18226
rect 4448 18086 4476 19858
rect 4540 19514 4568 20538
rect 4816 20466 4844 21082
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4540 19310 4568 19450
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4066 17504 4122 17513
rect 4066 17439 4122 17448
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3528 16794 3556 17138
rect 4080 17066 4108 17439
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 4172 16998 4200 17614
rect 4356 17134 4384 17682
rect 4448 17134 4476 18022
rect 4540 17882 4568 19246
rect 4724 18766 4752 19246
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4724 18358 4752 18702
rect 4712 18352 4764 18358
rect 4712 18294 4764 18300
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 4172 16590 4200 16934
rect 4356 16726 4384 17070
rect 4344 16720 4396 16726
rect 4344 16662 4396 16668
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3436 15570 3464 16186
rect 3804 15638 3832 16390
rect 4356 16114 4384 16662
rect 4724 16658 4752 18294
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4816 16522 4844 16934
rect 4804 16516 4856 16522
rect 4804 16458 4856 16464
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 4908 15162 4936 28750
rect 5276 28642 5304 28750
rect 5354 28739 5410 29539
rect 5920 28750 6224 28778
rect 5368 28642 5396 28739
rect 5276 28614 5396 28642
rect 5136 26684 5444 26704
rect 5136 26682 5142 26684
rect 5198 26682 5222 26684
rect 5278 26682 5302 26684
rect 5358 26682 5382 26684
rect 5438 26682 5444 26684
rect 5198 26630 5200 26682
rect 5380 26630 5382 26682
rect 5136 26628 5142 26630
rect 5198 26628 5222 26630
rect 5278 26628 5302 26630
rect 5358 26628 5382 26630
rect 5438 26628 5444 26630
rect 5136 26608 5444 26628
rect 5632 25900 5684 25906
rect 5632 25842 5684 25848
rect 5136 25596 5444 25616
rect 5136 25594 5142 25596
rect 5198 25594 5222 25596
rect 5278 25594 5302 25596
rect 5358 25594 5382 25596
rect 5438 25594 5444 25596
rect 5198 25542 5200 25594
rect 5380 25542 5382 25594
rect 5136 25540 5142 25542
rect 5198 25540 5222 25542
rect 5278 25540 5302 25542
rect 5358 25540 5382 25542
rect 5438 25540 5444 25542
rect 5136 25520 5444 25540
rect 5644 25430 5672 25842
rect 5816 25832 5868 25838
rect 5816 25774 5868 25780
rect 5632 25424 5684 25430
rect 5632 25366 5684 25372
rect 5828 25362 5856 25774
rect 5816 25356 5868 25362
rect 5816 25298 5868 25304
rect 5540 25288 5592 25294
rect 5592 25248 5672 25276
rect 5540 25230 5592 25236
rect 5644 24614 5672 25248
rect 5632 24608 5684 24614
rect 5632 24550 5684 24556
rect 5136 24508 5444 24528
rect 5136 24506 5142 24508
rect 5198 24506 5222 24508
rect 5278 24506 5302 24508
rect 5358 24506 5382 24508
rect 5438 24506 5444 24508
rect 5198 24454 5200 24506
rect 5380 24454 5382 24506
rect 5136 24452 5142 24454
rect 5198 24452 5222 24454
rect 5278 24452 5302 24454
rect 5358 24452 5382 24454
rect 5438 24452 5444 24454
rect 5136 24432 5444 24452
rect 5540 24404 5592 24410
rect 5540 24346 5592 24352
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 5276 23730 5304 24006
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5136 23420 5444 23440
rect 5136 23418 5142 23420
rect 5198 23418 5222 23420
rect 5278 23418 5302 23420
rect 5358 23418 5382 23420
rect 5438 23418 5444 23420
rect 5198 23366 5200 23418
rect 5380 23366 5382 23418
rect 5136 23364 5142 23366
rect 5198 23364 5222 23366
rect 5278 23364 5302 23366
rect 5358 23364 5382 23366
rect 5438 23364 5444 23366
rect 5136 23344 5444 23364
rect 5552 23186 5580 24346
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 5644 23118 5672 24550
rect 5724 24200 5776 24206
rect 5828 24154 5856 25298
rect 5776 24148 5856 24154
rect 5724 24142 5856 24148
rect 5736 24126 5856 24142
rect 5828 23798 5856 24126
rect 5816 23792 5868 23798
rect 5816 23734 5868 23740
rect 5828 23186 5856 23734
rect 5816 23180 5868 23186
rect 5816 23122 5868 23128
rect 5632 23112 5684 23118
rect 5632 23054 5684 23060
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5136 22332 5444 22352
rect 5136 22330 5142 22332
rect 5198 22330 5222 22332
rect 5278 22330 5302 22332
rect 5358 22330 5382 22332
rect 5438 22330 5444 22332
rect 5198 22278 5200 22330
rect 5380 22278 5382 22330
rect 5136 22276 5142 22278
rect 5198 22276 5222 22278
rect 5278 22276 5302 22278
rect 5358 22276 5382 22278
rect 5438 22276 5444 22278
rect 5136 22256 5444 22276
rect 5136 21244 5444 21264
rect 5136 21242 5142 21244
rect 5198 21242 5222 21244
rect 5278 21242 5302 21244
rect 5358 21242 5382 21244
rect 5438 21242 5444 21244
rect 5198 21190 5200 21242
rect 5380 21190 5382 21242
rect 5136 21188 5142 21190
rect 5198 21188 5222 21190
rect 5278 21188 5302 21190
rect 5358 21188 5382 21190
rect 5438 21188 5444 21190
rect 5136 21168 5444 21188
rect 5552 20942 5580 22714
rect 5644 22438 5672 23054
rect 5828 22778 5856 23122
rect 5816 22772 5868 22778
rect 5816 22714 5868 22720
rect 5632 22432 5684 22438
rect 5632 22374 5684 22380
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5448 20460 5500 20466
rect 5632 20460 5684 20466
rect 5500 20420 5580 20448
rect 5448 20402 5500 20408
rect 5276 20369 5304 20402
rect 5262 20360 5318 20369
rect 5262 20295 5318 20304
rect 5552 20262 5580 20420
rect 5920 20448 5948 28750
rect 6196 28642 6224 28750
rect 6274 28739 6330 29539
rect 7286 28739 7342 29539
rect 8298 28739 8354 29539
rect 9218 28739 9274 29539
rect 10230 28739 10286 29539
rect 11242 28739 11298 29539
rect 11624 28750 12112 28778
rect 6288 28642 6316 28739
rect 6196 28614 6316 28642
rect 7012 26512 7064 26518
rect 7012 26454 7064 26460
rect 7024 25226 7052 26454
rect 7104 26376 7156 26382
rect 7104 26318 7156 26324
rect 7288 26376 7340 26382
rect 7288 26318 7340 26324
rect 7116 26042 7144 26318
rect 7196 26240 7248 26246
rect 7196 26182 7248 26188
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 7208 25362 7236 26182
rect 7300 25498 7328 26318
rect 7840 26036 7892 26042
rect 7840 25978 7892 25984
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 7196 25356 7248 25362
rect 7196 25298 7248 25304
rect 6460 25220 6512 25226
rect 6460 25162 6512 25168
rect 7012 25220 7064 25226
rect 7012 25162 7064 25168
rect 6472 24954 6500 25162
rect 6460 24948 6512 24954
rect 6460 24890 6512 24896
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6000 24200 6052 24206
rect 6000 24142 6052 24148
rect 6932 24154 6960 24754
rect 7024 24750 7052 25162
rect 7208 24886 7236 25298
rect 7196 24880 7248 24886
rect 7196 24822 7248 24828
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 7024 24342 7052 24686
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7012 24336 7064 24342
rect 7012 24278 7064 24284
rect 7116 24274 7144 24550
rect 7104 24268 7156 24274
rect 7104 24210 7156 24216
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 7208 24154 7236 24210
rect 7300 24206 7328 25434
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 7760 24750 7788 25230
rect 7852 24818 7880 25978
rect 8024 25900 8076 25906
rect 8024 25842 8076 25848
rect 8036 25498 8064 25842
rect 8024 25492 8076 25498
rect 8024 25434 8076 25440
rect 7932 25288 7984 25294
rect 7932 25230 7984 25236
rect 8116 25288 8168 25294
rect 8116 25230 8168 25236
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 7748 24744 7800 24750
rect 7748 24686 7800 24692
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 6012 23866 6040 24142
rect 6932 24126 7236 24154
rect 7288 24200 7340 24206
rect 7288 24142 7340 24148
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 6828 23724 6880 23730
rect 6828 23666 6880 23672
rect 6840 23610 6868 23666
rect 6840 23582 7052 23610
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6092 22432 6144 22438
rect 6092 22374 6144 22380
rect 6104 22166 6132 22374
rect 6092 22160 6144 22166
rect 6092 22102 6144 22108
rect 6748 21978 6776 23462
rect 7024 23254 7052 23582
rect 7116 23322 7144 24006
rect 7300 23798 7328 24142
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7208 23322 7236 23666
rect 7392 23662 7420 24142
rect 7380 23656 7432 23662
rect 7380 23598 7432 23604
rect 7484 23526 7512 24346
rect 7564 24200 7616 24206
rect 7564 24142 7616 24148
rect 7472 23520 7524 23526
rect 7472 23462 7524 23468
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7012 23248 7064 23254
rect 7012 23190 7064 23196
rect 6920 23044 6972 23050
rect 6920 22986 6972 22992
rect 6932 22710 6960 22986
rect 6920 22704 6972 22710
rect 6920 22646 6972 22652
rect 6932 22098 6960 22646
rect 7024 22438 7052 23190
rect 7116 22642 7144 23258
rect 7208 22710 7236 23258
rect 7196 22704 7248 22710
rect 7196 22646 7248 22652
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 7116 22234 7144 22578
rect 7576 22506 7604 24142
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7668 22794 7696 24074
rect 7760 23526 7788 24686
rect 7852 24410 7880 24754
rect 7944 24614 7972 25230
rect 8128 24954 8156 25230
rect 8116 24948 8168 24954
rect 8116 24890 8168 24896
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 8024 24608 8076 24614
rect 8024 24550 8076 24556
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 8036 24274 8064 24550
rect 8024 24268 8076 24274
rect 8024 24210 8076 24216
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 7668 22766 7788 22794
rect 7852 22778 7880 23054
rect 7656 22704 7708 22710
rect 7656 22646 7708 22652
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 7668 22386 7696 22646
rect 7484 22358 7696 22386
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 6920 22092 6972 22098
rect 6920 22034 6972 22040
rect 6748 21950 6960 21978
rect 6932 20942 6960 21950
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 6000 20868 6052 20874
rect 6000 20810 6052 20816
rect 6092 20868 6144 20874
rect 6092 20810 6144 20816
rect 6276 20868 6328 20874
rect 6276 20810 6328 20816
rect 6012 20466 6040 20810
rect 6104 20602 6132 20810
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 6288 20534 6316 20810
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 6276 20528 6328 20534
rect 6276 20470 6328 20476
rect 5684 20420 5948 20448
rect 5632 20402 5684 20408
rect 5920 20346 5948 20420
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6380 20346 6408 20538
rect 6644 20528 6696 20534
rect 6644 20470 6696 20476
rect 6552 20460 6604 20466
rect 5920 20318 6408 20346
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5136 20156 5444 20176
rect 5136 20154 5142 20156
rect 5198 20154 5222 20156
rect 5278 20154 5302 20156
rect 5358 20154 5382 20156
rect 5438 20154 5444 20156
rect 5198 20102 5200 20154
rect 5380 20102 5382 20154
rect 5136 20100 5142 20102
rect 5198 20100 5222 20102
rect 5278 20100 5302 20102
rect 5358 20100 5382 20102
rect 5438 20100 5444 20102
rect 5136 20080 5444 20100
rect 5136 19068 5444 19088
rect 5136 19066 5142 19068
rect 5198 19066 5222 19068
rect 5278 19066 5302 19068
rect 5358 19066 5382 19068
rect 5438 19066 5444 19068
rect 5198 19014 5200 19066
rect 5380 19014 5382 19066
rect 5136 19012 5142 19014
rect 5198 19012 5222 19014
rect 5278 19012 5302 19014
rect 5358 19012 5382 19014
rect 5438 19012 5444 19014
rect 5136 18992 5444 19012
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5136 17980 5444 18000
rect 5136 17978 5142 17980
rect 5198 17978 5222 17980
rect 5278 17978 5302 17980
rect 5358 17978 5382 17980
rect 5438 17978 5444 17980
rect 5198 17926 5200 17978
rect 5380 17926 5382 17978
rect 5136 17924 5142 17926
rect 5198 17924 5222 17926
rect 5278 17924 5302 17926
rect 5358 17924 5382 17926
rect 5438 17924 5444 17926
rect 5136 17904 5444 17924
rect 5828 17202 5856 18022
rect 6380 17678 6408 20318
rect 6472 20420 6552 20448
rect 6472 20058 6500 20420
rect 6552 20402 6604 20408
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 6564 19854 6592 20198
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6656 19310 6684 20470
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6748 19378 6776 20334
rect 6840 19922 6868 20878
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7116 20330 7144 20402
rect 7104 20324 7156 20330
rect 7104 20266 7156 20272
rect 7288 20324 7340 20330
rect 7288 20266 7340 20272
rect 7116 20058 7144 20266
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 7300 19786 7328 20266
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7484 19718 7512 22358
rect 7760 22250 7788 22766
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 7576 22222 7788 22250
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6748 18970 6776 19314
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6932 18834 6960 19314
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 6564 18290 6592 18702
rect 7024 18290 7052 18702
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6104 17202 6132 17478
rect 6184 17332 6236 17338
rect 6236 17292 6408 17320
rect 6184 17274 6236 17280
rect 6182 17232 6238 17241
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 6092 17196 6144 17202
rect 6380 17202 6408 17292
rect 6748 17202 6776 18022
rect 6182 17167 6184 17176
rect 6092 17138 6144 17144
rect 6236 17167 6238 17176
rect 6368 17196 6420 17202
rect 6184 17138 6236 17144
rect 6368 17138 6420 17144
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 5000 16250 5028 17138
rect 5136 16892 5444 16912
rect 5136 16890 5142 16892
rect 5198 16890 5222 16892
rect 5278 16890 5302 16892
rect 5358 16890 5382 16892
rect 5438 16890 5444 16892
rect 5198 16838 5200 16890
rect 5380 16838 5382 16890
rect 5136 16836 5142 16838
rect 5198 16836 5222 16838
rect 5278 16836 5302 16838
rect 5358 16836 5382 16838
rect 5438 16836 5444 16838
rect 5136 16816 5444 16836
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5828 16046 5856 17138
rect 6840 17134 6868 18022
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6840 16794 6868 17070
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 6288 16250 6316 16458
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6380 16182 6408 16390
rect 6368 16176 6420 16182
rect 6368 16118 6420 16124
rect 6564 16114 6592 16730
rect 6840 16114 6868 16730
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 6932 15910 6960 16050
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 5136 15804 5444 15824
rect 5136 15802 5142 15804
rect 5198 15802 5222 15804
rect 5278 15802 5302 15804
rect 5358 15802 5382 15804
rect 5438 15802 5444 15804
rect 5198 15750 5200 15802
rect 5380 15750 5382 15802
rect 5136 15748 5142 15750
rect 5198 15748 5222 15750
rect 5278 15748 5302 15750
rect 5358 15748 5382 15750
rect 5438 15748 5444 15750
rect 5136 15728 5444 15748
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2884 14074 2912 14894
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4080 14414 4108 14758
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1504 13326 1532 13806
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1504 11830 1532 13262
rect 2136 13252 2188 13258
rect 2136 13194 2188 13200
rect 2148 12986 2176 13194
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2332 12442 2360 13874
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2516 12918 2544 13398
rect 2504 12912 2556 12918
rect 2884 12866 2912 14010
rect 3436 13938 3464 14350
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2976 12889 3004 12922
rect 2504 12854 2556 12860
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2700 12838 2912 12866
rect 2962 12880 3018 12889
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2608 12186 2636 12786
rect 2700 12306 2728 12838
rect 2962 12815 3018 12824
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12374 2912 12718
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2608 12170 2728 12186
rect 2608 12164 2740 12170
rect 2608 12158 2688 12164
rect 2688 12106 2740 12112
rect 1492 11824 1544 11830
rect 1492 11766 1544 11772
rect 1504 11694 1532 11766
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1504 10130 1532 11630
rect 2332 11354 2360 11698
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2700 11098 2728 12106
rect 2884 11898 2912 12310
rect 2976 12220 3004 12650
rect 3160 12442 3188 13126
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3252 12238 3280 13262
rect 3344 12850 3372 13466
rect 3436 13394 3464 13874
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 3436 12986 3464 13194
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3514 12880 3570 12889
rect 3332 12844 3384 12850
rect 3514 12815 3516 12824
rect 3332 12786 3384 12792
rect 3568 12815 3570 12824
rect 3792 12844 3844 12850
rect 3516 12786 3568 12792
rect 3792 12786 3844 12792
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3344 12442 3372 12582
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3056 12232 3108 12238
rect 2976 12192 3056 12220
rect 3056 12174 3108 12180
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2884 11354 2912 11834
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 3068 11218 3096 12174
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2780 11144 2832 11150
rect 2700 11092 2780 11098
rect 2700 11086 2832 11092
rect 2700 11070 2820 11086
rect 2884 10810 2912 11154
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2884 10266 2912 10542
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2516 9722 2544 9930
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2884 9654 2912 10202
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2792 9042 2820 9522
rect 2976 9518 3004 9862
rect 3068 9586 3096 11154
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3344 10198 3372 10610
rect 3332 10192 3384 10198
rect 3332 10134 3384 10140
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 3068 9178 3096 9522
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3160 9058 3188 10066
rect 3344 10062 3372 10134
rect 3436 10062 3464 12174
rect 3528 11218 3556 12786
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3252 9178 3280 9386
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2976 9030 3188 9058
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 8498 2728 8774
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2792 7818 2820 8978
rect 2976 8974 3004 9030
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 7886 2912 8774
rect 2976 8634 3004 8910
rect 3344 8838 3372 9522
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7410 3280 7686
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3436 7290 3464 9590
rect 3620 9586 3648 10134
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3712 9382 3740 11086
rect 3804 10606 3832 12786
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11830 3924 12174
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 3988 11218 4016 12922
rect 4356 12782 4384 14826
rect 4724 14822 4752 14962
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4816 14074 4844 14826
rect 4908 14550 4936 15098
rect 5552 15094 5580 15302
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5136 14716 5444 14736
rect 5136 14714 5142 14716
rect 5198 14714 5222 14716
rect 5278 14714 5302 14716
rect 5358 14714 5382 14716
rect 5438 14714 5444 14716
rect 5198 14662 5200 14714
rect 5380 14662 5382 14714
rect 5136 14660 5142 14662
rect 5198 14660 5222 14662
rect 5278 14660 5302 14662
rect 5358 14660 5382 14662
rect 5438 14660 5444 14662
rect 5136 14640 5444 14660
rect 5552 14618 5580 15030
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 4896 14544 4948 14550
rect 4896 14486 4948 14492
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4448 12918 4476 13874
rect 4816 12918 4844 14010
rect 5136 13628 5444 13648
rect 5136 13626 5142 13628
rect 5198 13626 5222 13628
rect 5278 13626 5302 13628
rect 5358 13626 5382 13628
rect 5438 13626 5444 13628
rect 5198 13574 5200 13626
rect 5380 13574 5382 13626
rect 5136 13572 5142 13574
rect 5198 13572 5222 13574
rect 5278 13572 5302 13574
rect 5358 13572 5382 13574
rect 5438 13572 5444 13574
rect 5136 13552 5444 13572
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4540 12646 4568 12786
rect 4908 12782 4936 12922
rect 5000 12850 5028 13262
rect 5170 12880 5226 12889
rect 4988 12844 5040 12850
rect 5170 12815 5172 12824
rect 4988 12786 5040 12792
rect 5224 12815 5226 12824
rect 5538 12880 5594 12889
rect 5538 12815 5594 12824
rect 5172 12786 5224 12792
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4172 12238 4200 12582
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4724 12170 4752 12650
rect 4816 12442 4844 12718
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 5000 12442 5028 12582
rect 5136 12540 5444 12560
rect 5136 12538 5142 12540
rect 5198 12538 5222 12540
rect 5278 12538 5302 12540
rect 5358 12538 5382 12540
rect 5438 12538 5444 12540
rect 5198 12486 5200 12538
rect 5380 12486 5382 12538
rect 5136 12484 5142 12486
rect 5198 12484 5222 12486
rect 5278 12484 5302 12486
rect 5358 12484 5382 12486
rect 5438 12484 5444 12486
rect 5136 12464 5444 12484
rect 5552 12442 5580 12815
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 4448 11150 4476 11834
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4540 11354 4568 11698
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 4080 10130 4108 11086
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4632 9586 4660 11154
rect 4816 10962 4844 11630
rect 4908 11150 4936 12242
rect 5644 12238 5672 14962
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 5828 12850 5856 14894
rect 6564 14414 6592 14894
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6840 14113 6868 14894
rect 6826 14104 6882 14113
rect 6826 14039 6882 14048
rect 6840 14006 6868 14039
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6472 12986 6500 13262
rect 6932 13190 6960 13874
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7024 13258 7052 13806
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5736 12238 5764 12786
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 4986 11928 5042 11937
rect 4986 11863 5042 11872
rect 5172 11892 5224 11898
rect 5000 11626 5028 11863
rect 5172 11834 5224 11840
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5184 11801 5212 11834
rect 5170 11792 5226 11801
rect 5170 11727 5226 11736
rect 5276 11694 5304 11834
rect 5828 11778 5856 12786
rect 5908 12436 5960 12442
rect 6472 12434 6500 12922
rect 5908 12378 5960 12384
rect 6380 12406 6500 12434
rect 5920 12170 5948 12378
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 5368 11762 5856 11778
rect 5356 11756 5856 11762
rect 5408 11750 5856 11756
rect 5356 11698 5408 11704
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 5136 11452 5444 11472
rect 5136 11450 5142 11452
rect 5198 11450 5222 11452
rect 5278 11450 5302 11452
rect 5358 11450 5382 11452
rect 5438 11450 5444 11452
rect 5198 11398 5200 11450
rect 5380 11398 5382 11450
rect 5136 11396 5142 11398
rect 5198 11396 5222 11398
rect 5278 11396 5302 11398
rect 5358 11396 5382 11398
rect 5438 11396 5444 11398
rect 5136 11376 5444 11396
rect 5552 11150 5580 11630
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 11218 5672 11494
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 4724 10934 4844 10962
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3620 8498 3648 8774
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3712 7886 3740 9318
rect 3896 9178 3924 9318
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3896 7410 3924 8434
rect 3988 8265 4016 9318
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 4080 8974 4108 9046
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3974 8256 4030 8265
rect 3974 8191 4030 8200
rect 4172 8022 4200 9454
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4172 7546 4200 7958
rect 4356 7886 4384 8978
rect 4632 8974 4660 9522
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4632 8634 4660 8910
rect 4620 8628 4672 8634
rect 4724 8616 4752 10934
rect 4908 10826 4936 11086
rect 4816 10810 4936 10826
rect 4804 10804 4936 10810
rect 4856 10798 4936 10804
rect 4804 10746 4856 10752
rect 5276 10674 5304 11086
rect 5552 10810 5580 11086
rect 5644 11082 5672 11154
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5644 10810 5672 11018
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5552 10690 5580 10746
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 5264 10668 5316 10674
rect 5552 10662 5764 10690
rect 5264 10610 5316 10616
rect 4816 9518 4844 10610
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5136 10364 5444 10384
rect 5136 10362 5142 10364
rect 5198 10362 5222 10364
rect 5278 10362 5302 10364
rect 5358 10362 5382 10364
rect 5438 10362 5444 10364
rect 5198 10310 5200 10362
rect 5380 10310 5382 10362
rect 5136 10308 5142 10310
rect 5198 10308 5222 10310
rect 5278 10308 5302 10310
rect 5358 10308 5382 10310
rect 5438 10308 5444 10310
rect 5136 10288 5444 10308
rect 5552 10266 5580 10474
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 5000 8974 5028 9998
rect 5644 9926 5672 10662
rect 5736 10606 5764 10662
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5724 10056 5776 10062
rect 5828 10044 5856 11750
rect 5776 10016 5856 10044
rect 5724 9998 5776 10004
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5136 9276 5444 9296
rect 5136 9274 5142 9276
rect 5198 9274 5222 9276
rect 5278 9274 5302 9276
rect 5358 9274 5382 9276
rect 5438 9274 5444 9276
rect 5198 9222 5200 9274
rect 5380 9222 5382 9274
rect 5136 9220 5142 9222
rect 5198 9220 5222 9222
rect 5278 9220 5302 9222
rect 5358 9220 5382 9222
rect 5438 9220 5444 9222
rect 5136 9200 5444 9220
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4724 8588 4844 8616
rect 4620 8570 4672 8576
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4724 8090 4752 8434
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3252 7262 3464 7290
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2976 3942 3004 4082
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 662 3496 718 3505
rect 662 3431 718 3440
rect 676 800 704 3431
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1964 800 1992 2790
rect 2976 921 3004 3878
rect 2962 912 3018 921
rect 2962 847 3018 856
rect 3252 800 3280 7262
rect 3896 5302 3924 7346
rect 4816 5914 4844 8588
rect 4908 7868 4936 8774
rect 5000 8090 5028 8910
rect 5136 8188 5444 8208
rect 5136 8186 5142 8188
rect 5198 8186 5222 8188
rect 5278 8186 5302 8188
rect 5358 8186 5382 8188
rect 5438 8186 5444 8188
rect 5198 8134 5200 8186
rect 5380 8134 5382 8186
rect 5136 8132 5142 8134
rect 5198 8132 5222 8134
rect 5278 8132 5302 8134
rect 5358 8132 5382 8134
rect 5438 8132 5444 8134
rect 5136 8112 5444 8132
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4988 7880 5040 7886
rect 4908 7840 4988 7868
rect 4988 7822 5040 7828
rect 5000 6361 5028 7822
rect 5552 7750 5580 9114
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5644 8362 5672 8842
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5736 7886 5764 8434
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5828 7750 5856 10016
rect 5920 7886 5948 12106
rect 6196 11762 6224 12174
rect 6288 12102 6316 12310
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6196 10742 6224 11018
rect 6184 10736 6236 10742
rect 6184 10678 6236 10684
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 6012 8634 6040 10474
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6104 9994 6132 10406
rect 6092 9988 6144 9994
rect 6092 9930 6144 9936
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 6104 9178 6132 9386
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6012 7954 6040 8570
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6196 7886 6224 8910
rect 6380 7970 6408 12406
rect 7116 11898 7144 19450
rect 7286 19408 7342 19417
rect 7286 19343 7288 19352
rect 7340 19343 7342 19352
rect 7288 19314 7340 19320
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7196 18896 7248 18902
rect 7196 18838 7248 18844
rect 7208 15706 7236 18838
rect 7392 18766 7420 19246
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 18358 7420 18566
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 7288 16516 7340 16522
rect 7288 16458 7340 16464
rect 7300 16250 7328 16458
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7288 16108 7340 16114
rect 7392 16096 7420 16186
rect 7340 16068 7420 16096
rect 7288 16050 7340 16056
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7300 14346 7328 14894
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7196 13932 7248 13938
rect 7300 13920 7328 14282
rect 7392 13977 7420 14962
rect 7248 13892 7328 13920
rect 7378 13968 7434 13977
rect 7378 13903 7434 13912
rect 7196 13874 7248 13880
rect 7392 13734 7420 13903
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 6828 11756 6880 11762
rect 7116 11744 7144 11834
rect 6880 11716 7144 11744
rect 6828 11698 6880 11704
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10674 6500 10950
rect 6932 10742 6960 11086
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6932 10062 6960 10678
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6564 8090 6592 8366
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6748 8022 6776 8434
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 8090 6960 8230
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6736 8016 6788 8022
rect 6380 7942 6500 7970
rect 6736 7958 6788 7964
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5736 7546 5764 7686
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5920 7478 5948 7822
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 5136 7100 5444 7120
rect 5136 7098 5142 7100
rect 5198 7098 5222 7100
rect 5278 7098 5302 7100
rect 5358 7098 5382 7100
rect 5438 7098 5444 7100
rect 5198 7046 5200 7098
rect 5380 7046 5382 7098
rect 5136 7044 5142 7046
rect 5198 7044 5222 7046
rect 5278 7044 5302 7046
rect 5358 7044 5382 7046
rect 5438 7044 5444 7046
rect 5136 7024 5444 7044
rect 6012 6798 6040 7754
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 4986 6352 5042 6361
rect 4986 6287 5042 6296
rect 5136 6012 5444 6032
rect 5136 6010 5142 6012
rect 5198 6010 5222 6012
rect 5278 6010 5302 6012
rect 5358 6010 5382 6012
rect 5438 6010 5444 6012
rect 5198 5958 5200 6010
rect 5380 5958 5382 6010
rect 5136 5956 5142 5958
rect 5198 5956 5222 5958
rect 5278 5956 5302 5958
rect 5358 5956 5382 5958
rect 5438 5956 5444 5958
rect 5136 5936 5444 5956
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3712 4826 3740 5170
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3896 4622 3924 5238
rect 5276 5234 5304 5782
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5368 5370 5396 5646
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5644 5166 5672 6394
rect 6196 6390 6224 7822
rect 6380 7478 6408 7822
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 6184 6384 6236 6390
rect 6090 6352 6146 6361
rect 6184 6326 6236 6332
rect 6090 6287 6146 6296
rect 5816 6180 5868 6186
rect 5816 6122 5868 6128
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4448 4622 4476 5034
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 3436 4214 3464 4558
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3896 3058 3924 4558
rect 5000 4146 5028 5102
rect 5136 4924 5444 4944
rect 5136 4922 5142 4924
rect 5198 4922 5222 4924
rect 5278 4922 5302 4924
rect 5358 4922 5382 4924
rect 5438 4922 5444 4924
rect 5198 4870 5200 4922
rect 5380 4870 5382 4922
rect 5136 4868 5142 4870
rect 5198 4868 5222 4870
rect 5278 4868 5302 4870
rect 5358 4868 5382 4870
rect 5438 4868 5444 4870
rect 5136 4848 5444 4868
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 4540 800 4568 3946
rect 5000 3738 5028 4082
rect 5644 3942 5672 5102
rect 5736 4622 5764 5850
rect 5828 5710 5856 6122
rect 6104 5710 6132 6287
rect 6196 5914 6224 6326
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6288 5370 6316 5646
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6380 5370 6408 5578
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 5920 4622 5948 5170
rect 6288 4826 6316 5170
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6380 4690 6408 5306
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5136 3836 5444 3856
rect 5136 3834 5142 3836
rect 5198 3834 5222 3836
rect 5278 3834 5302 3836
rect 5358 3834 5382 3836
rect 5438 3834 5444 3836
rect 5198 3782 5200 3834
rect 5380 3782 5382 3834
rect 5136 3780 5142 3782
rect 5198 3780 5222 3782
rect 5278 3780 5302 3782
rect 5358 3780 5382 3782
rect 5438 3780 5444 3782
rect 5136 3760 5444 3780
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5136 2748 5444 2768
rect 5136 2746 5142 2748
rect 5198 2746 5222 2748
rect 5278 2746 5302 2748
rect 5358 2746 5382 2748
rect 5438 2746 5444 2748
rect 5198 2694 5200 2746
rect 5380 2694 5382 2746
rect 5136 2692 5142 2694
rect 5198 2692 5222 2694
rect 5278 2692 5302 2694
rect 5358 2692 5382 2694
rect 5438 2692 5444 2694
rect 5136 2672 5444 2692
rect 5828 800 5856 3402
rect 6196 3126 6224 4014
rect 6472 4010 6500 7942
rect 6840 7954 7052 7970
rect 6840 7948 7064 7954
rect 6840 7942 7012 7948
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6748 7002 6776 7754
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 6840 6866 6868 7942
rect 7012 7890 7064 7896
rect 7208 7562 7236 13126
rect 7484 12434 7512 19654
rect 7392 12406 7512 12434
rect 7392 9654 7420 12406
rect 7576 12306 7604 22222
rect 7748 22160 7800 22166
rect 7748 22102 7800 22108
rect 7656 21956 7708 21962
rect 7656 21898 7708 21904
rect 7668 21350 7696 21898
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7668 18766 7696 21286
rect 7760 19666 7788 22102
rect 7944 21690 7972 23054
rect 8036 22094 8064 24210
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8128 23526 8156 23802
rect 8208 23588 8260 23594
rect 8208 23530 8260 23536
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 8128 23202 8156 23462
rect 8220 23338 8248 23530
rect 8312 23474 8340 28739
rect 9322 27228 9630 27248
rect 9322 27226 9328 27228
rect 9384 27226 9408 27228
rect 9464 27226 9488 27228
rect 9544 27226 9568 27228
rect 9624 27226 9630 27228
rect 9384 27174 9386 27226
rect 9566 27174 9568 27226
rect 9322 27172 9328 27174
rect 9384 27172 9408 27174
rect 9464 27172 9488 27174
rect 9544 27172 9568 27174
rect 9624 27172 9630 27174
rect 9322 27152 9630 27172
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9220 26512 9272 26518
rect 9220 26454 9272 26460
rect 9128 26308 9180 26314
rect 9128 26250 9180 26256
rect 8484 25424 8536 25430
rect 8484 25366 8536 25372
rect 8496 24954 8524 25366
rect 8484 24948 8536 24954
rect 8484 24890 8536 24896
rect 9140 24750 9168 26250
rect 9232 25430 9260 26454
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 9322 26140 9630 26160
rect 9322 26138 9328 26140
rect 9384 26138 9408 26140
rect 9464 26138 9488 26140
rect 9544 26138 9568 26140
rect 9624 26138 9630 26140
rect 9384 26086 9386 26138
rect 9566 26086 9568 26138
rect 9322 26084 9328 26086
rect 9384 26084 9408 26086
rect 9464 26084 9488 26086
rect 9544 26084 9568 26086
rect 9624 26084 9630 26086
rect 9322 26064 9630 26084
rect 9692 26042 9720 26318
rect 9680 26036 9732 26042
rect 9680 25978 9732 25984
rect 9588 25832 9640 25838
rect 9588 25774 9640 25780
rect 9220 25424 9272 25430
rect 9220 25366 9272 25372
rect 9600 25242 9628 25774
rect 9784 25498 9812 26930
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9876 25786 9904 26182
rect 9968 25974 9996 26726
rect 9956 25968 10008 25974
rect 9956 25910 10008 25916
rect 9876 25758 9996 25786
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 9772 25288 9824 25294
rect 9220 25220 9272 25226
rect 9600 25214 9720 25242
rect 9772 25230 9824 25236
rect 9220 25162 9272 25168
rect 9128 24744 9180 24750
rect 9128 24686 9180 24692
rect 9232 24410 9260 25162
rect 9322 25052 9630 25072
rect 9322 25050 9328 25052
rect 9384 25050 9408 25052
rect 9464 25050 9488 25052
rect 9544 25050 9568 25052
rect 9624 25050 9630 25052
rect 9384 24998 9386 25050
rect 9566 24998 9568 25050
rect 9322 24996 9328 24998
rect 9384 24996 9408 24998
rect 9464 24996 9488 24998
rect 9544 24996 9568 24998
rect 9624 24996 9630 24998
rect 9322 24976 9630 24996
rect 9312 24880 9364 24886
rect 9692 24834 9720 25214
rect 9312 24822 9364 24828
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9324 24342 9352 24822
rect 9600 24806 9720 24834
rect 9600 24750 9628 24806
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 9312 24336 9364 24342
rect 9312 24278 9364 24284
rect 9600 24274 9628 24686
rect 9784 24410 9812 25230
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9876 24290 9904 25298
rect 9968 25158 9996 25758
rect 9956 25152 10008 25158
rect 9956 25094 10008 25100
rect 9968 24886 9996 25094
rect 9956 24880 10008 24886
rect 9956 24822 10008 24828
rect 9220 24268 9272 24274
rect 9220 24210 9272 24216
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9692 24262 9904 24290
rect 8576 23724 8628 23730
rect 8576 23666 8628 23672
rect 8312 23446 8524 23474
rect 8220 23310 8340 23338
rect 8128 23186 8248 23202
rect 8128 23180 8260 23186
rect 8128 23174 8208 23180
rect 8128 22438 8156 23174
rect 8208 23122 8260 23128
rect 8312 22778 8340 23310
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8312 22642 8340 22714
rect 8300 22636 8352 22642
rect 8300 22578 8352 22584
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 8036 22066 8248 22094
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7852 19922 7880 20878
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7760 19638 7880 19666
rect 7746 19408 7802 19417
rect 7746 19343 7802 19352
rect 7760 18970 7788 19343
rect 7852 19174 7880 19638
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7656 18760 7708 18766
rect 7656 18702 7708 18708
rect 7668 18222 7696 18702
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7668 18086 7696 18158
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7668 12442 7696 18022
rect 7760 17241 7788 18906
rect 7746 17232 7802 17241
rect 7746 17167 7802 17176
rect 7760 16250 7788 17167
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7760 15094 7788 15642
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7760 12986 7788 13874
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7484 10810 7512 11290
rect 7576 11082 7604 12242
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7760 11082 7788 11222
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7760 10810 7788 11018
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7380 9648 7432 9654
rect 7432 9608 7604 9636
rect 7380 9590 7432 9596
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8498 7420 8774
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7484 8022 7512 8910
rect 7576 8634 7604 9608
rect 7852 9178 7880 19110
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 7944 17270 7972 17546
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7944 16794 7972 17002
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 8036 16590 8064 18702
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8128 17202 8156 17478
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 8220 16674 8248 22066
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 8312 21010 8340 21898
rect 8404 21894 8432 22510
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8404 19854 8432 20334
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8404 19446 8432 19790
rect 8392 19440 8444 19446
rect 8392 19382 8444 19388
rect 8392 18896 8444 18902
rect 8392 18838 8444 18844
rect 8404 18766 8432 18838
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8312 17338 8340 17682
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8128 16646 8248 16674
rect 8312 16658 8340 17274
rect 8300 16652 8352 16658
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 8036 15570 8064 15846
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7944 13394 7972 14350
rect 8022 14104 8078 14113
rect 8022 14039 8078 14048
rect 8036 13938 8064 14039
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7944 12850 7972 13330
rect 8036 13258 8064 13874
rect 8128 13462 8156 16646
rect 8300 16594 8352 16600
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8220 15910 8248 16526
rect 8298 16144 8354 16153
rect 8298 16079 8300 16088
rect 8352 16079 8354 16088
rect 8300 16050 8352 16056
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8220 13870 8248 14282
rect 8312 14006 8340 14282
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8298 13832 8354 13841
rect 8220 13734 8248 13806
rect 8298 13767 8300 13776
rect 8352 13767 8354 13776
rect 8300 13738 8352 13744
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 8220 13376 8248 13670
rect 8300 13388 8352 13394
rect 8220 13348 8300 13376
rect 8300 13330 8352 13336
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7944 12442 7972 12786
rect 8036 12442 8064 13194
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12918 8156 13126
rect 8404 12986 8432 17818
rect 8496 14618 8524 23446
rect 8588 22506 8616 23666
rect 9232 23050 9260 24210
rect 9692 24138 9720 24262
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9680 24132 9732 24138
rect 9680 24074 9732 24080
rect 9322 23964 9630 23984
rect 9322 23962 9328 23964
rect 9384 23962 9408 23964
rect 9464 23962 9488 23964
rect 9544 23962 9568 23964
rect 9624 23962 9630 23964
rect 9384 23910 9386 23962
rect 9566 23910 9568 23962
rect 9322 23908 9328 23910
rect 9384 23908 9408 23910
rect 9464 23908 9488 23910
rect 9544 23908 9568 23910
rect 9624 23908 9630 23910
rect 9322 23888 9630 23908
rect 9692 23746 9720 24074
rect 9784 23866 9812 24142
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9692 23718 9812 23746
rect 9784 23662 9812 23718
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9784 23322 9812 23598
rect 9772 23316 9824 23322
rect 9772 23258 9824 23264
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 9220 23044 9272 23050
rect 9220 22986 9272 22992
rect 8852 22772 8904 22778
rect 8852 22714 8904 22720
rect 8944 22772 8996 22778
rect 8944 22714 8996 22720
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8680 22506 8708 22578
rect 8576 22500 8628 22506
rect 8576 22442 8628 22448
rect 8668 22500 8720 22506
rect 8668 22442 8720 22448
rect 8680 21554 8708 22442
rect 8864 22030 8892 22714
rect 8956 22438 8984 22714
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 8864 21554 8892 21966
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8956 21350 8984 22374
rect 9140 22030 9168 22646
rect 9232 22080 9260 22986
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 9322 22876 9630 22896
rect 9322 22874 9328 22876
rect 9384 22874 9408 22876
rect 9464 22874 9488 22876
rect 9544 22874 9568 22876
rect 9624 22874 9630 22876
rect 9384 22822 9386 22874
rect 9566 22822 9568 22874
rect 9322 22820 9328 22822
rect 9384 22820 9408 22822
rect 9464 22820 9488 22822
rect 9544 22820 9568 22822
rect 9624 22820 9630 22822
rect 9322 22800 9630 22820
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9312 22092 9364 22098
rect 9232 22052 9312 22080
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8956 21128 8984 21286
rect 9048 21146 9076 21490
rect 9140 21418 9168 21830
rect 9128 21412 9180 21418
rect 9128 21354 9180 21360
rect 8864 21100 8984 21128
rect 9036 21140 9088 21146
rect 8864 20942 8892 21100
rect 9036 21082 9088 21088
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 8852 20936 8904 20942
rect 8852 20878 8904 20884
rect 8864 20602 8892 20878
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8588 16046 8616 20538
rect 8956 19990 8984 20946
rect 8944 19984 8996 19990
rect 8944 19926 8996 19932
rect 8852 19780 8904 19786
rect 8852 19722 8904 19728
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8680 19378 8708 19654
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8680 19174 8708 19314
rect 8864 19174 8892 19722
rect 8956 19446 8984 19926
rect 9048 19854 9076 21082
rect 9140 20398 9168 21354
rect 9232 21078 9260 22052
rect 9312 22034 9364 22040
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9322 21788 9630 21808
rect 9322 21786 9328 21788
rect 9384 21786 9408 21788
rect 9464 21786 9488 21788
rect 9544 21786 9568 21788
rect 9624 21786 9630 21788
rect 9384 21734 9386 21786
rect 9566 21734 9568 21786
rect 9322 21732 9328 21734
rect 9384 21732 9408 21734
rect 9464 21732 9488 21734
rect 9544 21732 9568 21734
rect 9624 21732 9630 21734
rect 9322 21712 9630 21732
rect 9692 21690 9720 21830
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9220 21072 9272 21078
rect 9220 21014 9272 21020
rect 9232 20534 9260 21014
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9322 20700 9630 20720
rect 9322 20698 9328 20700
rect 9384 20698 9408 20700
rect 9464 20698 9488 20700
rect 9544 20698 9568 20700
rect 9624 20698 9630 20700
rect 9384 20646 9386 20698
rect 9566 20646 9568 20698
rect 9322 20644 9328 20646
rect 9384 20644 9408 20646
rect 9464 20644 9488 20646
rect 9544 20644 9568 20646
rect 9624 20644 9630 20646
rect 9322 20624 9630 20644
rect 9220 20528 9272 20534
rect 9220 20470 9272 20476
rect 9692 20466 9720 20742
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9784 20448 9812 22170
rect 9876 21622 9904 22918
rect 9968 22778 9996 23054
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 10060 22642 10088 23598
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10060 21690 10088 21966
rect 10048 21684 10100 21690
rect 10244 21672 10272 28739
rect 10692 26512 10744 26518
rect 10692 26454 10744 26460
rect 10704 25498 10732 26454
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 10980 25974 11008 26318
rect 11256 26042 11284 26386
rect 11244 26036 11296 26042
rect 11244 25978 11296 25984
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 11336 25492 11388 25498
rect 11336 25434 11388 25440
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 10428 24886 10456 25094
rect 10416 24880 10468 24886
rect 10416 24822 10468 24828
rect 10704 24818 10732 25434
rect 11348 24954 11376 25434
rect 11428 25288 11480 25294
rect 11428 25230 11480 25236
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10704 24154 10732 24754
rect 11440 24410 11468 25230
rect 11520 25220 11572 25226
rect 11520 25162 11572 25168
rect 11532 24818 11560 25162
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11428 24404 11480 24410
rect 11428 24346 11480 24352
rect 10704 24126 10824 24154
rect 10796 23798 10824 24126
rect 10784 23792 10836 23798
rect 10784 23734 10836 23740
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10336 22030 10364 22578
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10244 21644 10364 21672
rect 10048 21626 10100 21632
rect 9864 21616 9916 21622
rect 9864 21558 9916 21564
rect 9876 20874 9904 21558
rect 10060 21418 10088 21626
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10048 21412 10100 21418
rect 10048 21354 10100 21360
rect 10060 21146 10088 21354
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 10244 20942 10272 21490
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 9864 20868 9916 20874
rect 9864 20810 9916 20816
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 9864 20460 9916 20466
rect 9784 20420 9864 20448
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 9140 20058 9168 20334
rect 9692 20330 9720 20402
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 9692 20058 9720 20266
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9784 19854 9812 20420
rect 9864 20402 9916 20408
rect 9862 20360 9918 20369
rect 9862 20295 9918 20304
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 8944 19440 8996 19446
rect 8944 19382 8996 19388
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8864 18970 8892 19110
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 8956 18766 8984 19246
rect 8944 18760 8996 18766
rect 8942 18728 8944 18737
rect 8996 18728 8998 18737
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8852 18692 8904 18698
rect 8942 18663 8998 18672
rect 8852 18634 8904 18640
rect 8680 18426 8708 18634
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8680 18290 8708 18362
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 8666 17232 8722 17241
rect 8666 17167 8668 17176
rect 8720 17167 8722 17176
rect 8668 17138 8720 17144
rect 8680 16794 8708 17138
rect 8772 17134 8800 17614
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8772 16794 8800 17070
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8680 16114 8708 16730
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8496 14006 8524 14554
rect 8484 14000 8536 14006
rect 8484 13942 8536 13948
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 13530 8524 13806
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8588 13326 8616 15574
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 8680 14074 8708 15030
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8772 14006 8800 15914
rect 8864 15094 8892 18634
rect 9140 18154 9168 19246
rect 9232 18766 9260 19722
rect 9322 19612 9630 19632
rect 9322 19610 9328 19612
rect 9384 19610 9408 19612
rect 9464 19610 9488 19612
rect 9544 19610 9568 19612
rect 9624 19610 9630 19612
rect 9384 19558 9386 19610
rect 9566 19558 9568 19610
rect 9322 19556 9328 19558
rect 9384 19556 9408 19558
rect 9464 19556 9488 19558
rect 9544 19556 9568 19558
rect 9624 19556 9630 19558
rect 9322 19536 9630 19556
rect 9680 18896 9732 18902
rect 9680 18838 9732 18844
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9322 18524 9630 18544
rect 9322 18522 9328 18524
rect 9384 18522 9408 18524
rect 9464 18522 9488 18524
rect 9544 18522 9568 18524
rect 9624 18522 9630 18524
rect 9384 18470 9386 18522
rect 9566 18470 9568 18522
rect 9322 18468 9328 18470
rect 9384 18468 9408 18470
rect 9464 18468 9488 18470
rect 9544 18468 9568 18470
rect 9624 18468 9630 18470
rect 9322 18448 9630 18468
rect 9692 18426 9720 18838
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9784 18290 9812 18702
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 9404 18148 9456 18154
rect 9404 18090 9456 18096
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9324 17678 9352 18022
rect 9416 17814 9444 18090
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9692 17610 9720 18226
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8852 15088 8904 15094
rect 8852 15030 8904 15036
rect 8760 14000 8812 14006
rect 8666 13968 8722 13977
rect 8956 13954 8984 17478
rect 8760 13942 8812 13948
rect 8666 13903 8722 13912
rect 8864 13926 8984 13954
rect 9048 13938 9076 17546
rect 9876 17524 9904 20295
rect 9968 20262 9996 20538
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10336 20346 10364 21644
rect 10428 20602 10456 22510
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10600 20596 10652 20602
rect 10600 20538 10652 20544
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 10244 19700 10272 20334
rect 10336 20318 10456 20346
rect 10324 20256 10376 20262
rect 10324 20198 10376 20204
rect 10336 19854 10364 20198
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10324 19712 10376 19718
rect 10244 19672 10324 19700
rect 10324 19654 10376 19660
rect 10232 19372 10284 19378
rect 10232 19314 10284 19320
rect 10244 18970 10272 19314
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10138 18864 10194 18873
rect 10138 18799 10194 18808
rect 10232 18828 10284 18834
rect 10152 18766 10180 18799
rect 10232 18770 10284 18776
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9968 17882 9996 18566
rect 10244 18290 10272 18770
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 10336 18086 10364 19654
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 9956 17536 10008 17542
rect 9876 17496 9956 17524
rect 9956 17478 10008 17484
rect 9322 17436 9630 17456
rect 9322 17434 9328 17436
rect 9384 17434 9408 17436
rect 9464 17434 9488 17436
rect 9544 17434 9568 17436
rect 9624 17434 9630 17436
rect 9384 17382 9386 17434
rect 9566 17382 9568 17434
rect 9322 17380 9328 17382
rect 9384 17380 9408 17382
rect 9464 17380 9488 17382
rect 9544 17380 9568 17382
rect 9624 17380 9630 17382
rect 9322 17360 9630 17380
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9140 17218 9168 17274
rect 9968 17270 9996 17478
rect 9496 17264 9548 17270
rect 9494 17232 9496 17241
rect 9956 17264 10008 17270
rect 9548 17232 9550 17241
rect 9140 17190 9352 17218
rect 9128 17128 9180 17134
rect 9180 17088 9260 17116
rect 9128 17070 9180 17076
rect 9232 16454 9260 17088
rect 9324 16794 9352 17190
rect 9404 17196 9456 17202
rect 9956 17206 10008 17212
rect 9494 17167 9550 17176
rect 9404 17138 9456 17144
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9416 16697 9444 17138
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9692 16810 9720 17002
rect 9508 16782 9720 16810
rect 9402 16688 9458 16697
rect 9402 16623 9458 16632
rect 9508 16522 9536 16782
rect 9586 16688 9642 16697
rect 9642 16646 9904 16674
rect 9586 16623 9642 16632
rect 9496 16516 9548 16522
rect 9496 16458 9548 16464
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9140 15366 9168 16050
rect 9232 16046 9260 16390
rect 9322 16348 9630 16368
rect 9322 16346 9328 16348
rect 9384 16346 9408 16348
rect 9464 16346 9488 16348
rect 9544 16346 9568 16348
rect 9624 16346 9630 16348
rect 9384 16294 9386 16346
rect 9566 16294 9568 16346
rect 9322 16292 9328 16294
rect 9384 16292 9408 16294
rect 9464 16292 9488 16294
rect 9544 16292 9568 16294
rect 9624 16292 9630 16294
rect 9322 16272 9630 16292
rect 9588 16176 9640 16182
rect 9586 16144 9588 16153
rect 9640 16144 9642 16153
rect 9784 16114 9812 16458
rect 9586 16079 9642 16088
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9232 14958 9260 15982
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9508 15706 9536 15914
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9600 15502 9628 15982
rect 9784 15570 9812 16050
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9322 15260 9630 15280
rect 9322 15258 9328 15260
rect 9384 15258 9408 15260
rect 9464 15258 9488 15260
rect 9544 15258 9568 15260
rect 9624 15258 9630 15260
rect 9384 15206 9386 15258
rect 9566 15206 9568 15258
rect 9322 15204 9328 15206
rect 9384 15204 9408 15206
rect 9464 15204 9488 15206
rect 9544 15204 9568 15206
rect 9624 15204 9630 15206
rect 9322 15184 9630 15204
rect 9692 15144 9720 15506
rect 9876 15162 9904 16646
rect 10152 16250 10180 17070
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 9864 15156 9916 15162
rect 9692 15116 9812 15144
rect 9496 15088 9548 15094
rect 9496 15030 9548 15036
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9508 14822 9536 15030
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9496 14816 9548 14822
rect 9494 14784 9496 14793
rect 9548 14784 9550 14793
rect 9494 14719 9550 14728
rect 9692 14618 9720 14962
rect 9784 14770 9812 15116
rect 9864 15098 9916 15104
rect 9784 14742 9904 14770
rect 9680 14612 9732 14618
rect 9732 14572 9812 14600
rect 9680 14554 9732 14560
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9036 13932 9088 13938
rect 8680 13818 8708 13903
rect 8680 13790 8800 13818
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8116 12912 8168 12918
rect 8404 12889 8432 12922
rect 8116 12854 8168 12860
rect 8390 12880 8446 12889
rect 8390 12815 8446 12824
rect 8680 12782 8708 13466
rect 8772 12850 8800 13790
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8496 12442 8524 12718
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8484 12436 8536 12442
rect 8864 12434 8892 13926
rect 9036 13874 9088 13880
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8956 13530 8984 13806
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 9048 13326 9076 13874
rect 9232 13394 9260 14350
rect 9322 14172 9630 14192
rect 9322 14170 9328 14172
rect 9384 14170 9408 14172
rect 9464 14170 9488 14172
rect 9544 14170 9568 14172
rect 9624 14170 9630 14172
rect 9384 14118 9386 14170
rect 9566 14118 9568 14170
rect 9322 14116 9328 14118
rect 9384 14116 9408 14118
rect 9464 14116 9488 14118
rect 9544 14116 9568 14118
rect 9624 14116 9630 14118
rect 9322 14096 9630 14116
rect 9312 14000 9364 14006
rect 9310 13968 9312 13977
rect 9364 13968 9366 13977
rect 9310 13903 9366 13912
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9036 13320 9088 13326
rect 9088 13280 9168 13308
rect 9036 13262 9088 13268
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8484 12378 8536 12384
rect 8588 12406 8892 12434
rect 7944 10674 7972 12378
rect 8496 12306 8524 12378
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8036 10674 8064 11630
rect 8496 11218 8524 12242
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8312 10266 8340 10950
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8312 9382 8340 9998
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8404 9194 8432 10134
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 8312 9166 8432 9194
rect 7852 8974 7880 9114
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 8312 8480 8340 9166
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8220 8452 8340 8480
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7116 7534 7236 7562
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6840 6458 6868 6802
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6656 5778 6684 6054
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6564 5409 6592 5578
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6550 5400 6606 5409
rect 6550 5335 6606 5344
rect 6656 5302 6684 5510
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6644 5160 6696 5166
rect 6642 5128 6644 5137
rect 6696 5128 6698 5137
rect 6642 5063 6698 5072
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4146 6684 4966
rect 6748 4826 6776 6258
rect 6840 5574 6868 6258
rect 6932 5778 6960 6598
rect 7024 6458 7052 7142
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5234 6868 5510
rect 6932 5302 6960 5714
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6748 4282 6776 4762
rect 6840 4622 6868 4762
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6932 4282 6960 5102
rect 7024 4826 7052 6394
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 7024 4010 7052 4490
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 7116 800 7144 7534
rect 7380 7472 7432 7478
rect 7208 7420 7380 7426
rect 7208 7414 7432 7420
rect 7208 7410 7420 7414
rect 7484 7410 7512 7822
rect 7760 7478 7788 7822
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7196 7404 7420 7410
rect 7248 7398 7420 7404
rect 7196 7346 7248 7352
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7208 5778 7236 6666
rect 7196 5772 7248 5778
rect 7248 5732 7328 5760
rect 7196 5714 7248 5720
rect 7194 5400 7250 5409
rect 7194 5335 7250 5344
rect 7208 5302 7236 5335
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7300 5166 7328 5732
rect 7392 5234 7420 7398
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7484 6798 7512 7346
rect 7760 7342 7788 7414
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7760 7002 7788 7278
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7576 6322 7604 6598
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7484 6118 7512 6258
rect 7852 6118 7880 6870
rect 8036 6458 8064 7278
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8128 6866 8156 7210
rect 8220 6905 8248 8452
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8206 6896 8262 6905
rect 8116 6860 8168 6866
rect 8206 6831 8262 6840
rect 8116 6802 8168 6808
rect 8128 6474 8156 6802
rect 8312 6730 8340 8298
rect 8404 8090 8432 8842
rect 8496 8566 8524 9590
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8404 7546 8432 8026
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8496 7478 8524 8502
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8300 6724 8352 6730
rect 8352 6684 8432 6712
rect 8300 6666 8352 6672
rect 8024 6452 8076 6458
rect 8128 6446 8248 6474
rect 8024 6394 8076 6400
rect 8220 6390 8248 6446
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7484 5846 7512 6054
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7576 5370 7604 5646
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7208 4622 7236 4762
rect 7392 4622 7420 5170
rect 7484 4865 7512 5170
rect 7470 4856 7526 4865
rect 7576 4826 7604 5306
rect 7852 5273 7880 6054
rect 7838 5264 7894 5273
rect 7656 5228 7708 5234
rect 7838 5199 7894 5208
rect 7656 5170 7708 5176
rect 7470 4791 7526 4800
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7380 4616 7432 4622
rect 7668 4604 7696 5170
rect 7748 5092 7800 5098
rect 7852 5080 7880 5199
rect 7944 5098 7972 6326
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8128 6118 8156 6258
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8128 5778 8156 6054
rect 8220 5846 8248 6326
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8220 5692 8248 5782
rect 8300 5704 8352 5710
rect 8220 5664 8300 5692
rect 8300 5646 8352 5652
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8022 5264 8078 5273
rect 8022 5199 8024 5208
rect 8076 5199 8078 5208
rect 8208 5228 8260 5234
rect 8024 5170 8076 5176
rect 8208 5170 8260 5176
rect 7800 5052 7880 5080
rect 7932 5092 7984 5098
rect 7748 5034 7800 5040
rect 7932 5034 7984 5040
rect 7840 4616 7892 4622
rect 7668 4576 7840 4604
rect 7380 4558 7432 4564
rect 7840 4558 7892 4564
rect 7392 4282 7420 4558
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7576 3738 7604 4082
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7760 3194 7788 4082
rect 7852 4010 7880 4558
rect 7944 4214 7972 5034
rect 8036 4826 8064 5170
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7840 4004 7892 4010
rect 7840 3946 7892 3952
rect 8128 3534 8156 4966
rect 8220 4622 8248 5170
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8220 4146 8248 4558
rect 8312 4486 8340 5510
rect 8404 5166 8432 6684
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8404 4622 8432 5102
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8496 3602 8524 7414
rect 8588 3738 8616 12406
rect 8956 12238 8984 13126
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9048 12050 9076 12650
rect 9140 12238 9168 13280
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9322 13084 9630 13104
rect 9322 13082 9328 13084
rect 9384 13082 9408 13084
rect 9464 13082 9488 13084
rect 9544 13082 9568 13084
rect 9624 13082 9630 13084
rect 9384 13030 9386 13082
rect 9566 13030 9568 13082
rect 9322 13028 9328 13030
rect 9384 13028 9408 13030
rect 9464 13028 9488 13030
rect 9544 13028 9568 13030
rect 9624 13028 9630 13030
rect 9322 13008 9630 13028
rect 9692 12986 9720 13194
rect 9784 12986 9812 14572
rect 9876 13190 9904 14742
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9784 12850 9812 12922
rect 9954 12880 10010 12889
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9772 12844 9824 12850
rect 9954 12815 9956 12824
rect 9772 12786 9824 12792
rect 10008 12815 10010 12824
rect 9956 12786 10008 12792
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9232 12102 9260 12718
rect 9416 12442 9444 12786
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9128 12096 9180 12102
rect 9048 12044 9128 12050
rect 9048 12038 9180 12044
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9048 12022 9168 12038
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 10062 8708 11494
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8772 10062 8800 10610
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8956 9586 8984 9862
rect 9048 9674 9076 11154
rect 9140 9994 9168 12022
rect 9232 10588 9260 12038
rect 9322 11996 9630 12016
rect 9322 11994 9328 11996
rect 9384 11994 9408 11996
rect 9464 11994 9488 11996
rect 9544 11994 9568 11996
rect 9624 11994 9630 11996
rect 9384 11942 9386 11994
rect 9566 11942 9568 11994
rect 9322 11940 9328 11942
rect 9384 11940 9408 11942
rect 9464 11940 9488 11942
rect 9544 11940 9568 11942
rect 9624 11940 9630 11942
rect 9322 11920 9630 11940
rect 9968 11830 9996 12038
rect 9588 11824 9640 11830
rect 9586 11792 9588 11801
rect 9956 11824 10008 11830
rect 9640 11792 9642 11801
rect 9496 11756 9548 11762
rect 9956 11766 10008 11772
rect 9586 11727 9642 11736
rect 9864 11756 9916 11762
rect 9496 11698 9548 11704
rect 9864 11698 9916 11704
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9416 11558 9444 11630
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9312 11348 9364 11354
rect 9508 11336 9536 11698
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9364 11308 9536 11336
rect 9312 11290 9364 11296
rect 9600 11218 9628 11494
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9322 10908 9630 10928
rect 9322 10906 9328 10908
rect 9384 10906 9408 10908
rect 9464 10906 9488 10908
rect 9544 10906 9568 10908
rect 9624 10906 9630 10908
rect 9384 10854 9386 10906
rect 9566 10854 9568 10906
rect 9322 10852 9328 10854
rect 9384 10852 9408 10854
rect 9464 10852 9488 10854
rect 9544 10852 9568 10854
rect 9624 10852 9630 10854
rect 9322 10832 9630 10852
rect 9692 10674 9720 10950
rect 9784 10810 9812 11630
rect 9876 11354 9904 11698
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9876 10810 9904 11290
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9404 10600 9456 10606
rect 9232 10560 9404 10588
rect 9864 10600 9916 10606
rect 9404 10542 9456 10548
rect 9600 10548 9864 10554
rect 9600 10542 9916 10548
rect 9416 10130 9444 10542
rect 9600 10526 9904 10542
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9600 9994 9628 10526
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9322 9820 9630 9840
rect 9322 9818 9328 9820
rect 9384 9818 9408 9820
rect 9464 9818 9488 9820
rect 9544 9818 9568 9820
rect 9624 9818 9630 9820
rect 9384 9766 9386 9818
rect 9566 9766 9568 9818
rect 9322 9764 9328 9766
rect 9384 9764 9408 9766
rect 9464 9764 9488 9766
rect 9544 9764 9568 9766
rect 9624 9764 9630 9766
rect 9322 9744 9630 9764
rect 9048 9646 9168 9674
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8772 8022 8800 8434
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8760 8016 8812 8022
rect 8666 7984 8722 7993
rect 8760 7958 8812 7964
rect 8666 7919 8722 7928
rect 8680 7886 8708 7919
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8680 7342 8708 7822
rect 8772 7410 8800 7958
rect 8864 7954 8892 8298
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8864 6798 8892 7890
rect 8956 7886 8984 8026
rect 9048 8022 9076 8230
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8956 7206 8984 7822
rect 9048 7449 9076 7822
rect 9034 7440 9090 7449
rect 9034 7375 9090 7384
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8956 6798 8984 7142
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8760 6656 8812 6662
rect 8956 6644 8984 6734
rect 8760 6598 8812 6604
rect 8864 6616 8984 6644
rect 8772 6361 8800 6598
rect 8758 6352 8814 6361
rect 8758 6287 8814 6296
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8680 4622 8708 5850
rect 8772 5846 8800 6122
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8772 4758 8800 5646
rect 8864 5642 8892 6616
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8850 5128 8906 5137
rect 8850 5063 8852 5072
rect 8904 5063 8906 5072
rect 8852 5034 8904 5040
rect 8760 4752 8812 4758
rect 8760 4694 8812 4700
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8956 4434 8984 6326
rect 9048 5370 9076 7278
rect 9140 7154 9168 9646
rect 10060 9330 10088 15302
rect 10152 15026 10180 16186
rect 10336 16182 10364 16934
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10244 14278 10272 14962
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10336 14482 10364 14758
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10244 12714 10272 14214
rect 10428 13530 10456 20318
rect 10520 18290 10548 20402
rect 10612 20330 10640 20538
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 10704 20058 10732 23666
rect 10796 23186 10824 23734
rect 10784 23180 10836 23186
rect 10784 23122 10836 23128
rect 11624 22094 11652 28750
rect 12084 28642 12112 28750
rect 12162 28739 12218 29539
rect 13174 28739 13230 29539
rect 14186 28739 14242 29539
rect 15106 28739 15162 29539
rect 16118 28739 16174 29539
rect 17038 28739 17094 29539
rect 18050 28739 18106 29539
rect 19062 28739 19118 29539
rect 19982 28739 20038 29539
rect 20088 28750 20392 28778
rect 12176 28642 12204 28739
rect 12084 28614 12204 28642
rect 11888 26308 11940 26314
rect 11888 26250 11940 26256
rect 12440 26308 12492 26314
rect 12440 26250 12492 26256
rect 11900 25974 11928 26250
rect 11888 25968 11940 25974
rect 11888 25910 11940 25916
rect 11900 25362 11928 25910
rect 12452 25838 12480 26250
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 12164 25356 12216 25362
rect 12164 25298 12216 25304
rect 11704 25152 11756 25158
rect 11704 25094 11756 25100
rect 11716 24614 11744 25094
rect 12176 24818 12204 25298
rect 12164 24812 12216 24818
rect 12164 24754 12216 24760
rect 12348 24676 12400 24682
rect 12348 24618 12400 24624
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11716 24206 11744 24550
rect 12360 24274 12388 24618
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 11808 23866 11836 24006
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 11900 23730 11928 24006
rect 12452 23866 12480 25774
rect 12624 25696 12676 25702
rect 12624 25638 12676 25644
rect 12636 25294 12664 25638
rect 13096 25498 13124 25842
rect 13188 25786 13216 28739
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 13508 26684 13816 26704
rect 13508 26682 13514 26684
rect 13570 26682 13594 26684
rect 13650 26682 13674 26684
rect 13730 26682 13754 26684
rect 13810 26682 13816 26684
rect 13570 26630 13572 26682
rect 13752 26630 13754 26682
rect 13508 26628 13514 26630
rect 13570 26628 13594 26630
rect 13650 26628 13674 26630
rect 13730 26628 13754 26630
rect 13810 26628 13816 26630
rect 13508 26608 13816 26628
rect 14108 26586 14136 26930
rect 14096 26580 14148 26586
rect 14096 26522 14148 26528
rect 13912 26512 13964 26518
rect 13912 26454 13964 26460
rect 13188 25758 13400 25786
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 13188 25498 13216 25638
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 13176 25492 13228 25498
rect 13176 25434 13228 25440
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 12624 24336 12676 24342
rect 12624 24278 12676 24284
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 12176 23526 12204 23666
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12176 23118 12204 23462
rect 12636 23322 12664 24278
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23866 13032 24074
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 11532 22066 11652 22094
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11164 21690 11192 21966
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10796 18834 10824 19110
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10520 17202 10548 18226
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10612 17678 10640 18090
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10520 14804 10548 17138
rect 10612 16590 10640 17614
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10612 15162 10640 16390
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10612 14958 10640 15098
rect 10704 15026 10732 15370
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10600 14816 10652 14822
rect 10520 14776 10600 14804
rect 10600 14758 10652 14764
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 10336 12442 10364 12786
rect 10428 12646 10456 13466
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10520 12850 10548 12922
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10336 12238 10364 12378
rect 10520 12238 10548 12786
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10232 12164 10284 12170
rect 10232 12106 10284 12112
rect 10244 11558 10272 12106
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10674 10548 10950
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10152 10062 10180 10406
rect 10244 10266 10272 10610
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10428 9586 10456 9998
rect 10612 9586 10640 14758
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12850 10732 13126
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10796 12434 10824 16050
rect 10704 12406 10824 12434
rect 10704 12102 10732 12406
rect 10980 12374 11008 20810
rect 11440 20398 11468 20878
rect 11428 20392 11480 20398
rect 11428 20334 11480 20340
rect 11440 19378 11468 20334
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11072 17542 11100 18566
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 11256 17338 11284 17546
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10704 9466 10732 12038
rect 10784 11756 10836 11762
rect 10980 11744 11008 12310
rect 11072 11898 11100 17138
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15434 11192 15846
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 11440 14890 11468 19314
rect 11532 16794 11560 22066
rect 11900 22030 11928 22578
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11900 21622 11928 21966
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 11992 21554 12020 21830
rect 12360 21690 12388 22034
rect 12452 21690 12480 22034
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12728 21622 12756 21830
rect 12716 21616 12768 21622
rect 12716 21558 12768 21564
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11992 21010 12020 21490
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12176 20262 12204 20878
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11716 19378 11744 19994
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11716 18834 11744 19314
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11164 12238 11192 12922
rect 11256 12782 11284 13194
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11256 12306 11284 12718
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11348 11898 11376 12786
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 10836 11716 11008 11744
rect 10784 11698 10836 11704
rect 11348 11150 11376 11834
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 10062 11008 10406
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10612 9438 10732 9466
rect 10784 9444 10836 9450
rect 10060 9302 10180 9330
rect 9322 8732 9630 8752
rect 9322 8730 9328 8732
rect 9384 8730 9408 8732
rect 9464 8730 9488 8732
rect 9544 8730 9568 8732
rect 9624 8730 9630 8732
rect 9384 8678 9386 8730
rect 9566 8678 9568 8730
rect 9322 8676 9328 8678
rect 9384 8676 9408 8678
rect 9464 8676 9488 8678
rect 9544 8676 9568 8678
rect 9624 8676 9630 8678
rect 9322 8656 9630 8676
rect 9220 8628 9272 8634
rect 9272 8588 9536 8616
rect 9220 8570 9272 8576
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9232 7970 9260 8434
rect 9232 7954 9444 7970
rect 9232 7948 9456 7954
rect 9232 7942 9404 7948
rect 9232 7546 9260 7942
rect 9404 7890 9456 7896
rect 9404 7812 9456 7818
rect 9508 7800 9536 8588
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9784 8090 9812 8502
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9864 8016 9916 8022
rect 9586 7984 9642 7993
rect 9864 7958 9916 7964
rect 9586 7919 9642 7928
rect 9600 7886 9628 7919
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9456 7772 9536 7800
rect 9680 7812 9732 7818
rect 9404 7754 9456 7760
rect 9680 7754 9732 7760
rect 9322 7644 9630 7664
rect 9322 7642 9328 7644
rect 9384 7642 9408 7644
rect 9464 7642 9488 7644
rect 9544 7642 9568 7644
rect 9624 7642 9630 7644
rect 9384 7590 9386 7642
rect 9566 7590 9568 7642
rect 9322 7588 9328 7590
rect 9384 7588 9408 7590
rect 9464 7588 9488 7590
rect 9544 7588 9568 7590
rect 9624 7588 9630 7590
rect 9322 7568 9630 7588
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9232 7342 9260 7482
rect 9692 7410 9720 7754
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9220 7336 9272 7342
rect 9876 7290 9904 7958
rect 9220 7278 9272 7284
rect 9784 7274 9904 7290
rect 9772 7268 9904 7274
rect 9824 7262 9904 7268
rect 9772 7210 9824 7216
rect 9140 7126 9260 7154
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9140 5710 9168 6394
rect 9232 6390 9260 7126
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 9322 6556 9630 6576
rect 9322 6554 9328 6556
rect 9384 6554 9408 6556
rect 9464 6554 9488 6556
rect 9544 6554 9568 6556
rect 9624 6554 9630 6556
rect 9384 6502 9386 6554
rect 9566 6502 9568 6554
rect 9322 6500 9328 6502
rect 9384 6500 9408 6502
rect 9464 6500 9488 6502
rect 9544 6500 9568 6502
rect 9624 6500 9630 6502
rect 9322 6480 9630 6500
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9232 5234 9260 6190
rect 10060 6118 10088 6666
rect 10152 6390 10180 9302
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10414 7440 10470 7449
rect 10414 7375 10416 7384
rect 10468 7375 10470 7384
rect 10416 7346 10468 7352
rect 10520 6662 10548 7958
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10520 6322 10548 6598
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9322 5468 9630 5488
rect 9322 5466 9328 5468
rect 9384 5466 9408 5468
rect 9464 5466 9488 5468
rect 9544 5466 9568 5468
rect 9624 5466 9630 5468
rect 9384 5414 9386 5466
rect 9566 5414 9568 5466
rect 9322 5412 9328 5414
rect 9384 5412 9408 5414
rect 9464 5412 9488 5414
rect 9544 5412 9568 5414
rect 9624 5412 9630 5414
rect 9322 5392 9630 5412
rect 10060 5234 10088 6054
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9034 4856 9090 4865
rect 9034 4791 9090 4800
rect 9048 4758 9076 4791
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 9140 4690 9168 5170
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 8680 4406 8984 4434
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8482 3360 8538 3369
rect 8482 3295 8538 3304
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 8496 800 8524 3295
rect 8588 3126 8616 3470
rect 8680 3398 8708 4406
rect 9232 4078 9260 4966
rect 9322 4380 9630 4400
rect 9322 4378 9328 4380
rect 9384 4378 9408 4380
rect 9464 4378 9488 4380
rect 9544 4378 9568 4380
rect 9624 4378 9630 4380
rect 9384 4326 9386 4378
rect 9566 4326 9568 4378
rect 9322 4324 9328 4326
rect 9384 4324 9408 4326
rect 9464 4324 9488 4326
rect 9544 4324 9568 4326
rect 9624 4324 9630 4326
rect 9322 4304 9630 4324
rect 10060 4214 10088 5170
rect 10152 4282 10180 5238
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10244 4826 10272 4966
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10428 4282 10456 5510
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8772 3194 8800 3674
rect 8850 3632 8906 3641
rect 8850 3567 8906 3576
rect 8864 3534 8892 3567
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8864 2990 8892 3470
rect 8956 3466 8984 3878
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 9048 3058 9076 3538
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9140 3126 9168 3334
rect 9232 3194 9260 3470
rect 9322 3292 9630 3312
rect 9322 3290 9328 3292
rect 9384 3290 9408 3292
rect 9464 3290 9488 3292
rect 9544 3290 9568 3292
rect 9624 3290 9630 3292
rect 9384 3238 9386 3290
rect 9566 3238 9568 3290
rect 9322 3236 9328 3238
rect 9384 3236 9408 3238
rect 9464 3236 9488 3238
rect 9544 3236 9568 3238
rect 9624 3236 9630 3238
rect 9322 3216 9630 3236
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 9232 1358 9260 3130
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9692 2650 9720 2994
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9876 2446 9904 3878
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9322 2204 9630 2224
rect 9322 2202 9328 2204
rect 9384 2202 9408 2204
rect 9464 2202 9488 2204
rect 9544 2202 9568 2204
rect 9624 2202 9630 2204
rect 9384 2150 9386 2202
rect 9566 2150 9568 2202
rect 9322 2148 9328 2150
rect 9384 2148 9408 2150
rect 9464 2148 9488 2150
rect 9544 2148 9568 2150
rect 9624 2148 9630 2150
rect 9322 2128 9630 2148
rect 10612 1442 10640 9438
rect 10784 9386 10836 9392
rect 10796 8634 10824 9386
rect 11164 8974 11192 9522
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 10888 6458 10916 7346
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10704 5710 10732 6258
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10704 5234 10732 5646
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10888 4622 10916 4966
rect 10980 4690 11008 6598
rect 11072 6458 11100 7142
rect 11164 6798 11192 7346
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11256 6322 11284 7210
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 6798 11376 7142
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11256 5250 11284 6258
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10980 4146 11008 4626
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11072 4078 11100 4694
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10968 3460 11020 3466
rect 10968 3402 11020 3408
rect 10980 3194 11008 3402
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 11164 3058 11192 5238
rect 11256 5222 11376 5250
rect 11348 5166 11376 5222
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11348 4214 11376 4558
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11256 3738 11284 4082
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11348 3602 11376 4150
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11348 3126 11376 3538
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 10244 1414 10640 1442
rect 9220 1352 9272 1358
rect 9220 1294 9272 1300
rect 9784 870 9904 898
rect 9784 800 9812 870
rect 662 0 718 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 8482 0 8538 800
rect 9770 0 9826 800
rect 9876 762 9904 870
rect 10244 762 10272 1414
rect 11072 870 11192 898
rect 11072 800 11100 870
rect 9876 734 10272 762
rect 11058 0 11114 800
rect 11164 762 11192 870
rect 11440 762 11468 13126
rect 11532 12918 11560 13670
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11624 11694 11652 18566
rect 11808 18222 11836 19790
rect 11900 19310 11928 20198
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12176 19514 12204 19722
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12452 19446 12480 21082
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12544 20466 12572 20810
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12636 19514 12664 19654
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11888 19304 11940 19310
rect 11888 19246 11940 19252
rect 11900 18834 11928 19246
rect 12084 18970 12112 19314
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11900 18426 11928 18770
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11716 17626 11744 18022
rect 11808 17882 11836 18158
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11716 17598 11836 17626
rect 12176 17610 12204 19178
rect 12452 19174 12480 19382
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12268 17678 12296 17818
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 16114 11744 16390
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11716 11830 11744 12922
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11624 10266 11652 10610
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 7274 11652 8230
rect 11716 7750 11744 8774
rect 11808 8498 11836 17598
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11900 13326 11928 16730
rect 12268 16522 12296 17478
rect 12360 17066 12388 18634
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12452 18358 12480 18566
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12348 17060 12400 17066
rect 12348 17002 12400 17008
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12072 14816 12124 14822
rect 12070 14784 12072 14793
rect 12124 14784 12126 14793
rect 12070 14719 12126 14728
rect 12176 14414 12204 16050
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 11992 13394 12020 13670
rect 12084 13394 12112 14214
rect 12268 13938 12296 16458
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12360 14346 12388 14962
rect 12544 14498 12572 18702
rect 12636 16250 12664 19314
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12728 17542 12756 17818
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12728 15638 12756 17070
rect 12820 16454 12848 22918
rect 13004 22710 13032 23802
rect 12992 22704 13044 22710
rect 12992 22646 13044 22652
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12912 19174 12940 20402
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 18766 12940 19110
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 13004 18698 13032 19790
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 13004 18408 13032 18634
rect 12912 18380 13032 18408
rect 12912 16794 12940 18380
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13004 16998 13032 18226
rect 13096 17678 13124 18702
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13096 17202 13124 17614
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12808 16040 12860 16046
rect 12912 16028 12940 16730
rect 12860 16000 12940 16028
rect 12808 15982 12860 15988
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12624 15496 12676 15502
rect 12820 15473 12848 15982
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12624 15438 12676 15444
rect 12806 15464 12862 15473
rect 12636 15162 12664 15438
rect 12806 15399 12862 15408
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12728 14618 12756 14962
rect 12820 14958 12848 15302
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12544 14470 12756 14498
rect 12532 14408 12584 14414
rect 12584 14368 12664 14396
rect 12532 14350 12584 14356
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12636 13938 12664 14368
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11900 13190 11928 13262
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11900 10674 11928 11698
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11808 7290 11836 8434
rect 11900 7546 11928 10610
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11992 8090 12020 8366
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11716 7262 11836 7290
rect 11624 7041 11652 7210
rect 11610 7032 11666 7041
rect 11520 6996 11572 7002
rect 11610 6967 11666 6976
rect 11520 6938 11572 6944
rect 11532 6186 11560 6938
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11716 5642 11744 7262
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11808 6730 11836 7142
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11900 5234 11928 7482
rect 12084 7410 12112 8842
rect 12176 8514 12204 13466
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12268 12986 12296 13262
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12268 11762 12296 12582
rect 12360 12442 12388 12582
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12452 12238 12480 12786
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12360 11082 12388 12038
rect 12452 11830 12480 12174
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12452 10606 12480 11766
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 9654 12480 10542
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12360 9110 12388 9522
rect 12544 9178 12572 9998
rect 12636 9654 12664 13874
rect 12728 12434 12756 14470
rect 12820 14414 12848 14894
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12912 13818 12940 15846
rect 12820 13790 12940 13818
rect 12820 13308 12848 13790
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 13462 12940 13670
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12820 13280 12940 13308
rect 12728 12406 12848 12434
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12728 10266 12756 10610
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12728 9110 12756 9454
rect 12820 9450 12848 12406
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12820 9110 12848 9386
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12452 8634 12480 8910
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12176 8498 12296 8514
rect 12176 8492 12308 8498
rect 12176 8486 12256 8492
rect 12256 8434 12308 8440
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12176 7886 12204 8366
rect 12256 8288 12308 8294
rect 12452 8242 12480 8570
rect 12256 8230 12308 8236
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 7206 12112 7346
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12176 5778 12204 7822
rect 12268 7818 12296 8230
rect 12360 8214 12480 8242
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12268 6798 12296 7278
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12360 6254 12388 8214
rect 12636 8022 12664 8910
rect 12820 8634 12848 8910
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12360 5574 12388 6190
rect 12544 6118 12572 6734
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 12360 4826 12388 5510
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11624 4146 11652 4558
rect 12452 4554 12480 4966
rect 12636 4622 12664 7686
rect 12912 7002 12940 13280
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12912 6746 12940 6938
rect 12820 6718 12940 6746
rect 12820 5710 12848 6718
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11532 2990 11560 3470
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11624 3126 11652 3334
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 11808 3058 11836 3878
rect 11900 3738 11928 3946
rect 12176 3942 12204 4422
rect 12452 4214 12480 4490
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 12820 3942 12848 5034
rect 13004 4026 13032 16934
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13096 15706 13124 16390
rect 13188 15978 13216 25094
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 13280 19718 13308 20538
rect 13268 19712 13320 19718
rect 13268 19654 13320 19660
rect 13280 17134 13308 19654
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13280 16794 13308 17070
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13372 16697 13400 25758
rect 13508 25596 13816 25616
rect 13508 25594 13514 25596
rect 13570 25594 13594 25596
rect 13650 25594 13674 25596
rect 13730 25594 13754 25596
rect 13810 25594 13816 25596
rect 13570 25542 13572 25594
rect 13752 25542 13754 25594
rect 13508 25540 13514 25542
rect 13570 25540 13594 25542
rect 13650 25540 13674 25542
rect 13730 25540 13754 25542
rect 13810 25540 13816 25542
rect 13508 25520 13816 25540
rect 13924 25498 13952 26454
rect 14200 26330 14228 28739
rect 14648 26784 14700 26790
rect 14648 26726 14700 26732
rect 14096 26308 14148 26314
rect 14200 26302 14320 26330
rect 14096 26250 14148 26256
rect 14004 25968 14056 25974
rect 14004 25910 14056 25916
rect 13912 25492 13964 25498
rect 13912 25434 13964 25440
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13508 24508 13816 24528
rect 13508 24506 13514 24508
rect 13570 24506 13594 24508
rect 13650 24506 13674 24508
rect 13730 24506 13754 24508
rect 13810 24506 13816 24508
rect 13570 24454 13572 24506
rect 13752 24454 13754 24506
rect 13508 24452 13514 24454
rect 13570 24452 13594 24454
rect 13650 24452 13674 24454
rect 13730 24452 13754 24454
rect 13810 24452 13816 24454
rect 13508 24432 13816 24452
rect 13924 24138 13952 24754
rect 13912 24132 13964 24138
rect 13912 24074 13964 24080
rect 13924 23866 13952 24074
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 14016 23730 14044 25910
rect 14108 25294 14136 26250
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 14292 24954 14320 26302
rect 14660 25974 14688 26726
rect 14740 26512 14792 26518
rect 15120 26466 15148 28739
rect 14740 26454 14792 26460
rect 14752 26246 14780 26454
rect 15028 26438 15148 26466
rect 14924 26308 14976 26314
rect 14924 26250 14976 26256
rect 14740 26240 14792 26246
rect 14740 26182 14792 26188
rect 14648 25968 14700 25974
rect 14648 25910 14700 25916
rect 14752 25702 14780 26182
rect 14740 25696 14792 25702
rect 14792 25644 14872 25650
rect 14740 25638 14872 25644
rect 14752 25622 14872 25638
rect 14740 25220 14792 25226
rect 14740 25162 14792 25168
rect 14280 24948 14332 24954
rect 14280 24890 14332 24896
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14648 24744 14700 24750
rect 14648 24686 14700 24692
rect 14108 24206 14136 24686
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 14384 24342 14412 24550
rect 14568 24410 14596 24686
rect 14556 24404 14608 24410
rect 14556 24346 14608 24352
rect 14372 24336 14424 24342
rect 14372 24278 14424 24284
rect 14660 24206 14688 24686
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14648 24064 14700 24070
rect 14648 24006 14700 24012
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 14096 23724 14148 23730
rect 14096 23666 14148 23672
rect 13508 23420 13816 23440
rect 13508 23418 13514 23420
rect 13570 23418 13594 23420
rect 13650 23418 13674 23420
rect 13730 23418 13754 23420
rect 13810 23418 13816 23420
rect 13570 23366 13572 23418
rect 13752 23366 13754 23418
rect 13508 23364 13514 23366
rect 13570 23364 13594 23366
rect 13650 23364 13674 23366
rect 13730 23364 13754 23366
rect 13810 23364 13816 23366
rect 13508 23344 13816 23364
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13832 22778 13860 23054
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 14016 22710 14044 23666
rect 14108 23322 14136 23666
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14004 22704 14056 22710
rect 14004 22646 14056 22652
rect 13508 22332 13816 22352
rect 13508 22330 13514 22332
rect 13570 22330 13594 22332
rect 13650 22330 13674 22332
rect 13730 22330 13754 22332
rect 13810 22330 13816 22332
rect 13570 22278 13572 22330
rect 13752 22278 13754 22330
rect 13508 22276 13514 22278
rect 13570 22276 13594 22278
rect 13650 22276 13674 22278
rect 13730 22276 13754 22278
rect 13810 22276 13816 22278
rect 13508 22256 13816 22276
rect 14016 22098 14044 22646
rect 14108 22506 14136 22918
rect 14096 22500 14148 22506
rect 14096 22442 14148 22448
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 14016 21554 14044 22034
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13508 21244 13816 21264
rect 13508 21242 13514 21244
rect 13570 21242 13594 21244
rect 13650 21242 13674 21244
rect 13730 21242 13754 21244
rect 13810 21242 13816 21244
rect 13570 21190 13572 21242
rect 13752 21190 13754 21242
rect 13508 21188 13514 21190
rect 13570 21188 13594 21190
rect 13650 21188 13674 21190
rect 13730 21188 13754 21190
rect 13810 21188 13816 21190
rect 13508 21168 13816 21188
rect 13636 20800 13688 20806
rect 13636 20742 13688 20748
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 13648 20602 13676 20742
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 14108 20466 14136 20742
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 13508 20156 13816 20176
rect 13508 20154 13514 20156
rect 13570 20154 13594 20156
rect 13650 20154 13674 20156
rect 13730 20154 13754 20156
rect 13810 20154 13816 20156
rect 13570 20102 13572 20154
rect 13752 20102 13754 20154
rect 13508 20100 13514 20102
rect 13570 20100 13594 20102
rect 13650 20100 13674 20102
rect 13730 20100 13754 20102
rect 13810 20100 13816 20102
rect 13508 20080 13816 20100
rect 14108 19922 14136 20402
rect 14200 20398 14228 21626
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 14384 20602 14412 20810
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 14004 19780 14056 19786
rect 14004 19722 14056 19728
rect 14016 19378 14044 19722
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 13508 19068 13816 19088
rect 13508 19066 13514 19068
rect 13570 19066 13594 19068
rect 13650 19066 13674 19068
rect 13730 19066 13754 19068
rect 13810 19066 13816 19068
rect 13570 19014 13572 19066
rect 13752 19014 13754 19066
rect 13508 19012 13514 19014
rect 13570 19012 13594 19014
rect 13650 19012 13674 19014
rect 13730 19012 13754 19014
rect 13810 19012 13816 19014
rect 13508 18992 13816 19012
rect 14200 18834 14228 19314
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14108 18222 14136 18702
rect 14200 18426 14228 18770
rect 14476 18630 14504 19314
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14004 18148 14056 18154
rect 14004 18090 14056 18096
rect 13508 17980 13816 18000
rect 13508 17978 13514 17980
rect 13570 17978 13594 17980
rect 13650 17978 13674 17980
rect 13730 17978 13754 17980
rect 13810 17978 13816 17980
rect 13570 17926 13572 17978
rect 13752 17926 13754 17978
rect 13508 17924 13514 17926
rect 13570 17924 13594 17926
rect 13650 17924 13674 17926
rect 13730 17924 13754 17926
rect 13810 17924 13816 17926
rect 13508 17904 13816 17924
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13556 17202 13584 17546
rect 13740 17218 13768 17614
rect 13740 17202 13952 17218
rect 13544 17196 13596 17202
rect 13740 17196 13964 17202
rect 13740 17190 13912 17196
rect 13544 17138 13596 17144
rect 13912 17138 13964 17144
rect 13924 16998 13952 17138
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13508 16892 13816 16912
rect 13508 16890 13514 16892
rect 13570 16890 13594 16892
rect 13650 16890 13674 16892
rect 13730 16890 13754 16892
rect 13810 16890 13816 16892
rect 13570 16838 13572 16890
rect 13752 16838 13754 16890
rect 13508 16836 13514 16838
rect 13570 16836 13594 16838
rect 13650 16836 13674 16838
rect 13730 16836 13754 16838
rect 13810 16836 13816 16838
rect 13508 16816 13816 16836
rect 13358 16688 13414 16697
rect 13358 16623 13414 16632
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13280 15858 13308 16390
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13188 15830 13308 15858
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13082 15464 13138 15473
rect 13082 15399 13138 15408
rect 13096 14618 13124 15399
rect 13188 15366 13216 15830
rect 13372 15638 13400 15982
rect 13508 15804 13816 15824
rect 13508 15802 13514 15804
rect 13570 15802 13594 15804
rect 13650 15802 13674 15804
rect 13730 15802 13754 15804
rect 13810 15802 13816 15804
rect 13570 15750 13572 15802
rect 13752 15750 13754 15802
rect 13508 15748 13514 15750
rect 13570 15748 13594 15750
rect 13650 15748 13674 15750
rect 13730 15748 13754 15750
rect 13810 15748 13816 15750
rect 13508 15728 13816 15748
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 13096 10742 13124 13398
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 13188 9654 13216 15302
rect 13280 13802 13308 15370
rect 13372 14498 13400 15574
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13508 14716 13816 14736
rect 13508 14714 13514 14716
rect 13570 14714 13594 14716
rect 13650 14714 13674 14716
rect 13730 14714 13754 14716
rect 13810 14714 13816 14716
rect 13570 14662 13572 14714
rect 13752 14662 13754 14714
rect 13508 14660 13514 14662
rect 13570 14660 13594 14662
rect 13650 14660 13674 14662
rect 13730 14660 13754 14662
rect 13810 14660 13816 14662
rect 13508 14640 13816 14660
rect 13924 14550 13952 15438
rect 14016 14958 14044 18090
rect 14108 17746 14136 18158
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 14292 17270 14320 18226
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13912 14544 13964 14550
rect 13372 14470 13584 14498
rect 13912 14486 13964 14492
rect 13372 14414 13400 14470
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13464 14006 13492 14350
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13556 13938 13584 14470
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13832 13938 13860 14418
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13728 13864 13780 13870
rect 13372 13812 13728 13818
rect 13372 13806 13780 13812
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13372 13790 13768 13806
rect 13372 13326 13400 13790
rect 13508 13628 13816 13648
rect 13508 13626 13514 13628
rect 13570 13626 13594 13628
rect 13650 13626 13674 13628
rect 13730 13626 13754 13628
rect 13810 13626 13816 13628
rect 13570 13574 13572 13626
rect 13752 13574 13754 13626
rect 13508 13572 13514 13574
rect 13570 13572 13594 13574
rect 13650 13572 13674 13574
rect 13730 13572 13754 13574
rect 13810 13572 13816 13574
rect 13508 13552 13816 13572
rect 14016 13530 14044 14350
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14016 13326 14044 13466
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13280 12918 13308 13194
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13508 12540 13816 12560
rect 13508 12538 13514 12540
rect 13570 12538 13594 12540
rect 13650 12538 13674 12540
rect 13730 12538 13754 12540
rect 13810 12538 13816 12540
rect 13570 12486 13572 12538
rect 13752 12486 13754 12538
rect 13508 12484 13514 12486
rect 13570 12484 13594 12486
rect 13650 12484 13674 12486
rect 13730 12484 13754 12486
rect 13810 12484 13816 12486
rect 13508 12464 13816 12484
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13508 11452 13816 11472
rect 13508 11450 13514 11452
rect 13570 11450 13594 11452
rect 13650 11450 13674 11452
rect 13730 11450 13754 11452
rect 13810 11450 13816 11452
rect 13570 11398 13572 11450
rect 13752 11398 13754 11450
rect 13508 11396 13514 11398
rect 13570 11396 13594 11398
rect 13650 11396 13674 11398
rect 13730 11396 13754 11398
rect 13810 11396 13816 11398
rect 13508 11376 13816 11396
rect 13924 11354 13952 11698
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14108 10810 14136 17070
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14384 16250 14412 17002
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14200 15366 14228 16050
rect 14292 15502 14320 16050
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14384 15570 14412 15982
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 13508 10364 13816 10384
rect 13508 10362 13514 10364
rect 13570 10362 13594 10364
rect 13650 10362 13674 10364
rect 13730 10362 13754 10364
rect 13810 10362 13816 10364
rect 13570 10310 13572 10362
rect 13752 10310 13754 10362
rect 13508 10308 13514 10310
rect 13570 10308 13594 10310
rect 13650 10308 13674 10310
rect 13730 10308 13754 10310
rect 13810 10308 13816 10310
rect 13508 10288 13816 10308
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13096 8634 13124 9454
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13188 8566 13216 9590
rect 13280 9058 13308 9862
rect 13556 9518 13584 9998
rect 14108 9994 14136 10066
rect 14200 10062 14228 15302
rect 14292 14074 14320 15438
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14384 14074 14412 14554
rect 14476 14414 14504 14758
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14384 13530 14412 14010
rect 14476 13938 14504 14214
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14384 13394 14412 13466
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14476 13326 14504 13738
rect 14568 13530 14596 23054
rect 14660 23050 14688 24006
rect 14648 23044 14700 23050
rect 14648 22986 14700 22992
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14660 19514 14688 20402
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14660 18698 14688 19110
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 14752 14618 14780 25162
rect 14844 24614 14872 25622
rect 14936 25362 14964 26250
rect 15028 26042 15056 26438
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 15016 26036 15068 26042
rect 15016 25978 15068 25984
rect 14924 25356 14976 25362
rect 14924 25298 14976 25304
rect 15016 25220 15068 25226
rect 15016 25162 15068 25168
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 14844 24410 14872 24550
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 14832 24132 14884 24138
rect 14832 24074 14884 24080
rect 14844 22982 14872 24074
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 14844 20058 14872 20402
rect 14936 20346 14964 24890
rect 15028 24698 15056 25162
rect 15120 24818 15148 26318
rect 16132 25974 16160 28739
rect 16120 25968 16172 25974
rect 16120 25910 16172 25916
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 16672 25832 16724 25838
rect 16672 25774 16724 25780
rect 15752 25696 15804 25702
rect 15752 25638 15804 25644
rect 15764 25362 15792 25638
rect 16684 25362 16712 25774
rect 16776 25498 16804 25842
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 15200 25356 15252 25362
rect 15200 25298 15252 25304
rect 15752 25356 15804 25362
rect 15752 25298 15804 25304
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 15212 24818 15240 25298
rect 15476 25288 15528 25294
rect 15476 25230 15528 25236
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 15488 24954 15516 25230
rect 16500 24954 16528 25230
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 15476 24948 15528 24954
rect 15476 24890 15528 24896
rect 16488 24948 16540 24954
rect 16488 24890 16540 24896
rect 15108 24812 15160 24818
rect 15108 24754 15160 24760
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15028 24670 15148 24698
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 15028 24206 15056 24550
rect 15120 24342 15148 24670
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15212 24410 15240 24550
rect 15200 24404 15252 24410
rect 15200 24346 15252 24352
rect 15108 24336 15160 24342
rect 15108 24278 15160 24284
rect 15016 24200 15068 24206
rect 15016 24142 15068 24148
rect 15120 23322 15148 24278
rect 15488 24274 15516 24890
rect 16592 24886 16620 25094
rect 16580 24880 16632 24886
rect 16580 24822 16632 24828
rect 16684 24818 16712 25298
rect 16856 25288 16908 25294
rect 16856 25230 16908 25236
rect 16764 25220 16816 25226
rect 16764 25162 16816 25168
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16212 24676 16264 24682
rect 16212 24618 16264 24624
rect 16224 24410 16252 24618
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15384 24200 15436 24206
rect 15384 24142 15436 24148
rect 15396 23866 15424 24142
rect 16592 24138 16620 24686
rect 16776 24274 16804 25162
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16868 24154 16896 25230
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16776 24126 16896 24154
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 16212 22568 16264 22574
rect 16212 22510 16264 22516
rect 15016 22092 15068 22098
rect 15016 22034 15068 22040
rect 15028 21486 15056 22034
rect 15304 22030 15332 22510
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15488 22030 15516 22374
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 16224 21622 16252 22510
rect 16212 21616 16264 21622
rect 16212 21558 16264 21564
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 15028 20942 15056 21422
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 20466 15240 20742
rect 15304 20602 15332 20810
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15396 20482 15424 20538
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15304 20454 15424 20482
rect 15304 20398 15332 20454
rect 15292 20392 15344 20398
rect 14936 20318 15148 20346
rect 15292 20334 15344 20340
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14936 19786 14964 20198
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14844 18873 14872 19110
rect 14830 18864 14886 18873
rect 14830 18799 14886 18808
rect 15120 18086 15148 20318
rect 15200 20324 15252 20330
rect 15200 20266 15252 20272
rect 15212 20058 15240 20266
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15304 19922 15332 20334
rect 15488 19922 15516 20878
rect 16040 20466 16068 21286
rect 16132 20602 16160 21490
rect 16224 21010 16252 21558
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 15764 20058 15792 20334
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15212 19514 15240 19790
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15304 19310 15332 19858
rect 15764 19446 15792 19994
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15304 18970 15332 19246
rect 15764 18970 15792 19382
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15660 18692 15712 18698
rect 15660 18634 15712 18640
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15384 17808 15436 17814
rect 15384 17750 15436 17756
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15212 15910 15240 15982
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15212 15609 15240 15846
rect 15304 15706 15332 16458
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15198 15600 15254 15609
rect 14832 15564 14884 15570
rect 15198 15535 15254 15544
rect 14832 15506 14884 15512
rect 14844 14822 14872 15506
rect 15396 15434 15424 17750
rect 15580 17338 15608 18362
rect 15672 18329 15700 18634
rect 15658 18320 15714 18329
rect 15658 18255 15714 18264
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 16454 15516 16594
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 14660 13802 14688 14486
rect 14844 14414 14872 14758
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14844 14006 14872 14214
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14292 10010 14320 13262
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 9586 13860 9862
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 14108 9518 14136 9930
rect 14200 9654 14228 9998
rect 14292 9994 14412 10010
rect 14292 9988 14424 9994
rect 14292 9982 14372 9988
rect 14372 9930 14424 9936
rect 14188 9648 14240 9654
rect 14240 9608 14320 9636
rect 14188 9590 14240 9596
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13372 9178 13400 9318
rect 13508 9276 13816 9296
rect 13508 9274 13514 9276
rect 13570 9274 13594 9276
rect 13650 9274 13674 9276
rect 13730 9274 13754 9276
rect 13810 9274 13816 9276
rect 13570 9222 13572 9274
rect 13752 9222 13754 9274
rect 13508 9220 13514 9222
rect 13570 9220 13594 9222
rect 13650 9220 13674 9222
rect 13730 9220 13754 9222
rect 13810 9220 13816 9222
rect 13508 9200 13816 9220
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13280 9030 13400 9058
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13096 8090 13124 8230
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13188 7954 13216 8502
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13280 6798 13308 8774
rect 13372 8294 13400 9030
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13740 8498 13768 8910
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13508 8188 13816 8208
rect 13508 8186 13514 8188
rect 13570 8186 13594 8188
rect 13650 8186 13674 8188
rect 13730 8186 13754 8188
rect 13810 8186 13816 8188
rect 13570 8134 13572 8186
rect 13752 8134 13754 8186
rect 13508 8132 13514 8134
rect 13570 8132 13594 8134
rect 13650 8132 13674 8134
rect 13730 8132 13754 8134
rect 13810 8132 13816 8134
rect 13508 8112 13816 8132
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13096 6458 13124 6734
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13372 5370 13400 7958
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13508 7100 13816 7120
rect 13508 7098 13514 7100
rect 13570 7098 13594 7100
rect 13650 7098 13674 7100
rect 13730 7098 13754 7100
rect 13810 7098 13816 7100
rect 13570 7046 13572 7098
rect 13752 7046 13754 7098
rect 13508 7044 13514 7046
rect 13570 7044 13594 7046
rect 13650 7044 13674 7046
rect 13730 7044 13754 7046
rect 13810 7044 13816 7046
rect 13508 7024 13816 7044
rect 13924 7002 13952 7346
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 14016 6866 14044 7346
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13508 6012 13816 6032
rect 13508 6010 13514 6012
rect 13570 6010 13594 6012
rect 13650 6010 13674 6012
rect 13730 6010 13754 6012
rect 13810 6010 13816 6012
rect 13570 5958 13572 6010
rect 13752 5958 13754 6010
rect 13508 5956 13514 5958
rect 13570 5956 13594 5958
rect 13650 5956 13674 5958
rect 13730 5956 13754 5958
rect 13810 5956 13816 5958
rect 13508 5936 13816 5956
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13832 5166 13860 5510
rect 14016 5250 14044 6802
rect 14108 5370 14136 8774
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14200 7886 14228 8230
rect 14292 7954 14320 9608
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14384 8498 14412 9318
rect 14476 8974 14504 9318
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 7206 14320 7346
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 13924 5222 14044 5250
rect 14096 5228 14148 5234
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13096 4690 13124 4966
rect 13508 4924 13816 4944
rect 13508 4922 13514 4924
rect 13570 4922 13594 4924
rect 13650 4922 13674 4924
rect 13730 4922 13754 4924
rect 13810 4922 13816 4924
rect 13570 4870 13572 4922
rect 13752 4870 13754 4922
rect 13508 4868 13514 4870
rect 13570 4868 13594 4870
rect 13650 4868 13674 4870
rect 13730 4868 13754 4870
rect 13810 4868 13816 4870
rect 13508 4848 13816 4868
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4282 13124 4422
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13924 4146 13952 5222
rect 14096 5170 14148 5176
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14016 4826 14044 4966
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14016 4146 14044 4422
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 12912 3998 13032 4026
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12452 3194 12480 3402
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 12544 2990 12572 3334
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12912 2854 12940 3998
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3466 13032 3878
rect 12992 3460 13044 3466
rect 12992 3402 13044 3408
rect 13188 3398 13216 4014
rect 13280 3398 13308 4014
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 13188 2446 13216 3334
rect 13280 2446 13308 3334
rect 13372 3194 13400 4082
rect 13508 3836 13816 3856
rect 13508 3834 13514 3836
rect 13570 3834 13594 3836
rect 13650 3834 13674 3836
rect 13730 3834 13754 3836
rect 13810 3834 13816 3836
rect 13570 3782 13572 3834
rect 13752 3782 13754 3834
rect 13508 3780 13514 3782
rect 13570 3780 13594 3782
rect 13650 3780 13674 3782
rect 13730 3780 13754 3782
rect 13810 3780 13816 3782
rect 13508 3760 13816 3780
rect 13924 3670 13952 4082
rect 14108 3670 14136 5170
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13372 2650 13400 3130
rect 13740 3058 13768 3334
rect 13924 3126 13952 3606
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13508 2748 13816 2768
rect 13508 2746 13514 2748
rect 13570 2746 13594 2748
rect 13650 2746 13674 2748
rect 13730 2746 13754 2748
rect 13810 2746 13816 2748
rect 13570 2694 13572 2746
rect 13752 2694 13754 2746
rect 13508 2692 13514 2694
rect 13570 2692 13594 2694
rect 13650 2692 13674 2694
rect 13730 2692 13754 2694
rect 13810 2692 13816 2694
rect 13508 2672 13816 2692
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 11164 734 11468 762
rect 12346 0 12402 800
rect 13634 0 13690 800
rect 14568 762 14596 12922
rect 14752 12374 14780 13806
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14844 12442 14872 13126
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14936 11286 14964 14894
rect 15120 14482 15148 14962
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15120 13410 15148 14282
rect 15212 14278 15240 14894
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15120 13382 15240 13410
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15120 12986 15148 13194
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15212 12866 15240 13382
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15028 12838 15240 12866
rect 15028 12306 15056 12838
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15304 12238 15332 13126
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15396 12238 15424 12582
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 15304 11218 15332 12174
rect 15396 11762 15424 12174
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15488 11558 15516 16390
rect 15580 16114 15608 16662
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15672 13394 15700 18255
rect 15856 18193 15884 18702
rect 15842 18184 15898 18193
rect 15842 18119 15898 18128
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15764 14958 15792 16526
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15856 13394 15884 18119
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16224 16590 16252 16730
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15948 16114 15976 16390
rect 16224 16250 16252 16526
rect 16408 16250 16436 16526
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 16224 16046 16252 16186
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15948 15434 15976 15846
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 16500 13530 16528 24006
rect 16592 23798 16620 24074
rect 16776 23866 16804 24126
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16580 23792 16632 23798
rect 16580 23734 16632 23740
rect 16868 23594 16896 24006
rect 16856 23588 16908 23594
rect 16856 23530 16908 23536
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16684 22710 16712 22918
rect 16672 22704 16724 22710
rect 16672 22646 16724 22652
rect 16672 22500 16724 22506
rect 16672 22442 16724 22448
rect 16684 21690 16712 22442
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16776 21690 16804 22374
rect 17052 22094 17080 28739
rect 17694 27228 18002 27248
rect 17694 27226 17700 27228
rect 17756 27226 17780 27228
rect 17836 27226 17860 27228
rect 17916 27226 17940 27228
rect 17996 27226 18002 27228
rect 17756 27174 17758 27226
rect 17938 27174 17940 27226
rect 17694 27172 17700 27174
rect 17756 27172 17780 27174
rect 17836 27172 17860 27174
rect 17916 27172 17940 27174
rect 17996 27172 18002 27174
rect 17694 27152 18002 27172
rect 17694 26140 18002 26160
rect 17694 26138 17700 26140
rect 17756 26138 17780 26140
rect 17836 26138 17860 26140
rect 17916 26138 17940 26140
rect 17996 26138 18002 26140
rect 17756 26086 17758 26138
rect 17938 26086 17940 26138
rect 17694 26084 17700 26086
rect 17756 26084 17780 26086
rect 17836 26084 17860 26086
rect 17916 26084 17940 26086
rect 17996 26084 18002 26086
rect 17694 26064 18002 26084
rect 17224 25968 17276 25974
rect 17224 25910 17276 25916
rect 17132 22704 17184 22710
rect 17132 22646 17184 22652
rect 17144 22234 17172 22646
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 16960 22066 17080 22094
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16684 19718 16712 19858
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16684 19378 16712 19654
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16776 18358 16804 19722
rect 16856 19712 16908 19718
rect 16854 19680 16856 19689
rect 16908 19680 16910 19689
rect 16854 19615 16910 19624
rect 16868 19514 16896 19615
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 16592 16182 16620 16662
rect 16580 16176 16632 16182
rect 16580 16118 16632 16124
rect 16684 16114 16712 17614
rect 16776 16454 16804 18294
rect 16960 17270 16988 22066
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 17052 18766 17080 19654
rect 17144 18970 17172 21490
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16948 17264 17000 17270
rect 16868 17224 16948 17252
rect 16868 16590 16896 17224
rect 16948 17206 17000 17212
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 17052 16590 17080 16730
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16592 15026 16620 15982
rect 16684 15502 16712 16050
rect 16776 15706 16804 16390
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16868 13394 16896 14010
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16040 12918 16068 13126
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 16408 12306 16436 12922
rect 16592 12322 16620 13194
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16684 12374 16712 12786
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16500 12294 16620 12322
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15948 11762 15976 12038
rect 16408 11898 16436 12242
rect 16500 12102 16528 12294
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15580 11150 15608 11562
rect 15856 11286 15884 11630
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 10674 15240 10950
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15212 10470 15240 10610
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 14740 9988 14792 9994
rect 14740 9930 14792 9936
rect 14752 9518 14780 9930
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14660 8294 14688 8978
rect 14752 8974 14780 9454
rect 15028 9042 15056 9454
rect 15212 9178 15240 10406
rect 15304 10130 15332 10406
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15304 9722 15332 9862
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 15396 8634 15424 11086
rect 15580 10674 15608 11086
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14660 7954 14688 8230
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 15396 7886 15424 8570
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14648 6928 14700 6934
rect 14648 6870 14700 6876
rect 14660 6730 14688 6870
rect 14844 6730 14872 7346
rect 14936 7002 14964 7686
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 15028 7342 15056 7414
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 15028 6458 15056 7278
rect 15120 7002 15148 7482
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15304 6798 15332 7142
rect 15396 6866 15424 7686
rect 15488 7546 15516 10474
rect 15672 10130 15700 10474
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15764 9994 15792 11154
rect 16592 11150 16620 12174
rect 16684 11830 16712 12310
rect 16776 12238 16804 12718
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 16776 11642 16804 12038
rect 16868 11898 16896 12582
rect 16960 12442 16988 13126
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 17052 11762 17080 12106
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16684 11614 16804 11642
rect 16948 11620 17000 11626
rect 16684 11558 16712 11614
rect 16948 11562 17000 11568
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16316 10130 16344 10406
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15752 9988 15804 9994
rect 15752 9930 15804 9936
rect 15764 9654 15792 9930
rect 16040 9654 16068 9998
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15764 9382 15792 9454
rect 16316 9382 16344 10066
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15488 6934 15516 7482
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15580 5370 15608 9318
rect 16316 9178 16344 9318
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16408 8838 16436 10678
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 7954 16160 8230
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16500 7818 16528 10406
rect 16592 9722 16620 10610
rect 16684 10062 16712 11494
rect 16960 11150 16988 11562
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16580 9716 16632 9722
rect 16776 9674 16804 11086
rect 17052 10810 17080 11698
rect 17144 11286 17172 18566
rect 17236 17338 17264 25910
rect 18064 25786 18092 28739
rect 19996 28642 20024 28739
rect 20088 28642 20116 28750
rect 19996 28614 20116 28642
rect 18064 25758 18276 25786
rect 18052 25696 18104 25702
rect 18052 25638 18104 25644
rect 18064 25294 18092 25638
rect 18144 25424 18196 25430
rect 18144 25366 18196 25372
rect 18156 25294 18184 25366
rect 17500 25288 17552 25294
rect 17500 25230 17552 25236
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 18052 25288 18104 25294
rect 18052 25230 18104 25236
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17328 24614 17356 24754
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17420 24274 17448 25094
rect 17512 24818 17540 25230
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17604 24614 17632 25230
rect 17694 25052 18002 25072
rect 17694 25050 17700 25052
rect 17756 25050 17780 25052
rect 17836 25050 17860 25052
rect 17916 25050 17940 25052
rect 17996 25050 18002 25052
rect 17756 24998 17758 25050
rect 17938 24998 17940 25050
rect 17694 24996 17700 24998
rect 17756 24996 17780 24998
rect 17836 24996 17860 24998
rect 17916 24996 17940 24998
rect 17996 24996 18002 24998
rect 17694 24976 18002 24996
rect 17592 24608 17644 24614
rect 17592 24550 17644 24556
rect 17604 24342 17632 24550
rect 17592 24336 17644 24342
rect 17592 24278 17644 24284
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17512 23866 17540 24210
rect 18064 24206 18092 25230
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18156 24954 18184 25094
rect 18144 24948 18196 24954
rect 18144 24890 18196 24896
rect 18052 24200 18104 24206
rect 18052 24142 18104 24148
rect 17694 23964 18002 23984
rect 17694 23962 17700 23964
rect 17756 23962 17780 23964
rect 17836 23962 17860 23964
rect 17916 23962 17940 23964
rect 17996 23962 18002 23964
rect 17756 23910 17758 23962
rect 17938 23910 17940 23962
rect 17694 23908 17700 23910
rect 17756 23908 17780 23910
rect 17836 23908 17860 23910
rect 17916 23908 17940 23910
rect 17996 23908 18002 23910
rect 17694 23888 18002 23908
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17316 22500 17368 22506
rect 17316 22442 17368 22448
rect 17328 22030 17356 22442
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17512 21894 17540 23802
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 17694 22876 18002 22896
rect 17694 22874 17700 22876
rect 17756 22874 17780 22876
rect 17836 22874 17860 22876
rect 17916 22874 17940 22876
rect 17996 22874 18002 22876
rect 17756 22822 17758 22874
rect 17938 22822 17940 22874
rect 17694 22820 17700 22822
rect 17756 22820 17780 22822
rect 17836 22820 17860 22822
rect 17916 22820 17940 22822
rect 17996 22820 18002 22822
rect 17694 22800 18002 22820
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17512 21486 17540 21830
rect 17694 21788 18002 21808
rect 17694 21786 17700 21788
rect 17756 21786 17780 21788
rect 17836 21786 17860 21788
rect 17916 21786 17940 21788
rect 17996 21786 18002 21788
rect 17756 21734 17758 21786
rect 17938 21734 17940 21786
rect 17694 21732 17700 21734
rect 17756 21732 17780 21734
rect 17836 21732 17860 21734
rect 17916 21732 17940 21734
rect 17996 21732 18002 21734
rect 17694 21712 18002 21732
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17512 21146 17540 21422
rect 17500 21140 17552 21146
rect 17500 21082 17552 21088
rect 17694 20700 18002 20720
rect 17694 20698 17700 20700
rect 17756 20698 17780 20700
rect 17836 20698 17860 20700
rect 17916 20698 17940 20700
rect 17996 20698 18002 20700
rect 17756 20646 17758 20698
rect 17938 20646 17940 20698
rect 17694 20644 17700 20646
rect 17756 20644 17780 20646
rect 17836 20644 17860 20646
rect 17916 20644 17940 20646
rect 17996 20644 18002 20646
rect 17694 20624 18002 20644
rect 17316 20324 17368 20330
rect 17316 20266 17368 20272
rect 17328 18766 17356 20266
rect 18064 19718 18092 22986
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17420 18630 17448 19654
rect 17694 19612 18002 19632
rect 17694 19610 17700 19612
rect 17756 19610 17780 19612
rect 17836 19610 17860 19612
rect 17916 19610 17940 19612
rect 17996 19610 18002 19612
rect 17756 19558 17758 19610
rect 17938 19558 17940 19610
rect 17694 19556 17700 19558
rect 17756 19556 17780 19558
rect 17836 19556 17860 19558
rect 17916 19556 17940 19558
rect 17996 19556 18002 19558
rect 17694 19536 18002 19556
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17972 19122 18000 19382
rect 17880 19094 18000 19122
rect 17880 18970 17908 19094
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17592 18760 17644 18766
rect 17960 18760 18012 18766
rect 17592 18702 17644 18708
rect 17958 18728 17960 18737
rect 18012 18728 18014 18737
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17512 18426 17540 18566
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 17420 17066 17448 17750
rect 17512 17134 17540 18226
rect 17604 17882 17632 18702
rect 17958 18663 18014 18672
rect 17694 18524 18002 18544
rect 17694 18522 17700 18524
rect 17756 18522 17780 18524
rect 17836 18522 17860 18524
rect 17916 18522 17940 18524
rect 17996 18522 18002 18524
rect 17756 18470 17758 18522
rect 17938 18470 17940 18522
rect 17694 18468 17700 18470
rect 17756 18468 17780 18470
rect 17836 18468 17860 18470
rect 17916 18468 17940 18470
rect 17996 18468 18002 18470
rect 17694 18448 18002 18468
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17880 17882 17908 18158
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17694 17436 18002 17456
rect 17694 17434 17700 17436
rect 17756 17434 17780 17436
rect 17836 17434 17860 17436
rect 17916 17434 17940 17436
rect 17996 17434 18002 17436
rect 17756 17382 17758 17434
rect 17938 17382 17940 17434
rect 17694 17380 17700 17382
rect 17756 17380 17780 17382
rect 17836 17380 17860 17382
rect 17916 17380 17940 17382
rect 17996 17380 18002 17382
rect 17694 17360 18002 17380
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17236 16590 17264 16934
rect 17604 16590 17632 17274
rect 17958 17232 18014 17241
rect 17776 17196 17828 17202
rect 17958 17167 18014 17176
rect 17776 17138 17828 17144
rect 17788 16998 17816 17138
rect 17972 17134 18000 17167
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17236 15502 17264 16390
rect 17512 15706 17540 16526
rect 17694 16348 18002 16368
rect 17694 16346 17700 16348
rect 17756 16346 17780 16348
rect 17836 16346 17860 16348
rect 17916 16346 17940 16348
rect 17996 16346 18002 16348
rect 17756 16294 17758 16346
rect 17938 16294 17940 16346
rect 17694 16292 17700 16294
rect 17756 16292 17780 16294
rect 17836 16292 17860 16294
rect 17916 16292 17940 16294
rect 17996 16292 18002 16294
rect 17694 16272 18002 16292
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17236 13326 17264 13738
rect 17224 13320 17276 13326
rect 17222 13288 17224 13297
rect 17276 13288 17278 13297
rect 17222 13223 17278 13232
rect 17328 13138 17356 15642
rect 17694 15260 18002 15280
rect 17694 15258 17700 15260
rect 17756 15258 17780 15260
rect 17836 15258 17860 15260
rect 17916 15258 17940 15260
rect 17996 15258 18002 15260
rect 17756 15206 17758 15258
rect 17938 15206 17940 15258
rect 17694 15204 17700 15206
rect 17756 15204 17780 15206
rect 17836 15204 17860 15206
rect 17916 15204 17940 15206
rect 17996 15204 18002 15206
rect 17694 15184 18002 15204
rect 18064 15094 18092 19654
rect 18248 19514 18276 25758
rect 19340 25356 19392 25362
rect 19340 25298 19392 25304
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 18616 24886 18644 25230
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 18524 24138 18552 24686
rect 18616 24206 18644 24822
rect 19248 24676 19300 24682
rect 19248 24618 19300 24624
rect 18880 24336 18932 24342
rect 18880 24278 18932 24284
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18604 24200 18656 24206
rect 18604 24142 18656 24148
rect 18512 24132 18564 24138
rect 18512 24074 18564 24080
rect 18328 23724 18380 23730
rect 18328 23666 18380 23672
rect 18340 22982 18368 23666
rect 18524 23594 18552 24074
rect 18512 23588 18564 23594
rect 18512 23530 18564 23536
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18328 22432 18380 22438
rect 18328 22374 18380 22380
rect 18340 21962 18368 22374
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18524 21690 18552 22578
rect 18512 21684 18564 21690
rect 18512 21626 18564 21632
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18156 18698 18184 18770
rect 18144 18692 18196 18698
rect 18144 18634 18196 18640
rect 18156 18222 18184 18634
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18156 17882 18184 18158
rect 18248 18154 18276 19314
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 18156 17202 18184 17818
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18340 16454 18368 21490
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18432 17882 18460 19654
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18524 18766 18552 18906
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18524 18426 18552 18702
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 18524 18136 18552 18362
rect 18616 18358 18644 19450
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18604 18148 18656 18154
rect 18524 18108 18604 18136
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 18432 17678 18460 17818
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18524 17524 18552 18108
rect 18604 18090 18656 18096
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18432 17496 18552 17524
rect 18432 17241 18460 17496
rect 18616 17338 18644 17546
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18418 17232 18474 17241
rect 18418 17167 18474 17176
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18524 16726 18552 17138
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18432 16250 18460 16390
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17420 13394 17448 14758
rect 17512 14618 17540 14894
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17512 13818 17540 14554
rect 18156 14414 18184 15846
rect 18248 15570 18276 16186
rect 18524 16130 18552 16662
rect 18432 16102 18552 16130
rect 18604 16108 18656 16114
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 18340 15026 18368 15370
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 17694 14172 18002 14192
rect 17694 14170 17700 14172
rect 17756 14170 17780 14172
rect 17836 14170 17860 14172
rect 17916 14170 17940 14172
rect 17996 14170 18002 14172
rect 17756 14118 17758 14170
rect 17938 14118 17940 14170
rect 17694 14116 17700 14118
rect 17756 14116 17780 14118
rect 17836 14116 17860 14118
rect 17916 14116 17940 14118
rect 17996 14116 18002 14118
rect 17694 14096 18002 14116
rect 18156 14074 18184 14350
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 17512 13790 17632 13818
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17512 13530 17540 13670
rect 17604 13530 17632 13790
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17236 13110 17356 13138
rect 17236 12238 17264 13110
rect 17604 13002 17632 13330
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17694 13084 18002 13104
rect 17694 13082 17700 13084
rect 17756 13082 17780 13084
rect 17836 13082 17860 13084
rect 17916 13082 17940 13084
rect 17996 13082 18002 13084
rect 17756 13030 17758 13082
rect 17938 13030 17940 13082
rect 17694 13028 17700 13030
rect 17756 13028 17780 13030
rect 17836 13028 17860 13030
rect 17916 13028 17940 13030
rect 17996 13028 18002 13030
rect 17694 13008 18002 13028
rect 17512 12986 17632 13002
rect 18064 12986 18092 13126
rect 17500 12980 17632 12986
rect 17328 12940 17500 12968
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17236 11762 17264 12174
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17328 11626 17356 12940
rect 17552 12974 17632 12980
rect 18052 12980 18104 12986
rect 17500 12922 17552 12928
rect 18052 12922 18104 12928
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 12434 17540 12718
rect 17420 12406 17540 12434
rect 17316 11620 17368 11626
rect 17316 11562 17368 11568
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 17052 10266 17080 10610
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17144 10130 17172 11018
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16580 9658 16632 9664
rect 16684 9646 16804 9674
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 15948 6866 15976 7686
rect 16224 7206 16252 7686
rect 16408 7478 16436 7686
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15948 6390 15976 6802
rect 15936 6384 15988 6390
rect 15936 6326 15988 6332
rect 16684 6186 16712 9646
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 7886 16896 9318
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 16776 6798 16804 6870
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 15028 4826 15056 4966
rect 15488 4826 15516 5034
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 16224 4758 16252 5102
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 16212 4752 16264 4758
rect 16212 4694 16264 4700
rect 14832 4548 14884 4554
rect 14832 4490 14884 4496
rect 14844 4282 14872 4490
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14660 3534 14688 3674
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14660 3194 14688 3470
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14752 3058 14780 3470
rect 14936 3466 14964 4694
rect 15108 4616 15160 4622
rect 15028 4576 15108 4604
rect 15028 3942 15056 4576
rect 15108 4558 15160 4564
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15304 4146 15332 4490
rect 15396 4214 15424 4558
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 15028 3534 15056 3878
rect 15396 3738 15424 4150
rect 16224 4078 16252 4694
rect 16408 4690 16436 4966
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16500 4214 16528 5034
rect 16960 4622 16988 9862
rect 17328 9586 17356 11562
rect 17420 11558 17448 12406
rect 17512 12374 17540 12406
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17512 11830 17540 12174
rect 17604 11898 17632 12854
rect 18052 12844 18104 12850
rect 18156 12832 18184 14010
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18248 12850 18276 13194
rect 18104 12804 18184 12832
rect 18236 12844 18288 12850
rect 18052 12786 18104 12792
rect 18236 12786 18288 12792
rect 17684 12368 17736 12374
rect 17684 12310 17736 12316
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 17696 12238 17724 12310
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 18248 12102 18276 12310
rect 18340 12306 18368 14962
rect 18432 13988 18460 16102
rect 18604 16050 18656 16056
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18524 15026 18552 15642
rect 18616 15366 18644 16050
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18512 14000 18564 14006
rect 18432 13960 18512 13988
rect 18512 13942 18564 13948
rect 18524 13394 18552 13942
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 17694 11996 18002 12016
rect 17694 11994 17700 11996
rect 17756 11994 17780 11996
rect 17836 11994 17860 11996
rect 17916 11994 17940 11996
rect 17996 11994 18002 11996
rect 17756 11942 17758 11994
rect 17938 11942 17940 11994
rect 17694 11940 17700 11942
rect 17756 11940 17780 11942
rect 17836 11940 17860 11942
rect 17916 11940 17940 11942
rect 17996 11940 18002 11942
rect 17694 11920 18002 11940
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 18064 11762 18092 12038
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17604 11354 17632 11698
rect 18340 11694 18368 12242
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17420 10062 17448 11222
rect 17694 10908 18002 10928
rect 17694 10906 17700 10908
rect 17756 10906 17780 10908
rect 17836 10906 17860 10908
rect 17916 10906 17940 10908
rect 17996 10906 18002 10908
rect 17756 10854 17758 10906
rect 17938 10854 17940 10906
rect 17694 10852 17700 10854
rect 17756 10852 17780 10854
rect 17836 10852 17860 10854
rect 17916 10852 17940 10854
rect 17996 10852 18002 10854
rect 17694 10832 18002 10852
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17604 10198 17632 10678
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17408 10056 17460 10062
rect 17592 10056 17644 10062
rect 17408 9998 17460 10004
rect 17512 10016 17592 10044
rect 17420 9722 17448 9998
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17512 9654 17540 10016
rect 17592 9998 17644 10004
rect 17696 9994 17724 10610
rect 17788 10130 17816 10610
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17880 10062 17908 10406
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17328 8974 17356 9522
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17420 9178 17448 9454
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17420 8634 17448 9114
rect 17604 8906 17632 9862
rect 17694 9820 18002 9840
rect 17694 9818 17700 9820
rect 17756 9818 17780 9820
rect 17836 9818 17860 9820
rect 17916 9818 17940 9820
rect 17996 9818 18002 9820
rect 17756 9766 17758 9818
rect 17938 9766 17940 9818
rect 17694 9764 17700 9766
rect 17756 9764 17780 9766
rect 17836 9764 17860 9766
rect 17916 9764 17940 9766
rect 17996 9764 18002 9766
rect 17694 9744 18002 9764
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18248 9518 18276 9658
rect 18616 9654 18644 15302
rect 18708 13530 18736 24210
rect 18892 23798 18920 24278
rect 18880 23792 18932 23798
rect 18880 23734 18932 23740
rect 19260 23594 19288 24618
rect 19352 24342 19380 25298
rect 19708 25220 19760 25226
rect 19708 25162 19760 25168
rect 19720 24954 19748 25162
rect 19708 24948 19760 24954
rect 19708 24890 19760 24896
rect 19708 24608 19760 24614
rect 19708 24550 19760 24556
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 19352 23866 19380 24278
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19248 23588 19300 23594
rect 19248 23530 19300 23536
rect 19156 22704 19208 22710
rect 19156 22646 19208 22652
rect 19064 21956 19116 21962
rect 19064 21898 19116 21904
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18892 21078 18920 21422
rect 19076 21078 19104 21898
rect 19168 21554 19196 22646
rect 19352 22094 19380 23802
rect 19444 23526 19472 24346
rect 19720 23866 19748 24550
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19708 23656 19760 23662
rect 19708 23598 19760 23604
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19720 23118 19748 23598
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19260 22066 19380 22094
rect 19260 22030 19288 22066
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 19260 21486 19288 21830
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19352 21350 19380 21830
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19444 21457 19472 21490
rect 19430 21448 19486 21457
rect 19430 21383 19486 21392
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 18880 21072 18932 21078
rect 18880 21014 18932 21020
rect 19064 21072 19116 21078
rect 19064 21014 19116 21020
rect 18892 20602 18920 21014
rect 19628 21010 19656 21286
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18786 18320 18842 18329
rect 18786 18255 18788 18264
rect 18840 18255 18842 18264
rect 18788 18226 18840 18232
rect 18786 18184 18842 18193
rect 18786 18119 18788 18128
rect 18840 18119 18842 18128
rect 18788 18090 18840 18096
rect 18892 17134 18920 18838
rect 18984 18766 19012 19246
rect 19352 18884 19380 19450
rect 19260 18856 19380 18884
rect 18972 18760 19024 18766
rect 19260 18737 19288 18856
rect 18972 18702 19024 18708
rect 19246 18728 19302 18737
rect 19246 18663 19302 18672
rect 19628 18426 19656 20742
rect 19720 20534 19748 21490
rect 19708 20528 19760 20534
rect 19708 20470 19760 20476
rect 19892 18692 19944 18698
rect 19892 18634 19944 18640
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19904 18290 19932 18634
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 19260 17882 19288 18226
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18800 16114 18828 16390
rect 18892 16250 18920 16934
rect 19076 16726 19104 17614
rect 19064 16720 19116 16726
rect 19064 16662 19116 16668
rect 19154 16688 19210 16697
rect 19154 16623 19210 16632
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 18800 15026 18828 15914
rect 18892 15706 18920 16186
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18892 15502 18920 15642
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18984 15178 19012 15438
rect 19076 15434 19104 16118
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 18892 15162 19012 15178
rect 18880 15156 19012 15162
rect 18932 15150 19012 15156
rect 18880 15098 18932 15104
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 19076 14958 19104 15370
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19168 14822 19196 16623
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19904 16114 19932 16526
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19352 15162 19380 16050
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19352 14550 19380 15098
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19996 14074 20024 23666
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 20088 21486 20116 21830
rect 20076 21480 20128 21486
rect 20168 21480 20220 21486
rect 20076 21422 20128 21428
rect 20166 21448 20168 21457
rect 20220 21448 20222 21457
rect 20088 20602 20116 21422
rect 20222 21406 20300 21434
rect 20166 21383 20222 21392
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 20180 19922 20208 20810
rect 20272 20466 20300 21406
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20364 19514 20392 28750
rect 20994 28739 21050 29539
rect 21652 28750 21956 28778
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20732 24886 20760 25094
rect 20720 24880 20772 24886
rect 20720 24822 20772 24828
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 21088 24336 21140 24342
rect 21088 24278 21140 24284
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 20548 23866 20576 24006
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 21100 23798 21128 24278
rect 21192 24274 21220 24754
rect 21180 24268 21232 24274
rect 21180 24210 21232 24216
rect 21192 23866 21220 24210
rect 21180 23860 21232 23866
rect 21180 23802 21232 23808
rect 21088 23792 21140 23798
rect 21088 23734 21140 23740
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20548 23118 20576 23598
rect 20628 23248 20680 23254
rect 20628 23190 20680 23196
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 20536 21004 20588 21010
rect 20536 20946 20588 20952
rect 20548 20602 20576 20946
rect 20640 20874 20668 23190
rect 20628 20868 20680 20874
rect 20628 20810 20680 20816
rect 20536 20596 20588 20602
rect 20536 20538 20588 20544
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20732 18766 20760 18838
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20352 18284 20404 18290
rect 20404 18244 20484 18272
rect 20352 18226 20404 18232
rect 20180 17882 20208 18226
rect 20456 18204 20484 18244
rect 20456 18176 20576 18204
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20272 17134 20300 17818
rect 20548 17542 20576 18176
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20536 17536 20588 17542
rect 20628 17536 20680 17542
rect 20536 17478 20588 17484
rect 20626 17504 20628 17513
rect 20680 17504 20682 17513
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 20272 16250 20300 17070
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 20076 15972 20128 15978
rect 20076 15914 20128 15920
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 19260 13394 19288 14010
rect 19628 13530 19656 14010
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19524 13456 19576 13462
rect 19524 13398 19576 13404
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19536 12374 19564 13398
rect 19904 13258 19932 13806
rect 19892 13252 19944 13258
rect 19892 13194 19944 13200
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19708 12708 19760 12714
rect 19708 12650 19760 12656
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19720 12238 19748 12650
rect 19812 12646 19840 13126
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19904 12102 19932 13194
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 19996 12238 20024 12786
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19904 11150 19932 12038
rect 19996 11898 20024 12174
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 18800 10266 18828 10610
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18984 9722 19012 10406
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18156 9178 18184 9454
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18616 8974 18644 9590
rect 19076 9586 19104 9998
rect 19444 9722 19472 10610
rect 19628 10606 19656 11086
rect 19904 10810 19932 11086
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19628 10266 19656 10542
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19628 10062 19656 10202
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19628 8974 19656 9318
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 17694 8732 18002 8752
rect 17694 8730 17700 8732
rect 17756 8730 17780 8732
rect 17836 8730 17860 8732
rect 17916 8730 17940 8732
rect 17996 8730 18002 8732
rect 17756 8678 17758 8730
rect 17938 8678 17940 8730
rect 17694 8676 17700 8678
rect 17756 8676 17780 8678
rect 17836 8676 17860 8678
rect 17916 8676 17940 8678
rect 17996 8676 18002 8678
rect 17694 8656 18002 8676
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17052 6798 17080 7142
rect 17236 6934 17264 7822
rect 17604 7206 17632 7822
rect 17694 7644 18002 7664
rect 17694 7642 17700 7644
rect 17756 7642 17780 7644
rect 17836 7642 17860 7644
rect 17916 7642 17940 7644
rect 17996 7642 18002 7644
rect 17756 7590 17758 7642
rect 17938 7590 17940 7642
rect 17694 7588 17700 7590
rect 17756 7588 17780 7590
rect 17836 7588 17860 7590
rect 17916 7588 17940 7590
rect 17996 7588 18002 7590
rect 17694 7568 18002 7588
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17144 6254 17172 6734
rect 17328 6662 17356 6938
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17328 6322 17356 6598
rect 17694 6556 18002 6576
rect 17694 6554 17700 6556
rect 17756 6554 17780 6556
rect 17836 6554 17860 6556
rect 17916 6554 17940 6556
rect 17996 6554 18002 6556
rect 17756 6502 17758 6554
rect 17938 6502 17940 6554
rect 17694 6500 17700 6502
rect 17756 6500 17780 6502
rect 17836 6500 17860 6502
rect 17916 6500 17940 6502
rect 17996 6500 18002 6502
rect 17694 6480 18002 6500
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17694 5468 18002 5488
rect 17694 5466 17700 5468
rect 17756 5466 17780 5468
rect 17836 5466 17860 5468
rect 17916 5466 17940 5468
rect 17996 5466 18002 5468
rect 17756 5414 17758 5466
rect 17938 5414 17940 5466
rect 17694 5412 17700 5414
rect 17756 5412 17780 5414
rect 17836 5412 17860 5414
rect 17916 5412 17940 5414
rect 17996 5412 18002 5414
rect 17694 5392 18002 5412
rect 18064 5370 18092 8774
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18248 7546 18276 8026
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18340 6322 18368 7822
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 6730 18460 7686
rect 19260 7546 19288 8774
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19444 7546 19472 7754
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 18524 6390 18552 7278
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18788 5568 18840 5574
rect 18788 5510 18840 5516
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 17236 4554 17264 5102
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 17512 4826 17540 4966
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 18432 4554 18460 4966
rect 18800 4554 18828 5510
rect 18892 5370 18920 7278
rect 19444 7002 19472 7482
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19260 5710 19288 6734
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 19248 5704 19300 5710
rect 19248 5646 19300 5652
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 19076 4826 19104 4966
rect 19064 4820 19116 4826
rect 19064 4762 19116 4768
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 18420 4548 18472 4554
rect 18420 4490 18472 4496
rect 18788 4548 18840 4554
rect 18788 4490 18840 4496
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16302 4040 16358 4049
rect 16302 3975 16358 3984
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15672 3534 15700 3878
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 14924 3460 14976 3466
rect 14924 3402 14976 3408
rect 14936 3126 14964 3402
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14936 870 15056 898
rect 14936 762 14964 870
rect 15028 800 15056 870
rect 16316 800 16344 3975
rect 16592 3942 16620 4422
rect 16960 3942 16988 4422
rect 17144 4282 17172 4422
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16684 3058 16712 3878
rect 17052 3738 17080 4014
rect 17236 3942 17264 4490
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 17694 4380 18002 4400
rect 17694 4378 17700 4380
rect 17756 4378 17780 4380
rect 17836 4378 17860 4380
rect 17916 4378 17940 4380
rect 17996 4378 18002 4380
rect 17756 4326 17758 4378
rect 17938 4326 17940 4378
rect 17694 4324 17700 4326
rect 17756 4324 17780 4326
rect 17836 4324 17860 4326
rect 17916 4324 17940 4326
rect 17996 4324 18002 4326
rect 17694 4304 18002 4324
rect 18064 4214 18092 4422
rect 18432 4214 18460 4490
rect 18800 4282 18828 4490
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18878 4040 18934 4049
rect 18878 3975 18934 3984
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17236 3670 17264 3878
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16868 3194 16896 3402
rect 17694 3292 18002 3312
rect 17694 3290 17700 3292
rect 17756 3290 17780 3292
rect 17836 3290 17860 3292
rect 17916 3290 17940 3292
rect 17996 3290 18002 3292
rect 17756 3238 17758 3290
rect 17938 3238 17940 3290
rect 17694 3236 17700 3238
rect 17756 3236 17780 3238
rect 17836 3236 17860 3238
rect 17916 3236 17940 3238
rect 17996 3236 18002 3238
rect 17694 3216 18002 3236
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 17694 2204 18002 2224
rect 17694 2202 17700 2204
rect 17756 2202 17780 2204
rect 17836 2202 17860 2204
rect 17916 2202 17940 2204
rect 17996 2202 18002 2204
rect 17756 2150 17758 2202
rect 17938 2150 17940 2202
rect 17694 2148 17700 2150
rect 17756 2148 17780 2150
rect 17836 2148 17860 2150
rect 17916 2148 17940 2150
rect 17996 2148 18002 2150
rect 17694 2128 18002 2148
rect 18892 800 18920 3975
rect 19352 3942 19380 6666
rect 19536 6322 19564 7142
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19628 6458 19656 6666
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19628 5250 19656 6258
rect 19812 5370 19840 10406
rect 19904 10062 19932 10746
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19996 10130 20024 10406
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 20088 9654 20116 15914
rect 20364 15706 20392 15982
rect 20548 15978 20576 17478
rect 20626 17439 20682 17448
rect 20732 17338 20760 17546
rect 20720 17332 20772 17338
rect 20640 17292 20720 17320
rect 20640 16590 20668 17292
rect 20720 17274 20772 17280
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20640 16266 20668 16526
rect 20732 16522 20760 17138
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20640 16238 20760 16266
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20548 15502 20576 15642
rect 20640 15570 20668 16050
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20732 15502 20760 16238
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20180 13870 20208 14214
rect 20824 14074 20852 23666
rect 21284 22094 21312 25978
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 21468 22710 21496 23122
rect 21456 22704 21508 22710
rect 21456 22646 21508 22652
rect 21192 22066 21312 22094
rect 20904 21072 20956 21078
rect 20904 21014 20956 21020
rect 20916 20602 20944 21014
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 21192 18970 21220 22066
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21272 21480 21324 21486
rect 21270 21448 21272 21457
rect 21324 21448 21326 21457
rect 21270 21383 21326 21392
rect 21376 20806 21404 21490
rect 21456 21412 21508 21418
rect 21456 21354 21508 21360
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21468 20602 21496 21354
rect 21652 21350 21680 28750
rect 21928 28642 21956 28750
rect 22006 28739 22062 29539
rect 22926 28739 22982 29539
rect 23938 28739 23994 29539
rect 24950 28739 25006 29539
rect 25870 28739 25926 29539
rect 26330 28792 26386 28801
rect 22020 28642 22048 28739
rect 21928 28614 22048 28642
rect 21880 26684 22188 26704
rect 21880 26682 21886 26684
rect 21942 26682 21966 26684
rect 22022 26682 22046 26684
rect 22102 26682 22126 26684
rect 22182 26682 22188 26684
rect 21942 26630 21944 26682
rect 22124 26630 22126 26682
rect 21880 26628 21886 26630
rect 21942 26628 21966 26630
rect 22022 26628 22046 26630
rect 22102 26628 22126 26630
rect 22182 26628 22188 26630
rect 21880 26608 22188 26628
rect 23952 25906 23980 28739
rect 24964 25906 24992 28739
rect 26882 28739 26938 29539
rect 26330 28727 26332 28736
rect 26384 28727 26386 28736
rect 26332 28698 26384 28704
rect 23940 25900 23992 25906
rect 23940 25842 23992 25848
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 26896 25838 26924 28739
rect 26884 25832 26936 25838
rect 26884 25774 26936 25780
rect 21880 25596 22188 25616
rect 21880 25594 21886 25596
rect 21942 25594 21966 25596
rect 22022 25594 22046 25596
rect 22102 25594 22126 25596
rect 22182 25594 22188 25596
rect 21942 25542 21944 25594
rect 22124 25542 22126 25594
rect 21880 25540 21886 25542
rect 21942 25540 21966 25542
rect 22022 25540 22046 25542
rect 22102 25540 22126 25542
rect 22182 25540 22188 25542
rect 21880 25520 22188 25540
rect 26330 24576 26386 24585
rect 21880 24508 22188 24528
rect 26330 24511 26332 24520
rect 21880 24506 21886 24508
rect 21942 24506 21966 24508
rect 22022 24506 22046 24508
rect 22102 24506 22126 24508
rect 22182 24506 22188 24508
rect 21942 24454 21944 24506
rect 22124 24454 22126 24506
rect 26384 24511 26386 24520
rect 26332 24482 26384 24488
rect 21880 24452 21886 24454
rect 21942 24452 21966 24454
rect 22022 24452 22046 24454
rect 22102 24452 22126 24454
rect 22182 24452 22188 24454
rect 21880 24432 22188 24452
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 21928 23798 21956 24142
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22560 24132 22612 24138
rect 22560 24074 22612 24080
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21744 23322 21772 23666
rect 22112 23662 22140 24074
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 21880 23420 22188 23440
rect 21880 23418 21886 23420
rect 21942 23418 21966 23420
rect 22022 23418 22046 23420
rect 22102 23418 22126 23420
rect 22182 23418 22188 23420
rect 21942 23366 21944 23418
rect 22124 23366 22126 23418
rect 21880 23364 21886 23366
rect 21942 23364 21966 23366
rect 22022 23364 22046 23366
rect 22102 23364 22126 23366
rect 22182 23364 22188 23366
rect 21880 23344 22188 23364
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 22572 23186 22600 24074
rect 23216 23866 23244 24142
rect 24032 24132 24084 24138
rect 24032 24074 24084 24080
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 24044 23798 24072 24074
rect 24032 23792 24084 23798
rect 24032 23734 24084 23740
rect 22744 23520 22796 23526
rect 22744 23462 22796 23468
rect 22560 23180 22612 23186
rect 22560 23122 22612 23128
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22284 22500 22336 22506
rect 22284 22442 22336 22448
rect 21880 22332 22188 22352
rect 21880 22330 21886 22332
rect 21942 22330 21966 22332
rect 22022 22330 22046 22332
rect 22102 22330 22126 22332
rect 22182 22330 22188 22332
rect 21942 22278 21944 22330
rect 22124 22278 22126 22330
rect 21880 22276 21886 22278
rect 21942 22276 21966 22278
rect 22022 22276 22046 22278
rect 22102 22276 22126 22278
rect 22182 22276 22188 22278
rect 21880 22256 22188 22276
rect 22296 22234 22324 22442
rect 22284 22228 22336 22234
rect 22284 22170 22336 22176
rect 22480 22137 22508 22918
rect 22756 22642 22784 23462
rect 24044 23186 24072 23734
rect 25134 23216 25190 23225
rect 24032 23180 24084 23186
rect 25134 23151 25136 23160
rect 24032 23122 24084 23128
rect 25188 23151 25190 23160
rect 25136 23122 25188 23128
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 23020 23044 23072 23050
rect 23020 22986 23072 22992
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 22744 22636 22796 22642
rect 22744 22578 22796 22584
rect 22466 22128 22522 22137
rect 22466 22063 22522 22072
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 22652 21888 22704 21894
rect 22282 21856 22338 21865
rect 22652 21830 22704 21836
rect 22282 21791 22338 21800
rect 22296 21622 22324 21791
rect 21824 21616 21876 21622
rect 21744 21576 21824 21604
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 21008 18222 21036 18362
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 20916 18068 20944 18158
rect 20916 18040 21036 18068
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20916 16794 20944 17682
rect 21008 17270 21036 18040
rect 21100 17678 21128 18226
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 21192 17542 21220 18906
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21192 17338 21220 17478
rect 21284 17338 21312 20402
rect 21652 18902 21680 20878
rect 21744 20874 21772 21576
rect 21824 21558 21876 21564
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 21880 21244 22188 21264
rect 21880 21242 21886 21244
rect 21942 21242 21966 21244
rect 22022 21242 22046 21244
rect 22102 21242 22126 21244
rect 22182 21242 22188 21244
rect 21942 21190 21944 21242
rect 22124 21190 22126 21242
rect 21880 21188 21886 21190
rect 21942 21188 21966 21190
rect 22022 21188 22046 21190
rect 22102 21188 22126 21190
rect 22182 21188 22188 21190
rect 21880 21168 22188 21188
rect 21732 20868 21784 20874
rect 21732 20810 21784 20816
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 21880 20156 22188 20176
rect 21880 20154 21886 20156
rect 21942 20154 21966 20156
rect 22022 20154 22046 20156
rect 22102 20154 22126 20156
rect 22182 20154 22188 20156
rect 21942 20102 21944 20154
rect 22124 20102 22126 20154
rect 21880 20100 21886 20102
rect 21942 20100 21966 20102
rect 22022 20100 22046 20102
rect 22102 20100 22126 20102
rect 22182 20100 22188 20102
rect 21880 20080 22188 20100
rect 22296 19990 22324 20198
rect 22388 20058 22416 20402
rect 22376 20052 22428 20058
rect 22376 19994 22428 20000
rect 22284 19984 22336 19990
rect 22284 19926 22336 19932
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22388 19514 22416 19858
rect 22572 19802 22600 21490
rect 22480 19774 22600 19802
rect 22480 19718 22508 19774
rect 22468 19712 22520 19718
rect 22468 19654 22520 19660
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22572 19514 22600 19654
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 22388 19174 22416 19450
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 21880 19068 22188 19088
rect 21880 19066 21886 19068
rect 21942 19066 21966 19068
rect 22022 19066 22046 19068
rect 22102 19066 22126 19068
rect 22182 19066 22188 19068
rect 21942 19014 21944 19066
rect 22124 19014 22126 19066
rect 21880 19012 21886 19014
rect 21942 19012 21966 19014
rect 22022 19012 22046 19014
rect 22102 19012 22126 19014
rect 22182 19012 22188 19014
rect 21880 18992 22188 19012
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21652 18766 21680 18838
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21376 17678 21404 18362
rect 21638 18320 21694 18329
rect 21638 18255 21694 18264
rect 21652 17746 21680 18255
rect 21744 18154 21772 18906
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22190 18184 22246 18193
rect 21732 18148 21784 18154
rect 22190 18119 22192 18128
rect 21732 18090 21784 18096
rect 22244 18119 22246 18128
rect 22192 18090 22244 18096
rect 21880 17980 22188 18000
rect 21880 17978 21886 17980
rect 21942 17978 21966 17980
rect 22022 17978 22046 17980
rect 22102 17978 22126 17980
rect 22182 17978 22188 17980
rect 21942 17926 21944 17978
rect 22124 17926 22126 17978
rect 21880 17924 21886 17926
rect 21942 17924 21966 17926
rect 22022 17924 22046 17926
rect 22102 17924 22126 17926
rect 22182 17924 22188 17926
rect 21880 17904 22188 17924
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 22296 17678 22324 18226
rect 22388 17882 22416 18634
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 21008 17066 21036 17206
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 21376 16590 21404 17614
rect 21928 17542 21956 17614
rect 22388 17542 22416 17682
rect 21916 17536 21968 17542
rect 21454 17504 21510 17513
rect 22284 17536 22336 17542
rect 21916 17478 21968 17484
rect 22282 17504 22284 17513
rect 22376 17536 22428 17542
rect 22336 17504 22338 17513
rect 21454 17439 21510 17448
rect 22376 17478 22428 17484
rect 22282 17439 22338 17448
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 15910 21312 16390
rect 21468 16046 21496 17439
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 21548 17128 21600 17134
rect 21548 17070 21600 17076
rect 21560 16454 21588 17070
rect 21880 16892 22188 16912
rect 21880 16890 21886 16892
rect 21942 16890 21966 16892
rect 22022 16890 22046 16892
rect 22102 16890 22126 16892
rect 22182 16890 22188 16892
rect 21942 16838 21944 16890
rect 22124 16838 22126 16890
rect 21880 16836 21886 16838
rect 21942 16836 21966 16838
rect 22022 16836 22046 16838
rect 22102 16836 22126 16838
rect 22182 16836 22188 16838
rect 21880 16816 22188 16836
rect 22296 16454 22324 17206
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22388 16794 22416 17070
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21100 15570 21128 15846
rect 21468 15706 21496 15982
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20180 12374 20208 13806
rect 20364 13326 20392 13806
rect 20456 13530 20484 13874
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20364 12442 20392 12718
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20168 12368 20220 12374
rect 20168 12310 20220 12316
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20364 11762 20392 12038
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20364 11150 20392 11698
rect 20640 11558 20668 13262
rect 20824 12850 20852 13874
rect 20916 13734 20944 14962
rect 21100 14414 21128 15506
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21284 15094 21312 15370
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21272 15088 21324 15094
rect 21272 15030 21324 15036
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21284 14618 21312 14894
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 20916 13326 20944 13670
rect 21008 13530 21036 13670
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21272 13456 21324 13462
rect 21272 13398 21324 13404
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 21284 12986 21312 13398
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 20824 11762 20852 12786
rect 21008 12306 21036 12786
rect 21284 12442 21312 12922
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20536 11008 20588 11014
rect 20536 10950 20588 10956
rect 20548 10810 20576 10950
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20640 10674 20668 11494
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 21192 10810 21220 11222
rect 21376 11150 21404 15302
rect 21468 13302 21496 15370
rect 21456 13296 21508 13302
rect 21456 13238 21508 13244
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21468 12374 21496 12718
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21560 11354 21588 16390
rect 22282 16144 22338 16153
rect 21732 16108 21784 16114
rect 22282 16079 22338 16088
rect 22376 16108 22428 16114
rect 21732 16050 21784 16056
rect 21744 15026 21772 16050
rect 21880 15804 22188 15824
rect 21880 15802 21886 15804
rect 21942 15802 21966 15804
rect 22022 15802 22046 15804
rect 22102 15802 22126 15804
rect 22182 15802 22188 15804
rect 21942 15750 21944 15802
rect 22124 15750 22126 15802
rect 21880 15748 21886 15750
rect 21942 15748 21966 15750
rect 22022 15748 22046 15750
rect 22102 15748 22126 15750
rect 22182 15748 22188 15750
rect 21880 15728 22188 15748
rect 22296 15638 22324 16079
rect 22376 16050 22428 16056
rect 22388 15706 22416 16050
rect 22376 15700 22428 15706
rect 22376 15642 22428 15648
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21836 14906 21864 15438
rect 21744 14878 21864 14906
rect 21744 14618 21772 14878
rect 21880 14716 22188 14736
rect 21880 14714 21886 14716
rect 21942 14714 21966 14716
rect 22022 14714 22046 14716
rect 22102 14714 22126 14716
rect 22182 14714 22188 14716
rect 21942 14662 21944 14714
rect 22124 14662 22126 14714
rect 21880 14660 21886 14662
rect 21942 14660 21966 14662
rect 22022 14660 22046 14662
rect 22102 14660 22126 14662
rect 22182 14660 22188 14662
rect 21880 14640 22188 14660
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 21652 13462 21680 13670
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 21744 13410 21772 14554
rect 22376 14544 22428 14550
rect 22376 14486 22428 14492
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 21928 14074 21956 14350
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 22020 13938 22048 14214
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 21880 13628 22188 13648
rect 21880 13626 21886 13628
rect 21942 13626 21966 13628
rect 22022 13626 22046 13628
rect 22102 13626 22126 13628
rect 22182 13626 22188 13628
rect 21942 13574 21944 13626
rect 22124 13574 22126 13626
rect 21880 13572 21886 13574
rect 21942 13572 21966 13574
rect 22022 13572 22046 13574
rect 22102 13572 22126 13574
rect 22182 13572 22188 13574
rect 21880 13552 22188 13572
rect 22296 13530 22324 13874
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 21744 13382 21864 13410
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21652 12850 21680 13126
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 21652 12442 21680 12786
rect 21744 12782 21772 13262
rect 21836 13258 21864 13382
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 21824 13252 21876 13258
rect 21824 13194 21876 13200
rect 22020 12918 22048 13262
rect 22008 12912 22060 12918
rect 22008 12854 22060 12860
rect 22192 12844 22244 12850
rect 22296 12832 22324 13466
rect 22388 12850 22416 14486
rect 22480 14346 22508 19314
rect 22558 19000 22614 19009
rect 22558 18935 22614 18944
rect 22572 18630 22600 18935
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 22572 16538 22600 18362
rect 22664 17338 22692 21830
rect 22848 21434 22876 22034
rect 23032 22030 23060 22986
rect 23492 22234 23520 22986
rect 23584 22778 23612 23054
rect 23572 22772 23624 22778
rect 23572 22714 23624 22720
rect 23480 22228 23532 22234
rect 23480 22170 23532 22176
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 23492 21554 23520 22170
rect 23584 22030 23612 22714
rect 24044 22030 24072 23122
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 23204 21548 23256 21554
rect 23204 21490 23256 21496
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 22756 21406 22876 21434
rect 22756 20398 22784 21406
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22928 21344 22980 21350
rect 22928 21286 22980 21292
rect 22848 20942 22876 21286
rect 22836 20936 22888 20942
rect 22836 20878 22888 20884
rect 22940 20602 22968 21286
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 23216 20534 23244 21490
rect 23296 21480 23348 21486
rect 23296 21422 23348 21428
rect 23308 21146 23336 21422
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23308 20534 23336 21082
rect 23492 20534 23520 21490
rect 23204 20528 23256 20534
rect 23204 20470 23256 20476
rect 23296 20528 23348 20534
rect 23296 20470 23348 20476
rect 23480 20528 23532 20534
rect 23480 20470 23532 20476
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22836 19712 22888 19718
rect 22836 19654 22888 19660
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 22848 19378 22876 19654
rect 23112 19440 23164 19446
rect 23112 19382 23164 19388
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 22836 18624 22888 18630
rect 22836 18566 22888 18572
rect 22744 18352 22796 18358
rect 22742 18320 22744 18329
rect 22796 18320 22798 18329
rect 22848 18290 22876 18566
rect 22742 18255 22798 18264
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22756 18034 22784 18158
rect 22848 18154 22876 18226
rect 22836 18148 22888 18154
rect 22836 18090 22888 18096
rect 22756 18006 22876 18034
rect 22848 17678 22876 18006
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22756 16658 22784 17614
rect 22848 17542 22876 17614
rect 22836 17536 22888 17542
rect 22836 17478 22888 17484
rect 22848 16726 22876 17478
rect 22836 16720 22888 16726
rect 22836 16662 22888 16668
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22836 16584 22888 16590
rect 22572 16510 22784 16538
rect 22836 16526 22888 16532
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22244 12804 22324 12832
rect 22376 12844 22428 12850
rect 22192 12786 22244 12792
rect 22376 12786 22428 12792
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21744 12238 21772 12718
rect 21880 12540 22188 12560
rect 21880 12538 21886 12540
rect 21942 12538 21966 12540
rect 22022 12538 22046 12540
rect 22102 12538 22126 12540
rect 22182 12538 22188 12540
rect 21942 12486 21944 12538
rect 22124 12486 22126 12538
rect 21880 12484 21886 12486
rect 21942 12484 21966 12486
rect 22022 12484 22046 12486
rect 22102 12484 22126 12486
rect 22182 12484 22188 12486
rect 21880 12464 22188 12484
rect 22480 12434 22508 14282
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22572 13326 22600 13806
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22480 12406 22600 12434
rect 22468 12368 22520 12374
rect 22466 12336 22468 12345
rect 22520 12336 22522 12345
rect 22466 12271 22522 12280
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21880 11452 22188 11472
rect 21880 11450 21886 11452
rect 21942 11450 21966 11452
rect 22022 11450 22046 11452
rect 22102 11450 22126 11452
rect 22182 11450 22188 11452
rect 21942 11398 21944 11450
rect 22124 11398 22126 11450
rect 21880 11396 21886 11398
rect 21942 11396 21966 11398
rect 22022 11396 22046 11398
rect 22102 11396 22126 11398
rect 22182 11396 22188 11398
rect 21880 11376 22188 11396
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 21192 10674 21220 10746
rect 21376 10674 21404 11086
rect 21732 11076 21784 11082
rect 21732 11018 21784 11024
rect 21456 11008 21508 11014
rect 21456 10950 21508 10956
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 20640 10130 20668 10610
rect 21468 10606 21496 10950
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 20088 9178 20116 9454
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 19904 8906 19932 8978
rect 20272 8974 20300 9590
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20364 9042 20392 9386
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 19904 8634 19932 8842
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 20364 7342 20392 7890
rect 20456 7546 20484 9318
rect 20732 7562 20760 9862
rect 20824 9722 20852 10406
rect 21744 10062 21772 11018
rect 22204 10810 22232 11222
rect 22572 11150 22600 12406
rect 22664 12238 22692 13670
rect 22756 12850 22784 16510
rect 22848 14550 22876 16526
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 22836 13932 22888 13938
rect 22836 13874 22888 13880
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22848 12730 22876 13874
rect 22940 12782 22968 18906
rect 23018 18320 23074 18329
rect 23018 18255 23074 18264
rect 23032 17814 23060 18255
rect 23124 18193 23152 19382
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23204 19168 23256 19174
rect 23204 19110 23256 19116
rect 23110 18184 23166 18193
rect 23110 18119 23166 18128
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 23216 17354 23244 19110
rect 23124 17326 23244 17354
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23032 15706 23060 17138
rect 23124 17134 23152 17326
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23124 15638 23152 16730
rect 23112 15632 23164 15638
rect 23112 15574 23164 15580
rect 23124 14600 23152 15574
rect 23216 15366 23244 17206
rect 23308 16794 23336 19246
rect 25056 19242 25084 19654
rect 25044 19236 25096 19242
rect 25044 19178 25096 19184
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23400 18358 23428 18634
rect 23388 18352 23440 18358
rect 23388 18294 23440 18300
rect 23478 18184 23534 18193
rect 23478 18119 23534 18128
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 23308 15450 23336 16458
rect 23400 15978 23428 16526
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 23492 15910 23520 18119
rect 24228 17746 24256 18702
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24136 16182 24164 16458
rect 24228 16250 24256 17682
rect 25778 17640 25834 17649
rect 25778 17575 25834 17584
rect 25792 17542 25820 17575
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 24124 16176 24176 16182
rect 24124 16118 24176 16124
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23492 15502 23520 15846
rect 23480 15496 23532 15502
rect 23308 15422 23428 15450
rect 23480 15438 23532 15444
rect 23204 15360 23256 15366
rect 23204 15302 23256 15308
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 23032 14572 23152 14600
rect 23032 13802 23060 14572
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 23020 13796 23072 13802
rect 23020 13738 23072 13744
rect 23124 13190 23152 14418
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 22756 12714 22876 12730
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 22744 12708 22876 12714
rect 22796 12702 22876 12708
rect 22744 12650 22796 12656
rect 22848 12374 22876 12702
rect 23020 12708 23072 12714
rect 23020 12650 23072 12656
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22388 10606 22416 11018
rect 22468 11008 22520 11014
rect 22468 10950 22520 10956
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 21880 10364 22188 10384
rect 21880 10362 21886 10364
rect 21942 10362 21966 10364
rect 22022 10362 22046 10364
rect 22102 10362 22126 10364
rect 22182 10362 22188 10364
rect 21942 10310 21944 10362
rect 22124 10310 22126 10362
rect 21880 10308 21886 10310
rect 21942 10308 21966 10310
rect 22022 10308 22046 10310
rect 22102 10308 22126 10310
rect 22182 10308 22188 10310
rect 21880 10288 22188 10308
rect 22296 10062 22324 10406
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 21008 9518 21036 9998
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 21008 8906 21036 9454
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 20444 7540 20496 7546
rect 20732 7534 20852 7562
rect 20444 7482 20496 7488
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20352 7336 20404 7342
rect 20352 7278 20404 7284
rect 20732 6458 20760 7346
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 19800 5364 19852 5370
rect 19800 5306 19852 5312
rect 19444 5234 19656 5250
rect 19432 5228 19656 5234
rect 19484 5222 19656 5228
rect 20628 5228 20680 5234
rect 19432 5170 19484 5176
rect 20628 5170 20680 5176
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19616 5160 19668 5166
rect 19616 5102 19668 5108
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19536 4826 19564 5102
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19628 4758 19656 5102
rect 19812 4758 19840 5102
rect 20352 5092 20404 5098
rect 20352 5034 20404 5040
rect 19616 4752 19668 4758
rect 19616 4694 19668 4700
rect 19800 4752 19852 4758
rect 19800 4694 19852 4700
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19352 3602 19380 3878
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 19076 3126 19104 3334
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 19352 3074 19380 3538
rect 19352 3058 19472 3074
rect 19352 3052 19484 3058
rect 19352 3046 19432 3052
rect 19432 2994 19484 3000
rect 19536 2990 19564 4558
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19628 3942 19656 4422
rect 19812 4010 19840 4694
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 20088 4010 20116 4422
rect 20364 4146 20392 5034
rect 20640 4690 20668 5170
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20456 4146 20484 4558
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 19800 4004 19852 4010
rect 19800 3946 19852 3952
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19812 3466 19840 3946
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20180 3534 20208 3878
rect 20364 3534 20392 4082
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 19616 3460 19668 3466
rect 19616 3402 19668 3408
rect 19800 3460 19852 3466
rect 19800 3402 19852 3408
rect 19628 3194 19656 3402
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 20456 2582 20484 4082
rect 20444 2576 20496 2582
rect 20444 2518 20496 2524
rect 20640 2446 20668 4626
rect 20732 4214 20760 6054
rect 20824 4554 20852 7534
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 21008 7410 21036 7482
rect 21652 7410 21680 7890
rect 21744 7886 21772 9318
rect 21880 9276 22188 9296
rect 21880 9274 21886 9276
rect 21942 9274 21966 9276
rect 22022 9274 22046 9276
rect 22102 9274 22126 9276
rect 22182 9274 22188 9276
rect 21942 9222 21944 9274
rect 22124 9222 22126 9274
rect 21880 9220 21886 9222
rect 21942 9220 21966 9222
rect 22022 9220 22046 9222
rect 22102 9220 22126 9222
rect 22182 9220 22188 9222
rect 21880 9200 22188 9220
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 21880 8188 22188 8208
rect 21880 8186 21886 8188
rect 21942 8186 21966 8188
rect 22022 8186 22046 8188
rect 22102 8186 22126 8188
rect 22182 8186 22188 8188
rect 21942 8134 21944 8186
rect 22124 8134 22126 8186
rect 21880 8132 21886 8134
rect 21942 8132 21966 8134
rect 22022 8132 22046 8134
rect 22102 8132 22126 8134
rect 22182 8132 22188 8134
rect 21880 8112 22188 8132
rect 22296 8022 22324 8230
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 22284 7812 22336 7818
rect 22284 7754 22336 7760
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21836 7410 21864 7482
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 20916 5930 20944 6258
rect 21008 6118 21036 7346
rect 22112 7274 22140 7686
rect 22204 7342 22232 7686
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 21880 7100 22188 7120
rect 21880 7098 21886 7100
rect 21942 7098 21966 7100
rect 22022 7098 22046 7100
rect 22102 7098 22126 7100
rect 22182 7098 22188 7100
rect 21942 7046 21944 7098
rect 22124 7046 22126 7098
rect 21880 7044 21886 7046
rect 21942 7044 21966 7046
rect 22022 7044 22046 7046
rect 22102 7044 22126 7046
rect 22182 7044 22188 7046
rect 21880 7024 22188 7044
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21192 6254 21220 6598
rect 21744 6458 21772 6598
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 20916 5902 21036 5930
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20916 4622 20944 5578
rect 21008 5370 21036 5902
rect 20996 5364 21048 5370
rect 20996 5306 21048 5312
rect 21192 4622 21220 6190
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 21284 4826 21312 5102
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 20904 4616 20956 4622
rect 21180 4616 21232 4622
rect 20956 4576 21128 4604
rect 20904 4558 20956 4564
rect 20812 4548 20864 4554
rect 20812 4490 20864 4496
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20916 3738 20944 4082
rect 21100 3738 21128 4576
rect 21376 4570 21404 5714
rect 21744 5710 21772 6394
rect 22100 6384 22152 6390
rect 22098 6352 22100 6361
rect 22152 6352 22154 6361
rect 22098 6287 22154 6296
rect 22296 6254 22324 7754
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 21880 6012 22188 6032
rect 21880 6010 21886 6012
rect 21942 6010 21966 6012
rect 22022 6010 22046 6012
rect 22102 6010 22126 6012
rect 22182 6010 22188 6012
rect 21942 5958 21944 6010
rect 22124 5958 22126 6010
rect 21880 5956 21886 5958
rect 21942 5956 21966 5958
rect 22022 5956 22046 5958
rect 22102 5956 22126 5958
rect 22182 5956 22188 5958
rect 21880 5936 22188 5956
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21468 5030 21496 5510
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21456 5024 21508 5030
rect 21456 4966 21508 4972
rect 21744 4826 21772 5034
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 21880 4924 22188 4944
rect 21880 4922 21886 4924
rect 21942 4922 21966 4924
rect 22022 4922 22046 4924
rect 22102 4922 22126 4924
rect 22182 4922 22188 4924
rect 21942 4870 21944 4922
rect 22124 4870 22126 4922
rect 21880 4868 21886 4870
rect 21942 4868 21966 4870
rect 22022 4868 22046 4870
rect 22102 4868 22126 4870
rect 22182 4868 22188 4870
rect 21880 4848 22188 4868
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 21180 4558 21232 4564
rect 21284 4542 21404 4570
rect 21640 4548 21692 4554
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 21100 3398 21128 3674
rect 21284 3602 21312 4542
rect 21640 4490 21692 4496
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21376 3942 21404 4422
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 20916 2446 20944 3334
rect 21284 3194 21312 3538
rect 21468 3194 21496 4014
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21560 3534 21588 3878
rect 21652 3738 21680 4490
rect 22204 4078 22232 4626
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 22296 3942 22324 4966
rect 22388 4622 22416 9862
rect 22480 9654 22508 10950
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22572 9722 22600 10746
rect 22652 10736 22704 10742
rect 22652 10678 22704 10684
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22468 9648 22520 9654
rect 22468 9590 22520 9596
rect 22664 9602 22692 10678
rect 22848 10554 22876 12310
rect 23032 11762 23060 12650
rect 23216 12434 23244 15302
rect 23308 15162 23336 15302
rect 23400 15162 23428 15422
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23308 14346 23336 15098
rect 23400 14822 23428 15098
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23400 13818 23428 14758
rect 23492 14414 23520 15438
rect 26332 15224 26384 15230
rect 26332 15166 26384 15172
rect 26344 14793 26372 15166
rect 26330 14784 26386 14793
rect 26330 14719 26386 14728
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23400 13790 23520 13818
rect 23386 13424 23442 13433
rect 23386 13359 23442 13368
rect 23400 13326 23428 13359
rect 23492 13326 23520 13790
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12850 23336 13126
rect 23492 12850 23520 13262
rect 23676 12850 23704 13262
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 23216 12406 23428 12434
rect 23400 11898 23428 12406
rect 25148 11937 25176 12582
rect 25134 11928 25190 11937
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 23388 11892 23440 11898
rect 25134 11863 25190 11872
rect 23388 11834 23440 11840
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 22928 11076 22980 11082
rect 22928 11018 22980 11024
rect 22756 10526 22876 10554
rect 22756 10130 22784 10526
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22756 9722 22784 9862
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 22664 9574 22784 9602
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22480 7886 22508 8774
rect 22468 7880 22520 7886
rect 22468 7822 22520 7828
rect 22664 5370 22692 9318
rect 22756 9217 22784 9574
rect 22742 9208 22798 9217
rect 22742 9143 22798 9152
rect 22848 8974 22876 10406
rect 22940 9178 22968 11018
rect 23032 10810 23060 11698
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 23124 10690 23152 11834
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23032 10674 23152 10690
rect 23020 10668 23152 10674
rect 23072 10662 23152 10668
rect 23020 10610 23072 10616
rect 23124 9722 23152 10662
rect 23112 9716 23164 9722
rect 23112 9658 23164 9664
rect 23216 9654 23244 11086
rect 23308 10606 23336 11154
rect 23296 10600 23348 10606
rect 23296 10542 23348 10548
rect 23308 10130 23336 10542
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 23308 9926 23336 10066
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 23216 8974 23244 9590
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23492 8974 23520 9318
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22756 6730 22784 7142
rect 22940 7002 22968 7686
rect 23216 7478 23244 7686
rect 23204 7472 23256 7478
rect 23204 7414 23256 7420
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 23032 6798 23060 7346
rect 23848 7200 23900 7206
rect 23848 7142 23900 7148
rect 23860 6914 23888 7142
rect 23768 6886 23888 6914
rect 23768 6798 23796 6886
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 22744 6724 22796 6730
rect 22744 6666 22796 6672
rect 22652 5364 22704 5370
rect 22652 5306 22704 5312
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22480 4690 22508 5102
rect 23032 4826 23060 6734
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23400 6322 23428 6598
rect 23492 6390 23520 6734
rect 23480 6384 23532 6390
rect 23480 6326 23532 6332
rect 23768 6322 23796 6734
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23400 5234 23428 6258
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23492 5914 23520 6054
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23848 5160 23900 5166
rect 23848 5102 23900 5108
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22664 4214 22692 4422
rect 22652 4208 22704 4214
rect 22652 4150 22704 4156
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 21880 3836 22188 3856
rect 21880 3834 21886 3836
rect 21942 3834 21966 3836
rect 22022 3834 22046 3836
rect 22102 3834 22126 3836
rect 22182 3834 22188 3836
rect 21942 3782 21944 3834
rect 22124 3782 22126 3834
rect 21880 3780 21886 3782
rect 21942 3780 21966 3782
rect 22022 3780 22046 3782
rect 22102 3780 22126 3782
rect 22182 3780 22188 3782
rect 21880 3760 22188 3780
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 21652 3602 21680 3674
rect 21640 3596 21692 3602
rect 21640 3538 21692 3544
rect 22756 3534 22784 4626
rect 23860 4214 23888 5102
rect 24124 5092 24176 5098
rect 24124 5034 24176 5040
rect 24136 4826 24164 5034
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 23848 4208 23900 4214
rect 23216 4146 23520 4162
rect 23848 4150 23900 4156
rect 23216 4140 23532 4146
rect 23216 4134 23480 4140
rect 23216 4078 23244 4134
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23308 3738 23336 4014
rect 23400 3738 23428 4134
rect 23480 4082 23532 4088
rect 24596 4010 24624 4558
rect 24584 4004 24636 4010
rect 24584 3946 24636 3952
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 21548 3528 21600 3534
rect 22744 3528 22796 3534
rect 21548 3470 21600 3476
rect 22098 3496 22154 3505
rect 22744 3470 22796 3476
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 22098 3431 22154 3440
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 22112 2922 22140 3431
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 22836 2848 22888 2854
rect 22836 2790 22888 2796
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 20180 800 20208 2382
rect 21560 800 21588 2790
rect 21880 2748 22188 2768
rect 21880 2746 21886 2748
rect 21942 2746 21966 2748
rect 22022 2746 22046 2748
rect 22102 2746 22126 2748
rect 22182 2746 22188 2748
rect 21942 2694 21944 2746
rect 22124 2694 22126 2746
rect 21880 2692 21886 2694
rect 21942 2692 21966 2694
rect 22022 2692 22046 2694
rect 22102 2692 22126 2694
rect 22182 2692 22188 2694
rect 21880 2672 22188 2692
rect 22100 1352 22152 1358
rect 22100 1294 22152 1300
rect 14568 734 14964 762
rect 15014 0 15070 800
rect 16302 0 16358 800
rect 17590 0 17646 800
rect 18878 0 18934 800
rect 20166 0 20222 800
rect 21546 0 21602 800
rect 22112 785 22140 1294
rect 22848 800 22876 2790
rect 24136 800 24164 3470
rect 26712 800 26740 3470
rect 22098 776 22154 785
rect 22098 711 22154 720
rect 22834 0 22890 800
rect 24122 0 24178 800
rect 25410 0 25466 800
rect 26698 0 26754 800
<< via2 >>
rect 4066 17448 4122 17504
rect 5142 26682 5198 26684
rect 5222 26682 5278 26684
rect 5302 26682 5358 26684
rect 5382 26682 5438 26684
rect 5142 26630 5188 26682
rect 5188 26630 5198 26682
rect 5222 26630 5252 26682
rect 5252 26630 5264 26682
rect 5264 26630 5278 26682
rect 5302 26630 5316 26682
rect 5316 26630 5328 26682
rect 5328 26630 5358 26682
rect 5382 26630 5392 26682
rect 5392 26630 5438 26682
rect 5142 26628 5198 26630
rect 5222 26628 5278 26630
rect 5302 26628 5358 26630
rect 5382 26628 5438 26630
rect 5142 25594 5198 25596
rect 5222 25594 5278 25596
rect 5302 25594 5358 25596
rect 5382 25594 5438 25596
rect 5142 25542 5188 25594
rect 5188 25542 5198 25594
rect 5222 25542 5252 25594
rect 5252 25542 5264 25594
rect 5264 25542 5278 25594
rect 5302 25542 5316 25594
rect 5316 25542 5328 25594
rect 5328 25542 5358 25594
rect 5382 25542 5392 25594
rect 5392 25542 5438 25594
rect 5142 25540 5198 25542
rect 5222 25540 5278 25542
rect 5302 25540 5358 25542
rect 5382 25540 5438 25542
rect 5142 24506 5198 24508
rect 5222 24506 5278 24508
rect 5302 24506 5358 24508
rect 5382 24506 5438 24508
rect 5142 24454 5188 24506
rect 5188 24454 5198 24506
rect 5222 24454 5252 24506
rect 5252 24454 5264 24506
rect 5264 24454 5278 24506
rect 5302 24454 5316 24506
rect 5316 24454 5328 24506
rect 5328 24454 5358 24506
rect 5382 24454 5392 24506
rect 5392 24454 5438 24506
rect 5142 24452 5198 24454
rect 5222 24452 5278 24454
rect 5302 24452 5358 24454
rect 5382 24452 5438 24454
rect 5142 23418 5198 23420
rect 5222 23418 5278 23420
rect 5302 23418 5358 23420
rect 5382 23418 5438 23420
rect 5142 23366 5188 23418
rect 5188 23366 5198 23418
rect 5222 23366 5252 23418
rect 5252 23366 5264 23418
rect 5264 23366 5278 23418
rect 5302 23366 5316 23418
rect 5316 23366 5328 23418
rect 5328 23366 5358 23418
rect 5382 23366 5392 23418
rect 5392 23366 5438 23418
rect 5142 23364 5198 23366
rect 5222 23364 5278 23366
rect 5302 23364 5358 23366
rect 5382 23364 5438 23366
rect 5142 22330 5198 22332
rect 5222 22330 5278 22332
rect 5302 22330 5358 22332
rect 5382 22330 5438 22332
rect 5142 22278 5188 22330
rect 5188 22278 5198 22330
rect 5222 22278 5252 22330
rect 5252 22278 5264 22330
rect 5264 22278 5278 22330
rect 5302 22278 5316 22330
rect 5316 22278 5328 22330
rect 5328 22278 5358 22330
rect 5382 22278 5392 22330
rect 5392 22278 5438 22330
rect 5142 22276 5198 22278
rect 5222 22276 5278 22278
rect 5302 22276 5358 22278
rect 5382 22276 5438 22278
rect 5142 21242 5198 21244
rect 5222 21242 5278 21244
rect 5302 21242 5358 21244
rect 5382 21242 5438 21244
rect 5142 21190 5188 21242
rect 5188 21190 5198 21242
rect 5222 21190 5252 21242
rect 5252 21190 5264 21242
rect 5264 21190 5278 21242
rect 5302 21190 5316 21242
rect 5316 21190 5328 21242
rect 5328 21190 5358 21242
rect 5382 21190 5392 21242
rect 5392 21190 5438 21242
rect 5142 21188 5198 21190
rect 5222 21188 5278 21190
rect 5302 21188 5358 21190
rect 5382 21188 5438 21190
rect 5262 20304 5318 20360
rect 5142 20154 5198 20156
rect 5222 20154 5278 20156
rect 5302 20154 5358 20156
rect 5382 20154 5438 20156
rect 5142 20102 5188 20154
rect 5188 20102 5198 20154
rect 5222 20102 5252 20154
rect 5252 20102 5264 20154
rect 5264 20102 5278 20154
rect 5302 20102 5316 20154
rect 5316 20102 5328 20154
rect 5328 20102 5358 20154
rect 5382 20102 5392 20154
rect 5392 20102 5438 20154
rect 5142 20100 5198 20102
rect 5222 20100 5278 20102
rect 5302 20100 5358 20102
rect 5382 20100 5438 20102
rect 5142 19066 5198 19068
rect 5222 19066 5278 19068
rect 5302 19066 5358 19068
rect 5382 19066 5438 19068
rect 5142 19014 5188 19066
rect 5188 19014 5198 19066
rect 5222 19014 5252 19066
rect 5252 19014 5264 19066
rect 5264 19014 5278 19066
rect 5302 19014 5316 19066
rect 5316 19014 5328 19066
rect 5328 19014 5358 19066
rect 5382 19014 5392 19066
rect 5392 19014 5438 19066
rect 5142 19012 5198 19014
rect 5222 19012 5278 19014
rect 5302 19012 5358 19014
rect 5382 19012 5438 19014
rect 5142 17978 5198 17980
rect 5222 17978 5278 17980
rect 5302 17978 5358 17980
rect 5382 17978 5438 17980
rect 5142 17926 5188 17978
rect 5188 17926 5198 17978
rect 5222 17926 5252 17978
rect 5252 17926 5264 17978
rect 5264 17926 5278 17978
rect 5302 17926 5316 17978
rect 5316 17926 5328 17978
rect 5328 17926 5358 17978
rect 5382 17926 5392 17978
rect 5392 17926 5438 17978
rect 5142 17924 5198 17926
rect 5222 17924 5278 17926
rect 5302 17924 5358 17926
rect 5382 17924 5438 17926
rect 6182 17196 6238 17232
rect 6182 17176 6184 17196
rect 6184 17176 6236 17196
rect 6236 17176 6238 17196
rect 5142 16890 5198 16892
rect 5222 16890 5278 16892
rect 5302 16890 5358 16892
rect 5382 16890 5438 16892
rect 5142 16838 5188 16890
rect 5188 16838 5198 16890
rect 5222 16838 5252 16890
rect 5252 16838 5264 16890
rect 5264 16838 5278 16890
rect 5302 16838 5316 16890
rect 5316 16838 5328 16890
rect 5328 16838 5358 16890
rect 5382 16838 5392 16890
rect 5392 16838 5438 16890
rect 5142 16836 5198 16838
rect 5222 16836 5278 16838
rect 5302 16836 5358 16838
rect 5382 16836 5438 16838
rect 5142 15802 5198 15804
rect 5222 15802 5278 15804
rect 5302 15802 5358 15804
rect 5382 15802 5438 15804
rect 5142 15750 5188 15802
rect 5188 15750 5198 15802
rect 5222 15750 5252 15802
rect 5252 15750 5264 15802
rect 5264 15750 5278 15802
rect 5302 15750 5316 15802
rect 5316 15750 5328 15802
rect 5328 15750 5358 15802
rect 5382 15750 5392 15802
rect 5392 15750 5438 15802
rect 5142 15748 5198 15750
rect 5222 15748 5278 15750
rect 5302 15748 5358 15750
rect 5382 15748 5438 15750
rect 2962 12824 3018 12880
rect 3514 12844 3570 12880
rect 3514 12824 3516 12844
rect 3516 12824 3568 12844
rect 3568 12824 3570 12844
rect 5142 14714 5198 14716
rect 5222 14714 5278 14716
rect 5302 14714 5358 14716
rect 5382 14714 5438 14716
rect 5142 14662 5188 14714
rect 5188 14662 5198 14714
rect 5222 14662 5252 14714
rect 5252 14662 5264 14714
rect 5264 14662 5278 14714
rect 5302 14662 5316 14714
rect 5316 14662 5328 14714
rect 5328 14662 5358 14714
rect 5382 14662 5392 14714
rect 5392 14662 5438 14714
rect 5142 14660 5198 14662
rect 5222 14660 5278 14662
rect 5302 14660 5358 14662
rect 5382 14660 5438 14662
rect 5142 13626 5198 13628
rect 5222 13626 5278 13628
rect 5302 13626 5358 13628
rect 5382 13626 5438 13628
rect 5142 13574 5188 13626
rect 5188 13574 5198 13626
rect 5222 13574 5252 13626
rect 5252 13574 5264 13626
rect 5264 13574 5278 13626
rect 5302 13574 5316 13626
rect 5316 13574 5328 13626
rect 5328 13574 5358 13626
rect 5382 13574 5392 13626
rect 5392 13574 5438 13626
rect 5142 13572 5198 13574
rect 5222 13572 5278 13574
rect 5302 13572 5358 13574
rect 5382 13572 5438 13574
rect 5170 12844 5226 12880
rect 5170 12824 5172 12844
rect 5172 12824 5224 12844
rect 5224 12824 5226 12844
rect 5538 12824 5594 12880
rect 5142 12538 5198 12540
rect 5222 12538 5278 12540
rect 5302 12538 5358 12540
rect 5382 12538 5438 12540
rect 5142 12486 5188 12538
rect 5188 12486 5198 12538
rect 5222 12486 5252 12538
rect 5252 12486 5264 12538
rect 5264 12486 5278 12538
rect 5302 12486 5316 12538
rect 5316 12486 5328 12538
rect 5328 12486 5358 12538
rect 5382 12486 5392 12538
rect 5392 12486 5438 12538
rect 5142 12484 5198 12486
rect 5222 12484 5278 12486
rect 5302 12484 5358 12486
rect 5382 12484 5438 12486
rect 6826 14048 6882 14104
rect 4986 11872 5042 11928
rect 5170 11736 5226 11792
rect 5142 11450 5198 11452
rect 5222 11450 5278 11452
rect 5302 11450 5358 11452
rect 5382 11450 5438 11452
rect 5142 11398 5188 11450
rect 5188 11398 5198 11450
rect 5222 11398 5252 11450
rect 5252 11398 5264 11450
rect 5264 11398 5278 11450
rect 5302 11398 5316 11450
rect 5316 11398 5328 11450
rect 5328 11398 5358 11450
rect 5382 11398 5392 11450
rect 5392 11398 5438 11450
rect 5142 11396 5198 11398
rect 5222 11396 5278 11398
rect 5302 11396 5358 11398
rect 5382 11396 5438 11398
rect 3974 8200 4030 8256
rect 5142 10362 5198 10364
rect 5222 10362 5278 10364
rect 5302 10362 5358 10364
rect 5382 10362 5438 10364
rect 5142 10310 5188 10362
rect 5188 10310 5198 10362
rect 5222 10310 5252 10362
rect 5252 10310 5264 10362
rect 5264 10310 5278 10362
rect 5302 10310 5316 10362
rect 5316 10310 5328 10362
rect 5328 10310 5358 10362
rect 5382 10310 5392 10362
rect 5392 10310 5438 10362
rect 5142 10308 5198 10310
rect 5222 10308 5278 10310
rect 5302 10308 5358 10310
rect 5382 10308 5438 10310
rect 5142 9274 5198 9276
rect 5222 9274 5278 9276
rect 5302 9274 5358 9276
rect 5382 9274 5438 9276
rect 5142 9222 5188 9274
rect 5188 9222 5198 9274
rect 5222 9222 5252 9274
rect 5252 9222 5264 9274
rect 5264 9222 5278 9274
rect 5302 9222 5316 9274
rect 5316 9222 5328 9274
rect 5328 9222 5358 9274
rect 5382 9222 5392 9274
rect 5392 9222 5438 9274
rect 5142 9220 5198 9222
rect 5222 9220 5278 9222
rect 5302 9220 5358 9222
rect 5382 9220 5438 9222
rect 662 3440 718 3496
rect 2962 856 3018 912
rect 5142 8186 5198 8188
rect 5222 8186 5278 8188
rect 5302 8186 5358 8188
rect 5382 8186 5438 8188
rect 5142 8134 5188 8186
rect 5188 8134 5198 8186
rect 5222 8134 5252 8186
rect 5252 8134 5264 8186
rect 5264 8134 5278 8186
rect 5302 8134 5316 8186
rect 5316 8134 5328 8186
rect 5328 8134 5358 8186
rect 5382 8134 5392 8186
rect 5392 8134 5438 8186
rect 5142 8132 5198 8134
rect 5222 8132 5278 8134
rect 5302 8132 5358 8134
rect 5382 8132 5438 8134
rect 7286 19372 7342 19408
rect 7286 19352 7288 19372
rect 7288 19352 7340 19372
rect 7340 19352 7342 19372
rect 7378 13912 7434 13968
rect 5142 7098 5198 7100
rect 5222 7098 5278 7100
rect 5302 7098 5358 7100
rect 5382 7098 5438 7100
rect 5142 7046 5188 7098
rect 5188 7046 5198 7098
rect 5222 7046 5252 7098
rect 5252 7046 5264 7098
rect 5264 7046 5278 7098
rect 5302 7046 5316 7098
rect 5316 7046 5328 7098
rect 5328 7046 5358 7098
rect 5382 7046 5392 7098
rect 5392 7046 5438 7098
rect 5142 7044 5198 7046
rect 5222 7044 5278 7046
rect 5302 7044 5358 7046
rect 5382 7044 5438 7046
rect 4986 6296 5042 6352
rect 5142 6010 5198 6012
rect 5222 6010 5278 6012
rect 5302 6010 5358 6012
rect 5382 6010 5438 6012
rect 5142 5958 5188 6010
rect 5188 5958 5198 6010
rect 5222 5958 5252 6010
rect 5252 5958 5264 6010
rect 5264 5958 5278 6010
rect 5302 5958 5316 6010
rect 5316 5958 5328 6010
rect 5328 5958 5358 6010
rect 5382 5958 5392 6010
rect 5392 5958 5438 6010
rect 5142 5956 5198 5958
rect 5222 5956 5278 5958
rect 5302 5956 5358 5958
rect 5382 5956 5438 5958
rect 6090 6296 6146 6352
rect 5142 4922 5198 4924
rect 5222 4922 5278 4924
rect 5302 4922 5358 4924
rect 5382 4922 5438 4924
rect 5142 4870 5188 4922
rect 5188 4870 5198 4922
rect 5222 4870 5252 4922
rect 5252 4870 5264 4922
rect 5264 4870 5278 4922
rect 5302 4870 5316 4922
rect 5316 4870 5328 4922
rect 5328 4870 5358 4922
rect 5382 4870 5392 4922
rect 5392 4870 5438 4922
rect 5142 4868 5198 4870
rect 5222 4868 5278 4870
rect 5302 4868 5358 4870
rect 5382 4868 5438 4870
rect 5142 3834 5198 3836
rect 5222 3834 5278 3836
rect 5302 3834 5358 3836
rect 5382 3834 5438 3836
rect 5142 3782 5188 3834
rect 5188 3782 5198 3834
rect 5222 3782 5252 3834
rect 5252 3782 5264 3834
rect 5264 3782 5278 3834
rect 5302 3782 5316 3834
rect 5316 3782 5328 3834
rect 5328 3782 5358 3834
rect 5382 3782 5392 3834
rect 5392 3782 5438 3834
rect 5142 3780 5198 3782
rect 5222 3780 5278 3782
rect 5302 3780 5358 3782
rect 5382 3780 5438 3782
rect 5142 2746 5198 2748
rect 5222 2746 5278 2748
rect 5302 2746 5358 2748
rect 5382 2746 5438 2748
rect 5142 2694 5188 2746
rect 5188 2694 5198 2746
rect 5222 2694 5252 2746
rect 5252 2694 5264 2746
rect 5264 2694 5278 2746
rect 5302 2694 5316 2746
rect 5316 2694 5328 2746
rect 5328 2694 5358 2746
rect 5382 2694 5392 2746
rect 5392 2694 5438 2746
rect 5142 2692 5198 2694
rect 5222 2692 5278 2694
rect 5302 2692 5358 2694
rect 5382 2692 5438 2694
rect 9328 27226 9384 27228
rect 9408 27226 9464 27228
rect 9488 27226 9544 27228
rect 9568 27226 9624 27228
rect 9328 27174 9374 27226
rect 9374 27174 9384 27226
rect 9408 27174 9438 27226
rect 9438 27174 9450 27226
rect 9450 27174 9464 27226
rect 9488 27174 9502 27226
rect 9502 27174 9514 27226
rect 9514 27174 9544 27226
rect 9568 27174 9578 27226
rect 9578 27174 9624 27226
rect 9328 27172 9384 27174
rect 9408 27172 9464 27174
rect 9488 27172 9544 27174
rect 9568 27172 9624 27174
rect 9328 26138 9384 26140
rect 9408 26138 9464 26140
rect 9488 26138 9544 26140
rect 9568 26138 9624 26140
rect 9328 26086 9374 26138
rect 9374 26086 9384 26138
rect 9408 26086 9438 26138
rect 9438 26086 9450 26138
rect 9450 26086 9464 26138
rect 9488 26086 9502 26138
rect 9502 26086 9514 26138
rect 9514 26086 9544 26138
rect 9568 26086 9578 26138
rect 9578 26086 9624 26138
rect 9328 26084 9384 26086
rect 9408 26084 9464 26086
rect 9488 26084 9544 26086
rect 9568 26084 9624 26086
rect 9328 25050 9384 25052
rect 9408 25050 9464 25052
rect 9488 25050 9544 25052
rect 9568 25050 9624 25052
rect 9328 24998 9374 25050
rect 9374 24998 9384 25050
rect 9408 24998 9438 25050
rect 9438 24998 9450 25050
rect 9450 24998 9464 25050
rect 9488 24998 9502 25050
rect 9502 24998 9514 25050
rect 9514 24998 9544 25050
rect 9568 24998 9578 25050
rect 9578 24998 9624 25050
rect 9328 24996 9384 24998
rect 9408 24996 9464 24998
rect 9488 24996 9544 24998
rect 9568 24996 9624 24998
rect 7746 19352 7802 19408
rect 7746 17176 7802 17232
rect 8022 14048 8078 14104
rect 8298 16108 8354 16144
rect 8298 16088 8300 16108
rect 8300 16088 8352 16108
rect 8352 16088 8354 16108
rect 8298 13796 8354 13832
rect 8298 13776 8300 13796
rect 8300 13776 8352 13796
rect 8352 13776 8354 13796
rect 9328 23962 9384 23964
rect 9408 23962 9464 23964
rect 9488 23962 9544 23964
rect 9568 23962 9624 23964
rect 9328 23910 9374 23962
rect 9374 23910 9384 23962
rect 9408 23910 9438 23962
rect 9438 23910 9450 23962
rect 9450 23910 9464 23962
rect 9488 23910 9502 23962
rect 9502 23910 9514 23962
rect 9514 23910 9544 23962
rect 9568 23910 9578 23962
rect 9578 23910 9624 23962
rect 9328 23908 9384 23910
rect 9408 23908 9464 23910
rect 9488 23908 9544 23910
rect 9568 23908 9624 23910
rect 9328 22874 9384 22876
rect 9408 22874 9464 22876
rect 9488 22874 9544 22876
rect 9568 22874 9624 22876
rect 9328 22822 9374 22874
rect 9374 22822 9384 22874
rect 9408 22822 9438 22874
rect 9438 22822 9450 22874
rect 9450 22822 9464 22874
rect 9488 22822 9502 22874
rect 9502 22822 9514 22874
rect 9514 22822 9544 22874
rect 9568 22822 9578 22874
rect 9578 22822 9624 22874
rect 9328 22820 9384 22822
rect 9408 22820 9464 22822
rect 9488 22820 9544 22822
rect 9568 22820 9624 22822
rect 9328 21786 9384 21788
rect 9408 21786 9464 21788
rect 9488 21786 9544 21788
rect 9568 21786 9624 21788
rect 9328 21734 9374 21786
rect 9374 21734 9384 21786
rect 9408 21734 9438 21786
rect 9438 21734 9450 21786
rect 9450 21734 9464 21786
rect 9488 21734 9502 21786
rect 9502 21734 9514 21786
rect 9514 21734 9544 21786
rect 9568 21734 9578 21786
rect 9578 21734 9624 21786
rect 9328 21732 9384 21734
rect 9408 21732 9464 21734
rect 9488 21732 9544 21734
rect 9568 21732 9624 21734
rect 9328 20698 9384 20700
rect 9408 20698 9464 20700
rect 9488 20698 9544 20700
rect 9568 20698 9624 20700
rect 9328 20646 9374 20698
rect 9374 20646 9384 20698
rect 9408 20646 9438 20698
rect 9438 20646 9450 20698
rect 9450 20646 9464 20698
rect 9488 20646 9502 20698
rect 9502 20646 9514 20698
rect 9514 20646 9544 20698
rect 9568 20646 9578 20698
rect 9578 20646 9624 20698
rect 9328 20644 9384 20646
rect 9408 20644 9464 20646
rect 9488 20644 9544 20646
rect 9568 20644 9624 20646
rect 9862 20304 9918 20360
rect 8942 18708 8944 18728
rect 8944 18708 8996 18728
rect 8996 18708 8998 18728
rect 8942 18672 8998 18708
rect 8666 17196 8722 17232
rect 8666 17176 8668 17196
rect 8668 17176 8720 17196
rect 8720 17176 8722 17196
rect 9328 19610 9384 19612
rect 9408 19610 9464 19612
rect 9488 19610 9544 19612
rect 9568 19610 9624 19612
rect 9328 19558 9374 19610
rect 9374 19558 9384 19610
rect 9408 19558 9438 19610
rect 9438 19558 9450 19610
rect 9450 19558 9464 19610
rect 9488 19558 9502 19610
rect 9502 19558 9514 19610
rect 9514 19558 9544 19610
rect 9568 19558 9578 19610
rect 9578 19558 9624 19610
rect 9328 19556 9384 19558
rect 9408 19556 9464 19558
rect 9488 19556 9544 19558
rect 9568 19556 9624 19558
rect 9328 18522 9384 18524
rect 9408 18522 9464 18524
rect 9488 18522 9544 18524
rect 9568 18522 9624 18524
rect 9328 18470 9374 18522
rect 9374 18470 9384 18522
rect 9408 18470 9438 18522
rect 9438 18470 9450 18522
rect 9450 18470 9464 18522
rect 9488 18470 9502 18522
rect 9502 18470 9514 18522
rect 9514 18470 9544 18522
rect 9568 18470 9578 18522
rect 9578 18470 9624 18522
rect 9328 18468 9384 18470
rect 9408 18468 9464 18470
rect 9488 18468 9544 18470
rect 9568 18468 9624 18470
rect 8666 13912 8722 13968
rect 10138 18808 10194 18864
rect 9328 17434 9384 17436
rect 9408 17434 9464 17436
rect 9488 17434 9544 17436
rect 9568 17434 9624 17436
rect 9328 17382 9374 17434
rect 9374 17382 9384 17434
rect 9408 17382 9438 17434
rect 9438 17382 9450 17434
rect 9450 17382 9464 17434
rect 9488 17382 9502 17434
rect 9502 17382 9514 17434
rect 9514 17382 9544 17434
rect 9568 17382 9578 17434
rect 9578 17382 9624 17434
rect 9328 17380 9384 17382
rect 9408 17380 9464 17382
rect 9488 17380 9544 17382
rect 9568 17380 9624 17382
rect 9494 17212 9496 17232
rect 9496 17212 9548 17232
rect 9548 17212 9550 17232
rect 9494 17176 9550 17212
rect 9402 16632 9458 16688
rect 9586 16632 9642 16688
rect 9328 16346 9384 16348
rect 9408 16346 9464 16348
rect 9488 16346 9544 16348
rect 9568 16346 9624 16348
rect 9328 16294 9374 16346
rect 9374 16294 9384 16346
rect 9408 16294 9438 16346
rect 9438 16294 9450 16346
rect 9450 16294 9464 16346
rect 9488 16294 9502 16346
rect 9502 16294 9514 16346
rect 9514 16294 9544 16346
rect 9568 16294 9578 16346
rect 9578 16294 9624 16346
rect 9328 16292 9384 16294
rect 9408 16292 9464 16294
rect 9488 16292 9544 16294
rect 9568 16292 9624 16294
rect 9586 16124 9588 16144
rect 9588 16124 9640 16144
rect 9640 16124 9642 16144
rect 9586 16088 9642 16124
rect 9328 15258 9384 15260
rect 9408 15258 9464 15260
rect 9488 15258 9544 15260
rect 9568 15258 9624 15260
rect 9328 15206 9374 15258
rect 9374 15206 9384 15258
rect 9408 15206 9438 15258
rect 9438 15206 9450 15258
rect 9450 15206 9464 15258
rect 9488 15206 9502 15258
rect 9502 15206 9514 15258
rect 9514 15206 9544 15258
rect 9568 15206 9578 15258
rect 9578 15206 9624 15258
rect 9328 15204 9384 15206
rect 9408 15204 9464 15206
rect 9488 15204 9544 15206
rect 9568 15204 9624 15206
rect 9494 14764 9496 14784
rect 9496 14764 9548 14784
rect 9548 14764 9550 14784
rect 9494 14728 9550 14764
rect 8390 12824 8446 12880
rect 9328 14170 9384 14172
rect 9408 14170 9464 14172
rect 9488 14170 9544 14172
rect 9568 14170 9624 14172
rect 9328 14118 9374 14170
rect 9374 14118 9384 14170
rect 9408 14118 9438 14170
rect 9438 14118 9450 14170
rect 9450 14118 9464 14170
rect 9488 14118 9502 14170
rect 9502 14118 9514 14170
rect 9514 14118 9544 14170
rect 9568 14118 9578 14170
rect 9578 14118 9624 14170
rect 9328 14116 9384 14118
rect 9408 14116 9464 14118
rect 9488 14116 9544 14118
rect 9568 14116 9624 14118
rect 9310 13948 9312 13968
rect 9312 13948 9364 13968
rect 9364 13948 9366 13968
rect 9310 13912 9366 13948
rect 6550 5344 6606 5400
rect 6642 5108 6644 5128
rect 6644 5108 6696 5128
rect 6696 5108 6698 5128
rect 6642 5072 6698 5108
rect 7194 5344 7250 5400
rect 8206 6840 8262 6896
rect 7470 4800 7526 4856
rect 7838 5208 7894 5264
rect 8022 5228 8078 5264
rect 8022 5208 8024 5228
rect 8024 5208 8076 5228
rect 8076 5208 8078 5228
rect 9328 13082 9384 13084
rect 9408 13082 9464 13084
rect 9488 13082 9544 13084
rect 9568 13082 9624 13084
rect 9328 13030 9374 13082
rect 9374 13030 9384 13082
rect 9408 13030 9438 13082
rect 9438 13030 9450 13082
rect 9450 13030 9464 13082
rect 9488 13030 9502 13082
rect 9502 13030 9514 13082
rect 9514 13030 9544 13082
rect 9568 13030 9578 13082
rect 9578 13030 9624 13082
rect 9328 13028 9384 13030
rect 9408 13028 9464 13030
rect 9488 13028 9544 13030
rect 9568 13028 9624 13030
rect 9954 12844 10010 12880
rect 9954 12824 9956 12844
rect 9956 12824 10008 12844
rect 10008 12824 10010 12844
rect 9328 11994 9384 11996
rect 9408 11994 9464 11996
rect 9488 11994 9544 11996
rect 9568 11994 9624 11996
rect 9328 11942 9374 11994
rect 9374 11942 9384 11994
rect 9408 11942 9438 11994
rect 9438 11942 9450 11994
rect 9450 11942 9464 11994
rect 9488 11942 9502 11994
rect 9502 11942 9514 11994
rect 9514 11942 9544 11994
rect 9568 11942 9578 11994
rect 9578 11942 9624 11994
rect 9328 11940 9384 11942
rect 9408 11940 9464 11942
rect 9488 11940 9544 11942
rect 9568 11940 9624 11942
rect 9586 11772 9588 11792
rect 9588 11772 9640 11792
rect 9640 11772 9642 11792
rect 9586 11736 9642 11772
rect 9328 10906 9384 10908
rect 9408 10906 9464 10908
rect 9488 10906 9544 10908
rect 9568 10906 9624 10908
rect 9328 10854 9374 10906
rect 9374 10854 9384 10906
rect 9408 10854 9438 10906
rect 9438 10854 9450 10906
rect 9450 10854 9464 10906
rect 9488 10854 9502 10906
rect 9502 10854 9514 10906
rect 9514 10854 9544 10906
rect 9568 10854 9578 10906
rect 9578 10854 9624 10906
rect 9328 10852 9384 10854
rect 9408 10852 9464 10854
rect 9488 10852 9544 10854
rect 9568 10852 9624 10854
rect 9328 9818 9384 9820
rect 9408 9818 9464 9820
rect 9488 9818 9544 9820
rect 9568 9818 9624 9820
rect 9328 9766 9374 9818
rect 9374 9766 9384 9818
rect 9408 9766 9438 9818
rect 9438 9766 9450 9818
rect 9450 9766 9464 9818
rect 9488 9766 9502 9818
rect 9502 9766 9514 9818
rect 9514 9766 9544 9818
rect 9568 9766 9578 9818
rect 9578 9766 9624 9818
rect 9328 9764 9384 9766
rect 9408 9764 9464 9766
rect 9488 9764 9544 9766
rect 9568 9764 9624 9766
rect 8666 7928 8722 7984
rect 9034 7384 9090 7440
rect 8758 6296 8814 6352
rect 8850 5092 8906 5128
rect 8850 5072 8852 5092
rect 8852 5072 8904 5092
rect 8904 5072 8906 5092
rect 13514 26682 13570 26684
rect 13594 26682 13650 26684
rect 13674 26682 13730 26684
rect 13754 26682 13810 26684
rect 13514 26630 13560 26682
rect 13560 26630 13570 26682
rect 13594 26630 13624 26682
rect 13624 26630 13636 26682
rect 13636 26630 13650 26682
rect 13674 26630 13688 26682
rect 13688 26630 13700 26682
rect 13700 26630 13730 26682
rect 13754 26630 13764 26682
rect 13764 26630 13810 26682
rect 13514 26628 13570 26630
rect 13594 26628 13650 26630
rect 13674 26628 13730 26630
rect 13754 26628 13810 26630
rect 9328 8730 9384 8732
rect 9408 8730 9464 8732
rect 9488 8730 9544 8732
rect 9568 8730 9624 8732
rect 9328 8678 9374 8730
rect 9374 8678 9384 8730
rect 9408 8678 9438 8730
rect 9438 8678 9450 8730
rect 9450 8678 9464 8730
rect 9488 8678 9502 8730
rect 9502 8678 9514 8730
rect 9514 8678 9544 8730
rect 9568 8678 9578 8730
rect 9578 8678 9624 8730
rect 9328 8676 9384 8678
rect 9408 8676 9464 8678
rect 9488 8676 9544 8678
rect 9568 8676 9624 8678
rect 9586 7928 9642 7984
rect 9328 7642 9384 7644
rect 9408 7642 9464 7644
rect 9488 7642 9544 7644
rect 9568 7642 9624 7644
rect 9328 7590 9374 7642
rect 9374 7590 9384 7642
rect 9408 7590 9438 7642
rect 9438 7590 9450 7642
rect 9450 7590 9464 7642
rect 9488 7590 9502 7642
rect 9502 7590 9514 7642
rect 9514 7590 9544 7642
rect 9568 7590 9578 7642
rect 9578 7590 9624 7642
rect 9328 7588 9384 7590
rect 9408 7588 9464 7590
rect 9488 7588 9544 7590
rect 9568 7588 9624 7590
rect 9328 6554 9384 6556
rect 9408 6554 9464 6556
rect 9488 6554 9544 6556
rect 9568 6554 9624 6556
rect 9328 6502 9374 6554
rect 9374 6502 9384 6554
rect 9408 6502 9438 6554
rect 9438 6502 9450 6554
rect 9450 6502 9464 6554
rect 9488 6502 9502 6554
rect 9502 6502 9514 6554
rect 9514 6502 9544 6554
rect 9568 6502 9578 6554
rect 9578 6502 9624 6554
rect 9328 6500 9384 6502
rect 9408 6500 9464 6502
rect 9488 6500 9544 6502
rect 9568 6500 9624 6502
rect 10414 7404 10470 7440
rect 10414 7384 10416 7404
rect 10416 7384 10468 7404
rect 10468 7384 10470 7404
rect 9328 5466 9384 5468
rect 9408 5466 9464 5468
rect 9488 5466 9544 5468
rect 9568 5466 9624 5468
rect 9328 5414 9374 5466
rect 9374 5414 9384 5466
rect 9408 5414 9438 5466
rect 9438 5414 9450 5466
rect 9450 5414 9464 5466
rect 9488 5414 9502 5466
rect 9502 5414 9514 5466
rect 9514 5414 9544 5466
rect 9568 5414 9578 5466
rect 9578 5414 9624 5466
rect 9328 5412 9384 5414
rect 9408 5412 9464 5414
rect 9488 5412 9544 5414
rect 9568 5412 9624 5414
rect 9034 4800 9090 4856
rect 8482 3304 8538 3360
rect 9328 4378 9384 4380
rect 9408 4378 9464 4380
rect 9488 4378 9544 4380
rect 9568 4378 9624 4380
rect 9328 4326 9374 4378
rect 9374 4326 9384 4378
rect 9408 4326 9438 4378
rect 9438 4326 9450 4378
rect 9450 4326 9464 4378
rect 9488 4326 9502 4378
rect 9502 4326 9514 4378
rect 9514 4326 9544 4378
rect 9568 4326 9578 4378
rect 9578 4326 9624 4378
rect 9328 4324 9384 4326
rect 9408 4324 9464 4326
rect 9488 4324 9544 4326
rect 9568 4324 9624 4326
rect 8850 3576 8906 3632
rect 9328 3290 9384 3292
rect 9408 3290 9464 3292
rect 9488 3290 9544 3292
rect 9568 3290 9624 3292
rect 9328 3238 9374 3290
rect 9374 3238 9384 3290
rect 9408 3238 9438 3290
rect 9438 3238 9450 3290
rect 9450 3238 9464 3290
rect 9488 3238 9502 3290
rect 9502 3238 9514 3290
rect 9514 3238 9544 3290
rect 9568 3238 9578 3290
rect 9578 3238 9624 3290
rect 9328 3236 9384 3238
rect 9408 3236 9464 3238
rect 9488 3236 9544 3238
rect 9568 3236 9624 3238
rect 9328 2202 9384 2204
rect 9408 2202 9464 2204
rect 9488 2202 9544 2204
rect 9568 2202 9624 2204
rect 9328 2150 9374 2202
rect 9374 2150 9384 2202
rect 9408 2150 9438 2202
rect 9438 2150 9450 2202
rect 9450 2150 9464 2202
rect 9488 2150 9502 2202
rect 9502 2150 9514 2202
rect 9514 2150 9544 2202
rect 9568 2150 9578 2202
rect 9578 2150 9624 2202
rect 9328 2148 9384 2150
rect 9408 2148 9464 2150
rect 9488 2148 9544 2150
rect 9568 2148 9624 2150
rect 12070 14764 12072 14784
rect 12072 14764 12124 14784
rect 12124 14764 12126 14784
rect 12070 14728 12126 14764
rect 12806 15408 12862 15464
rect 11610 6976 11666 7032
rect 13514 25594 13570 25596
rect 13594 25594 13650 25596
rect 13674 25594 13730 25596
rect 13754 25594 13810 25596
rect 13514 25542 13560 25594
rect 13560 25542 13570 25594
rect 13594 25542 13624 25594
rect 13624 25542 13636 25594
rect 13636 25542 13650 25594
rect 13674 25542 13688 25594
rect 13688 25542 13700 25594
rect 13700 25542 13730 25594
rect 13754 25542 13764 25594
rect 13764 25542 13810 25594
rect 13514 25540 13570 25542
rect 13594 25540 13650 25542
rect 13674 25540 13730 25542
rect 13754 25540 13810 25542
rect 13514 24506 13570 24508
rect 13594 24506 13650 24508
rect 13674 24506 13730 24508
rect 13754 24506 13810 24508
rect 13514 24454 13560 24506
rect 13560 24454 13570 24506
rect 13594 24454 13624 24506
rect 13624 24454 13636 24506
rect 13636 24454 13650 24506
rect 13674 24454 13688 24506
rect 13688 24454 13700 24506
rect 13700 24454 13730 24506
rect 13754 24454 13764 24506
rect 13764 24454 13810 24506
rect 13514 24452 13570 24454
rect 13594 24452 13650 24454
rect 13674 24452 13730 24454
rect 13754 24452 13810 24454
rect 13514 23418 13570 23420
rect 13594 23418 13650 23420
rect 13674 23418 13730 23420
rect 13754 23418 13810 23420
rect 13514 23366 13560 23418
rect 13560 23366 13570 23418
rect 13594 23366 13624 23418
rect 13624 23366 13636 23418
rect 13636 23366 13650 23418
rect 13674 23366 13688 23418
rect 13688 23366 13700 23418
rect 13700 23366 13730 23418
rect 13754 23366 13764 23418
rect 13764 23366 13810 23418
rect 13514 23364 13570 23366
rect 13594 23364 13650 23366
rect 13674 23364 13730 23366
rect 13754 23364 13810 23366
rect 13514 22330 13570 22332
rect 13594 22330 13650 22332
rect 13674 22330 13730 22332
rect 13754 22330 13810 22332
rect 13514 22278 13560 22330
rect 13560 22278 13570 22330
rect 13594 22278 13624 22330
rect 13624 22278 13636 22330
rect 13636 22278 13650 22330
rect 13674 22278 13688 22330
rect 13688 22278 13700 22330
rect 13700 22278 13730 22330
rect 13754 22278 13764 22330
rect 13764 22278 13810 22330
rect 13514 22276 13570 22278
rect 13594 22276 13650 22278
rect 13674 22276 13730 22278
rect 13754 22276 13810 22278
rect 13514 21242 13570 21244
rect 13594 21242 13650 21244
rect 13674 21242 13730 21244
rect 13754 21242 13810 21244
rect 13514 21190 13560 21242
rect 13560 21190 13570 21242
rect 13594 21190 13624 21242
rect 13624 21190 13636 21242
rect 13636 21190 13650 21242
rect 13674 21190 13688 21242
rect 13688 21190 13700 21242
rect 13700 21190 13730 21242
rect 13754 21190 13764 21242
rect 13764 21190 13810 21242
rect 13514 21188 13570 21190
rect 13594 21188 13650 21190
rect 13674 21188 13730 21190
rect 13754 21188 13810 21190
rect 13514 20154 13570 20156
rect 13594 20154 13650 20156
rect 13674 20154 13730 20156
rect 13754 20154 13810 20156
rect 13514 20102 13560 20154
rect 13560 20102 13570 20154
rect 13594 20102 13624 20154
rect 13624 20102 13636 20154
rect 13636 20102 13650 20154
rect 13674 20102 13688 20154
rect 13688 20102 13700 20154
rect 13700 20102 13730 20154
rect 13754 20102 13764 20154
rect 13764 20102 13810 20154
rect 13514 20100 13570 20102
rect 13594 20100 13650 20102
rect 13674 20100 13730 20102
rect 13754 20100 13810 20102
rect 13514 19066 13570 19068
rect 13594 19066 13650 19068
rect 13674 19066 13730 19068
rect 13754 19066 13810 19068
rect 13514 19014 13560 19066
rect 13560 19014 13570 19066
rect 13594 19014 13624 19066
rect 13624 19014 13636 19066
rect 13636 19014 13650 19066
rect 13674 19014 13688 19066
rect 13688 19014 13700 19066
rect 13700 19014 13730 19066
rect 13754 19014 13764 19066
rect 13764 19014 13810 19066
rect 13514 19012 13570 19014
rect 13594 19012 13650 19014
rect 13674 19012 13730 19014
rect 13754 19012 13810 19014
rect 13514 17978 13570 17980
rect 13594 17978 13650 17980
rect 13674 17978 13730 17980
rect 13754 17978 13810 17980
rect 13514 17926 13560 17978
rect 13560 17926 13570 17978
rect 13594 17926 13624 17978
rect 13624 17926 13636 17978
rect 13636 17926 13650 17978
rect 13674 17926 13688 17978
rect 13688 17926 13700 17978
rect 13700 17926 13730 17978
rect 13754 17926 13764 17978
rect 13764 17926 13810 17978
rect 13514 17924 13570 17926
rect 13594 17924 13650 17926
rect 13674 17924 13730 17926
rect 13754 17924 13810 17926
rect 13514 16890 13570 16892
rect 13594 16890 13650 16892
rect 13674 16890 13730 16892
rect 13754 16890 13810 16892
rect 13514 16838 13560 16890
rect 13560 16838 13570 16890
rect 13594 16838 13624 16890
rect 13624 16838 13636 16890
rect 13636 16838 13650 16890
rect 13674 16838 13688 16890
rect 13688 16838 13700 16890
rect 13700 16838 13730 16890
rect 13754 16838 13764 16890
rect 13764 16838 13810 16890
rect 13514 16836 13570 16838
rect 13594 16836 13650 16838
rect 13674 16836 13730 16838
rect 13754 16836 13810 16838
rect 13358 16632 13414 16688
rect 13082 15408 13138 15464
rect 13514 15802 13570 15804
rect 13594 15802 13650 15804
rect 13674 15802 13730 15804
rect 13754 15802 13810 15804
rect 13514 15750 13560 15802
rect 13560 15750 13570 15802
rect 13594 15750 13624 15802
rect 13624 15750 13636 15802
rect 13636 15750 13650 15802
rect 13674 15750 13688 15802
rect 13688 15750 13700 15802
rect 13700 15750 13730 15802
rect 13754 15750 13764 15802
rect 13764 15750 13810 15802
rect 13514 15748 13570 15750
rect 13594 15748 13650 15750
rect 13674 15748 13730 15750
rect 13754 15748 13810 15750
rect 13514 14714 13570 14716
rect 13594 14714 13650 14716
rect 13674 14714 13730 14716
rect 13754 14714 13810 14716
rect 13514 14662 13560 14714
rect 13560 14662 13570 14714
rect 13594 14662 13624 14714
rect 13624 14662 13636 14714
rect 13636 14662 13650 14714
rect 13674 14662 13688 14714
rect 13688 14662 13700 14714
rect 13700 14662 13730 14714
rect 13754 14662 13764 14714
rect 13764 14662 13810 14714
rect 13514 14660 13570 14662
rect 13594 14660 13650 14662
rect 13674 14660 13730 14662
rect 13754 14660 13810 14662
rect 13514 13626 13570 13628
rect 13594 13626 13650 13628
rect 13674 13626 13730 13628
rect 13754 13626 13810 13628
rect 13514 13574 13560 13626
rect 13560 13574 13570 13626
rect 13594 13574 13624 13626
rect 13624 13574 13636 13626
rect 13636 13574 13650 13626
rect 13674 13574 13688 13626
rect 13688 13574 13700 13626
rect 13700 13574 13730 13626
rect 13754 13574 13764 13626
rect 13764 13574 13810 13626
rect 13514 13572 13570 13574
rect 13594 13572 13650 13574
rect 13674 13572 13730 13574
rect 13754 13572 13810 13574
rect 13514 12538 13570 12540
rect 13594 12538 13650 12540
rect 13674 12538 13730 12540
rect 13754 12538 13810 12540
rect 13514 12486 13560 12538
rect 13560 12486 13570 12538
rect 13594 12486 13624 12538
rect 13624 12486 13636 12538
rect 13636 12486 13650 12538
rect 13674 12486 13688 12538
rect 13688 12486 13700 12538
rect 13700 12486 13730 12538
rect 13754 12486 13764 12538
rect 13764 12486 13810 12538
rect 13514 12484 13570 12486
rect 13594 12484 13650 12486
rect 13674 12484 13730 12486
rect 13754 12484 13810 12486
rect 13514 11450 13570 11452
rect 13594 11450 13650 11452
rect 13674 11450 13730 11452
rect 13754 11450 13810 11452
rect 13514 11398 13560 11450
rect 13560 11398 13570 11450
rect 13594 11398 13624 11450
rect 13624 11398 13636 11450
rect 13636 11398 13650 11450
rect 13674 11398 13688 11450
rect 13688 11398 13700 11450
rect 13700 11398 13730 11450
rect 13754 11398 13764 11450
rect 13764 11398 13810 11450
rect 13514 11396 13570 11398
rect 13594 11396 13650 11398
rect 13674 11396 13730 11398
rect 13754 11396 13810 11398
rect 13514 10362 13570 10364
rect 13594 10362 13650 10364
rect 13674 10362 13730 10364
rect 13754 10362 13810 10364
rect 13514 10310 13560 10362
rect 13560 10310 13570 10362
rect 13594 10310 13624 10362
rect 13624 10310 13636 10362
rect 13636 10310 13650 10362
rect 13674 10310 13688 10362
rect 13688 10310 13700 10362
rect 13700 10310 13730 10362
rect 13754 10310 13764 10362
rect 13764 10310 13810 10362
rect 13514 10308 13570 10310
rect 13594 10308 13650 10310
rect 13674 10308 13730 10310
rect 13754 10308 13810 10310
rect 14830 18808 14886 18864
rect 15198 15544 15254 15600
rect 15658 18264 15714 18320
rect 13514 9274 13570 9276
rect 13594 9274 13650 9276
rect 13674 9274 13730 9276
rect 13754 9274 13810 9276
rect 13514 9222 13560 9274
rect 13560 9222 13570 9274
rect 13594 9222 13624 9274
rect 13624 9222 13636 9274
rect 13636 9222 13650 9274
rect 13674 9222 13688 9274
rect 13688 9222 13700 9274
rect 13700 9222 13730 9274
rect 13754 9222 13764 9274
rect 13764 9222 13810 9274
rect 13514 9220 13570 9222
rect 13594 9220 13650 9222
rect 13674 9220 13730 9222
rect 13754 9220 13810 9222
rect 13514 8186 13570 8188
rect 13594 8186 13650 8188
rect 13674 8186 13730 8188
rect 13754 8186 13810 8188
rect 13514 8134 13560 8186
rect 13560 8134 13570 8186
rect 13594 8134 13624 8186
rect 13624 8134 13636 8186
rect 13636 8134 13650 8186
rect 13674 8134 13688 8186
rect 13688 8134 13700 8186
rect 13700 8134 13730 8186
rect 13754 8134 13764 8186
rect 13764 8134 13810 8186
rect 13514 8132 13570 8134
rect 13594 8132 13650 8134
rect 13674 8132 13730 8134
rect 13754 8132 13810 8134
rect 13514 7098 13570 7100
rect 13594 7098 13650 7100
rect 13674 7098 13730 7100
rect 13754 7098 13810 7100
rect 13514 7046 13560 7098
rect 13560 7046 13570 7098
rect 13594 7046 13624 7098
rect 13624 7046 13636 7098
rect 13636 7046 13650 7098
rect 13674 7046 13688 7098
rect 13688 7046 13700 7098
rect 13700 7046 13730 7098
rect 13754 7046 13764 7098
rect 13764 7046 13810 7098
rect 13514 7044 13570 7046
rect 13594 7044 13650 7046
rect 13674 7044 13730 7046
rect 13754 7044 13810 7046
rect 13514 6010 13570 6012
rect 13594 6010 13650 6012
rect 13674 6010 13730 6012
rect 13754 6010 13810 6012
rect 13514 5958 13560 6010
rect 13560 5958 13570 6010
rect 13594 5958 13624 6010
rect 13624 5958 13636 6010
rect 13636 5958 13650 6010
rect 13674 5958 13688 6010
rect 13688 5958 13700 6010
rect 13700 5958 13730 6010
rect 13754 5958 13764 6010
rect 13764 5958 13810 6010
rect 13514 5956 13570 5958
rect 13594 5956 13650 5958
rect 13674 5956 13730 5958
rect 13754 5956 13810 5958
rect 13514 4922 13570 4924
rect 13594 4922 13650 4924
rect 13674 4922 13730 4924
rect 13754 4922 13810 4924
rect 13514 4870 13560 4922
rect 13560 4870 13570 4922
rect 13594 4870 13624 4922
rect 13624 4870 13636 4922
rect 13636 4870 13650 4922
rect 13674 4870 13688 4922
rect 13688 4870 13700 4922
rect 13700 4870 13730 4922
rect 13754 4870 13764 4922
rect 13764 4870 13810 4922
rect 13514 4868 13570 4870
rect 13594 4868 13650 4870
rect 13674 4868 13730 4870
rect 13754 4868 13810 4870
rect 13514 3834 13570 3836
rect 13594 3834 13650 3836
rect 13674 3834 13730 3836
rect 13754 3834 13810 3836
rect 13514 3782 13560 3834
rect 13560 3782 13570 3834
rect 13594 3782 13624 3834
rect 13624 3782 13636 3834
rect 13636 3782 13650 3834
rect 13674 3782 13688 3834
rect 13688 3782 13700 3834
rect 13700 3782 13730 3834
rect 13754 3782 13764 3834
rect 13764 3782 13810 3834
rect 13514 3780 13570 3782
rect 13594 3780 13650 3782
rect 13674 3780 13730 3782
rect 13754 3780 13810 3782
rect 13514 2746 13570 2748
rect 13594 2746 13650 2748
rect 13674 2746 13730 2748
rect 13754 2746 13810 2748
rect 13514 2694 13560 2746
rect 13560 2694 13570 2746
rect 13594 2694 13624 2746
rect 13624 2694 13636 2746
rect 13636 2694 13650 2746
rect 13674 2694 13688 2746
rect 13688 2694 13700 2746
rect 13700 2694 13730 2746
rect 13754 2694 13764 2746
rect 13764 2694 13810 2746
rect 13514 2692 13570 2694
rect 13594 2692 13650 2694
rect 13674 2692 13730 2694
rect 13754 2692 13810 2694
rect 15842 18128 15898 18184
rect 17700 27226 17756 27228
rect 17780 27226 17836 27228
rect 17860 27226 17916 27228
rect 17940 27226 17996 27228
rect 17700 27174 17746 27226
rect 17746 27174 17756 27226
rect 17780 27174 17810 27226
rect 17810 27174 17822 27226
rect 17822 27174 17836 27226
rect 17860 27174 17874 27226
rect 17874 27174 17886 27226
rect 17886 27174 17916 27226
rect 17940 27174 17950 27226
rect 17950 27174 17996 27226
rect 17700 27172 17756 27174
rect 17780 27172 17836 27174
rect 17860 27172 17916 27174
rect 17940 27172 17996 27174
rect 17700 26138 17756 26140
rect 17780 26138 17836 26140
rect 17860 26138 17916 26140
rect 17940 26138 17996 26140
rect 17700 26086 17746 26138
rect 17746 26086 17756 26138
rect 17780 26086 17810 26138
rect 17810 26086 17822 26138
rect 17822 26086 17836 26138
rect 17860 26086 17874 26138
rect 17874 26086 17886 26138
rect 17886 26086 17916 26138
rect 17940 26086 17950 26138
rect 17950 26086 17996 26138
rect 17700 26084 17756 26086
rect 17780 26084 17836 26086
rect 17860 26084 17916 26086
rect 17940 26084 17996 26086
rect 16854 19660 16856 19680
rect 16856 19660 16908 19680
rect 16908 19660 16910 19680
rect 16854 19624 16910 19660
rect 17700 25050 17756 25052
rect 17780 25050 17836 25052
rect 17860 25050 17916 25052
rect 17940 25050 17996 25052
rect 17700 24998 17746 25050
rect 17746 24998 17756 25050
rect 17780 24998 17810 25050
rect 17810 24998 17822 25050
rect 17822 24998 17836 25050
rect 17860 24998 17874 25050
rect 17874 24998 17886 25050
rect 17886 24998 17916 25050
rect 17940 24998 17950 25050
rect 17950 24998 17996 25050
rect 17700 24996 17756 24998
rect 17780 24996 17836 24998
rect 17860 24996 17916 24998
rect 17940 24996 17996 24998
rect 17700 23962 17756 23964
rect 17780 23962 17836 23964
rect 17860 23962 17916 23964
rect 17940 23962 17996 23964
rect 17700 23910 17746 23962
rect 17746 23910 17756 23962
rect 17780 23910 17810 23962
rect 17810 23910 17822 23962
rect 17822 23910 17836 23962
rect 17860 23910 17874 23962
rect 17874 23910 17886 23962
rect 17886 23910 17916 23962
rect 17940 23910 17950 23962
rect 17950 23910 17996 23962
rect 17700 23908 17756 23910
rect 17780 23908 17836 23910
rect 17860 23908 17916 23910
rect 17940 23908 17996 23910
rect 17700 22874 17756 22876
rect 17780 22874 17836 22876
rect 17860 22874 17916 22876
rect 17940 22874 17996 22876
rect 17700 22822 17746 22874
rect 17746 22822 17756 22874
rect 17780 22822 17810 22874
rect 17810 22822 17822 22874
rect 17822 22822 17836 22874
rect 17860 22822 17874 22874
rect 17874 22822 17886 22874
rect 17886 22822 17916 22874
rect 17940 22822 17950 22874
rect 17950 22822 17996 22874
rect 17700 22820 17756 22822
rect 17780 22820 17836 22822
rect 17860 22820 17916 22822
rect 17940 22820 17996 22822
rect 17700 21786 17756 21788
rect 17780 21786 17836 21788
rect 17860 21786 17916 21788
rect 17940 21786 17996 21788
rect 17700 21734 17746 21786
rect 17746 21734 17756 21786
rect 17780 21734 17810 21786
rect 17810 21734 17822 21786
rect 17822 21734 17836 21786
rect 17860 21734 17874 21786
rect 17874 21734 17886 21786
rect 17886 21734 17916 21786
rect 17940 21734 17950 21786
rect 17950 21734 17996 21786
rect 17700 21732 17756 21734
rect 17780 21732 17836 21734
rect 17860 21732 17916 21734
rect 17940 21732 17996 21734
rect 17700 20698 17756 20700
rect 17780 20698 17836 20700
rect 17860 20698 17916 20700
rect 17940 20698 17996 20700
rect 17700 20646 17746 20698
rect 17746 20646 17756 20698
rect 17780 20646 17810 20698
rect 17810 20646 17822 20698
rect 17822 20646 17836 20698
rect 17860 20646 17874 20698
rect 17874 20646 17886 20698
rect 17886 20646 17916 20698
rect 17940 20646 17950 20698
rect 17950 20646 17996 20698
rect 17700 20644 17756 20646
rect 17780 20644 17836 20646
rect 17860 20644 17916 20646
rect 17940 20644 17996 20646
rect 17700 19610 17756 19612
rect 17780 19610 17836 19612
rect 17860 19610 17916 19612
rect 17940 19610 17996 19612
rect 17700 19558 17746 19610
rect 17746 19558 17756 19610
rect 17780 19558 17810 19610
rect 17810 19558 17822 19610
rect 17822 19558 17836 19610
rect 17860 19558 17874 19610
rect 17874 19558 17886 19610
rect 17886 19558 17916 19610
rect 17940 19558 17950 19610
rect 17950 19558 17996 19610
rect 17700 19556 17756 19558
rect 17780 19556 17836 19558
rect 17860 19556 17916 19558
rect 17940 19556 17996 19558
rect 17958 18708 17960 18728
rect 17960 18708 18012 18728
rect 18012 18708 18014 18728
rect 17958 18672 18014 18708
rect 17700 18522 17756 18524
rect 17780 18522 17836 18524
rect 17860 18522 17916 18524
rect 17940 18522 17996 18524
rect 17700 18470 17746 18522
rect 17746 18470 17756 18522
rect 17780 18470 17810 18522
rect 17810 18470 17822 18522
rect 17822 18470 17836 18522
rect 17860 18470 17874 18522
rect 17874 18470 17886 18522
rect 17886 18470 17916 18522
rect 17940 18470 17950 18522
rect 17950 18470 17996 18522
rect 17700 18468 17756 18470
rect 17780 18468 17836 18470
rect 17860 18468 17916 18470
rect 17940 18468 17996 18470
rect 17700 17434 17756 17436
rect 17780 17434 17836 17436
rect 17860 17434 17916 17436
rect 17940 17434 17996 17436
rect 17700 17382 17746 17434
rect 17746 17382 17756 17434
rect 17780 17382 17810 17434
rect 17810 17382 17822 17434
rect 17822 17382 17836 17434
rect 17860 17382 17874 17434
rect 17874 17382 17886 17434
rect 17886 17382 17916 17434
rect 17940 17382 17950 17434
rect 17950 17382 17996 17434
rect 17700 17380 17756 17382
rect 17780 17380 17836 17382
rect 17860 17380 17916 17382
rect 17940 17380 17996 17382
rect 17958 17176 18014 17232
rect 17700 16346 17756 16348
rect 17780 16346 17836 16348
rect 17860 16346 17916 16348
rect 17940 16346 17996 16348
rect 17700 16294 17746 16346
rect 17746 16294 17756 16346
rect 17780 16294 17810 16346
rect 17810 16294 17822 16346
rect 17822 16294 17836 16346
rect 17860 16294 17874 16346
rect 17874 16294 17886 16346
rect 17886 16294 17916 16346
rect 17940 16294 17950 16346
rect 17950 16294 17996 16346
rect 17700 16292 17756 16294
rect 17780 16292 17836 16294
rect 17860 16292 17916 16294
rect 17940 16292 17996 16294
rect 17222 13268 17224 13288
rect 17224 13268 17276 13288
rect 17276 13268 17278 13288
rect 17222 13232 17278 13268
rect 17700 15258 17756 15260
rect 17780 15258 17836 15260
rect 17860 15258 17916 15260
rect 17940 15258 17996 15260
rect 17700 15206 17746 15258
rect 17746 15206 17756 15258
rect 17780 15206 17810 15258
rect 17810 15206 17822 15258
rect 17822 15206 17836 15258
rect 17860 15206 17874 15258
rect 17874 15206 17886 15258
rect 17886 15206 17916 15258
rect 17940 15206 17950 15258
rect 17950 15206 17996 15258
rect 17700 15204 17756 15206
rect 17780 15204 17836 15206
rect 17860 15204 17916 15206
rect 17940 15204 17996 15206
rect 18418 17176 18474 17232
rect 17700 14170 17756 14172
rect 17780 14170 17836 14172
rect 17860 14170 17916 14172
rect 17940 14170 17996 14172
rect 17700 14118 17746 14170
rect 17746 14118 17756 14170
rect 17780 14118 17810 14170
rect 17810 14118 17822 14170
rect 17822 14118 17836 14170
rect 17860 14118 17874 14170
rect 17874 14118 17886 14170
rect 17886 14118 17916 14170
rect 17940 14118 17950 14170
rect 17950 14118 17996 14170
rect 17700 14116 17756 14118
rect 17780 14116 17836 14118
rect 17860 14116 17916 14118
rect 17940 14116 17996 14118
rect 17700 13082 17756 13084
rect 17780 13082 17836 13084
rect 17860 13082 17916 13084
rect 17940 13082 17996 13084
rect 17700 13030 17746 13082
rect 17746 13030 17756 13082
rect 17780 13030 17810 13082
rect 17810 13030 17822 13082
rect 17822 13030 17836 13082
rect 17860 13030 17874 13082
rect 17874 13030 17886 13082
rect 17886 13030 17916 13082
rect 17940 13030 17950 13082
rect 17950 13030 17996 13082
rect 17700 13028 17756 13030
rect 17780 13028 17836 13030
rect 17860 13028 17916 13030
rect 17940 13028 17996 13030
rect 17700 11994 17756 11996
rect 17780 11994 17836 11996
rect 17860 11994 17916 11996
rect 17940 11994 17996 11996
rect 17700 11942 17746 11994
rect 17746 11942 17756 11994
rect 17780 11942 17810 11994
rect 17810 11942 17822 11994
rect 17822 11942 17836 11994
rect 17860 11942 17874 11994
rect 17874 11942 17886 11994
rect 17886 11942 17916 11994
rect 17940 11942 17950 11994
rect 17950 11942 17996 11994
rect 17700 11940 17756 11942
rect 17780 11940 17836 11942
rect 17860 11940 17916 11942
rect 17940 11940 17996 11942
rect 17700 10906 17756 10908
rect 17780 10906 17836 10908
rect 17860 10906 17916 10908
rect 17940 10906 17996 10908
rect 17700 10854 17746 10906
rect 17746 10854 17756 10906
rect 17780 10854 17810 10906
rect 17810 10854 17822 10906
rect 17822 10854 17836 10906
rect 17860 10854 17874 10906
rect 17874 10854 17886 10906
rect 17886 10854 17916 10906
rect 17940 10854 17950 10906
rect 17950 10854 17996 10906
rect 17700 10852 17756 10854
rect 17780 10852 17836 10854
rect 17860 10852 17916 10854
rect 17940 10852 17996 10854
rect 17700 9818 17756 9820
rect 17780 9818 17836 9820
rect 17860 9818 17916 9820
rect 17940 9818 17996 9820
rect 17700 9766 17746 9818
rect 17746 9766 17756 9818
rect 17780 9766 17810 9818
rect 17810 9766 17822 9818
rect 17822 9766 17836 9818
rect 17860 9766 17874 9818
rect 17874 9766 17886 9818
rect 17886 9766 17916 9818
rect 17940 9766 17950 9818
rect 17950 9766 17996 9818
rect 17700 9764 17756 9766
rect 17780 9764 17836 9766
rect 17860 9764 17916 9766
rect 17940 9764 17996 9766
rect 19430 21392 19486 21448
rect 18786 18284 18842 18320
rect 18786 18264 18788 18284
rect 18788 18264 18840 18284
rect 18840 18264 18842 18284
rect 18786 18148 18842 18184
rect 18786 18128 18788 18148
rect 18788 18128 18840 18148
rect 18840 18128 18842 18148
rect 19246 18672 19302 18728
rect 19154 16632 19210 16688
rect 20166 21428 20168 21448
rect 20168 21428 20220 21448
rect 20220 21428 20222 21448
rect 20166 21392 20222 21428
rect 20626 17484 20628 17504
rect 20628 17484 20680 17504
rect 20680 17484 20682 17504
rect 17700 8730 17756 8732
rect 17780 8730 17836 8732
rect 17860 8730 17916 8732
rect 17940 8730 17996 8732
rect 17700 8678 17746 8730
rect 17746 8678 17756 8730
rect 17780 8678 17810 8730
rect 17810 8678 17822 8730
rect 17822 8678 17836 8730
rect 17860 8678 17874 8730
rect 17874 8678 17886 8730
rect 17886 8678 17916 8730
rect 17940 8678 17950 8730
rect 17950 8678 17996 8730
rect 17700 8676 17756 8678
rect 17780 8676 17836 8678
rect 17860 8676 17916 8678
rect 17940 8676 17996 8678
rect 17700 7642 17756 7644
rect 17780 7642 17836 7644
rect 17860 7642 17916 7644
rect 17940 7642 17996 7644
rect 17700 7590 17746 7642
rect 17746 7590 17756 7642
rect 17780 7590 17810 7642
rect 17810 7590 17822 7642
rect 17822 7590 17836 7642
rect 17860 7590 17874 7642
rect 17874 7590 17886 7642
rect 17886 7590 17916 7642
rect 17940 7590 17950 7642
rect 17950 7590 17996 7642
rect 17700 7588 17756 7590
rect 17780 7588 17836 7590
rect 17860 7588 17916 7590
rect 17940 7588 17996 7590
rect 17700 6554 17756 6556
rect 17780 6554 17836 6556
rect 17860 6554 17916 6556
rect 17940 6554 17996 6556
rect 17700 6502 17746 6554
rect 17746 6502 17756 6554
rect 17780 6502 17810 6554
rect 17810 6502 17822 6554
rect 17822 6502 17836 6554
rect 17860 6502 17874 6554
rect 17874 6502 17886 6554
rect 17886 6502 17916 6554
rect 17940 6502 17950 6554
rect 17950 6502 17996 6554
rect 17700 6500 17756 6502
rect 17780 6500 17836 6502
rect 17860 6500 17916 6502
rect 17940 6500 17996 6502
rect 17700 5466 17756 5468
rect 17780 5466 17836 5468
rect 17860 5466 17916 5468
rect 17940 5466 17996 5468
rect 17700 5414 17746 5466
rect 17746 5414 17756 5466
rect 17780 5414 17810 5466
rect 17810 5414 17822 5466
rect 17822 5414 17836 5466
rect 17860 5414 17874 5466
rect 17874 5414 17886 5466
rect 17886 5414 17916 5466
rect 17940 5414 17950 5466
rect 17950 5414 17996 5466
rect 17700 5412 17756 5414
rect 17780 5412 17836 5414
rect 17860 5412 17916 5414
rect 17940 5412 17996 5414
rect 16302 3984 16358 4040
rect 17700 4378 17756 4380
rect 17780 4378 17836 4380
rect 17860 4378 17916 4380
rect 17940 4378 17996 4380
rect 17700 4326 17746 4378
rect 17746 4326 17756 4378
rect 17780 4326 17810 4378
rect 17810 4326 17822 4378
rect 17822 4326 17836 4378
rect 17860 4326 17874 4378
rect 17874 4326 17886 4378
rect 17886 4326 17916 4378
rect 17940 4326 17950 4378
rect 17950 4326 17996 4378
rect 17700 4324 17756 4326
rect 17780 4324 17836 4326
rect 17860 4324 17916 4326
rect 17940 4324 17996 4326
rect 18878 3984 18934 4040
rect 17700 3290 17756 3292
rect 17780 3290 17836 3292
rect 17860 3290 17916 3292
rect 17940 3290 17996 3292
rect 17700 3238 17746 3290
rect 17746 3238 17756 3290
rect 17780 3238 17810 3290
rect 17810 3238 17822 3290
rect 17822 3238 17836 3290
rect 17860 3238 17874 3290
rect 17874 3238 17886 3290
rect 17886 3238 17916 3290
rect 17940 3238 17950 3290
rect 17950 3238 17996 3290
rect 17700 3236 17756 3238
rect 17780 3236 17836 3238
rect 17860 3236 17916 3238
rect 17940 3236 17996 3238
rect 17700 2202 17756 2204
rect 17780 2202 17836 2204
rect 17860 2202 17916 2204
rect 17940 2202 17996 2204
rect 17700 2150 17746 2202
rect 17746 2150 17756 2202
rect 17780 2150 17810 2202
rect 17810 2150 17822 2202
rect 17822 2150 17836 2202
rect 17860 2150 17874 2202
rect 17874 2150 17886 2202
rect 17886 2150 17916 2202
rect 17940 2150 17950 2202
rect 17950 2150 17996 2202
rect 17700 2148 17756 2150
rect 17780 2148 17836 2150
rect 17860 2148 17916 2150
rect 17940 2148 17996 2150
rect 20626 17448 20682 17484
rect 21270 21428 21272 21448
rect 21272 21428 21324 21448
rect 21324 21428 21326 21448
rect 21270 21392 21326 21428
rect 26330 28756 26386 28792
rect 21886 26682 21942 26684
rect 21966 26682 22022 26684
rect 22046 26682 22102 26684
rect 22126 26682 22182 26684
rect 21886 26630 21932 26682
rect 21932 26630 21942 26682
rect 21966 26630 21996 26682
rect 21996 26630 22008 26682
rect 22008 26630 22022 26682
rect 22046 26630 22060 26682
rect 22060 26630 22072 26682
rect 22072 26630 22102 26682
rect 22126 26630 22136 26682
rect 22136 26630 22182 26682
rect 21886 26628 21942 26630
rect 21966 26628 22022 26630
rect 22046 26628 22102 26630
rect 22126 26628 22182 26630
rect 26330 28736 26332 28756
rect 26332 28736 26384 28756
rect 26384 28736 26386 28756
rect 21886 25594 21942 25596
rect 21966 25594 22022 25596
rect 22046 25594 22102 25596
rect 22126 25594 22182 25596
rect 21886 25542 21932 25594
rect 21932 25542 21942 25594
rect 21966 25542 21996 25594
rect 21996 25542 22008 25594
rect 22008 25542 22022 25594
rect 22046 25542 22060 25594
rect 22060 25542 22072 25594
rect 22072 25542 22102 25594
rect 22126 25542 22136 25594
rect 22136 25542 22182 25594
rect 21886 25540 21942 25542
rect 21966 25540 22022 25542
rect 22046 25540 22102 25542
rect 22126 25540 22182 25542
rect 26330 24540 26386 24576
rect 26330 24520 26332 24540
rect 26332 24520 26384 24540
rect 26384 24520 26386 24540
rect 21886 24506 21942 24508
rect 21966 24506 22022 24508
rect 22046 24506 22102 24508
rect 22126 24506 22182 24508
rect 21886 24454 21932 24506
rect 21932 24454 21942 24506
rect 21966 24454 21996 24506
rect 21996 24454 22008 24506
rect 22008 24454 22022 24506
rect 22046 24454 22060 24506
rect 22060 24454 22072 24506
rect 22072 24454 22102 24506
rect 22126 24454 22136 24506
rect 22136 24454 22182 24506
rect 21886 24452 21942 24454
rect 21966 24452 22022 24454
rect 22046 24452 22102 24454
rect 22126 24452 22182 24454
rect 21886 23418 21942 23420
rect 21966 23418 22022 23420
rect 22046 23418 22102 23420
rect 22126 23418 22182 23420
rect 21886 23366 21932 23418
rect 21932 23366 21942 23418
rect 21966 23366 21996 23418
rect 21996 23366 22008 23418
rect 22008 23366 22022 23418
rect 22046 23366 22060 23418
rect 22060 23366 22072 23418
rect 22072 23366 22102 23418
rect 22126 23366 22136 23418
rect 22136 23366 22182 23418
rect 21886 23364 21942 23366
rect 21966 23364 22022 23366
rect 22046 23364 22102 23366
rect 22126 23364 22182 23366
rect 21886 22330 21942 22332
rect 21966 22330 22022 22332
rect 22046 22330 22102 22332
rect 22126 22330 22182 22332
rect 21886 22278 21932 22330
rect 21932 22278 21942 22330
rect 21966 22278 21996 22330
rect 21996 22278 22008 22330
rect 22008 22278 22022 22330
rect 22046 22278 22060 22330
rect 22060 22278 22072 22330
rect 22072 22278 22102 22330
rect 22126 22278 22136 22330
rect 22136 22278 22182 22330
rect 21886 22276 21942 22278
rect 21966 22276 22022 22278
rect 22046 22276 22102 22278
rect 22126 22276 22182 22278
rect 25134 23180 25190 23216
rect 25134 23160 25136 23180
rect 25136 23160 25188 23180
rect 25188 23160 25190 23180
rect 22466 22072 22522 22128
rect 22282 21800 22338 21856
rect 21886 21242 21942 21244
rect 21966 21242 22022 21244
rect 22046 21242 22102 21244
rect 22126 21242 22182 21244
rect 21886 21190 21932 21242
rect 21932 21190 21942 21242
rect 21966 21190 21996 21242
rect 21996 21190 22008 21242
rect 22008 21190 22022 21242
rect 22046 21190 22060 21242
rect 22060 21190 22072 21242
rect 22072 21190 22102 21242
rect 22126 21190 22136 21242
rect 22136 21190 22182 21242
rect 21886 21188 21942 21190
rect 21966 21188 22022 21190
rect 22046 21188 22102 21190
rect 22126 21188 22182 21190
rect 21886 20154 21942 20156
rect 21966 20154 22022 20156
rect 22046 20154 22102 20156
rect 22126 20154 22182 20156
rect 21886 20102 21932 20154
rect 21932 20102 21942 20154
rect 21966 20102 21996 20154
rect 21996 20102 22008 20154
rect 22008 20102 22022 20154
rect 22046 20102 22060 20154
rect 22060 20102 22072 20154
rect 22072 20102 22102 20154
rect 22126 20102 22136 20154
rect 22136 20102 22182 20154
rect 21886 20100 21942 20102
rect 21966 20100 22022 20102
rect 22046 20100 22102 20102
rect 22126 20100 22182 20102
rect 21886 19066 21942 19068
rect 21966 19066 22022 19068
rect 22046 19066 22102 19068
rect 22126 19066 22182 19068
rect 21886 19014 21932 19066
rect 21932 19014 21942 19066
rect 21966 19014 21996 19066
rect 21996 19014 22008 19066
rect 22008 19014 22022 19066
rect 22046 19014 22060 19066
rect 22060 19014 22072 19066
rect 22072 19014 22102 19066
rect 22126 19014 22136 19066
rect 22136 19014 22182 19066
rect 21886 19012 21942 19014
rect 21966 19012 22022 19014
rect 22046 19012 22102 19014
rect 22126 19012 22182 19014
rect 21638 18264 21694 18320
rect 22190 18148 22246 18184
rect 22190 18128 22192 18148
rect 22192 18128 22244 18148
rect 22244 18128 22246 18148
rect 21886 17978 21942 17980
rect 21966 17978 22022 17980
rect 22046 17978 22102 17980
rect 22126 17978 22182 17980
rect 21886 17926 21932 17978
rect 21932 17926 21942 17978
rect 21966 17926 21996 17978
rect 21996 17926 22008 17978
rect 22008 17926 22022 17978
rect 22046 17926 22060 17978
rect 22060 17926 22072 17978
rect 22072 17926 22102 17978
rect 22126 17926 22136 17978
rect 22136 17926 22182 17978
rect 21886 17924 21942 17926
rect 21966 17924 22022 17926
rect 22046 17924 22102 17926
rect 22126 17924 22182 17926
rect 21454 17448 21510 17504
rect 22282 17484 22284 17504
rect 22284 17484 22336 17504
rect 22336 17484 22338 17504
rect 22282 17448 22338 17484
rect 21886 16890 21942 16892
rect 21966 16890 22022 16892
rect 22046 16890 22102 16892
rect 22126 16890 22182 16892
rect 21886 16838 21932 16890
rect 21932 16838 21942 16890
rect 21966 16838 21996 16890
rect 21996 16838 22008 16890
rect 22008 16838 22022 16890
rect 22046 16838 22060 16890
rect 22060 16838 22072 16890
rect 22072 16838 22102 16890
rect 22126 16838 22136 16890
rect 22136 16838 22182 16890
rect 21886 16836 21942 16838
rect 21966 16836 22022 16838
rect 22046 16836 22102 16838
rect 22126 16836 22182 16838
rect 22282 16088 22338 16144
rect 21886 15802 21942 15804
rect 21966 15802 22022 15804
rect 22046 15802 22102 15804
rect 22126 15802 22182 15804
rect 21886 15750 21932 15802
rect 21932 15750 21942 15802
rect 21966 15750 21996 15802
rect 21996 15750 22008 15802
rect 22008 15750 22022 15802
rect 22046 15750 22060 15802
rect 22060 15750 22072 15802
rect 22072 15750 22102 15802
rect 22126 15750 22136 15802
rect 22136 15750 22182 15802
rect 21886 15748 21942 15750
rect 21966 15748 22022 15750
rect 22046 15748 22102 15750
rect 22126 15748 22182 15750
rect 21886 14714 21942 14716
rect 21966 14714 22022 14716
rect 22046 14714 22102 14716
rect 22126 14714 22182 14716
rect 21886 14662 21932 14714
rect 21932 14662 21942 14714
rect 21966 14662 21996 14714
rect 21996 14662 22008 14714
rect 22008 14662 22022 14714
rect 22046 14662 22060 14714
rect 22060 14662 22072 14714
rect 22072 14662 22102 14714
rect 22126 14662 22136 14714
rect 22136 14662 22182 14714
rect 21886 14660 21942 14662
rect 21966 14660 22022 14662
rect 22046 14660 22102 14662
rect 22126 14660 22182 14662
rect 21886 13626 21942 13628
rect 21966 13626 22022 13628
rect 22046 13626 22102 13628
rect 22126 13626 22182 13628
rect 21886 13574 21932 13626
rect 21932 13574 21942 13626
rect 21966 13574 21996 13626
rect 21996 13574 22008 13626
rect 22008 13574 22022 13626
rect 22046 13574 22060 13626
rect 22060 13574 22072 13626
rect 22072 13574 22102 13626
rect 22126 13574 22136 13626
rect 22136 13574 22182 13626
rect 21886 13572 21942 13574
rect 21966 13572 22022 13574
rect 22046 13572 22102 13574
rect 22126 13572 22182 13574
rect 22558 18944 22614 19000
rect 22742 18300 22744 18320
rect 22744 18300 22796 18320
rect 22796 18300 22798 18320
rect 22742 18264 22798 18300
rect 21886 12538 21942 12540
rect 21966 12538 22022 12540
rect 22046 12538 22102 12540
rect 22126 12538 22182 12540
rect 21886 12486 21932 12538
rect 21932 12486 21942 12538
rect 21966 12486 21996 12538
rect 21996 12486 22008 12538
rect 22008 12486 22022 12538
rect 22046 12486 22060 12538
rect 22060 12486 22072 12538
rect 22072 12486 22102 12538
rect 22126 12486 22136 12538
rect 22136 12486 22182 12538
rect 21886 12484 21942 12486
rect 21966 12484 22022 12486
rect 22046 12484 22102 12486
rect 22126 12484 22182 12486
rect 22466 12316 22468 12336
rect 22468 12316 22520 12336
rect 22520 12316 22522 12336
rect 22466 12280 22522 12316
rect 21886 11450 21942 11452
rect 21966 11450 22022 11452
rect 22046 11450 22102 11452
rect 22126 11450 22182 11452
rect 21886 11398 21932 11450
rect 21932 11398 21942 11450
rect 21966 11398 21996 11450
rect 21996 11398 22008 11450
rect 22008 11398 22022 11450
rect 22046 11398 22060 11450
rect 22060 11398 22072 11450
rect 22072 11398 22102 11450
rect 22126 11398 22136 11450
rect 22136 11398 22182 11450
rect 21886 11396 21942 11398
rect 21966 11396 22022 11398
rect 22046 11396 22102 11398
rect 22126 11396 22182 11398
rect 23018 18264 23074 18320
rect 23110 18128 23166 18184
rect 23478 18128 23534 18184
rect 25778 17584 25834 17640
rect 21886 10362 21942 10364
rect 21966 10362 22022 10364
rect 22046 10362 22102 10364
rect 22126 10362 22182 10364
rect 21886 10310 21932 10362
rect 21932 10310 21942 10362
rect 21966 10310 21996 10362
rect 21996 10310 22008 10362
rect 22008 10310 22022 10362
rect 22046 10310 22060 10362
rect 22060 10310 22072 10362
rect 22072 10310 22102 10362
rect 22126 10310 22136 10362
rect 22136 10310 22182 10362
rect 21886 10308 21942 10310
rect 21966 10308 22022 10310
rect 22046 10308 22102 10310
rect 22126 10308 22182 10310
rect 21886 9274 21942 9276
rect 21966 9274 22022 9276
rect 22046 9274 22102 9276
rect 22126 9274 22182 9276
rect 21886 9222 21932 9274
rect 21932 9222 21942 9274
rect 21966 9222 21996 9274
rect 21996 9222 22008 9274
rect 22008 9222 22022 9274
rect 22046 9222 22060 9274
rect 22060 9222 22072 9274
rect 22072 9222 22102 9274
rect 22126 9222 22136 9274
rect 22136 9222 22182 9274
rect 21886 9220 21942 9222
rect 21966 9220 22022 9222
rect 22046 9220 22102 9222
rect 22126 9220 22182 9222
rect 21886 8186 21942 8188
rect 21966 8186 22022 8188
rect 22046 8186 22102 8188
rect 22126 8186 22182 8188
rect 21886 8134 21932 8186
rect 21932 8134 21942 8186
rect 21966 8134 21996 8186
rect 21996 8134 22008 8186
rect 22008 8134 22022 8186
rect 22046 8134 22060 8186
rect 22060 8134 22072 8186
rect 22072 8134 22102 8186
rect 22126 8134 22136 8186
rect 22136 8134 22182 8186
rect 21886 8132 21942 8134
rect 21966 8132 22022 8134
rect 22046 8132 22102 8134
rect 22126 8132 22182 8134
rect 21886 7098 21942 7100
rect 21966 7098 22022 7100
rect 22046 7098 22102 7100
rect 22126 7098 22182 7100
rect 21886 7046 21932 7098
rect 21932 7046 21942 7098
rect 21966 7046 21996 7098
rect 21996 7046 22008 7098
rect 22008 7046 22022 7098
rect 22046 7046 22060 7098
rect 22060 7046 22072 7098
rect 22072 7046 22102 7098
rect 22126 7046 22136 7098
rect 22136 7046 22182 7098
rect 21886 7044 21942 7046
rect 21966 7044 22022 7046
rect 22046 7044 22102 7046
rect 22126 7044 22182 7046
rect 22098 6332 22100 6352
rect 22100 6332 22152 6352
rect 22152 6332 22154 6352
rect 22098 6296 22154 6332
rect 21886 6010 21942 6012
rect 21966 6010 22022 6012
rect 22046 6010 22102 6012
rect 22126 6010 22182 6012
rect 21886 5958 21932 6010
rect 21932 5958 21942 6010
rect 21966 5958 21996 6010
rect 21996 5958 22008 6010
rect 22008 5958 22022 6010
rect 22046 5958 22060 6010
rect 22060 5958 22072 6010
rect 22072 5958 22102 6010
rect 22126 5958 22136 6010
rect 22136 5958 22182 6010
rect 21886 5956 21942 5958
rect 21966 5956 22022 5958
rect 22046 5956 22102 5958
rect 22126 5956 22182 5958
rect 21886 4922 21942 4924
rect 21966 4922 22022 4924
rect 22046 4922 22102 4924
rect 22126 4922 22182 4924
rect 21886 4870 21932 4922
rect 21932 4870 21942 4922
rect 21966 4870 21996 4922
rect 21996 4870 22008 4922
rect 22008 4870 22022 4922
rect 22046 4870 22060 4922
rect 22060 4870 22072 4922
rect 22072 4870 22102 4922
rect 22126 4870 22136 4922
rect 22136 4870 22182 4922
rect 21886 4868 21942 4870
rect 21966 4868 22022 4870
rect 22046 4868 22102 4870
rect 22126 4868 22182 4870
rect 26330 14728 26386 14784
rect 23386 13368 23442 13424
rect 25134 11872 25190 11928
rect 22742 9152 22798 9208
rect 21886 3834 21942 3836
rect 21966 3834 22022 3836
rect 22046 3834 22102 3836
rect 22126 3834 22182 3836
rect 21886 3782 21932 3834
rect 21932 3782 21942 3834
rect 21966 3782 21996 3834
rect 21996 3782 22008 3834
rect 22008 3782 22022 3834
rect 22046 3782 22060 3834
rect 22060 3782 22072 3834
rect 22072 3782 22102 3834
rect 22126 3782 22136 3834
rect 22136 3782 22182 3834
rect 21886 3780 21942 3782
rect 21966 3780 22022 3782
rect 22046 3780 22102 3782
rect 22126 3780 22182 3782
rect 22098 3440 22154 3496
rect 21886 2746 21942 2748
rect 21966 2746 22022 2748
rect 22046 2746 22102 2748
rect 22126 2746 22182 2748
rect 21886 2694 21932 2746
rect 21932 2694 21942 2746
rect 21966 2694 21996 2746
rect 21996 2694 22008 2746
rect 22008 2694 22022 2746
rect 22046 2694 22060 2746
rect 22060 2694 22072 2746
rect 22072 2694 22102 2746
rect 22126 2694 22136 2746
rect 22136 2694 22182 2746
rect 21886 2692 21942 2694
rect 21966 2692 22022 2694
rect 22046 2692 22102 2694
rect 22126 2692 22182 2694
rect 22098 720 22154 776
<< metal3 >>
rect 26325 28794 26391 28797
rect 26595 28794 27395 28824
rect 26325 28792 27395 28794
rect 26325 28736 26330 28792
rect 26386 28736 27395 28792
rect 26325 28734 27395 28736
rect 26325 28731 26391 28734
rect 26595 28704 27395 28734
rect 0 28432 800 28552
rect 26595 27344 27395 27464
rect 9316 27232 9636 27233
rect 9316 27168 9324 27232
rect 9388 27168 9404 27232
rect 9468 27168 9484 27232
rect 9548 27168 9564 27232
rect 9628 27168 9636 27232
rect 9316 27167 9636 27168
rect 17688 27232 18008 27233
rect 17688 27168 17696 27232
rect 17760 27168 17776 27232
rect 17840 27168 17856 27232
rect 17920 27168 17936 27232
rect 18000 27168 18008 27232
rect 17688 27167 18008 27168
rect 5130 26688 5450 26689
rect 0 26528 800 26648
rect 5130 26624 5138 26688
rect 5202 26624 5218 26688
rect 5282 26624 5298 26688
rect 5362 26624 5378 26688
rect 5442 26624 5450 26688
rect 5130 26623 5450 26624
rect 13502 26688 13822 26689
rect 13502 26624 13510 26688
rect 13574 26624 13590 26688
rect 13654 26624 13670 26688
rect 13734 26624 13750 26688
rect 13814 26624 13822 26688
rect 13502 26623 13822 26624
rect 21874 26688 22194 26689
rect 21874 26624 21882 26688
rect 21946 26624 21962 26688
rect 22026 26624 22042 26688
rect 22106 26624 22122 26688
rect 22186 26624 22194 26688
rect 21874 26623 22194 26624
rect 9316 26144 9636 26145
rect 9316 26080 9324 26144
rect 9388 26080 9404 26144
rect 9468 26080 9484 26144
rect 9548 26080 9564 26144
rect 9628 26080 9636 26144
rect 9316 26079 9636 26080
rect 17688 26144 18008 26145
rect 17688 26080 17696 26144
rect 17760 26080 17776 26144
rect 17840 26080 17856 26144
rect 17920 26080 17936 26144
rect 18000 26080 18008 26144
rect 17688 26079 18008 26080
rect 26595 25984 27395 26104
rect 5130 25600 5450 25601
rect 5130 25536 5138 25600
rect 5202 25536 5218 25600
rect 5282 25536 5298 25600
rect 5362 25536 5378 25600
rect 5442 25536 5450 25600
rect 5130 25535 5450 25536
rect 13502 25600 13822 25601
rect 13502 25536 13510 25600
rect 13574 25536 13590 25600
rect 13654 25536 13670 25600
rect 13734 25536 13750 25600
rect 13814 25536 13822 25600
rect 13502 25535 13822 25536
rect 21874 25600 22194 25601
rect 21874 25536 21882 25600
rect 21946 25536 21962 25600
rect 22026 25536 22042 25600
rect 22106 25536 22122 25600
rect 22186 25536 22194 25600
rect 21874 25535 22194 25536
rect 9316 25056 9636 25057
rect 9316 24992 9324 25056
rect 9388 24992 9404 25056
rect 9468 24992 9484 25056
rect 9548 24992 9564 25056
rect 9628 24992 9636 25056
rect 9316 24991 9636 24992
rect 17688 25056 18008 25057
rect 17688 24992 17696 25056
rect 17760 24992 17776 25056
rect 17840 24992 17856 25056
rect 17920 24992 17936 25056
rect 18000 24992 18008 25056
rect 17688 24991 18008 24992
rect 0 24760 800 24880
rect 26325 24578 26391 24581
rect 26595 24578 27395 24608
rect 26325 24576 27395 24578
rect 26325 24520 26330 24576
rect 26386 24520 27395 24576
rect 26325 24518 27395 24520
rect 26325 24515 26391 24518
rect 5130 24512 5450 24513
rect 5130 24448 5138 24512
rect 5202 24448 5218 24512
rect 5282 24448 5298 24512
rect 5362 24448 5378 24512
rect 5442 24448 5450 24512
rect 5130 24447 5450 24448
rect 13502 24512 13822 24513
rect 13502 24448 13510 24512
rect 13574 24448 13590 24512
rect 13654 24448 13670 24512
rect 13734 24448 13750 24512
rect 13814 24448 13822 24512
rect 13502 24447 13822 24448
rect 21874 24512 22194 24513
rect 21874 24448 21882 24512
rect 21946 24448 21962 24512
rect 22026 24448 22042 24512
rect 22106 24448 22122 24512
rect 22186 24448 22194 24512
rect 26595 24488 27395 24518
rect 21874 24447 22194 24448
rect 9316 23968 9636 23969
rect 9316 23904 9324 23968
rect 9388 23904 9404 23968
rect 9468 23904 9484 23968
rect 9548 23904 9564 23968
rect 9628 23904 9636 23968
rect 9316 23903 9636 23904
rect 17688 23968 18008 23969
rect 17688 23904 17696 23968
rect 17760 23904 17776 23968
rect 17840 23904 17856 23968
rect 17920 23904 17936 23968
rect 18000 23904 18008 23968
rect 17688 23903 18008 23904
rect 5130 23424 5450 23425
rect 5130 23360 5138 23424
rect 5202 23360 5218 23424
rect 5282 23360 5298 23424
rect 5362 23360 5378 23424
rect 5442 23360 5450 23424
rect 5130 23359 5450 23360
rect 13502 23424 13822 23425
rect 13502 23360 13510 23424
rect 13574 23360 13590 23424
rect 13654 23360 13670 23424
rect 13734 23360 13750 23424
rect 13814 23360 13822 23424
rect 13502 23359 13822 23360
rect 21874 23424 22194 23425
rect 21874 23360 21882 23424
rect 21946 23360 21962 23424
rect 22026 23360 22042 23424
rect 22106 23360 22122 23424
rect 22186 23360 22194 23424
rect 21874 23359 22194 23360
rect 25129 23218 25195 23221
rect 26595 23218 27395 23248
rect 25129 23216 27395 23218
rect 25129 23160 25134 23216
rect 25190 23160 27395 23216
rect 25129 23158 27395 23160
rect 25129 23155 25195 23158
rect 26595 23128 27395 23158
rect 0 22856 800 22976
rect 9316 22880 9636 22881
rect 9316 22816 9324 22880
rect 9388 22816 9404 22880
rect 9468 22816 9484 22880
rect 9548 22816 9564 22880
rect 9628 22816 9636 22880
rect 9316 22815 9636 22816
rect 17688 22880 18008 22881
rect 17688 22816 17696 22880
rect 17760 22816 17776 22880
rect 17840 22816 17856 22880
rect 17920 22816 17936 22880
rect 18000 22816 18008 22880
rect 17688 22815 18008 22816
rect 5130 22336 5450 22337
rect 5130 22272 5138 22336
rect 5202 22272 5218 22336
rect 5282 22272 5298 22336
rect 5362 22272 5378 22336
rect 5442 22272 5450 22336
rect 5130 22271 5450 22272
rect 13502 22336 13822 22337
rect 13502 22272 13510 22336
rect 13574 22272 13590 22336
rect 13654 22272 13670 22336
rect 13734 22272 13750 22336
rect 13814 22272 13822 22336
rect 13502 22271 13822 22272
rect 21874 22336 22194 22337
rect 21874 22272 21882 22336
rect 21946 22272 21962 22336
rect 22026 22272 22042 22336
rect 22106 22272 22122 22336
rect 22186 22272 22194 22336
rect 21874 22271 22194 22272
rect 22461 22132 22527 22133
rect 22461 22128 22508 22132
rect 22572 22130 22578 22132
rect 22461 22072 22466 22128
rect 22461 22068 22508 22072
rect 22572 22070 22618 22130
rect 22572 22068 22578 22070
rect 22461 22067 22527 22068
rect 22277 21858 22343 21861
rect 26595 21858 27395 21888
rect 22277 21856 27395 21858
rect 22277 21800 22282 21856
rect 22338 21800 27395 21856
rect 22277 21798 27395 21800
rect 22277 21795 22343 21798
rect 9316 21792 9636 21793
rect 9316 21728 9324 21792
rect 9388 21728 9404 21792
rect 9468 21728 9484 21792
rect 9548 21728 9564 21792
rect 9628 21728 9636 21792
rect 9316 21727 9636 21728
rect 17688 21792 18008 21793
rect 17688 21728 17696 21792
rect 17760 21728 17776 21792
rect 17840 21728 17856 21792
rect 17920 21728 17936 21792
rect 18000 21728 18008 21792
rect 26595 21768 27395 21798
rect 17688 21727 18008 21728
rect 19425 21450 19491 21453
rect 20161 21450 20227 21453
rect 21265 21450 21331 21453
rect 19425 21448 21331 21450
rect 19425 21392 19430 21448
rect 19486 21392 20166 21448
rect 20222 21392 21270 21448
rect 21326 21392 21331 21448
rect 19425 21390 21331 21392
rect 19425 21387 19491 21390
rect 20161 21387 20227 21390
rect 21265 21387 21331 21390
rect 5130 21248 5450 21249
rect 0 21088 800 21208
rect 5130 21184 5138 21248
rect 5202 21184 5218 21248
rect 5282 21184 5298 21248
rect 5362 21184 5378 21248
rect 5442 21184 5450 21248
rect 5130 21183 5450 21184
rect 13502 21248 13822 21249
rect 13502 21184 13510 21248
rect 13574 21184 13590 21248
rect 13654 21184 13670 21248
rect 13734 21184 13750 21248
rect 13814 21184 13822 21248
rect 13502 21183 13822 21184
rect 21874 21248 22194 21249
rect 21874 21184 21882 21248
rect 21946 21184 21962 21248
rect 22026 21184 22042 21248
rect 22106 21184 22122 21248
rect 22186 21184 22194 21248
rect 21874 21183 22194 21184
rect 9316 20704 9636 20705
rect 9316 20640 9324 20704
rect 9388 20640 9404 20704
rect 9468 20640 9484 20704
rect 9548 20640 9564 20704
rect 9628 20640 9636 20704
rect 9316 20639 9636 20640
rect 17688 20704 18008 20705
rect 17688 20640 17696 20704
rect 17760 20640 17776 20704
rect 17840 20640 17856 20704
rect 17920 20640 17936 20704
rect 18000 20640 18008 20704
rect 17688 20639 18008 20640
rect 5257 20362 5323 20365
rect 9857 20362 9923 20365
rect 5257 20360 9923 20362
rect 5257 20304 5262 20360
rect 5318 20304 9862 20360
rect 9918 20304 9923 20360
rect 5257 20302 9923 20304
rect 5257 20299 5323 20302
rect 9857 20299 9923 20302
rect 26595 20272 27395 20392
rect 5130 20160 5450 20161
rect 5130 20096 5138 20160
rect 5202 20096 5218 20160
rect 5282 20096 5298 20160
rect 5362 20096 5378 20160
rect 5442 20096 5450 20160
rect 5130 20095 5450 20096
rect 13502 20160 13822 20161
rect 13502 20096 13510 20160
rect 13574 20096 13590 20160
rect 13654 20096 13670 20160
rect 13734 20096 13750 20160
rect 13814 20096 13822 20160
rect 13502 20095 13822 20096
rect 21874 20160 22194 20161
rect 21874 20096 21882 20160
rect 21946 20096 21962 20160
rect 22026 20096 22042 20160
rect 22106 20096 22122 20160
rect 22186 20096 22194 20160
rect 21874 20095 22194 20096
rect 16849 19682 16915 19685
rect 16982 19682 16988 19684
rect 16849 19680 16988 19682
rect 16849 19624 16854 19680
rect 16910 19624 16988 19680
rect 16849 19622 16988 19624
rect 16849 19619 16915 19622
rect 16982 19620 16988 19622
rect 17052 19620 17058 19684
rect 9316 19616 9636 19617
rect 9316 19552 9324 19616
rect 9388 19552 9404 19616
rect 9468 19552 9484 19616
rect 9548 19552 9564 19616
rect 9628 19552 9636 19616
rect 9316 19551 9636 19552
rect 17688 19616 18008 19617
rect 17688 19552 17696 19616
rect 17760 19552 17776 19616
rect 17840 19552 17856 19616
rect 17920 19552 17936 19616
rect 18000 19552 18008 19616
rect 17688 19551 18008 19552
rect 7281 19410 7347 19413
rect 7741 19410 7807 19413
rect 7281 19408 7807 19410
rect 7281 19352 7286 19408
rect 7342 19352 7746 19408
rect 7802 19352 7807 19408
rect 7281 19350 7807 19352
rect 7281 19347 7347 19350
rect 7741 19347 7807 19350
rect 0 19184 800 19304
rect 5130 19072 5450 19073
rect 5130 19008 5138 19072
rect 5202 19008 5218 19072
rect 5282 19008 5298 19072
rect 5362 19008 5378 19072
rect 5442 19008 5450 19072
rect 5130 19007 5450 19008
rect 13502 19072 13822 19073
rect 13502 19008 13510 19072
rect 13574 19008 13590 19072
rect 13654 19008 13670 19072
rect 13734 19008 13750 19072
rect 13814 19008 13822 19072
rect 13502 19007 13822 19008
rect 21874 19072 22194 19073
rect 21874 19008 21882 19072
rect 21946 19008 21962 19072
rect 22026 19008 22042 19072
rect 22106 19008 22122 19072
rect 22186 19008 22194 19072
rect 21874 19007 22194 19008
rect 22553 19002 22619 19005
rect 26595 19002 27395 19032
rect 22553 19000 27395 19002
rect 22553 18944 22558 19000
rect 22614 18944 27395 19000
rect 22553 18942 27395 18944
rect 22553 18939 22619 18942
rect 26595 18912 27395 18942
rect 10133 18866 10199 18869
rect 14825 18866 14891 18869
rect 10133 18864 14891 18866
rect 10133 18808 10138 18864
rect 10194 18808 14830 18864
rect 14886 18808 14891 18864
rect 10133 18806 14891 18808
rect 10133 18803 10199 18806
rect 14825 18803 14891 18806
rect 8937 18732 9003 18733
rect 8886 18668 8892 18732
rect 8956 18730 9003 18732
rect 17953 18730 18019 18733
rect 19241 18730 19307 18733
rect 8956 18728 9048 18730
rect 8998 18672 9048 18728
rect 8956 18670 9048 18672
rect 17953 18728 19307 18730
rect 17953 18672 17958 18728
rect 18014 18672 19246 18728
rect 19302 18672 19307 18728
rect 17953 18670 19307 18672
rect 8956 18668 9003 18670
rect 8937 18667 9003 18668
rect 17953 18667 18019 18670
rect 19241 18667 19307 18670
rect 9316 18528 9636 18529
rect 9316 18464 9324 18528
rect 9388 18464 9404 18528
rect 9468 18464 9484 18528
rect 9548 18464 9564 18528
rect 9628 18464 9636 18528
rect 9316 18463 9636 18464
rect 17688 18528 18008 18529
rect 17688 18464 17696 18528
rect 17760 18464 17776 18528
rect 17840 18464 17856 18528
rect 17920 18464 17936 18528
rect 18000 18464 18008 18528
rect 17688 18463 18008 18464
rect 15653 18322 15719 18325
rect 18781 18322 18847 18325
rect 15653 18320 18847 18322
rect 15653 18264 15658 18320
rect 15714 18264 18786 18320
rect 18842 18264 18847 18320
rect 15653 18262 18847 18264
rect 15653 18259 15719 18262
rect 18781 18259 18847 18262
rect 21633 18322 21699 18325
rect 22737 18322 22803 18325
rect 23013 18322 23079 18325
rect 21633 18320 23079 18322
rect 21633 18264 21638 18320
rect 21694 18264 22742 18320
rect 22798 18264 23018 18320
rect 23074 18264 23079 18320
rect 21633 18262 23079 18264
rect 21633 18259 21699 18262
rect 22737 18259 22803 18262
rect 23013 18259 23079 18262
rect 15837 18186 15903 18189
rect 18781 18186 18847 18189
rect 15837 18184 18847 18186
rect 15837 18128 15842 18184
rect 15898 18128 18786 18184
rect 18842 18128 18847 18184
rect 15837 18126 18847 18128
rect 15837 18123 15903 18126
rect 18781 18123 18847 18126
rect 22185 18186 22251 18189
rect 23105 18186 23171 18189
rect 23473 18186 23539 18189
rect 22185 18184 23539 18186
rect 22185 18128 22190 18184
rect 22246 18128 23110 18184
rect 23166 18128 23478 18184
rect 23534 18128 23539 18184
rect 22185 18126 23539 18128
rect 22185 18123 22251 18126
rect 23105 18123 23171 18126
rect 23473 18123 23539 18126
rect 5130 17984 5450 17985
rect 5130 17920 5138 17984
rect 5202 17920 5218 17984
rect 5282 17920 5298 17984
rect 5362 17920 5378 17984
rect 5442 17920 5450 17984
rect 5130 17919 5450 17920
rect 13502 17984 13822 17985
rect 13502 17920 13510 17984
rect 13574 17920 13590 17984
rect 13654 17920 13670 17984
rect 13734 17920 13750 17984
rect 13814 17920 13822 17984
rect 13502 17919 13822 17920
rect 21874 17984 22194 17985
rect 21874 17920 21882 17984
rect 21946 17920 21962 17984
rect 22026 17920 22042 17984
rect 22106 17920 22122 17984
rect 22186 17920 22194 17984
rect 21874 17919 22194 17920
rect 25773 17642 25839 17645
rect 26595 17642 27395 17672
rect 25773 17640 27395 17642
rect 25773 17584 25778 17640
rect 25834 17584 27395 17640
rect 25773 17582 27395 17584
rect 25773 17579 25839 17582
rect 26595 17552 27395 17582
rect 0 17506 800 17536
rect 4061 17506 4127 17509
rect 0 17504 4127 17506
rect 0 17448 4066 17504
rect 4122 17448 4127 17504
rect 0 17446 4127 17448
rect 0 17416 800 17446
rect 4061 17443 4127 17446
rect 20621 17506 20687 17509
rect 21449 17506 21515 17509
rect 22277 17506 22343 17509
rect 20621 17504 22343 17506
rect 20621 17448 20626 17504
rect 20682 17448 21454 17504
rect 21510 17448 22282 17504
rect 22338 17448 22343 17504
rect 20621 17446 22343 17448
rect 20621 17443 20687 17446
rect 21449 17443 21515 17446
rect 22277 17443 22343 17446
rect 9316 17440 9636 17441
rect 9316 17376 9324 17440
rect 9388 17376 9404 17440
rect 9468 17376 9484 17440
rect 9548 17376 9564 17440
rect 9628 17376 9636 17440
rect 9316 17375 9636 17376
rect 17688 17440 18008 17441
rect 17688 17376 17696 17440
rect 17760 17376 17776 17440
rect 17840 17376 17856 17440
rect 17920 17376 17936 17440
rect 18000 17376 18008 17440
rect 17688 17375 18008 17376
rect 6177 17234 6243 17237
rect 7741 17234 7807 17237
rect 6177 17232 7807 17234
rect 6177 17176 6182 17232
rect 6238 17176 7746 17232
rect 7802 17176 7807 17232
rect 6177 17174 7807 17176
rect 6177 17171 6243 17174
rect 7741 17171 7807 17174
rect 8661 17234 8727 17237
rect 9489 17234 9555 17237
rect 8661 17232 9555 17234
rect 8661 17176 8666 17232
rect 8722 17176 9494 17232
rect 9550 17176 9555 17232
rect 8661 17174 9555 17176
rect 8661 17171 8727 17174
rect 9489 17171 9555 17174
rect 17953 17234 18019 17237
rect 18413 17234 18479 17237
rect 17953 17232 18479 17234
rect 17953 17176 17958 17232
rect 18014 17176 18418 17232
rect 18474 17176 18479 17232
rect 17953 17174 18479 17176
rect 17953 17171 18019 17174
rect 18413 17171 18479 17174
rect 5130 16896 5450 16897
rect 5130 16832 5138 16896
rect 5202 16832 5218 16896
rect 5282 16832 5298 16896
rect 5362 16832 5378 16896
rect 5442 16832 5450 16896
rect 5130 16831 5450 16832
rect 13502 16896 13822 16897
rect 13502 16832 13510 16896
rect 13574 16832 13590 16896
rect 13654 16832 13670 16896
rect 13734 16832 13750 16896
rect 13814 16832 13822 16896
rect 13502 16831 13822 16832
rect 21874 16896 22194 16897
rect 21874 16832 21882 16896
rect 21946 16832 21962 16896
rect 22026 16832 22042 16896
rect 22106 16832 22122 16896
rect 22186 16832 22194 16896
rect 21874 16831 22194 16832
rect 9397 16690 9463 16693
rect 9581 16690 9647 16693
rect 9397 16688 9647 16690
rect 9397 16632 9402 16688
rect 9458 16632 9586 16688
rect 9642 16632 9647 16688
rect 9397 16630 9647 16632
rect 9397 16627 9463 16630
rect 9581 16627 9647 16630
rect 13353 16690 13419 16693
rect 19149 16690 19215 16693
rect 13353 16688 19215 16690
rect 13353 16632 13358 16688
rect 13414 16632 19154 16688
rect 19210 16632 19215 16688
rect 13353 16630 19215 16632
rect 13353 16627 13419 16630
rect 19149 16627 19215 16630
rect 9316 16352 9636 16353
rect 9316 16288 9324 16352
rect 9388 16288 9404 16352
rect 9468 16288 9484 16352
rect 9548 16288 9564 16352
rect 9628 16288 9636 16352
rect 9316 16287 9636 16288
rect 17688 16352 18008 16353
rect 17688 16288 17696 16352
rect 17760 16288 17776 16352
rect 17840 16288 17856 16352
rect 17920 16288 17936 16352
rect 18000 16288 18008 16352
rect 17688 16287 18008 16288
rect 8293 16146 8359 16149
rect 9581 16146 9647 16149
rect 8293 16144 9647 16146
rect 8293 16088 8298 16144
rect 8354 16088 9586 16144
rect 9642 16088 9647 16144
rect 8293 16086 9647 16088
rect 8293 16083 8359 16086
rect 9581 16083 9647 16086
rect 22277 16146 22343 16149
rect 26595 16146 27395 16176
rect 22277 16144 27395 16146
rect 22277 16088 22282 16144
rect 22338 16088 27395 16144
rect 22277 16086 27395 16088
rect 22277 16083 22343 16086
rect 26595 16056 27395 16086
rect 5130 15808 5450 15809
rect 5130 15744 5138 15808
rect 5202 15744 5218 15808
rect 5282 15744 5298 15808
rect 5362 15744 5378 15808
rect 5442 15744 5450 15808
rect 5130 15743 5450 15744
rect 13502 15808 13822 15809
rect 13502 15744 13510 15808
rect 13574 15744 13590 15808
rect 13654 15744 13670 15808
rect 13734 15744 13750 15808
rect 13814 15744 13822 15808
rect 13502 15743 13822 15744
rect 21874 15808 22194 15809
rect 21874 15744 21882 15808
rect 21946 15744 21962 15808
rect 22026 15744 22042 15808
rect 22106 15744 22122 15808
rect 22186 15744 22194 15808
rect 21874 15743 22194 15744
rect 0 15602 800 15632
rect 15193 15602 15259 15605
rect 0 15600 15259 15602
rect 0 15544 15198 15600
rect 15254 15544 15259 15600
rect 0 15542 15259 15544
rect 0 15512 800 15542
rect 15193 15539 15259 15542
rect 12801 15466 12867 15469
rect 13077 15466 13143 15469
rect 12801 15464 13143 15466
rect 12801 15408 12806 15464
rect 12862 15408 13082 15464
rect 13138 15408 13143 15464
rect 12801 15406 13143 15408
rect 12801 15403 12867 15406
rect 13077 15403 13143 15406
rect 9316 15264 9636 15265
rect 9316 15200 9324 15264
rect 9388 15200 9404 15264
rect 9468 15200 9484 15264
rect 9548 15200 9564 15264
rect 9628 15200 9636 15264
rect 9316 15199 9636 15200
rect 17688 15264 18008 15265
rect 17688 15200 17696 15264
rect 17760 15200 17776 15264
rect 17840 15200 17856 15264
rect 17920 15200 17936 15264
rect 18000 15200 18008 15264
rect 17688 15199 18008 15200
rect 9070 14724 9076 14788
rect 9140 14786 9146 14788
rect 9489 14786 9555 14789
rect 12065 14788 12131 14789
rect 9140 14784 9555 14786
rect 9140 14728 9494 14784
rect 9550 14728 9555 14784
rect 9140 14726 9555 14728
rect 9140 14724 9146 14726
rect 9489 14723 9555 14726
rect 12014 14724 12020 14788
rect 12084 14786 12131 14788
rect 26325 14786 26391 14789
rect 26595 14786 27395 14816
rect 12084 14784 12176 14786
rect 12126 14728 12176 14784
rect 12084 14726 12176 14728
rect 26325 14784 27395 14786
rect 26325 14728 26330 14784
rect 26386 14728 27395 14784
rect 26325 14726 27395 14728
rect 12084 14724 12131 14726
rect 12065 14723 12131 14724
rect 26325 14723 26391 14726
rect 5130 14720 5450 14721
rect 5130 14656 5138 14720
rect 5202 14656 5218 14720
rect 5282 14656 5298 14720
rect 5362 14656 5378 14720
rect 5442 14656 5450 14720
rect 5130 14655 5450 14656
rect 13502 14720 13822 14721
rect 13502 14656 13510 14720
rect 13574 14656 13590 14720
rect 13654 14656 13670 14720
rect 13734 14656 13750 14720
rect 13814 14656 13822 14720
rect 13502 14655 13822 14656
rect 21874 14720 22194 14721
rect 21874 14656 21882 14720
rect 21946 14656 21962 14720
rect 22026 14656 22042 14720
rect 22106 14656 22122 14720
rect 22186 14656 22194 14720
rect 26595 14696 27395 14726
rect 21874 14655 22194 14656
rect 9316 14176 9636 14177
rect 9316 14112 9324 14176
rect 9388 14112 9404 14176
rect 9468 14112 9484 14176
rect 9548 14112 9564 14176
rect 9628 14112 9636 14176
rect 9316 14111 9636 14112
rect 17688 14176 18008 14177
rect 17688 14112 17696 14176
rect 17760 14112 17776 14176
rect 17840 14112 17856 14176
rect 17920 14112 17936 14176
rect 18000 14112 18008 14176
rect 17688 14111 18008 14112
rect 6821 14106 6887 14109
rect 8017 14106 8083 14109
rect 6821 14104 8083 14106
rect 6821 14048 6826 14104
rect 6882 14048 8022 14104
rect 8078 14048 8083 14104
rect 6821 14046 8083 14048
rect 6821 14043 6887 14046
rect 8017 14043 8083 14046
rect 7373 13970 7439 13973
rect 8661 13970 8727 13973
rect 9305 13970 9371 13973
rect 7373 13968 9371 13970
rect 7373 13912 7378 13968
rect 7434 13912 8666 13968
rect 8722 13912 9310 13968
rect 9366 13912 9371 13968
rect 7373 13910 9371 13912
rect 7373 13907 7439 13910
rect 8661 13907 8727 13910
rect 9305 13907 9371 13910
rect 8293 13834 8359 13837
rect 4846 13832 8359 13834
rect 4846 13776 8298 13832
rect 8354 13776 8359 13832
rect 4846 13774 8359 13776
rect 0 13698 800 13728
rect 4846 13698 4906 13774
rect 8293 13771 8359 13774
rect 0 13638 4906 13698
rect 0 13608 800 13638
rect 5130 13632 5450 13633
rect 5130 13568 5138 13632
rect 5202 13568 5218 13632
rect 5282 13568 5298 13632
rect 5362 13568 5378 13632
rect 5442 13568 5450 13632
rect 5130 13567 5450 13568
rect 13502 13632 13822 13633
rect 13502 13568 13510 13632
rect 13574 13568 13590 13632
rect 13654 13568 13670 13632
rect 13734 13568 13750 13632
rect 13814 13568 13822 13632
rect 13502 13567 13822 13568
rect 21874 13632 22194 13633
rect 21874 13568 21882 13632
rect 21946 13568 21962 13632
rect 22026 13568 22042 13632
rect 22106 13568 22122 13632
rect 22186 13568 22194 13632
rect 21874 13567 22194 13568
rect 23381 13426 23447 13429
rect 26595 13426 27395 13456
rect 23381 13424 27395 13426
rect 23381 13368 23386 13424
rect 23442 13368 27395 13424
rect 23381 13366 27395 13368
rect 23381 13363 23447 13366
rect 26595 13336 27395 13366
rect 16798 13228 16804 13292
rect 16868 13290 16874 13292
rect 17217 13290 17283 13293
rect 16868 13288 17283 13290
rect 16868 13232 17222 13288
rect 17278 13232 17283 13288
rect 16868 13230 17283 13232
rect 16868 13228 16874 13230
rect 17217 13227 17283 13230
rect 9316 13088 9636 13089
rect 9316 13024 9324 13088
rect 9388 13024 9404 13088
rect 9468 13024 9484 13088
rect 9548 13024 9564 13088
rect 9628 13024 9636 13088
rect 9316 13023 9636 13024
rect 17688 13088 18008 13089
rect 17688 13024 17696 13088
rect 17760 13024 17776 13088
rect 17840 13024 17856 13088
rect 17920 13024 17936 13088
rect 18000 13024 18008 13088
rect 17688 13023 18008 13024
rect 2957 12882 3023 12885
rect 3509 12882 3575 12885
rect 5165 12882 5231 12885
rect 5533 12882 5599 12885
rect 2957 12880 5599 12882
rect 2957 12824 2962 12880
rect 3018 12824 3514 12880
rect 3570 12824 5170 12880
rect 5226 12824 5538 12880
rect 5594 12824 5599 12880
rect 2957 12822 5599 12824
rect 2957 12819 3023 12822
rect 3509 12819 3575 12822
rect 5165 12819 5231 12822
rect 5533 12819 5599 12822
rect 8385 12882 8451 12885
rect 8702 12882 8708 12884
rect 8385 12880 8708 12882
rect 8385 12824 8390 12880
rect 8446 12824 8708 12880
rect 8385 12822 8708 12824
rect 8385 12819 8451 12822
rect 8702 12820 8708 12822
rect 8772 12882 8778 12884
rect 9949 12882 10015 12885
rect 8772 12880 10015 12882
rect 8772 12824 9954 12880
rect 10010 12824 10015 12880
rect 8772 12822 10015 12824
rect 8772 12820 8778 12822
rect 9949 12819 10015 12822
rect 5130 12544 5450 12545
rect 5130 12480 5138 12544
rect 5202 12480 5218 12544
rect 5282 12480 5298 12544
rect 5362 12480 5378 12544
rect 5442 12480 5450 12544
rect 5130 12479 5450 12480
rect 13502 12544 13822 12545
rect 13502 12480 13510 12544
rect 13574 12480 13590 12544
rect 13654 12480 13670 12544
rect 13734 12480 13750 12544
rect 13814 12480 13822 12544
rect 13502 12479 13822 12480
rect 21874 12544 22194 12545
rect 21874 12480 21882 12544
rect 21946 12480 21962 12544
rect 22026 12480 22042 12544
rect 22106 12480 22122 12544
rect 22186 12480 22194 12544
rect 21874 12479 22194 12480
rect 22461 12340 22527 12341
rect 22461 12338 22508 12340
rect 22416 12336 22508 12338
rect 22416 12280 22466 12336
rect 22416 12278 22508 12280
rect 22461 12276 22508 12278
rect 22572 12276 22578 12340
rect 22461 12275 22527 12276
rect 9316 12000 9636 12001
rect 0 11930 800 11960
rect 9316 11936 9324 12000
rect 9388 11936 9404 12000
rect 9468 11936 9484 12000
rect 9548 11936 9564 12000
rect 9628 11936 9636 12000
rect 9316 11935 9636 11936
rect 17688 12000 18008 12001
rect 17688 11936 17696 12000
rect 17760 11936 17776 12000
rect 17840 11936 17856 12000
rect 17920 11936 17936 12000
rect 18000 11936 18008 12000
rect 17688 11935 18008 11936
rect 4981 11930 5047 11933
rect 0 11928 5047 11930
rect 0 11872 4986 11928
rect 5042 11872 5047 11928
rect 0 11870 5047 11872
rect 0 11840 800 11870
rect 4981 11867 5047 11870
rect 25129 11930 25195 11933
rect 26595 11930 27395 11960
rect 25129 11928 27395 11930
rect 25129 11872 25134 11928
rect 25190 11872 27395 11928
rect 25129 11870 27395 11872
rect 25129 11867 25195 11870
rect 26595 11840 27395 11870
rect 5165 11794 5231 11797
rect 9581 11794 9647 11797
rect 5165 11792 9647 11794
rect 5165 11736 5170 11792
rect 5226 11736 9586 11792
rect 9642 11736 9647 11792
rect 5165 11734 9647 11736
rect 5165 11731 5231 11734
rect 9581 11731 9647 11734
rect 5130 11456 5450 11457
rect 5130 11392 5138 11456
rect 5202 11392 5218 11456
rect 5282 11392 5298 11456
rect 5362 11392 5378 11456
rect 5442 11392 5450 11456
rect 5130 11391 5450 11392
rect 13502 11456 13822 11457
rect 13502 11392 13510 11456
rect 13574 11392 13590 11456
rect 13654 11392 13670 11456
rect 13734 11392 13750 11456
rect 13814 11392 13822 11456
rect 13502 11391 13822 11392
rect 21874 11456 22194 11457
rect 21874 11392 21882 11456
rect 21946 11392 21962 11456
rect 22026 11392 22042 11456
rect 22106 11392 22122 11456
rect 22186 11392 22194 11456
rect 21874 11391 22194 11392
rect 9316 10912 9636 10913
rect 9316 10848 9324 10912
rect 9388 10848 9404 10912
rect 9468 10848 9484 10912
rect 9548 10848 9564 10912
rect 9628 10848 9636 10912
rect 9316 10847 9636 10848
rect 17688 10912 18008 10913
rect 17688 10848 17696 10912
rect 17760 10848 17776 10912
rect 17840 10848 17856 10912
rect 17920 10848 17936 10912
rect 18000 10848 18008 10912
rect 17688 10847 18008 10848
rect 26595 10480 27395 10600
rect 5130 10368 5450 10369
rect 5130 10304 5138 10368
rect 5202 10304 5218 10368
rect 5282 10304 5298 10368
rect 5362 10304 5378 10368
rect 5442 10304 5450 10368
rect 5130 10303 5450 10304
rect 13502 10368 13822 10369
rect 13502 10304 13510 10368
rect 13574 10304 13590 10368
rect 13654 10304 13670 10368
rect 13734 10304 13750 10368
rect 13814 10304 13822 10368
rect 13502 10303 13822 10304
rect 21874 10368 22194 10369
rect 21874 10304 21882 10368
rect 21946 10304 21962 10368
rect 22026 10304 22042 10368
rect 22106 10304 22122 10368
rect 22186 10304 22194 10368
rect 21874 10303 22194 10304
rect 0 9936 800 10056
rect 9316 9824 9636 9825
rect 9316 9760 9324 9824
rect 9388 9760 9404 9824
rect 9468 9760 9484 9824
rect 9548 9760 9564 9824
rect 9628 9760 9636 9824
rect 9316 9759 9636 9760
rect 17688 9824 18008 9825
rect 17688 9760 17696 9824
rect 17760 9760 17776 9824
rect 17840 9760 17856 9824
rect 17920 9760 17936 9824
rect 18000 9760 18008 9824
rect 17688 9759 18008 9760
rect 5130 9280 5450 9281
rect 5130 9216 5138 9280
rect 5202 9216 5218 9280
rect 5282 9216 5298 9280
rect 5362 9216 5378 9280
rect 5442 9216 5450 9280
rect 5130 9215 5450 9216
rect 13502 9280 13822 9281
rect 13502 9216 13510 9280
rect 13574 9216 13590 9280
rect 13654 9216 13670 9280
rect 13734 9216 13750 9280
rect 13814 9216 13822 9280
rect 13502 9215 13822 9216
rect 21874 9280 22194 9281
rect 21874 9216 21882 9280
rect 21946 9216 21962 9280
rect 22026 9216 22042 9280
rect 22106 9216 22122 9280
rect 22186 9216 22194 9280
rect 21874 9215 22194 9216
rect 22737 9210 22803 9213
rect 26595 9210 27395 9240
rect 22737 9208 27395 9210
rect 22737 9152 22742 9208
rect 22798 9152 27395 9208
rect 22737 9150 27395 9152
rect 22737 9147 22803 9150
rect 26595 9120 27395 9150
rect 9316 8736 9636 8737
rect 9316 8672 9324 8736
rect 9388 8672 9404 8736
rect 9468 8672 9484 8736
rect 9548 8672 9564 8736
rect 9628 8672 9636 8736
rect 9316 8671 9636 8672
rect 17688 8736 18008 8737
rect 17688 8672 17696 8736
rect 17760 8672 17776 8736
rect 17840 8672 17856 8736
rect 17920 8672 17936 8736
rect 18000 8672 18008 8736
rect 17688 8671 18008 8672
rect 0 8258 800 8288
rect 3969 8258 4035 8261
rect 0 8256 4035 8258
rect 0 8200 3974 8256
rect 4030 8200 4035 8256
rect 0 8198 4035 8200
rect 0 8168 800 8198
rect 3969 8195 4035 8198
rect 5130 8192 5450 8193
rect 5130 8128 5138 8192
rect 5202 8128 5218 8192
rect 5282 8128 5298 8192
rect 5362 8128 5378 8192
rect 5442 8128 5450 8192
rect 5130 8127 5450 8128
rect 13502 8192 13822 8193
rect 13502 8128 13510 8192
rect 13574 8128 13590 8192
rect 13654 8128 13670 8192
rect 13734 8128 13750 8192
rect 13814 8128 13822 8192
rect 13502 8127 13822 8128
rect 21874 8192 22194 8193
rect 21874 8128 21882 8192
rect 21946 8128 21962 8192
rect 22026 8128 22042 8192
rect 22106 8128 22122 8192
rect 22186 8128 22194 8192
rect 21874 8127 22194 8128
rect 8661 7986 8727 7989
rect 9581 7986 9647 7989
rect 8661 7984 9647 7986
rect 8661 7928 8666 7984
rect 8722 7928 9586 7984
rect 9642 7928 9647 7984
rect 8661 7926 9647 7928
rect 8661 7923 8727 7926
rect 9581 7923 9647 7926
rect 9316 7648 9636 7649
rect 9316 7584 9324 7648
rect 9388 7584 9404 7648
rect 9468 7584 9484 7648
rect 9548 7584 9564 7648
rect 9628 7584 9636 7648
rect 9316 7583 9636 7584
rect 17688 7648 18008 7649
rect 17688 7584 17696 7648
rect 17760 7584 17776 7648
rect 17840 7584 17856 7648
rect 17920 7584 17936 7648
rect 18000 7584 18008 7648
rect 26595 7624 27395 7744
rect 17688 7583 18008 7584
rect 9029 7442 9095 7445
rect 10409 7442 10475 7445
rect 9029 7440 10475 7442
rect 9029 7384 9034 7440
rect 9090 7384 10414 7440
rect 10470 7384 10475 7440
rect 9029 7382 10475 7384
rect 9029 7379 9095 7382
rect 10409 7379 10475 7382
rect 5130 7104 5450 7105
rect 5130 7040 5138 7104
rect 5202 7040 5218 7104
rect 5282 7040 5298 7104
rect 5362 7040 5378 7104
rect 5442 7040 5450 7104
rect 5130 7039 5450 7040
rect 13502 7104 13822 7105
rect 13502 7040 13510 7104
rect 13574 7040 13590 7104
rect 13654 7040 13670 7104
rect 13734 7040 13750 7104
rect 13814 7040 13822 7104
rect 13502 7039 13822 7040
rect 21874 7104 22194 7105
rect 21874 7040 21882 7104
rect 21946 7040 21962 7104
rect 22026 7040 22042 7104
rect 22106 7040 22122 7104
rect 22186 7040 22194 7104
rect 21874 7039 22194 7040
rect 11094 6972 11100 7036
rect 11164 7034 11170 7036
rect 11605 7034 11671 7037
rect 11164 7032 11671 7034
rect 11164 6976 11610 7032
rect 11666 6976 11671 7032
rect 11164 6974 11671 6976
rect 11164 6972 11170 6974
rect 11605 6971 11671 6974
rect 8201 6898 8267 6901
rect 614 6896 8267 6898
rect 614 6840 8206 6896
rect 8262 6840 8267 6896
rect 614 6838 8267 6840
rect 614 6626 674 6838
rect 8201 6835 8267 6838
rect 614 6566 858 6626
rect 798 6384 858 6566
rect 9316 6560 9636 6561
rect 9316 6496 9324 6560
rect 9388 6496 9404 6560
rect 9468 6496 9484 6560
rect 9548 6496 9564 6560
rect 9628 6496 9636 6560
rect 9316 6495 9636 6496
rect 17688 6560 18008 6561
rect 17688 6496 17696 6560
rect 17760 6496 17776 6560
rect 17840 6496 17856 6560
rect 17920 6496 17936 6560
rect 18000 6496 18008 6560
rect 17688 6495 18008 6496
rect 0 6294 858 6384
rect 4981 6354 5047 6357
rect 6085 6354 6151 6357
rect 8753 6354 8819 6357
rect 4981 6352 8819 6354
rect 4981 6296 4986 6352
rect 5042 6296 6090 6352
rect 6146 6296 8758 6352
rect 8814 6296 8819 6352
rect 4981 6294 8819 6296
rect 0 6264 800 6294
rect 4981 6291 5047 6294
rect 6085 6291 6151 6294
rect 8753 6291 8819 6294
rect 22093 6354 22159 6357
rect 26595 6354 27395 6384
rect 22093 6352 27395 6354
rect 22093 6296 22098 6352
rect 22154 6296 27395 6352
rect 22093 6294 27395 6296
rect 22093 6291 22159 6294
rect 26595 6264 27395 6294
rect 5130 6016 5450 6017
rect 5130 5952 5138 6016
rect 5202 5952 5218 6016
rect 5282 5952 5298 6016
rect 5362 5952 5378 6016
rect 5442 5952 5450 6016
rect 5130 5951 5450 5952
rect 13502 6016 13822 6017
rect 13502 5952 13510 6016
rect 13574 5952 13590 6016
rect 13654 5952 13670 6016
rect 13734 5952 13750 6016
rect 13814 5952 13822 6016
rect 13502 5951 13822 5952
rect 21874 6016 22194 6017
rect 21874 5952 21882 6016
rect 21946 5952 21962 6016
rect 22026 5952 22042 6016
rect 22106 5952 22122 6016
rect 22186 5952 22194 6016
rect 21874 5951 22194 5952
rect 9316 5472 9636 5473
rect 9316 5408 9324 5472
rect 9388 5408 9404 5472
rect 9468 5408 9484 5472
rect 9548 5408 9564 5472
rect 9628 5408 9636 5472
rect 9316 5407 9636 5408
rect 17688 5472 18008 5473
rect 17688 5408 17696 5472
rect 17760 5408 17776 5472
rect 17840 5408 17856 5472
rect 17920 5408 17936 5472
rect 18000 5408 18008 5472
rect 17688 5407 18008 5408
rect 6545 5402 6611 5405
rect 7189 5402 7255 5405
rect 6545 5400 7255 5402
rect 6545 5344 6550 5400
rect 6606 5344 7194 5400
rect 7250 5344 7255 5400
rect 6545 5342 7255 5344
rect 6545 5339 6611 5342
rect 7189 5339 7255 5342
rect 7833 5266 7899 5269
rect 8017 5266 8083 5269
rect 7833 5264 8083 5266
rect 7833 5208 7838 5264
rect 7894 5208 8022 5264
rect 8078 5208 8083 5264
rect 7833 5206 8083 5208
rect 7833 5203 7899 5206
rect 8017 5203 8083 5206
rect 6637 5130 6703 5133
rect 8845 5130 8911 5133
rect 6637 5128 8911 5130
rect 6637 5072 6642 5128
rect 6698 5072 8850 5128
rect 8906 5072 8911 5128
rect 6637 5070 8911 5072
rect 6637 5067 6703 5070
rect 8845 5067 8911 5070
rect 5130 4928 5450 4929
rect 5130 4864 5138 4928
rect 5202 4864 5218 4928
rect 5282 4864 5298 4928
rect 5362 4864 5378 4928
rect 5442 4864 5450 4928
rect 5130 4863 5450 4864
rect 13502 4928 13822 4929
rect 13502 4864 13510 4928
rect 13574 4864 13590 4928
rect 13654 4864 13670 4928
rect 13734 4864 13750 4928
rect 13814 4864 13822 4928
rect 13502 4863 13822 4864
rect 21874 4928 22194 4929
rect 21874 4864 21882 4928
rect 21946 4864 21962 4928
rect 22026 4864 22042 4928
rect 22106 4864 22122 4928
rect 22186 4864 22194 4928
rect 26595 4904 27395 5024
rect 21874 4863 22194 4864
rect 7465 4858 7531 4861
rect 9029 4858 9095 4861
rect 11094 4858 11100 4860
rect 7465 4856 11100 4858
rect 7465 4800 7470 4856
rect 7526 4800 9034 4856
rect 9090 4800 11100 4856
rect 7465 4798 11100 4800
rect 7465 4795 7531 4798
rect 9029 4795 9095 4798
rect 11094 4796 11100 4798
rect 11164 4796 11170 4860
rect 0 4586 800 4616
rect 9070 4586 9076 4588
rect 0 4526 9076 4586
rect 0 4496 800 4526
rect 9070 4524 9076 4526
rect 9140 4524 9146 4588
rect 9316 4384 9636 4385
rect 9316 4320 9324 4384
rect 9388 4320 9404 4384
rect 9468 4320 9484 4384
rect 9548 4320 9564 4384
rect 9628 4320 9636 4384
rect 9316 4319 9636 4320
rect 17688 4384 18008 4385
rect 17688 4320 17696 4384
rect 17760 4320 17776 4384
rect 17840 4320 17856 4384
rect 17920 4320 17936 4384
rect 18000 4320 18008 4384
rect 17688 4319 18008 4320
rect 16297 4042 16363 4045
rect 16798 4042 16804 4044
rect 16297 4040 16804 4042
rect 16297 3984 16302 4040
rect 16358 3984 16804 4040
rect 16297 3982 16804 3984
rect 16297 3979 16363 3982
rect 16798 3980 16804 3982
rect 16868 3980 16874 4044
rect 16982 3980 16988 4044
rect 17052 4042 17058 4044
rect 18873 4042 18939 4045
rect 17052 4040 18939 4042
rect 17052 3984 18878 4040
rect 18934 3984 18939 4040
rect 17052 3982 18939 3984
rect 17052 3980 17058 3982
rect 18873 3979 18939 3982
rect 5130 3840 5450 3841
rect 5130 3776 5138 3840
rect 5202 3776 5218 3840
rect 5282 3776 5298 3840
rect 5362 3776 5378 3840
rect 5442 3776 5450 3840
rect 5130 3775 5450 3776
rect 13502 3840 13822 3841
rect 13502 3776 13510 3840
rect 13574 3776 13590 3840
rect 13654 3776 13670 3840
rect 13734 3776 13750 3840
rect 13814 3776 13822 3840
rect 13502 3775 13822 3776
rect 21874 3840 22194 3841
rect 21874 3776 21882 3840
rect 21946 3776 21962 3840
rect 22026 3776 22042 3840
rect 22106 3776 22122 3840
rect 22186 3776 22194 3840
rect 21874 3775 22194 3776
rect 8845 3636 8911 3637
rect 8845 3634 8892 3636
rect 8800 3632 8892 3634
rect 8800 3576 8850 3632
rect 8800 3574 8892 3576
rect 8845 3572 8892 3574
rect 8956 3572 8962 3636
rect 8845 3571 8911 3572
rect 657 3498 723 3501
rect 12014 3498 12020 3500
rect 657 3496 12020 3498
rect 657 3440 662 3496
rect 718 3440 12020 3496
rect 657 3438 12020 3440
rect 657 3435 723 3438
rect 12014 3436 12020 3438
rect 12084 3436 12090 3500
rect 22093 3498 22159 3501
rect 26595 3498 27395 3528
rect 22093 3496 27395 3498
rect 22093 3440 22098 3496
rect 22154 3440 27395 3496
rect 22093 3438 27395 3440
rect 22093 3435 22159 3438
rect 26595 3408 27395 3438
rect 8477 3362 8543 3365
rect 8702 3362 8708 3364
rect 8477 3360 8708 3362
rect 8477 3304 8482 3360
rect 8538 3304 8708 3360
rect 8477 3302 8708 3304
rect 8477 3299 8543 3302
rect 8702 3300 8708 3302
rect 8772 3300 8778 3364
rect 9316 3296 9636 3297
rect 9316 3232 9324 3296
rect 9388 3232 9404 3296
rect 9468 3232 9484 3296
rect 9548 3232 9564 3296
rect 9628 3232 9636 3296
rect 9316 3231 9636 3232
rect 17688 3296 18008 3297
rect 17688 3232 17696 3296
rect 17760 3232 17776 3296
rect 17840 3232 17856 3296
rect 17920 3232 17936 3296
rect 18000 3232 18008 3296
rect 17688 3231 18008 3232
rect 5130 2752 5450 2753
rect 0 2592 800 2712
rect 5130 2688 5138 2752
rect 5202 2688 5218 2752
rect 5282 2688 5298 2752
rect 5362 2688 5378 2752
rect 5442 2688 5450 2752
rect 5130 2687 5450 2688
rect 13502 2752 13822 2753
rect 13502 2688 13510 2752
rect 13574 2688 13590 2752
rect 13654 2688 13670 2752
rect 13734 2688 13750 2752
rect 13814 2688 13822 2752
rect 13502 2687 13822 2688
rect 21874 2752 22194 2753
rect 21874 2688 21882 2752
rect 21946 2688 21962 2752
rect 22026 2688 22042 2752
rect 22106 2688 22122 2752
rect 22186 2688 22194 2752
rect 21874 2687 22194 2688
rect 9316 2208 9636 2209
rect 9316 2144 9324 2208
rect 9388 2144 9404 2208
rect 9468 2144 9484 2208
rect 9548 2144 9564 2208
rect 9628 2144 9636 2208
rect 9316 2143 9636 2144
rect 17688 2208 18008 2209
rect 17688 2144 17696 2208
rect 17760 2144 17776 2208
rect 17840 2144 17856 2208
rect 17920 2144 17936 2208
rect 18000 2144 18008 2208
rect 17688 2143 18008 2144
rect 26595 2048 27395 2168
rect 0 914 800 944
rect 2957 914 3023 917
rect 0 912 3023 914
rect 0 856 2962 912
rect 3018 856 3023 912
rect 0 854 3023 856
rect 0 824 800 854
rect 2957 851 3023 854
rect 22093 778 22159 781
rect 26595 778 27395 808
rect 22093 776 27395 778
rect 22093 720 22098 776
rect 22154 720 27395 776
rect 22093 718 27395 720
rect 22093 715 22159 718
rect 26595 688 27395 718
<< via3 >>
rect 9324 27228 9388 27232
rect 9324 27172 9328 27228
rect 9328 27172 9384 27228
rect 9384 27172 9388 27228
rect 9324 27168 9388 27172
rect 9404 27228 9468 27232
rect 9404 27172 9408 27228
rect 9408 27172 9464 27228
rect 9464 27172 9468 27228
rect 9404 27168 9468 27172
rect 9484 27228 9548 27232
rect 9484 27172 9488 27228
rect 9488 27172 9544 27228
rect 9544 27172 9548 27228
rect 9484 27168 9548 27172
rect 9564 27228 9628 27232
rect 9564 27172 9568 27228
rect 9568 27172 9624 27228
rect 9624 27172 9628 27228
rect 9564 27168 9628 27172
rect 17696 27228 17760 27232
rect 17696 27172 17700 27228
rect 17700 27172 17756 27228
rect 17756 27172 17760 27228
rect 17696 27168 17760 27172
rect 17776 27228 17840 27232
rect 17776 27172 17780 27228
rect 17780 27172 17836 27228
rect 17836 27172 17840 27228
rect 17776 27168 17840 27172
rect 17856 27228 17920 27232
rect 17856 27172 17860 27228
rect 17860 27172 17916 27228
rect 17916 27172 17920 27228
rect 17856 27168 17920 27172
rect 17936 27228 18000 27232
rect 17936 27172 17940 27228
rect 17940 27172 17996 27228
rect 17996 27172 18000 27228
rect 17936 27168 18000 27172
rect 5138 26684 5202 26688
rect 5138 26628 5142 26684
rect 5142 26628 5198 26684
rect 5198 26628 5202 26684
rect 5138 26624 5202 26628
rect 5218 26684 5282 26688
rect 5218 26628 5222 26684
rect 5222 26628 5278 26684
rect 5278 26628 5282 26684
rect 5218 26624 5282 26628
rect 5298 26684 5362 26688
rect 5298 26628 5302 26684
rect 5302 26628 5358 26684
rect 5358 26628 5362 26684
rect 5298 26624 5362 26628
rect 5378 26684 5442 26688
rect 5378 26628 5382 26684
rect 5382 26628 5438 26684
rect 5438 26628 5442 26684
rect 5378 26624 5442 26628
rect 13510 26684 13574 26688
rect 13510 26628 13514 26684
rect 13514 26628 13570 26684
rect 13570 26628 13574 26684
rect 13510 26624 13574 26628
rect 13590 26684 13654 26688
rect 13590 26628 13594 26684
rect 13594 26628 13650 26684
rect 13650 26628 13654 26684
rect 13590 26624 13654 26628
rect 13670 26684 13734 26688
rect 13670 26628 13674 26684
rect 13674 26628 13730 26684
rect 13730 26628 13734 26684
rect 13670 26624 13734 26628
rect 13750 26684 13814 26688
rect 13750 26628 13754 26684
rect 13754 26628 13810 26684
rect 13810 26628 13814 26684
rect 13750 26624 13814 26628
rect 21882 26684 21946 26688
rect 21882 26628 21886 26684
rect 21886 26628 21942 26684
rect 21942 26628 21946 26684
rect 21882 26624 21946 26628
rect 21962 26684 22026 26688
rect 21962 26628 21966 26684
rect 21966 26628 22022 26684
rect 22022 26628 22026 26684
rect 21962 26624 22026 26628
rect 22042 26684 22106 26688
rect 22042 26628 22046 26684
rect 22046 26628 22102 26684
rect 22102 26628 22106 26684
rect 22042 26624 22106 26628
rect 22122 26684 22186 26688
rect 22122 26628 22126 26684
rect 22126 26628 22182 26684
rect 22182 26628 22186 26684
rect 22122 26624 22186 26628
rect 9324 26140 9388 26144
rect 9324 26084 9328 26140
rect 9328 26084 9384 26140
rect 9384 26084 9388 26140
rect 9324 26080 9388 26084
rect 9404 26140 9468 26144
rect 9404 26084 9408 26140
rect 9408 26084 9464 26140
rect 9464 26084 9468 26140
rect 9404 26080 9468 26084
rect 9484 26140 9548 26144
rect 9484 26084 9488 26140
rect 9488 26084 9544 26140
rect 9544 26084 9548 26140
rect 9484 26080 9548 26084
rect 9564 26140 9628 26144
rect 9564 26084 9568 26140
rect 9568 26084 9624 26140
rect 9624 26084 9628 26140
rect 9564 26080 9628 26084
rect 17696 26140 17760 26144
rect 17696 26084 17700 26140
rect 17700 26084 17756 26140
rect 17756 26084 17760 26140
rect 17696 26080 17760 26084
rect 17776 26140 17840 26144
rect 17776 26084 17780 26140
rect 17780 26084 17836 26140
rect 17836 26084 17840 26140
rect 17776 26080 17840 26084
rect 17856 26140 17920 26144
rect 17856 26084 17860 26140
rect 17860 26084 17916 26140
rect 17916 26084 17920 26140
rect 17856 26080 17920 26084
rect 17936 26140 18000 26144
rect 17936 26084 17940 26140
rect 17940 26084 17996 26140
rect 17996 26084 18000 26140
rect 17936 26080 18000 26084
rect 5138 25596 5202 25600
rect 5138 25540 5142 25596
rect 5142 25540 5198 25596
rect 5198 25540 5202 25596
rect 5138 25536 5202 25540
rect 5218 25596 5282 25600
rect 5218 25540 5222 25596
rect 5222 25540 5278 25596
rect 5278 25540 5282 25596
rect 5218 25536 5282 25540
rect 5298 25596 5362 25600
rect 5298 25540 5302 25596
rect 5302 25540 5358 25596
rect 5358 25540 5362 25596
rect 5298 25536 5362 25540
rect 5378 25596 5442 25600
rect 5378 25540 5382 25596
rect 5382 25540 5438 25596
rect 5438 25540 5442 25596
rect 5378 25536 5442 25540
rect 13510 25596 13574 25600
rect 13510 25540 13514 25596
rect 13514 25540 13570 25596
rect 13570 25540 13574 25596
rect 13510 25536 13574 25540
rect 13590 25596 13654 25600
rect 13590 25540 13594 25596
rect 13594 25540 13650 25596
rect 13650 25540 13654 25596
rect 13590 25536 13654 25540
rect 13670 25596 13734 25600
rect 13670 25540 13674 25596
rect 13674 25540 13730 25596
rect 13730 25540 13734 25596
rect 13670 25536 13734 25540
rect 13750 25596 13814 25600
rect 13750 25540 13754 25596
rect 13754 25540 13810 25596
rect 13810 25540 13814 25596
rect 13750 25536 13814 25540
rect 21882 25596 21946 25600
rect 21882 25540 21886 25596
rect 21886 25540 21942 25596
rect 21942 25540 21946 25596
rect 21882 25536 21946 25540
rect 21962 25596 22026 25600
rect 21962 25540 21966 25596
rect 21966 25540 22022 25596
rect 22022 25540 22026 25596
rect 21962 25536 22026 25540
rect 22042 25596 22106 25600
rect 22042 25540 22046 25596
rect 22046 25540 22102 25596
rect 22102 25540 22106 25596
rect 22042 25536 22106 25540
rect 22122 25596 22186 25600
rect 22122 25540 22126 25596
rect 22126 25540 22182 25596
rect 22182 25540 22186 25596
rect 22122 25536 22186 25540
rect 9324 25052 9388 25056
rect 9324 24996 9328 25052
rect 9328 24996 9384 25052
rect 9384 24996 9388 25052
rect 9324 24992 9388 24996
rect 9404 25052 9468 25056
rect 9404 24996 9408 25052
rect 9408 24996 9464 25052
rect 9464 24996 9468 25052
rect 9404 24992 9468 24996
rect 9484 25052 9548 25056
rect 9484 24996 9488 25052
rect 9488 24996 9544 25052
rect 9544 24996 9548 25052
rect 9484 24992 9548 24996
rect 9564 25052 9628 25056
rect 9564 24996 9568 25052
rect 9568 24996 9624 25052
rect 9624 24996 9628 25052
rect 9564 24992 9628 24996
rect 17696 25052 17760 25056
rect 17696 24996 17700 25052
rect 17700 24996 17756 25052
rect 17756 24996 17760 25052
rect 17696 24992 17760 24996
rect 17776 25052 17840 25056
rect 17776 24996 17780 25052
rect 17780 24996 17836 25052
rect 17836 24996 17840 25052
rect 17776 24992 17840 24996
rect 17856 25052 17920 25056
rect 17856 24996 17860 25052
rect 17860 24996 17916 25052
rect 17916 24996 17920 25052
rect 17856 24992 17920 24996
rect 17936 25052 18000 25056
rect 17936 24996 17940 25052
rect 17940 24996 17996 25052
rect 17996 24996 18000 25052
rect 17936 24992 18000 24996
rect 5138 24508 5202 24512
rect 5138 24452 5142 24508
rect 5142 24452 5198 24508
rect 5198 24452 5202 24508
rect 5138 24448 5202 24452
rect 5218 24508 5282 24512
rect 5218 24452 5222 24508
rect 5222 24452 5278 24508
rect 5278 24452 5282 24508
rect 5218 24448 5282 24452
rect 5298 24508 5362 24512
rect 5298 24452 5302 24508
rect 5302 24452 5358 24508
rect 5358 24452 5362 24508
rect 5298 24448 5362 24452
rect 5378 24508 5442 24512
rect 5378 24452 5382 24508
rect 5382 24452 5438 24508
rect 5438 24452 5442 24508
rect 5378 24448 5442 24452
rect 13510 24508 13574 24512
rect 13510 24452 13514 24508
rect 13514 24452 13570 24508
rect 13570 24452 13574 24508
rect 13510 24448 13574 24452
rect 13590 24508 13654 24512
rect 13590 24452 13594 24508
rect 13594 24452 13650 24508
rect 13650 24452 13654 24508
rect 13590 24448 13654 24452
rect 13670 24508 13734 24512
rect 13670 24452 13674 24508
rect 13674 24452 13730 24508
rect 13730 24452 13734 24508
rect 13670 24448 13734 24452
rect 13750 24508 13814 24512
rect 13750 24452 13754 24508
rect 13754 24452 13810 24508
rect 13810 24452 13814 24508
rect 13750 24448 13814 24452
rect 21882 24508 21946 24512
rect 21882 24452 21886 24508
rect 21886 24452 21942 24508
rect 21942 24452 21946 24508
rect 21882 24448 21946 24452
rect 21962 24508 22026 24512
rect 21962 24452 21966 24508
rect 21966 24452 22022 24508
rect 22022 24452 22026 24508
rect 21962 24448 22026 24452
rect 22042 24508 22106 24512
rect 22042 24452 22046 24508
rect 22046 24452 22102 24508
rect 22102 24452 22106 24508
rect 22042 24448 22106 24452
rect 22122 24508 22186 24512
rect 22122 24452 22126 24508
rect 22126 24452 22182 24508
rect 22182 24452 22186 24508
rect 22122 24448 22186 24452
rect 9324 23964 9388 23968
rect 9324 23908 9328 23964
rect 9328 23908 9384 23964
rect 9384 23908 9388 23964
rect 9324 23904 9388 23908
rect 9404 23964 9468 23968
rect 9404 23908 9408 23964
rect 9408 23908 9464 23964
rect 9464 23908 9468 23964
rect 9404 23904 9468 23908
rect 9484 23964 9548 23968
rect 9484 23908 9488 23964
rect 9488 23908 9544 23964
rect 9544 23908 9548 23964
rect 9484 23904 9548 23908
rect 9564 23964 9628 23968
rect 9564 23908 9568 23964
rect 9568 23908 9624 23964
rect 9624 23908 9628 23964
rect 9564 23904 9628 23908
rect 17696 23964 17760 23968
rect 17696 23908 17700 23964
rect 17700 23908 17756 23964
rect 17756 23908 17760 23964
rect 17696 23904 17760 23908
rect 17776 23964 17840 23968
rect 17776 23908 17780 23964
rect 17780 23908 17836 23964
rect 17836 23908 17840 23964
rect 17776 23904 17840 23908
rect 17856 23964 17920 23968
rect 17856 23908 17860 23964
rect 17860 23908 17916 23964
rect 17916 23908 17920 23964
rect 17856 23904 17920 23908
rect 17936 23964 18000 23968
rect 17936 23908 17940 23964
rect 17940 23908 17996 23964
rect 17996 23908 18000 23964
rect 17936 23904 18000 23908
rect 5138 23420 5202 23424
rect 5138 23364 5142 23420
rect 5142 23364 5198 23420
rect 5198 23364 5202 23420
rect 5138 23360 5202 23364
rect 5218 23420 5282 23424
rect 5218 23364 5222 23420
rect 5222 23364 5278 23420
rect 5278 23364 5282 23420
rect 5218 23360 5282 23364
rect 5298 23420 5362 23424
rect 5298 23364 5302 23420
rect 5302 23364 5358 23420
rect 5358 23364 5362 23420
rect 5298 23360 5362 23364
rect 5378 23420 5442 23424
rect 5378 23364 5382 23420
rect 5382 23364 5438 23420
rect 5438 23364 5442 23420
rect 5378 23360 5442 23364
rect 13510 23420 13574 23424
rect 13510 23364 13514 23420
rect 13514 23364 13570 23420
rect 13570 23364 13574 23420
rect 13510 23360 13574 23364
rect 13590 23420 13654 23424
rect 13590 23364 13594 23420
rect 13594 23364 13650 23420
rect 13650 23364 13654 23420
rect 13590 23360 13654 23364
rect 13670 23420 13734 23424
rect 13670 23364 13674 23420
rect 13674 23364 13730 23420
rect 13730 23364 13734 23420
rect 13670 23360 13734 23364
rect 13750 23420 13814 23424
rect 13750 23364 13754 23420
rect 13754 23364 13810 23420
rect 13810 23364 13814 23420
rect 13750 23360 13814 23364
rect 21882 23420 21946 23424
rect 21882 23364 21886 23420
rect 21886 23364 21942 23420
rect 21942 23364 21946 23420
rect 21882 23360 21946 23364
rect 21962 23420 22026 23424
rect 21962 23364 21966 23420
rect 21966 23364 22022 23420
rect 22022 23364 22026 23420
rect 21962 23360 22026 23364
rect 22042 23420 22106 23424
rect 22042 23364 22046 23420
rect 22046 23364 22102 23420
rect 22102 23364 22106 23420
rect 22042 23360 22106 23364
rect 22122 23420 22186 23424
rect 22122 23364 22126 23420
rect 22126 23364 22182 23420
rect 22182 23364 22186 23420
rect 22122 23360 22186 23364
rect 9324 22876 9388 22880
rect 9324 22820 9328 22876
rect 9328 22820 9384 22876
rect 9384 22820 9388 22876
rect 9324 22816 9388 22820
rect 9404 22876 9468 22880
rect 9404 22820 9408 22876
rect 9408 22820 9464 22876
rect 9464 22820 9468 22876
rect 9404 22816 9468 22820
rect 9484 22876 9548 22880
rect 9484 22820 9488 22876
rect 9488 22820 9544 22876
rect 9544 22820 9548 22876
rect 9484 22816 9548 22820
rect 9564 22876 9628 22880
rect 9564 22820 9568 22876
rect 9568 22820 9624 22876
rect 9624 22820 9628 22876
rect 9564 22816 9628 22820
rect 17696 22876 17760 22880
rect 17696 22820 17700 22876
rect 17700 22820 17756 22876
rect 17756 22820 17760 22876
rect 17696 22816 17760 22820
rect 17776 22876 17840 22880
rect 17776 22820 17780 22876
rect 17780 22820 17836 22876
rect 17836 22820 17840 22876
rect 17776 22816 17840 22820
rect 17856 22876 17920 22880
rect 17856 22820 17860 22876
rect 17860 22820 17916 22876
rect 17916 22820 17920 22876
rect 17856 22816 17920 22820
rect 17936 22876 18000 22880
rect 17936 22820 17940 22876
rect 17940 22820 17996 22876
rect 17996 22820 18000 22876
rect 17936 22816 18000 22820
rect 5138 22332 5202 22336
rect 5138 22276 5142 22332
rect 5142 22276 5198 22332
rect 5198 22276 5202 22332
rect 5138 22272 5202 22276
rect 5218 22332 5282 22336
rect 5218 22276 5222 22332
rect 5222 22276 5278 22332
rect 5278 22276 5282 22332
rect 5218 22272 5282 22276
rect 5298 22332 5362 22336
rect 5298 22276 5302 22332
rect 5302 22276 5358 22332
rect 5358 22276 5362 22332
rect 5298 22272 5362 22276
rect 5378 22332 5442 22336
rect 5378 22276 5382 22332
rect 5382 22276 5438 22332
rect 5438 22276 5442 22332
rect 5378 22272 5442 22276
rect 13510 22332 13574 22336
rect 13510 22276 13514 22332
rect 13514 22276 13570 22332
rect 13570 22276 13574 22332
rect 13510 22272 13574 22276
rect 13590 22332 13654 22336
rect 13590 22276 13594 22332
rect 13594 22276 13650 22332
rect 13650 22276 13654 22332
rect 13590 22272 13654 22276
rect 13670 22332 13734 22336
rect 13670 22276 13674 22332
rect 13674 22276 13730 22332
rect 13730 22276 13734 22332
rect 13670 22272 13734 22276
rect 13750 22332 13814 22336
rect 13750 22276 13754 22332
rect 13754 22276 13810 22332
rect 13810 22276 13814 22332
rect 13750 22272 13814 22276
rect 21882 22332 21946 22336
rect 21882 22276 21886 22332
rect 21886 22276 21942 22332
rect 21942 22276 21946 22332
rect 21882 22272 21946 22276
rect 21962 22332 22026 22336
rect 21962 22276 21966 22332
rect 21966 22276 22022 22332
rect 22022 22276 22026 22332
rect 21962 22272 22026 22276
rect 22042 22332 22106 22336
rect 22042 22276 22046 22332
rect 22046 22276 22102 22332
rect 22102 22276 22106 22332
rect 22042 22272 22106 22276
rect 22122 22332 22186 22336
rect 22122 22276 22126 22332
rect 22126 22276 22182 22332
rect 22182 22276 22186 22332
rect 22122 22272 22186 22276
rect 22508 22128 22572 22132
rect 22508 22072 22522 22128
rect 22522 22072 22572 22128
rect 22508 22068 22572 22072
rect 9324 21788 9388 21792
rect 9324 21732 9328 21788
rect 9328 21732 9384 21788
rect 9384 21732 9388 21788
rect 9324 21728 9388 21732
rect 9404 21788 9468 21792
rect 9404 21732 9408 21788
rect 9408 21732 9464 21788
rect 9464 21732 9468 21788
rect 9404 21728 9468 21732
rect 9484 21788 9548 21792
rect 9484 21732 9488 21788
rect 9488 21732 9544 21788
rect 9544 21732 9548 21788
rect 9484 21728 9548 21732
rect 9564 21788 9628 21792
rect 9564 21732 9568 21788
rect 9568 21732 9624 21788
rect 9624 21732 9628 21788
rect 9564 21728 9628 21732
rect 17696 21788 17760 21792
rect 17696 21732 17700 21788
rect 17700 21732 17756 21788
rect 17756 21732 17760 21788
rect 17696 21728 17760 21732
rect 17776 21788 17840 21792
rect 17776 21732 17780 21788
rect 17780 21732 17836 21788
rect 17836 21732 17840 21788
rect 17776 21728 17840 21732
rect 17856 21788 17920 21792
rect 17856 21732 17860 21788
rect 17860 21732 17916 21788
rect 17916 21732 17920 21788
rect 17856 21728 17920 21732
rect 17936 21788 18000 21792
rect 17936 21732 17940 21788
rect 17940 21732 17996 21788
rect 17996 21732 18000 21788
rect 17936 21728 18000 21732
rect 5138 21244 5202 21248
rect 5138 21188 5142 21244
rect 5142 21188 5198 21244
rect 5198 21188 5202 21244
rect 5138 21184 5202 21188
rect 5218 21244 5282 21248
rect 5218 21188 5222 21244
rect 5222 21188 5278 21244
rect 5278 21188 5282 21244
rect 5218 21184 5282 21188
rect 5298 21244 5362 21248
rect 5298 21188 5302 21244
rect 5302 21188 5358 21244
rect 5358 21188 5362 21244
rect 5298 21184 5362 21188
rect 5378 21244 5442 21248
rect 5378 21188 5382 21244
rect 5382 21188 5438 21244
rect 5438 21188 5442 21244
rect 5378 21184 5442 21188
rect 13510 21244 13574 21248
rect 13510 21188 13514 21244
rect 13514 21188 13570 21244
rect 13570 21188 13574 21244
rect 13510 21184 13574 21188
rect 13590 21244 13654 21248
rect 13590 21188 13594 21244
rect 13594 21188 13650 21244
rect 13650 21188 13654 21244
rect 13590 21184 13654 21188
rect 13670 21244 13734 21248
rect 13670 21188 13674 21244
rect 13674 21188 13730 21244
rect 13730 21188 13734 21244
rect 13670 21184 13734 21188
rect 13750 21244 13814 21248
rect 13750 21188 13754 21244
rect 13754 21188 13810 21244
rect 13810 21188 13814 21244
rect 13750 21184 13814 21188
rect 21882 21244 21946 21248
rect 21882 21188 21886 21244
rect 21886 21188 21942 21244
rect 21942 21188 21946 21244
rect 21882 21184 21946 21188
rect 21962 21244 22026 21248
rect 21962 21188 21966 21244
rect 21966 21188 22022 21244
rect 22022 21188 22026 21244
rect 21962 21184 22026 21188
rect 22042 21244 22106 21248
rect 22042 21188 22046 21244
rect 22046 21188 22102 21244
rect 22102 21188 22106 21244
rect 22042 21184 22106 21188
rect 22122 21244 22186 21248
rect 22122 21188 22126 21244
rect 22126 21188 22182 21244
rect 22182 21188 22186 21244
rect 22122 21184 22186 21188
rect 9324 20700 9388 20704
rect 9324 20644 9328 20700
rect 9328 20644 9384 20700
rect 9384 20644 9388 20700
rect 9324 20640 9388 20644
rect 9404 20700 9468 20704
rect 9404 20644 9408 20700
rect 9408 20644 9464 20700
rect 9464 20644 9468 20700
rect 9404 20640 9468 20644
rect 9484 20700 9548 20704
rect 9484 20644 9488 20700
rect 9488 20644 9544 20700
rect 9544 20644 9548 20700
rect 9484 20640 9548 20644
rect 9564 20700 9628 20704
rect 9564 20644 9568 20700
rect 9568 20644 9624 20700
rect 9624 20644 9628 20700
rect 9564 20640 9628 20644
rect 17696 20700 17760 20704
rect 17696 20644 17700 20700
rect 17700 20644 17756 20700
rect 17756 20644 17760 20700
rect 17696 20640 17760 20644
rect 17776 20700 17840 20704
rect 17776 20644 17780 20700
rect 17780 20644 17836 20700
rect 17836 20644 17840 20700
rect 17776 20640 17840 20644
rect 17856 20700 17920 20704
rect 17856 20644 17860 20700
rect 17860 20644 17916 20700
rect 17916 20644 17920 20700
rect 17856 20640 17920 20644
rect 17936 20700 18000 20704
rect 17936 20644 17940 20700
rect 17940 20644 17996 20700
rect 17996 20644 18000 20700
rect 17936 20640 18000 20644
rect 5138 20156 5202 20160
rect 5138 20100 5142 20156
rect 5142 20100 5198 20156
rect 5198 20100 5202 20156
rect 5138 20096 5202 20100
rect 5218 20156 5282 20160
rect 5218 20100 5222 20156
rect 5222 20100 5278 20156
rect 5278 20100 5282 20156
rect 5218 20096 5282 20100
rect 5298 20156 5362 20160
rect 5298 20100 5302 20156
rect 5302 20100 5358 20156
rect 5358 20100 5362 20156
rect 5298 20096 5362 20100
rect 5378 20156 5442 20160
rect 5378 20100 5382 20156
rect 5382 20100 5438 20156
rect 5438 20100 5442 20156
rect 5378 20096 5442 20100
rect 13510 20156 13574 20160
rect 13510 20100 13514 20156
rect 13514 20100 13570 20156
rect 13570 20100 13574 20156
rect 13510 20096 13574 20100
rect 13590 20156 13654 20160
rect 13590 20100 13594 20156
rect 13594 20100 13650 20156
rect 13650 20100 13654 20156
rect 13590 20096 13654 20100
rect 13670 20156 13734 20160
rect 13670 20100 13674 20156
rect 13674 20100 13730 20156
rect 13730 20100 13734 20156
rect 13670 20096 13734 20100
rect 13750 20156 13814 20160
rect 13750 20100 13754 20156
rect 13754 20100 13810 20156
rect 13810 20100 13814 20156
rect 13750 20096 13814 20100
rect 21882 20156 21946 20160
rect 21882 20100 21886 20156
rect 21886 20100 21942 20156
rect 21942 20100 21946 20156
rect 21882 20096 21946 20100
rect 21962 20156 22026 20160
rect 21962 20100 21966 20156
rect 21966 20100 22022 20156
rect 22022 20100 22026 20156
rect 21962 20096 22026 20100
rect 22042 20156 22106 20160
rect 22042 20100 22046 20156
rect 22046 20100 22102 20156
rect 22102 20100 22106 20156
rect 22042 20096 22106 20100
rect 22122 20156 22186 20160
rect 22122 20100 22126 20156
rect 22126 20100 22182 20156
rect 22182 20100 22186 20156
rect 22122 20096 22186 20100
rect 16988 19620 17052 19684
rect 9324 19612 9388 19616
rect 9324 19556 9328 19612
rect 9328 19556 9384 19612
rect 9384 19556 9388 19612
rect 9324 19552 9388 19556
rect 9404 19612 9468 19616
rect 9404 19556 9408 19612
rect 9408 19556 9464 19612
rect 9464 19556 9468 19612
rect 9404 19552 9468 19556
rect 9484 19612 9548 19616
rect 9484 19556 9488 19612
rect 9488 19556 9544 19612
rect 9544 19556 9548 19612
rect 9484 19552 9548 19556
rect 9564 19612 9628 19616
rect 9564 19556 9568 19612
rect 9568 19556 9624 19612
rect 9624 19556 9628 19612
rect 9564 19552 9628 19556
rect 17696 19612 17760 19616
rect 17696 19556 17700 19612
rect 17700 19556 17756 19612
rect 17756 19556 17760 19612
rect 17696 19552 17760 19556
rect 17776 19612 17840 19616
rect 17776 19556 17780 19612
rect 17780 19556 17836 19612
rect 17836 19556 17840 19612
rect 17776 19552 17840 19556
rect 17856 19612 17920 19616
rect 17856 19556 17860 19612
rect 17860 19556 17916 19612
rect 17916 19556 17920 19612
rect 17856 19552 17920 19556
rect 17936 19612 18000 19616
rect 17936 19556 17940 19612
rect 17940 19556 17996 19612
rect 17996 19556 18000 19612
rect 17936 19552 18000 19556
rect 5138 19068 5202 19072
rect 5138 19012 5142 19068
rect 5142 19012 5198 19068
rect 5198 19012 5202 19068
rect 5138 19008 5202 19012
rect 5218 19068 5282 19072
rect 5218 19012 5222 19068
rect 5222 19012 5278 19068
rect 5278 19012 5282 19068
rect 5218 19008 5282 19012
rect 5298 19068 5362 19072
rect 5298 19012 5302 19068
rect 5302 19012 5358 19068
rect 5358 19012 5362 19068
rect 5298 19008 5362 19012
rect 5378 19068 5442 19072
rect 5378 19012 5382 19068
rect 5382 19012 5438 19068
rect 5438 19012 5442 19068
rect 5378 19008 5442 19012
rect 13510 19068 13574 19072
rect 13510 19012 13514 19068
rect 13514 19012 13570 19068
rect 13570 19012 13574 19068
rect 13510 19008 13574 19012
rect 13590 19068 13654 19072
rect 13590 19012 13594 19068
rect 13594 19012 13650 19068
rect 13650 19012 13654 19068
rect 13590 19008 13654 19012
rect 13670 19068 13734 19072
rect 13670 19012 13674 19068
rect 13674 19012 13730 19068
rect 13730 19012 13734 19068
rect 13670 19008 13734 19012
rect 13750 19068 13814 19072
rect 13750 19012 13754 19068
rect 13754 19012 13810 19068
rect 13810 19012 13814 19068
rect 13750 19008 13814 19012
rect 21882 19068 21946 19072
rect 21882 19012 21886 19068
rect 21886 19012 21942 19068
rect 21942 19012 21946 19068
rect 21882 19008 21946 19012
rect 21962 19068 22026 19072
rect 21962 19012 21966 19068
rect 21966 19012 22022 19068
rect 22022 19012 22026 19068
rect 21962 19008 22026 19012
rect 22042 19068 22106 19072
rect 22042 19012 22046 19068
rect 22046 19012 22102 19068
rect 22102 19012 22106 19068
rect 22042 19008 22106 19012
rect 22122 19068 22186 19072
rect 22122 19012 22126 19068
rect 22126 19012 22182 19068
rect 22182 19012 22186 19068
rect 22122 19008 22186 19012
rect 8892 18728 8956 18732
rect 8892 18672 8942 18728
rect 8942 18672 8956 18728
rect 8892 18668 8956 18672
rect 9324 18524 9388 18528
rect 9324 18468 9328 18524
rect 9328 18468 9384 18524
rect 9384 18468 9388 18524
rect 9324 18464 9388 18468
rect 9404 18524 9468 18528
rect 9404 18468 9408 18524
rect 9408 18468 9464 18524
rect 9464 18468 9468 18524
rect 9404 18464 9468 18468
rect 9484 18524 9548 18528
rect 9484 18468 9488 18524
rect 9488 18468 9544 18524
rect 9544 18468 9548 18524
rect 9484 18464 9548 18468
rect 9564 18524 9628 18528
rect 9564 18468 9568 18524
rect 9568 18468 9624 18524
rect 9624 18468 9628 18524
rect 9564 18464 9628 18468
rect 17696 18524 17760 18528
rect 17696 18468 17700 18524
rect 17700 18468 17756 18524
rect 17756 18468 17760 18524
rect 17696 18464 17760 18468
rect 17776 18524 17840 18528
rect 17776 18468 17780 18524
rect 17780 18468 17836 18524
rect 17836 18468 17840 18524
rect 17776 18464 17840 18468
rect 17856 18524 17920 18528
rect 17856 18468 17860 18524
rect 17860 18468 17916 18524
rect 17916 18468 17920 18524
rect 17856 18464 17920 18468
rect 17936 18524 18000 18528
rect 17936 18468 17940 18524
rect 17940 18468 17996 18524
rect 17996 18468 18000 18524
rect 17936 18464 18000 18468
rect 5138 17980 5202 17984
rect 5138 17924 5142 17980
rect 5142 17924 5198 17980
rect 5198 17924 5202 17980
rect 5138 17920 5202 17924
rect 5218 17980 5282 17984
rect 5218 17924 5222 17980
rect 5222 17924 5278 17980
rect 5278 17924 5282 17980
rect 5218 17920 5282 17924
rect 5298 17980 5362 17984
rect 5298 17924 5302 17980
rect 5302 17924 5358 17980
rect 5358 17924 5362 17980
rect 5298 17920 5362 17924
rect 5378 17980 5442 17984
rect 5378 17924 5382 17980
rect 5382 17924 5438 17980
rect 5438 17924 5442 17980
rect 5378 17920 5442 17924
rect 13510 17980 13574 17984
rect 13510 17924 13514 17980
rect 13514 17924 13570 17980
rect 13570 17924 13574 17980
rect 13510 17920 13574 17924
rect 13590 17980 13654 17984
rect 13590 17924 13594 17980
rect 13594 17924 13650 17980
rect 13650 17924 13654 17980
rect 13590 17920 13654 17924
rect 13670 17980 13734 17984
rect 13670 17924 13674 17980
rect 13674 17924 13730 17980
rect 13730 17924 13734 17980
rect 13670 17920 13734 17924
rect 13750 17980 13814 17984
rect 13750 17924 13754 17980
rect 13754 17924 13810 17980
rect 13810 17924 13814 17980
rect 13750 17920 13814 17924
rect 21882 17980 21946 17984
rect 21882 17924 21886 17980
rect 21886 17924 21942 17980
rect 21942 17924 21946 17980
rect 21882 17920 21946 17924
rect 21962 17980 22026 17984
rect 21962 17924 21966 17980
rect 21966 17924 22022 17980
rect 22022 17924 22026 17980
rect 21962 17920 22026 17924
rect 22042 17980 22106 17984
rect 22042 17924 22046 17980
rect 22046 17924 22102 17980
rect 22102 17924 22106 17980
rect 22042 17920 22106 17924
rect 22122 17980 22186 17984
rect 22122 17924 22126 17980
rect 22126 17924 22182 17980
rect 22182 17924 22186 17980
rect 22122 17920 22186 17924
rect 9324 17436 9388 17440
rect 9324 17380 9328 17436
rect 9328 17380 9384 17436
rect 9384 17380 9388 17436
rect 9324 17376 9388 17380
rect 9404 17436 9468 17440
rect 9404 17380 9408 17436
rect 9408 17380 9464 17436
rect 9464 17380 9468 17436
rect 9404 17376 9468 17380
rect 9484 17436 9548 17440
rect 9484 17380 9488 17436
rect 9488 17380 9544 17436
rect 9544 17380 9548 17436
rect 9484 17376 9548 17380
rect 9564 17436 9628 17440
rect 9564 17380 9568 17436
rect 9568 17380 9624 17436
rect 9624 17380 9628 17436
rect 9564 17376 9628 17380
rect 17696 17436 17760 17440
rect 17696 17380 17700 17436
rect 17700 17380 17756 17436
rect 17756 17380 17760 17436
rect 17696 17376 17760 17380
rect 17776 17436 17840 17440
rect 17776 17380 17780 17436
rect 17780 17380 17836 17436
rect 17836 17380 17840 17436
rect 17776 17376 17840 17380
rect 17856 17436 17920 17440
rect 17856 17380 17860 17436
rect 17860 17380 17916 17436
rect 17916 17380 17920 17436
rect 17856 17376 17920 17380
rect 17936 17436 18000 17440
rect 17936 17380 17940 17436
rect 17940 17380 17996 17436
rect 17996 17380 18000 17436
rect 17936 17376 18000 17380
rect 5138 16892 5202 16896
rect 5138 16836 5142 16892
rect 5142 16836 5198 16892
rect 5198 16836 5202 16892
rect 5138 16832 5202 16836
rect 5218 16892 5282 16896
rect 5218 16836 5222 16892
rect 5222 16836 5278 16892
rect 5278 16836 5282 16892
rect 5218 16832 5282 16836
rect 5298 16892 5362 16896
rect 5298 16836 5302 16892
rect 5302 16836 5358 16892
rect 5358 16836 5362 16892
rect 5298 16832 5362 16836
rect 5378 16892 5442 16896
rect 5378 16836 5382 16892
rect 5382 16836 5438 16892
rect 5438 16836 5442 16892
rect 5378 16832 5442 16836
rect 13510 16892 13574 16896
rect 13510 16836 13514 16892
rect 13514 16836 13570 16892
rect 13570 16836 13574 16892
rect 13510 16832 13574 16836
rect 13590 16892 13654 16896
rect 13590 16836 13594 16892
rect 13594 16836 13650 16892
rect 13650 16836 13654 16892
rect 13590 16832 13654 16836
rect 13670 16892 13734 16896
rect 13670 16836 13674 16892
rect 13674 16836 13730 16892
rect 13730 16836 13734 16892
rect 13670 16832 13734 16836
rect 13750 16892 13814 16896
rect 13750 16836 13754 16892
rect 13754 16836 13810 16892
rect 13810 16836 13814 16892
rect 13750 16832 13814 16836
rect 21882 16892 21946 16896
rect 21882 16836 21886 16892
rect 21886 16836 21942 16892
rect 21942 16836 21946 16892
rect 21882 16832 21946 16836
rect 21962 16892 22026 16896
rect 21962 16836 21966 16892
rect 21966 16836 22022 16892
rect 22022 16836 22026 16892
rect 21962 16832 22026 16836
rect 22042 16892 22106 16896
rect 22042 16836 22046 16892
rect 22046 16836 22102 16892
rect 22102 16836 22106 16892
rect 22042 16832 22106 16836
rect 22122 16892 22186 16896
rect 22122 16836 22126 16892
rect 22126 16836 22182 16892
rect 22182 16836 22186 16892
rect 22122 16832 22186 16836
rect 9324 16348 9388 16352
rect 9324 16292 9328 16348
rect 9328 16292 9384 16348
rect 9384 16292 9388 16348
rect 9324 16288 9388 16292
rect 9404 16348 9468 16352
rect 9404 16292 9408 16348
rect 9408 16292 9464 16348
rect 9464 16292 9468 16348
rect 9404 16288 9468 16292
rect 9484 16348 9548 16352
rect 9484 16292 9488 16348
rect 9488 16292 9544 16348
rect 9544 16292 9548 16348
rect 9484 16288 9548 16292
rect 9564 16348 9628 16352
rect 9564 16292 9568 16348
rect 9568 16292 9624 16348
rect 9624 16292 9628 16348
rect 9564 16288 9628 16292
rect 17696 16348 17760 16352
rect 17696 16292 17700 16348
rect 17700 16292 17756 16348
rect 17756 16292 17760 16348
rect 17696 16288 17760 16292
rect 17776 16348 17840 16352
rect 17776 16292 17780 16348
rect 17780 16292 17836 16348
rect 17836 16292 17840 16348
rect 17776 16288 17840 16292
rect 17856 16348 17920 16352
rect 17856 16292 17860 16348
rect 17860 16292 17916 16348
rect 17916 16292 17920 16348
rect 17856 16288 17920 16292
rect 17936 16348 18000 16352
rect 17936 16292 17940 16348
rect 17940 16292 17996 16348
rect 17996 16292 18000 16348
rect 17936 16288 18000 16292
rect 5138 15804 5202 15808
rect 5138 15748 5142 15804
rect 5142 15748 5198 15804
rect 5198 15748 5202 15804
rect 5138 15744 5202 15748
rect 5218 15804 5282 15808
rect 5218 15748 5222 15804
rect 5222 15748 5278 15804
rect 5278 15748 5282 15804
rect 5218 15744 5282 15748
rect 5298 15804 5362 15808
rect 5298 15748 5302 15804
rect 5302 15748 5358 15804
rect 5358 15748 5362 15804
rect 5298 15744 5362 15748
rect 5378 15804 5442 15808
rect 5378 15748 5382 15804
rect 5382 15748 5438 15804
rect 5438 15748 5442 15804
rect 5378 15744 5442 15748
rect 13510 15804 13574 15808
rect 13510 15748 13514 15804
rect 13514 15748 13570 15804
rect 13570 15748 13574 15804
rect 13510 15744 13574 15748
rect 13590 15804 13654 15808
rect 13590 15748 13594 15804
rect 13594 15748 13650 15804
rect 13650 15748 13654 15804
rect 13590 15744 13654 15748
rect 13670 15804 13734 15808
rect 13670 15748 13674 15804
rect 13674 15748 13730 15804
rect 13730 15748 13734 15804
rect 13670 15744 13734 15748
rect 13750 15804 13814 15808
rect 13750 15748 13754 15804
rect 13754 15748 13810 15804
rect 13810 15748 13814 15804
rect 13750 15744 13814 15748
rect 21882 15804 21946 15808
rect 21882 15748 21886 15804
rect 21886 15748 21942 15804
rect 21942 15748 21946 15804
rect 21882 15744 21946 15748
rect 21962 15804 22026 15808
rect 21962 15748 21966 15804
rect 21966 15748 22022 15804
rect 22022 15748 22026 15804
rect 21962 15744 22026 15748
rect 22042 15804 22106 15808
rect 22042 15748 22046 15804
rect 22046 15748 22102 15804
rect 22102 15748 22106 15804
rect 22042 15744 22106 15748
rect 22122 15804 22186 15808
rect 22122 15748 22126 15804
rect 22126 15748 22182 15804
rect 22182 15748 22186 15804
rect 22122 15744 22186 15748
rect 9324 15260 9388 15264
rect 9324 15204 9328 15260
rect 9328 15204 9384 15260
rect 9384 15204 9388 15260
rect 9324 15200 9388 15204
rect 9404 15260 9468 15264
rect 9404 15204 9408 15260
rect 9408 15204 9464 15260
rect 9464 15204 9468 15260
rect 9404 15200 9468 15204
rect 9484 15260 9548 15264
rect 9484 15204 9488 15260
rect 9488 15204 9544 15260
rect 9544 15204 9548 15260
rect 9484 15200 9548 15204
rect 9564 15260 9628 15264
rect 9564 15204 9568 15260
rect 9568 15204 9624 15260
rect 9624 15204 9628 15260
rect 9564 15200 9628 15204
rect 17696 15260 17760 15264
rect 17696 15204 17700 15260
rect 17700 15204 17756 15260
rect 17756 15204 17760 15260
rect 17696 15200 17760 15204
rect 17776 15260 17840 15264
rect 17776 15204 17780 15260
rect 17780 15204 17836 15260
rect 17836 15204 17840 15260
rect 17776 15200 17840 15204
rect 17856 15260 17920 15264
rect 17856 15204 17860 15260
rect 17860 15204 17916 15260
rect 17916 15204 17920 15260
rect 17856 15200 17920 15204
rect 17936 15260 18000 15264
rect 17936 15204 17940 15260
rect 17940 15204 17996 15260
rect 17996 15204 18000 15260
rect 17936 15200 18000 15204
rect 9076 14724 9140 14788
rect 12020 14784 12084 14788
rect 12020 14728 12070 14784
rect 12070 14728 12084 14784
rect 12020 14724 12084 14728
rect 5138 14716 5202 14720
rect 5138 14660 5142 14716
rect 5142 14660 5198 14716
rect 5198 14660 5202 14716
rect 5138 14656 5202 14660
rect 5218 14716 5282 14720
rect 5218 14660 5222 14716
rect 5222 14660 5278 14716
rect 5278 14660 5282 14716
rect 5218 14656 5282 14660
rect 5298 14716 5362 14720
rect 5298 14660 5302 14716
rect 5302 14660 5358 14716
rect 5358 14660 5362 14716
rect 5298 14656 5362 14660
rect 5378 14716 5442 14720
rect 5378 14660 5382 14716
rect 5382 14660 5438 14716
rect 5438 14660 5442 14716
rect 5378 14656 5442 14660
rect 13510 14716 13574 14720
rect 13510 14660 13514 14716
rect 13514 14660 13570 14716
rect 13570 14660 13574 14716
rect 13510 14656 13574 14660
rect 13590 14716 13654 14720
rect 13590 14660 13594 14716
rect 13594 14660 13650 14716
rect 13650 14660 13654 14716
rect 13590 14656 13654 14660
rect 13670 14716 13734 14720
rect 13670 14660 13674 14716
rect 13674 14660 13730 14716
rect 13730 14660 13734 14716
rect 13670 14656 13734 14660
rect 13750 14716 13814 14720
rect 13750 14660 13754 14716
rect 13754 14660 13810 14716
rect 13810 14660 13814 14716
rect 13750 14656 13814 14660
rect 21882 14716 21946 14720
rect 21882 14660 21886 14716
rect 21886 14660 21942 14716
rect 21942 14660 21946 14716
rect 21882 14656 21946 14660
rect 21962 14716 22026 14720
rect 21962 14660 21966 14716
rect 21966 14660 22022 14716
rect 22022 14660 22026 14716
rect 21962 14656 22026 14660
rect 22042 14716 22106 14720
rect 22042 14660 22046 14716
rect 22046 14660 22102 14716
rect 22102 14660 22106 14716
rect 22042 14656 22106 14660
rect 22122 14716 22186 14720
rect 22122 14660 22126 14716
rect 22126 14660 22182 14716
rect 22182 14660 22186 14716
rect 22122 14656 22186 14660
rect 9324 14172 9388 14176
rect 9324 14116 9328 14172
rect 9328 14116 9384 14172
rect 9384 14116 9388 14172
rect 9324 14112 9388 14116
rect 9404 14172 9468 14176
rect 9404 14116 9408 14172
rect 9408 14116 9464 14172
rect 9464 14116 9468 14172
rect 9404 14112 9468 14116
rect 9484 14172 9548 14176
rect 9484 14116 9488 14172
rect 9488 14116 9544 14172
rect 9544 14116 9548 14172
rect 9484 14112 9548 14116
rect 9564 14172 9628 14176
rect 9564 14116 9568 14172
rect 9568 14116 9624 14172
rect 9624 14116 9628 14172
rect 9564 14112 9628 14116
rect 17696 14172 17760 14176
rect 17696 14116 17700 14172
rect 17700 14116 17756 14172
rect 17756 14116 17760 14172
rect 17696 14112 17760 14116
rect 17776 14172 17840 14176
rect 17776 14116 17780 14172
rect 17780 14116 17836 14172
rect 17836 14116 17840 14172
rect 17776 14112 17840 14116
rect 17856 14172 17920 14176
rect 17856 14116 17860 14172
rect 17860 14116 17916 14172
rect 17916 14116 17920 14172
rect 17856 14112 17920 14116
rect 17936 14172 18000 14176
rect 17936 14116 17940 14172
rect 17940 14116 17996 14172
rect 17996 14116 18000 14172
rect 17936 14112 18000 14116
rect 5138 13628 5202 13632
rect 5138 13572 5142 13628
rect 5142 13572 5198 13628
rect 5198 13572 5202 13628
rect 5138 13568 5202 13572
rect 5218 13628 5282 13632
rect 5218 13572 5222 13628
rect 5222 13572 5278 13628
rect 5278 13572 5282 13628
rect 5218 13568 5282 13572
rect 5298 13628 5362 13632
rect 5298 13572 5302 13628
rect 5302 13572 5358 13628
rect 5358 13572 5362 13628
rect 5298 13568 5362 13572
rect 5378 13628 5442 13632
rect 5378 13572 5382 13628
rect 5382 13572 5438 13628
rect 5438 13572 5442 13628
rect 5378 13568 5442 13572
rect 13510 13628 13574 13632
rect 13510 13572 13514 13628
rect 13514 13572 13570 13628
rect 13570 13572 13574 13628
rect 13510 13568 13574 13572
rect 13590 13628 13654 13632
rect 13590 13572 13594 13628
rect 13594 13572 13650 13628
rect 13650 13572 13654 13628
rect 13590 13568 13654 13572
rect 13670 13628 13734 13632
rect 13670 13572 13674 13628
rect 13674 13572 13730 13628
rect 13730 13572 13734 13628
rect 13670 13568 13734 13572
rect 13750 13628 13814 13632
rect 13750 13572 13754 13628
rect 13754 13572 13810 13628
rect 13810 13572 13814 13628
rect 13750 13568 13814 13572
rect 21882 13628 21946 13632
rect 21882 13572 21886 13628
rect 21886 13572 21942 13628
rect 21942 13572 21946 13628
rect 21882 13568 21946 13572
rect 21962 13628 22026 13632
rect 21962 13572 21966 13628
rect 21966 13572 22022 13628
rect 22022 13572 22026 13628
rect 21962 13568 22026 13572
rect 22042 13628 22106 13632
rect 22042 13572 22046 13628
rect 22046 13572 22102 13628
rect 22102 13572 22106 13628
rect 22042 13568 22106 13572
rect 22122 13628 22186 13632
rect 22122 13572 22126 13628
rect 22126 13572 22182 13628
rect 22182 13572 22186 13628
rect 22122 13568 22186 13572
rect 16804 13228 16868 13292
rect 9324 13084 9388 13088
rect 9324 13028 9328 13084
rect 9328 13028 9384 13084
rect 9384 13028 9388 13084
rect 9324 13024 9388 13028
rect 9404 13084 9468 13088
rect 9404 13028 9408 13084
rect 9408 13028 9464 13084
rect 9464 13028 9468 13084
rect 9404 13024 9468 13028
rect 9484 13084 9548 13088
rect 9484 13028 9488 13084
rect 9488 13028 9544 13084
rect 9544 13028 9548 13084
rect 9484 13024 9548 13028
rect 9564 13084 9628 13088
rect 9564 13028 9568 13084
rect 9568 13028 9624 13084
rect 9624 13028 9628 13084
rect 9564 13024 9628 13028
rect 17696 13084 17760 13088
rect 17696 13028 17700 13084
rect 17700 13028 17756 13084
rect 17756 13028 17760 13084
rect 17696 13024 17760 13028
rect 17776 13084 17840 13088
rect 17776 13028 17780 13084
rect 17780 13028 17836 13084
rect 17836 13028 17840 13084
rect 17776 13024 17840 13028
rect 17856 13084 17920 13088
rect 17856 13028 17860 13084
rect 17860 13028 17916 13084
rect 17916 13028 17920 13084
rect 17856 13024 17920 13028
rect 17936 13084 18000 13088
rect 17936 13028 17940 13084
rect 17940 13028 17996 13084
rect 17996 13028 18000 13084
rect 17936 13024 18000 13028
rect 8708 12820 8772 12884
rect 5138 12540 5202 12544
rect 5138 12484 5142 12540
rect 5142 12484 5198 12540
rect 5198 12484 5202 12540
rect 5138 12480 5202 12484
rect 5218 12540 5282 12544
rect 5218 12484 5222 12540
rect 5222 12484 5278 12540
rect 5278 12484 5282 12540
rect 5218 12480 5282 12484
rect 5298 12540 5362 12544
rect 5298 12484 5302 12540
rect 5302 12484 5358 12540
rect 5358 12484 5362 12540
rect 5298 12480 5362 12484
rect 5378 12540 5442 12544
rect 5378 12484 5382 12540
rect 5382 12484 5438 12540
rect 5438 12484 5442 12540
rect 5378 12480 5442 12484
rect 13510 12540 13574 12544
rect 13510 12484 13514 12540
rect 13514 12484 13570 12540
rect 13570 12484 13574 12540
rect 13510 12480 13574 12484
rect 13590 12540 13654 12544
rect 13590 12484 13594 12540
rect 13594 12484 13650 12540
rect 13650 12484 13654 12540
rect 13590 12480 13654 12484
rect 13670 12540 13734 12544
rect 13670 12484 13674 12540
rect 13674 12484 13730 12540
rect 13730 12484 13734 12540
rect 13670 12480 13734 12484
rect 13750 12540 13814 12544
rect 13750 12484 13754 12540
rect 13754 12484 13810 12540
rect 13810 12484 13814 12540
rect 13750 12480 13814 12484
rect 21882 12540 21946 12544
rect 21882 12484 21886 12540
rect 21886 12484 21942 12540
rect 21942 12484 21946 12540
rect 21882 12480 21946 12484
rect 21962 12540 22026 12544
rect 21962 12484 21966 12540
rect 21966 12484 22022 12540
rect 22022 12484 22026 12540
rect 21962 12480 22026 12484
rect 22042 12540 22106 12544
rect 22042 12484 22046 12540
rect 22046 12484 22102 12540
rect 22102 12484 22106 12540
rect 22042 12480 22106 12484
rect 22122 12540 22186 12544
rect 22122 12484 22126 12540
rect 22126 12484 22182 12540
rect 22182 12484 22186 12540
rect 22122 12480 22186 12484
rect 22508 12336 22572 12340
rect 22508 12280 22522 12336
rect 22522 12280 22572 12336
rect 22508 12276 22572 12280
rect 9324 11996 9388 12000
rect 9324 11940 9328 11996
rect 9328 11940 9384 11996
rect 9384 11940 9388 11996
rect 9324 11936 9388 11940
rect 9404 11996 9468 12000
rect 9404 11940 9408 11996
rect 9408 11940 9464 11996
rect 9464 11940 9468 11996
rect 9404 11936 9468 11940
rect 9484 11996 9548 12000
rect 9484 11940 9488 11996
rect 9488 11940 9544 11996
rect 9544 11940 9548 11996
rect 9484 11936 9548 11940
rect 9564 11996 9628 12000
rect 9564 11940 9568 11996
rect 9568 11940 9624 11996
rect 9624 11940 9628 11996
rect 9564 11936 9628 11940
rect 17696 11996 17760 12000
rect 17696 11940 17700 11996
rect 17700 11940 17756 11996
rect 17756 11940 17760 11996
rect 17696 11936 17760 11940
rect 17776 11996 17840 12000
rect 17776 11940 17780 11996
rect 17780 11940 17836 11996
rect 17836 11940 17840 11996
rect 17776 11936 17840 11940
rect 17856 11996 17920 12000
rect 17856 11940 17860 11996
rect 17860 11940 17916 11996
rect 17916 11940 17920 11996
rect 17856 11936 17920 11940
rect 17936 11996 18000 12000
rect 17936 11940 17940 11996
rect 17940 11940 17996 11996
rect 17996 11940 18000 11996
rect 17936 11936 18000 11940
rect 5138 11452 5202 11456
rect 5138 11396 5142 11452
rect 5142 11396 5198 11452
rect 5198 11396 5202 11452
rect 5138 11392 5202 11396
rect 5218 11452 5282 11456
rect 5218 11396 5222 11452
rect 5222 11396 5278 11452
rect 5278 11396 5282 11452
rect 5218 11392 5282 11396
rect 5298 11452 5362 11456
rect 5298 11396 5302 11452
rect 5302 11396 5358 11452
rect 5358 11396 5362 11452
rect 5298 11392 5362 11396
rect 5378 11452 5442 11456
rect 5378 11396 5382 11452
rect 5382 11396 5438 11452
rect 5438 11396 5442 11452
rect 5378 11392 5442 11396
rect 13510 11452 13574 11456
rect 13510 11396 13514 11452
rect 13514 11396 13570 11452
rect 13570 11396 13574 11452
rect 13510 11392 13574 11396
rect 13590 11452 13654 11456
rect 13590 11396 13594 11452
rect 13594 11396 13650 11452
rect 13650 11396 13654 11452
rect 13590 11392 13654 11396
rect 13670 11452 13734 11456
rect 13670 11396 13674 11452
rect 13674 11396 13730 11452
rect 13730 11396 13734 11452
rect 13670 11392 13734 11396
rect 13750 11452 13814 11456
rect 13750 11396 13754 11452
rect 13754 11396 13810 11452
rect 13810 11396 13814 11452
rect 13750 11392 13814 11396
rect 21882 11452 21946 11456
rect 21882 11396 21886 11452
rect 21886 11396 21942 11452
rect 21942 11396 21946 11452
rect 21882 11392 21946 11396
rect 21962 11452 22026 11456
rect 21962 11396 21966 11452
rect 21966 11396 22022 11452
rect 22022 11396 22026 11452
rect 21962 11392 22026 11396
rect 22042 11452 22106 11456
rect 22042 11396 22046 11452
rect 22046 11396 22102 11452
rect 22102 11396 22106 11452
rect 22042 11392 22106 11396
rect 22122 11452 22186 11456
rect 22122 11396 22126 11452
rect 22126 11396 22182 11452
rect 22182 11396 22186 11452
rect 22122 11392 22186 11396
rect 9324 10908 9388 10912
rect 9324 10852 9328 10908
rect 9328 10852 9384 10908
rect 9384 10852 9388 10908
rect 9324 10848 9388 10852
rect 9404 10908 9468 10912
rect 9404 10852 9408 10908
rect 9408 10852 9464 10908
rect 9464 10852 9468 10908
rect 9404 10848 9468 10852
rect 9484 10908 9548 10912
rect 9484 10852 9488 10908
rect 9488 10852 9544 10908
rect 9544 10852 9548 10908
rect 9484 10848 9548 10852
rect 9564 10908 9628 10912
rect 9564 10852 9568 10908
rect 9568 10852 9624 10908
rect 9624 10852 9628 10908
rect 9564 10848 9628 10852
rect 17696 10908 17760 10912
rect 17696 10852 17700 10908
rect 17700 10852 17756 10908
rect 17756 10852 17760 10908
rect 17696 10848 17760 10852
rect 17776 10908 17840 10912
rect 17776 10852 17780 10908
rect 17780 10852 17836 10908
rect 17836 10852 17840 10908
rect 17776 10848 17840 10852
rect 17856 10908 17920 10912
rect 17856 10852 17860 10908
rect 17860 10852 17916 10908
rect 17916 10852 17920 10908
rect 17856 10848 17920 10852
rect 17936 10908 18000 10912
rect 17936 10852 17940 10908
rect 17940 10852 17996 10908
rect 17996 10852 18000 10908
rect 17936 10848 18000 10852
rect 5138 10364 5202 10368
rect 5138 10308 5142 10364
rect 5142 10308 5198 10364
rect 5198 10308 5202 10364
rect 5138 10304 5202 10308
rect 5218 10364 5282 10368
rect 5218 10308 5222 10364
rect 5222 10308 5278 10364
rect 5278 10308 5282 10364
rect 5218 10304 5282 10308
rect 5298 10364 5362 10368
rect 5298 10308 5302 10364
rect 5302 10308 5358 10364
rect 5358 10308 5362 10364
rect 5298 10304 5362 10308
rect 5378 10364 5442 10368
rect 5378 10308 5382 10364
rect 5382 10308 5438 10364
rect 5438 10308 5442 10364
rect 5378 10304 5442 10308
rect 13510 10364 13574 10368
rect 13510 10308 13514 10364
rect 13514 10308 13570 10364
rect 13570 10308 13574 10364
rect 13510 10304 13574 10308
rect 13590 10364 13654 10368
rect 13590 10308 13594 10364
rect 13594 10308 13650 10364
rect 13650 10308 13654 10364
rect 13590 10304 13654 10308
rect 13670 10364 13734 10368
rect 13670 10308 13674 10364
rect 13674 10308 13730 10364
rect 13730 10308 13734 10364
rect 13670 10304 13734 10308
rect 13750 10364 13814 10368
rect 13750 10308 13754 10364
rect 13754 10308 13810 10364
rect 13810 10308 13814 10364
rect 13750 10304 13814 10308
rect 21882 10364 21946 10368
rect 21882 10308 21886 10364
rect 21886 10308 21942 10364
rect 21942 10308 21946 10364
rect 21882 10304 21946 10308
rect 21962 10364 22026 10368
rect 21962 10308 21966 10364
rect 21966 10308 22022 10364
rect 22022 10308 22026 10364
rect 21962 10304 22026 10308
rect 22042 10364 22106 10368
rect 22042 10308 22046 10364
rect 22046 10308 22102 10364
rect 22102 10308 22106 10364
rect 22042 10304 22106 10308
rect 22122 10364 22186 10368
rect 22122 10308 22126 10364
rect 22126 10308 22182 10364
rect 22182 10308 22186 10364
rect 22122 10304 22186 10308
rect 9324 9820 9388 9824
rect 9324 9764 9328 9820
rect 9328 9764 9384 9820
rect 9384 9764 9388 9820
rect 9324 9760 9388 9764
rect 9404 9820 9468 9824
rect 9404 9764 9408 9820
rect 9408 9764 9464 9820
rect 9464 9764 9468 9820
rect 9404 9760 9468 9764
rect 9484 9820 9548 9824
rect 9484 9764 9488 9820
rect 9488 9764 9544 9820
rect 9544 9764 9548 9820
rect 9484 9760 9548 9764
rect 9564 9820 9628 9824
rect 9564 9764 9568 9820
rect 9568 9764 9624 9820
rect 9624 9764 9628 9820
rect 9564 9760 9628 9764
rect 17696 9820 17760 9824
rect 17696 9764 17700 9820
rect 17700 9764 17756 9820
rect 17756 9764 17760 9820
rect 17696 9760 17760 9764
rect 17776 9820 17840 9824
rect 17776 9764 17780 9820
rect 17780 9764 17836 9820
rect 17836 9764 17840 9820
rect 17776 9760 17840 9764
rect 17856 9820 17920 9824
rect 17856 9764 17860 9820
rect 17860 9764 17916 9820
rect 17916 9764 17920 9820
rect 17856 9760 17920 9764
rect 17936 9820 18000 9824
rect 17936 9764 17940 9820
rect 17940 9764 17996 9820
rect 17996 9764 18000 9820
rect 17936 9760 18000 9764
rect 5138 9276 5202 9280
rect 5138 9220 5142 9276
rect 5142 9220 5198 9276
rect 5198 9220 5202 9276
rect 5138 9216 5202 9220
rect 5218 9276 5282 9280
rect 5218 9220 5222 9276
rect 5222 9220 5278 9276
rect 5278 9220 5282 9276
rect 5218 9216 5282 9220
rect 5298 9276 5362 9280
rect 5298 9220 5302 9276
rect 5302 9220 5358 9276
rect 5358 9220 5362 9276
rect 5298 9216 5362 9220
rect 5378 9276 5442 9280
rect 5378 9220 5382 9276
rect 5382 9220 5438 9276
rect 5438 9220 5442 9276
rect 5378 9216 5442 9220
rect 13510 9276 13574 9280
rect 13510 9220 13514 9276
rect 13514 9220 13570 9276
rect 13570 9220 13574 9276
rect 13510 9216 13574 9220
rect 13590 9276 13654 9280
rect 13590 9220 13594 9276
rect 13594 9220 13650 9276
rect 13650 9220 13654 9276
rect 13590 9216 13654 9220
rect 13670 9276 13734 9280
rect 13670 9220 13674 9276
rect 13674 9220 13730 9276
rect 13730 9220 13734 9276
rect 13670 9216 13734 9220
rect 13750 9276 13814 9280
rect 13750 9220 13754 9276
rect 13754 9220 13810 9276
rect 13810 9220 13814 9276
rect 13750 9216 13814 9220
rect 21882 9276 21946 9280
rect 21882 9220 21886 9276
rect 21886 9220 21942 9276
rect 21942 9220 21946 9276
rect 21882 9216 21946 9220
rect 21962 9276 22026 9280
rect 21962 9220 21966 9276
rect 21966 9220 22022 9276
rect 22022 9220 22026 9276
rect 21962 9216 22026 9220
rect 22042 9276 22106 9280
rect 22042 9220 22046 9276
rect 22046 9220 22102 9276
rect 22102 9220 22106 9276
rect 22042 9216 22106 9220
rect 22122 9276 22186 9280
rect 22122 9220 22126 9276
rect 22126 9220 22182 9276
rect 22182 9220 22186 9276
rect 22122 9216 22186 9220
rect 9324 8732 9388 8736
rect 9324 8676 9328 8732
rect 9328 8676 9384 8732
rect 9384 8676 9388 8732
rect 9324 8672 9388 8676
rect 9404 8732 9468 8736
rect 9404 8676 9408 8732
rect 9408 8676 9464 8732
rect 9464 8676 9468 8732
rect 9404 8672 9468 8676
rect 9484 8732 9548 8736
rect 9484 8676 9488 8732
rect 9488 8676 9544 8732
rect 9544 8676 9548 8732
rect 9484 8672 9548 8676
rect 9564 8732 9628 8736
rect 9564 8676 9568 8732
rect 9568 8676 9624 8732
rect 9624 8676 9628 8732
rect 9564 8672 9628 8676
rect 17696 8732 17760 8736
rect 17696 8676 17700 8732
rect 17700 8676 17756 8732
rect 17756 8676 17760 8732
rect 17696 8672 17760 8676
rect 17776 8732 17840 8736
rect 17776 8676 17780 8732
rect 17780 8676 17836 8732
rect 17836 8676 17840 8732
rect 17776 8672 17840 8676
rect 17856 8732 17920 8736
rect 17856 8676 17860 8732
rect 17860 8676 17916 8732
rect 17916 8676 17920 8732
rect 17856 8672 17920 8676
rect 17936 8732 18000 8736
rect 17936 8676 17940 8732
rect 17940 8676 17996 8732
rect 17996 8676 18000 8732
rect 17936 8672 18000 8676
rect 5138 8188 5202 8192
rect 5138 8132 5142 8188
rect 5142 8132 5198 8188
rect 5198 8132 5202 8188
rect 5138 8128 5202 8132
rect 5218 8188 5282 8192
rect 5218 8132 5222 8188
rect 5222 8132 5278 8188
rect 5278 8132 5282 8188
rect 5218 8128 5282 8132
rect 5298 8188 5362 8192
rect 5298 8132 5302 8188
rect 5302 8132 5358 8188
rect 5358 8132 5362 8188
rect 5298 8128 5362 8132
rect 5378 8188 5442 8192
rect 5378 8132 5382 8188
rect 5382 8132 5438 8188
rect 5438 8132 5442 8188
rect 5378 8128 5442 8132
rect 13510 8188 13574 8192
rect 13510 8132 13514 8188
rect 13514 8132 13570 8188
rect 13570 8132 13574 8188
rect 13510 8128 13574 8132
rect 13590 8188 13654 8192
rect 13590 8132 13594 8188
rect 13594 8132 13650 8188
rect 13650 8132 13654 8188
rect 13590 8128 13654 8132
rect 13670 8188 13734 8192
rect 13670 8132 13674 8188
rect 13674 8132 13730 8188
rect 13730 8132 13734 8188
rect 13670 8128 13734 8132
rect 13750 8188 13814 8192
rect 13750 8132 13754 8188
rect 13754 8132 13810 8188
rect 13810 8132 13814 8188
rect 13750 8128 13814 8132
rect 21882 8188 21946 8192
rect 21882 8132 21886 8188
rect 21886 8132 21942 8188
rect 21942 8132 21946 8188
rect 21882 8128 21946 8132
rect 21962 8188 22026 8192
rect 21962 8132 21966 8188
rect 21966 8132 22022 8188
rect 22022 8132 22026 8188
rect 21962 8128 22026 8132
rect 22042 8188 22106 8192
rect 22042 8132 22046 8188
rect 22046 8132 22102 8188
rect 22102 8132 22106 8188
rect 22042 8128 22106 8132
rect 22122 8188 22186 8192
rect 22122 8132 22126 8188
rect 22126 8132 22182 8188
rect 22182 8132 22186 8188
rect 22122 8128 22186 8132
rect 9324 7644 9388 7648
rect 9324 7588 9328 7644
rect 9328 7588 9384 7644
rect 9384 7588 9388 7644
rect 9324 7584 9388 7588
rect 9404 7644 9468 7648
rect 9404 7588 9408 7644
rect 9408 7588 9464 7644
rect 9464 7588 9468 7644
rect 9404 7584 9468 7588
rect 9484 7644 9548 7648
rect 9484 7588 9488 7644
rect 9488 7588 9544 7644
rect 9544 7588 9548 7644
rect 9484 7584 9548 7588
rect 9564 7644 9628 7648
rect 9564 7588 9568 7644
rect 9568 7588 9624 7644
rect 9624 7588 9628 7644
rect 9564 7584 9628 7588
rect 17696 7644 17760 7648
rect 17696 7588 17700 7644
rect 17700 7588 17756 7644
rect 17756 7588 17760 7644
rect 17696 7584 17760 7588
rect 17776 7644 17840 7648
rect 17776 7588 17780 7644
rect 17780 7588 17836 7644
rect 17836 7588 17840 7644
rect 17776 7584 17840 7588
rect 17856 7644 17920 7648
rect 17856 7588 17860 7644
rect 17860 7588 17916 7644
rect 17916 7588 17920 7644
rect 17856 7584 17920 7588
rect 17936 7644 18000 7648
rect 17936 7588 17940 7644
rect 17940 7588 17996 7644
rect 17996 7588 18000 7644
rect 17936 7584 18000 7588
rect 5138 7100 5202 7104
rect 5138 7044 5142 7100
rect 5142 7044 5198 7100
rect 5198 7044 5202 7100
rect 5138 7040 5202 7044
rect 5218 7100 5282 7104
rect 5218 7044 5222 7100
rect 5222 7044 5278 7100
rect 5278 7044 5282 7100
rect 5218 7040 5282 7044
rect 5298 7100 5362 7104
rect 5298 7044 5302 7100
rect 5302 7044 5358 7100
rect 5358 7044 5362 7100
rect 5298 7040 5362 7044
rect 5378 7100 5442 7104
rect 5378 7044 5382 7100
rect 5382 7044 5438 7100
rect 5438 7044 5442 7100
rect 5378 7040 5442 7044
rect 13510 7100 13574 7104
rect 13510 7044 13514 7100
rect 13514 7044 13570 7100
rect 13570 7044 13574 7100
rect 13510 7040 13574 7044
rect 13590 7100 13654 7104
rect 13590 7044 13594 7100
rect 13594 7044 13650 7100
rect 13650 7044 13654 7100
rect 13590 7040 13654 7044
rect 13670 7100 13734 7104
rect 13670 7044 13674 7100
rect 13674 7044 13730 7100
rect 13730 7044 13734 7100
rect 13670 7040 13734 7044
rect 13750 7100 13814 7104
rect 13750 7044 13754 7100
rect 13754 7044 13810 7100
rect 13810 7044 13814 7100
rect 13750 7040 13814 7044
rect 21882 7100 21946 7104
rect 21882 7044 21886 7100
rect 21886 7044 21942 7100
rect 21942 7044 21946 7100
rect 21882 7040 21946 7044
rect 21962 7100 22026 7104
rect 21962 7044 21966 7100
rect 21966 7044 22022 7100
rect 22022 7044 22026 7100
rect 21962 7040 22026 7044
rect 22042 7100 22106 7104
rect 22042 7044 22046 7100
rect 22046 7044 22102 7100
rect 22102 7044 22106 7100
rect 22042 7040 22106 7044
rect 22122 7100 22186 7104
rect 22122 7044 22126 7100
rect 22126 7044 22182 7100
rect 22182 7044 22186 7100
rect 22122 7040 22186 7044
rect 11100 6972 11164 7036
rect 9324 6556 9388 6560
rect 9324 6500 9328 6556
rect 9328 6500 9384 6556
rect 9384 6500 9388 6556
rect 9324 6496 9388 6500
rect 9404 6556 9468 6560
rect 9404 6500 9408 6556
rect 9408 6500 9464 6556
rect 9464 6500 9468 6556
rect 9404 6496 9468 6500
rect 9484 6556 9548 6560
rect 9484 6500 9488 6556
rect 9488 6500 9544 6556
rect 9544 6500 9548 6556
rect 9484 6496 9548 6500
rect 9564 6556 9628 6560
rect 9564 6500 9568 6556
rect 9568 6500 9624 6556
rect 9624 6500 9628 6556
rect 9564 6496 9628 6500
rect 17696 6556 17760 6560
rect 17696 6500 17700 6556
rect 17700 6500 17756 6556
rect 17756 6500 17760 6556
rect 17696 6496 17760 6500
rect 17776 6556 17840 6560
rect 17776 6500 17780 6556
rect 17780 6500 17836 6556
rect 17836 6500 17840 6556
rect 17776 6496 17840 6500
rect 17856 6556 17920 6560
rect 17856 6500 17860 6556
rect 17860 6500 17916 6556
rect 17916 6500 17920 6556
rect 17856 6496 17920 6500
rect 17936 6556 18000 6560
rect 17936 6500 17940 6556
rect 17940 6500 17996 6556
rect 17996 6500 18000 6556
rect 17936 6496 18000 6500
rect 5138 6012 5202 6016
rect 5138 5956 5142 6012
rect 5142 5956 5198 6012
rect 5198 5956 5202 6012
rect 5138 5952 5202 5956
rect 5218 6012 5282 6016
rect 5218 5956 5222 6012
rect 5222 5956 5278 6012
rect 5278 5956 5282 6012
rect 5218 5952 5282 5956
rect 5298 6012 5362 6016
rect 5298 5956 5302 6012
rect 5302 5956 5358 6012
rect 5358 5956 5362 6012
rect 5298 5952 5362 5956
rect 5378 6012 5442 6016
rect 5378 5956 5382 6012
rect 5382 5956 5438 6012
rect 5438 5956 5442 6012
rect 5378 5952 5442 5956
rect 13510 6012 13574 6016
rect 13510 5956 13514 6012
rect 13514 5956 13570 6012
rect 13570 5956 13574 6012
rect 13510 5952 13574 5956
rect 13590 6012 13654 6016
rect 13590 5956 13594 6012
rect 13594 5956 13650 6012
rect 13650 5956 13654 6012
rect 13590 5952 13654 5956
rect 13670 6012 13734 6016
rect 13670 5956 13674 6012
rect 13674 5956 13730 6012
rect 13730 5956 13734 6012
rect 13670 5952 13734 5956
rect 13750 6012 13814 6016
rect 13750 5956 13754 6012
rect 13754 5956 13810 6012
rect 13810 5956 13814 6012
rect 13750 5952 13814 5956
rect 21882 6012 21946 6016
rect 21882 5956 21886 6012
rect 21886 5956 21942 6012
rect 21942 5956 21946 6012
rect 21882 5952 21946 5956
rect 21962 6012 22026 6016
rect 21962 5956 21966 6012
rect 21966 5956 22022 6012
rect 22022 5956 22026 6012
rect 21962 5952 22026 5956
rect 22042 6012 22106 6016
rect 22042 5956 22046 6012
rect 22046 5956 22102 6012
rect 22102 5956 22106 6012
rect 22042 5952 22106 5956
rect 22122 6012 22186 6016
rect 22122 5956 22126 6012
rect 22126 5956 22182 6012
rect 22182 5956 22186 6012
rect 22122 5952 22186 5956
rect 9324 5468 9388 5472
rect 9324 5412 9328 5468
rect 9328 5412 9384 5468
rect 9384 5412 9388 5468
rect 9324 5408 9388 5412
rect 9404 5468 9468 5472
rect 9404 5412 9408 5468
rect 9408 5412 9464 5468
rect 9464 5412 9468 5468
rect 9404 5408 9468 5412
rect 9484 5468 9548 5472
rect 9484 5412 9488 5468
rect 9488 5412 9544 5468
rect 9544 5412 9548 5468
rect 9484 5408 9548 5412
rect 9564 5468 9628 5472
rect 9564 5412 9568 5468
rect 9568 5412 9624 5468
rect 9624 5412 9628 5468
rect 9564 5408 9628 5412
rect 17696 5468 17760 5472
rect 17696 5412 17700 5468
rect 17700 5412 17756 5468
rect 17756 5412 17760 5468
rect 17696 5408 17760 5412
rect 17776 5468 17840 5472
rect 17776 5412 17780 5468
rect 17780 5412 17836 5468
rect 17836 5412 17840 5468
rect 17776 5408 17840 5412
rect 17856 5468 17920 5472
rect 17856 5412 17860 5468
rect 17860 5412 17916 5468
rect 17916 5412 17920 5468
rect 17856 5408 17920 5412
rect 17936 5468 18000 5472
rect 17936 5412 17940 5468
rect 17940 5412 17996 5468
rect 17996 5412 18000 5468
rect 17936 5408 18000 5412
rect 5138 4924 5202 4928
rect 5138 4868 5142 4924
rect 5142 4868 5198 4924
rect 5198 4868 5202 4924
rect 5138 4864 5202 4868
rect 5218 4924 5282 4928
rect 5218 4868 5222 4924
rect 5222 4868 5278 4924
rect 5278 4868 5282 4924
rect 5218 4864 5282 4868
rect 5298 4924 5362 4928
rect 5298 4868 5302 4924
rect 5302 4868 5358 4924
rect 5358 4868 5362 4924
rect 5298 4864 5362 4868
rect 5378 4924 5442 4928
rect 5378 4868 5382 4924
rect 5382 4868 5438 4924
rect 5438 4868 5442 4924
rect 5378 4864 5442 4868
rect 13510 4924 13574 4928
rect 13510 4868 13514 4924
rect 13514 4868 13570 4924
rect 13570 4868 13574 4924
rect 13510 4864 13574 4868
rect 13590 4924 13654 4928
rect 13590 4868 13594 4924
rect 13594 4868 13650 4924
rect 13650 4868 13654 4924
rect 13590 4864 13654 4868
rect 13670 4924 13734 4928
rect 13670 4868 13674 4924
rect 13674 4868 13730 4924
rect 13730 4868 13734 4924
rect 13670 4864 13734 4868
rect 13750 4924 13814 4928
rect 13750 4868 13754 4924
rect 13754 4868 13810 4924
rect 13810 4868 13814 4924
rect 13750 4864 13814 4868
rect 21882 4924 21946 4928
rect 21882 4868 21886 4924
rect 21886 4868 21942 4924
rect 21942 4868 21946 4924
rect 21882 4864 21946 4868
rect 21962 4924 22026 4928
rect 21962 4868 21966 4924
rect 21966 4868 22022 4924
rect 22022 4868 22026 4924
rect 21962 4864 22026 4868
rect 22042 4924 22106 4928
rect 22042 4868 22046 4924
rect 22046 4868 22102 4924
rect 22102 4868 22106 4924
rect 22042 4864 22106 4868
rect 22122 4924 22186 4928
rect 22122 4868 22126 4924
rect 22126 4868 22182 4924
rect 22182 4868 22186 4924
rect 22122 4864 22186 4868
rect 11100 4796 11164 4860
rect 9076 4524 9140 4588
rect 9324 4380 9388 4384
rect 9324 4324 9328 4380
rect 9328 4324 9384 4380
rect 9384 4324 9388 4380
rect 9324 4320 9388 4324
rect 9404 4380 9468 4384
rect 9404 4324 9408 4380
rect 9408 4324 9464 4380
rect 9464 4324 9468 4380
rect 9404 4320 9468 4324
rect 9484 4380 9548 4384
rect 9484 4324 9488 4380
rect 9488 4324 9544 4380
rect 9544 4324 9548 4380
rect 9484 4320 9548 4324
rect 9564 4380 9628 4384
rect 9564 4324 9568 4380
rect 9568 4324 9624 4380
rect 9624 4324 9628 4380
rect 9564 4320 9628 4324
rect 17696 4380 17760 4384
rect 17696 4324 17700 4380
rect 17700 4324 17756 4380
rect 17756 4324 17760 4380
rect 17696 4320 17760 4324
rect 17776 4380 17840 4384
rect 17776 4324 17780 4380
rect 17780 4324 17836 4380
rect 17836 4324 17840 4380
rect 17776 4320 17840 4324
rect 17856 4380 17920 4384
rect 17856 4324 17860 4380
rect 17860 4324 17916 4380
rect 17916 4324 17920 4380
rect 17856 4320 17920 4324
rect 17936 4380 18000 4384
rect 17936 4324 17940 4380
rect 17940 4324 17996 4380
rect 17996 4324 18000 4380
rect 17936 4320 18000 4324
rect 16804 3980 16868 4044
rect 16988 3980 17052 4044
rect 5138 3836 5202 3840
rect 5138 3780 5142 3836
rect 5142 3780 5198 3836
rect 5198 3780 5202 3836
rect 5138 3776 5202 3780
rect 5218 3836 5282 3840
rect 5218 3780 5222 3836
rect 5222 3780 5278 3836
rect 5278 3780 5282 3836
rect 5218 3776 5282 3780
rect 5298 3836 5362 3840
rect 5298 3780 5302 3836
rect 5302 3780 5358 3836
rect 5358 3780 5362 3836
rect 5298 3776 5362 3780
rect 5378 3836 5442 3840
rect 5378 3780 5382 3836
rect 5382 3780 5438 3836
rect 5438 3780 5442 3836
rect 5378 3776 5442 3780
rect 13510 3836 13574 3840
rect 13510 3780 13514 3836
rect 13514 3780 13570 3836
rect 13570 3780 13574 3836
rect 13510 3776 13574 3780
rect 13590 3836 13654 3840
rect 13590 3780 13594 3836
rect 13594 3780 13650 3836
rect 13650 3780 13654 3836
rect 13590 3776 13654 3780
rect 13670 3836 13734 3840
rect 13670 3780 13674 3836
rect 13674 3780 13730 3836
rect 13730 3780 13734 3836
rect 13670 3776 13734 3780
rect 13750 3836 13814 3840
rect 13750 3780 13754 3836
rect 13754 3780 13810 3836
rect 13810 3780 13814 3836
rect 13750 3776 13814 3780
rect 21882 3836 21946 3840
rect 21882 3780 21886 3836
rect 21886 3780 21942 3836
rect 21942 3780 21946 3836
rect 21882 3776 21946 3780
rect 21962 3836 22026 3840
rect 21962 3780 21966 3836
rect 21966 3780 22022 3836
rect 22022 3780 22026 3836
rect 21962 3776 22026 3780
rect 22042 3836 22106 3840
rect 22042 3780 22046 3836
rect 22046 3780 22102 3836
rect 22102 3780 22106 3836
rect 22042 3776 22106 3780
rect 22122 3836 22186 3840
rect 22122 3780 22126 3836
rect 22126 3780 22182 3836
rect 22182 3780 22186 3836
rect 22122 3776 22186 3780
rect 8892 3632 8956 3636
rect 8892 3576 8906 3632
rect 8906 3576 8956 3632
rect 8892 3572 8956 3576
rect 12020 3436 12084 3500
rect 8708 3300 8772 3364
rect 9324 3292 9388 3296
rect 9324 3236 9328 3292
rect 9328 3236 9384 3292
rect 9384 3236 9388 3292
rect 9324 3232 9388 3236
rect 9404 3292 9468 3296
rect 9404 3236 9408 3292
rect 9408 3236 9464 3292
rect 9464 3236 9468 3292
rect 9404 3232 9468 3236
rect 9484 3292 9548 3296
rect 9484 3236 9488 3292
rect 9488 3236 9544 3292
rect 9544 3236 9548 3292
rect 9484 3232 9548 3236
rect 9564 3292 9628 3296
rect 9564 3236 9568 3292
rect 9568 3236 9624 3292
rect 9624 3236 9628 3292
rect 9564 3232 9628 3236
rect 17696 3292 17760 3296
rect 17696 3236 17700 3292
rect 17700 3236 17756 3292
rect 17756 3236 17760 3292
rect 17696 3232 17760 3236
rect 17776 3292 17840 3296
rect 17776 3236 17780 3292
rect 17780 3236 17836 3292
rect 17836 3236 17840 3292
rect 17776 3232 17840 3236
rect 17856 3292 17920 3296
rect 17856 3236 17860 3292
rect 17860 3236 17916 3292
rect 17916 3236 17920 3292
rect 17856 3232 17920 3236
rect 17936 3292 18000 3296
rect 17936 3236 17940 3292
rect 17940 3236 17996 3292
rect 17996 3236 18000 3292
rect 17936 3232 18000 3236
rect 5138 2748 5202 2752
rect 5138 2692 5142 2748
rect 5142 2692 5198 2748
rect 5198 2692 5202 2748
rect 5138 2688 5202 2692
rect 5218 2748 5282 2752
rect 5218 2692 5222 2748
rect 5222 2692 5278 2748
rect 5278 2692 5282 2748
rect 5218 2688 5282 2692
rect 5298 2748 5362 2752
rect 5298 2692 5302 2748
rect 5302 2692 5358 2748
rect 5358 2692 5362 2748
rect 5298 2688 5362 2692
rect 5378 2748 5442 2752
rect 5378 2692 5382 2748
rect 5382 2692 5438 2748
rect 5438 2692 5442 2748
rect 5378 2688 5442 2692
rect 13510 2748 13574 2752
rect 13510 2692 13514 2748
rect 13514 2692 13570 2748
rect 13570 2692 13574 2748
rect 13510 2688 13574 2692
rect 13590 2748 13654 2752
rect 13590 2692 13594 2748
rect 13594 2692 13650 2748
rect 13650 2692 13654 2748
rect 13590 2688 13654 2692
rect 13670 2748 13734 2752
rect 13670 2692 13674 2748
rect 13674 2692 13730 2748
rect 13730 2692 13734 2748
rect 13670 2688 13734 2692
rect 13750 2748 13814 2752
rect 13750 2692 13754 2748
rect 13754 2692 13810 2748
rect 13810 2692 13814 2748
rect 13750 2688 13814 2692
rect 21882 2748 21946 2752
rect 21882 2692 21886 2748
rect 21886 2692 21942 2748
rect 21942 2692 21946 2748
rect 21882 2688 21946 2692
rect 21962 2748 22026 2752
rect 21962 2692 21966 2748
rect 21966 2692 22022 2748
rect 22022 2692 22026 2748
rect 21962 2688 22026 2692
rect 22042 2748 22106 2752
rect 22042 2692 22046 2748
rect 22046 2692 22102 2748
rect 22102 2692 22106 2748
rect 22042 2688 22106 2692
rect 22122 2748 22186 2752
rect 22122 2692 22126 2748
rect 22126 2692 22182 2748
rect 22182 2692 22186 2748
rect 22122 2688 22186 2692
rect 9324 2204 9388 2208
rect 9324 2148 9328 2204
rect 9328 2148 9384 2204
rect 9384 2148 9388 2204
rect 9324 2144 9388 2148
rect 9404 2204 9468 2208
rect 9404 2148 9408 2204
rect 9408 2148 9464 2204
rect 9464 2148 9468 2204
rect 9404 2144 9468 2148
rect 9484 2204 9548 2208
rect 9484 2148 9488 2204
rect 9488 2148 9544 2204
rect 9544 2148 9548 2204
rect 9484 2144 9548 2148
rect 9564 2204 9628 2208
rect 9564 2148 9568 2204
rect 9568 2148 9624 2204
rect 9624 2148 9628 2204
rect 9564 2144 9628 2148
rect 17696 2204 17760 2208
rect 17696 2148 17700 2204
rect 17700 2148 17756 2204
rect 17756 2148 17760 2204
rect 17696 2144 17760 2148
rect 17776 2204 17840 2208
rect 17776 2148 17780 2204
rect 17780 2148 17836 2204
rect 17836 2148 17840 2204
rect 17776 2144 17840 2148
rect 17856 2204 17920 2208
rect 17856 2148 17860 2204
rect 17860 2148 17916 2204
rect 17916 2148 17920 2204
rect 17856 2144 17920 2148
rect 17936 2204 18000 2208
rect 17936 2148 17940 2204
rect 17940 2148 17996 2204
rect 17996 2148 18000 2204
rect 17936 2144 18000 2148
<< metal4 >>
rect 5130 26688 5450 27248
rect 5130 26624 5138 26688
rect 5202 26624 5218 26688
rect 5282 26624 5298 26688
rect 5362 26624 5378 26688
rect 5442 26624 5450 26688
rect 5130 25600 5450 26624
rect 5130 25536 5138 25600
rect 5202 25536 5218 25600
rect 5282 25536 5298 25600
rect 5362 25536 5378 25600
rect 5442 25536 5450 25600
rect 5130 24512 5450 25536
rect 5130 24448 5138 24512
rect 5202 24448 5218 24512
rect 5282 24448 5298 24512
rect 5362 24448 5378 24512
rect 5442 24448 5450 24512
rect 5130 23424 5450 24448
rect 5130 23360 5138 23424
rect 5202 23360 5218 23424
rect 5282 23360 5298 23424
rect 5362 23360 5378 23424
rect 5442 23360 5450 23424
rect 5130 22336 5450 23360
rect 5130 22272 5138 22336
rect 5202 22272 5218 22336
rect 5282 22272 5298 22336
rect 5362 22272 5378 22336
rect 5442 22272 5450 22336
rect 5130 21248 5450 22272
rect 5130 21184 5138 21248
rect 5202 21184 5218 21248
rect 5282 21184 5298 21248
rect 5362 21184 5378 21248
rect 5442 21184 5450 21248
rect 5130 20160 5450 21184
rect 5130 20096 5138 20160
rect 5202 20096 5218 20160
rect 5282 20096 5298 20160
rect 5362 20096 5378 20160
rect 5442 20096 5450 20160
rect 5130 19072 5450 20096
rect 5130 19008 5138 19072
rect 5202 19008 5218 19072
rect 5282 19008 5298 19072
rect 5362 19008 5378 19072
rect 5442 19008 5450 19072
rect 5130 17984 5450 19008
rect 9316 27232 9636 27248
rect 9316 27168 9324 27232
rect 9388 27168 9404 27232
rect 9468 27168 9484 27232
rect 9548 27168 9564 27232
rect 9628 27168 9636 27232
rect 9316 26144 9636 27168
rect 9316 26080 9324 26144
rect 9388 26080 9404 26144
rect 9468 26080 9484 26144
rect 9548 26080 9564 26144
rect 9628 26080 9636 26144
rect 9316 25056 9636 26080
rect 9316 24992 9324 25056
rect 9388 24992 9404 25056
rect 9468 24992 9484 25056
rect 9548 24992 9564 25056
rect 9628 24992 9636 25056
rect 9316 23968 9636 24992
rect 9316 23904 9324 23968
rect 9388 23904 9404 23968
rect 9468 23904 9484 23968
rect 9548 23904 9564 23968
rect 9628 23904 9636 23968
rect 9316 22880 9636 23904
rect 9316 22816 9324 22880
rect 9388 22816 9404 22880
rect 9468 22816 9484 22880
rect 9548 22816 9564 22880
rect 9628 22816 9636 22880
rect 9316 21792 9636 22816
rect 9316 21728 9324 21792
rect 9388 21728 9404 21792
rect 9468 21728 9484 21792
rect 9548 21728 9564 21792
rect 9628 21728 9636 21792
rect 9316 20704 9636 21728
rect 9316 20640 9324 20704
rect 9388 20640 9404 20704
rect 9468 20640 9484 20704
rect 9548 20640 9564 20704
rect 9628 20640 9636 20704
rect 9316 19616 9636 20640
rect 9316 19552 9324 19616
rect 9388 19552 9404 19616
rect 9468 19552 9484 19616
rect 9548 19552 9564 19616
rect 9628 19552 9636 19616
rect 8891 18732 8957 18733
rect 8891 18668 8892 18732
rect 8956 18668 8957 18732
rect 8891 18667 8957 18668
rect 5130 17920 5138 17984
rect 5202 17920 5218 17984
rect 5282 17920 5298 17984
rect 5362 17920 5378 17984
rect 5442 17920 5450 17984
rect 5130 16896 5450 17920
rect 5130 16832 5138 16896
rect 5202 16832 5218 16896
rect 5282 16832 5298 16896
rect 5362 16832 5378 16896
rect 5442 16832 5450 16896
rect 5130 15808 5450 16832
rect 5130 15744 5138 15808
rect 5202 15744 5218 15808
rect 5282 15744 5298 15808
rect 5362 15744 5378 15808
rect 5442 15744 5450 15808
rect 5130 14720 5450 15744
rect 5130 14656 5138 14720
rect 5202 14656 5218 14720
rect 5282 14656 5298 14720
rect 5362 14656 5378 14720
rect 5442 14656 5450 14720
rect 5130 13632 5450 14656
rect 5130 13568 5138 13632
rect 5202 13568 5218 13632
rect 5282 13568 5298 13632
rect 5362 13568 5378 13632
rect 5442 13568 5450 13632
rect 5130 12544 5450 13568
rect 8707 12884 8773 12885
rect 8707 12820 8708 12884
rect 8772 12820 8773 12884
rect 8707 12819 8773 12820
rect 5130 12480 5138 12544
rect 5202 12480 5218 12544
rect 5282 12480 5298 12544
rect 5362 12480 5378 12544
rect 5442 12480 5450 12544
rect 5130 11456 5450 12480
rect 5130 11392 5138 11456
rect 5202 11392 5218 11456
rect 5282 11392 5298 11456
rect 5362 11392 5378 11456
rect 5442 11392 5450 11456
rect 5130 10368 5450 11392
rect 5130 10304 5138 10368
rect 5202 10304 5218 10368
rect 5282 10304 5298 10368
rect 5362 10304 5378 10368
rect 5442 10304 5450 10368
rect 5130 9280 5450 10304
rect 5130 9216 5138 9280
rect 5202 9216 5218 9280
rect 5282 9216 5298 9280
rect 5362 9216 5378 9280
rect 5442 9216 5450 9280
rect 5130 8192 5450 9216
rect 5130 8128 5138 8192
rect 5202 8128 5218 8192
rect 5282 8128 5298 8192
rect 5362 8128 5378 8192
rect 5442 8128 5450 8192
rect 5130 7104 5450 8128
rect 5130 7040 5138 7104
rect 5202 7040 5218 7104
rect 5282 7040 5298 7104
rect 5362 7040 5378 7104
rect 5442 7040 5450 7104
rect 5130 6016 5450 7040
rect 5130 5952 5138 6016
rect 5202 5952 5218 6016
rect 5282 5952 5298 6016
rect 5362 5952 5378 6016
rect 5442 5952 5450 6016
rect 5130 4928 5450 5952
rect 5130 4864 5138 4928
rect 5202 4864 5218 4928
rect 5282 4864 5298 4928
rect 5362 4864 5378 4928
rect 5442 4864 5450 4928
rect 5130 3840 5450 4864
rect 5130 3776 5138 3840
rect 5202 3776 5218 3840
rect 5282 3776 5298 3840
rect 5362 3776 5378 3840
rect 5442 3776 5450 3840
rect 5130 2752 5450 3776
rect 8710 3365 8770 12819
rect 8894 3637 8954 18667
rect 9316 18528 9636 19552
rect 9316 18464 9324 18528
rect 9388 18464 9404 18528
rect 9468 18464 9484 18528
rect 9548 18464 9564 18528
rect 9628 18464 9636 18528
rect 9316 17440 9636 18464
rect 9316 17376 9324 17440
rect 9388 17376 9404 17440
rect 9468 17376 9484 17440
rect 9548 17376 9564 17440
rect 9628 17376 9636 17440
rect 9316 16352 9636 17376
rect 9316 16288 9324 16352
rect 9388 16288 9404 16352
rect 9468 16288 9484 16352
rect 9548 16288 9564 16352
rect 9628 16288 9636 16352
rect 9316 15264 9636 16288
rect 9316 15200 9324 15264
rect 9388 15200 9404 15264
rect 9468 15200 9484 15264
rect 9548 15200 9564 15264
rect 9628 15200 9636 15264
rect 9075 14788 9141 14789
rect 9075 14724 9076 14788
rect 9140 14724 9141 14788
rect 9075 14723 9141 14724
rect 9078 4589 9138 14723
rect 9316 14176 9636 15200
rect 13502 26688 13822 27248
rect 13502 26624 13510 26688
rect 13574 26624 13590 26688
rect 13654 26624 13670 26688
rect 13734 26624 13750 26688
rect 13814 26624 13822 26688
rect 13502 25600 13822 26624
rect 13502 25536 13510 25600
rect 13574 25536 13590 25600
rect 13654 25536 13670 25600
rect 13734 25536 13750 25600
rect 13814 25536 13822 25600
rect 13502 24512 13822 25536
rect 13502 24448 13510 24512
rect 13574 24448 13590 24512
rect 13654 24448 13670 24512
rect 13734 24448 13750 24512
rect 13814 24448 13822 24512
rect 13502 23424 13822 24448
rect 13502 23360 13510 23424
rect 13574 23360 13590 23424
rect 13654 23360 13670 23424
rect 13734 23360 13750 23424
rect 13814 23360 13822 23424
rect 13502 22336 13822 23360
rect 13502 22272 13510 22336
rect 13574 22272 13590 22336
rect 13654 22272 13670 22336
rect 13734 22272 13750 22336
rect 13814 22272 13822 22336
rect 13502 21248 13822 22272
rect 13502 21184 13510 21248
rect 13574 21184 13590 21248
rect 13654 21184 13670 21248
rect 13734 21184 13750 21248
rect 13814 21184 13822 21248
rect 13502 20160 13822 21184
rect 13502 20096 13510 20160
rect 13574 20096 13590 20160
rect 13654 20096 13670 20160
rect 13734 20096 13750 20160
rect 13814 20096 13822 20160
rect 13502 19072 13822 20096
rect 17688 27232 18008 27248
rect 17688 27168 17696 27232
rect 17760 27168 17776 27232
rect 17840 27168 17856 27232
rect 17920 27168 17936 27232
rect 18000 27168 18008 27232
rect 17688 26144 18008 27168
rect 17688 26080 17696 26144
rect 17760 26080 17776 26144
rect 17840 26080 17856 26144
rect 17920 26080 17936 26144
rect 18000 26080 18008 26144
rect 17688 25056 18008 26080
rect 17688 24992 17696 25056
rect 17760 24992 17776 25056
rect 17840 24992 17856 25056
rect 17920 24992 17936 25056
rect 18000 24992 18008 25056
rect 17688 23968 18008 24992
rect 17688 23904 17696 23968
rect 17760 23904 17776 23968
rect 17840 23904 17856 23968
rect 17920 23904 17936 23968
rect 18000 23904 18008 23968
rect 17688 22880 18008 23904
rect 17688 22816 17696 22880
rect 17760 22816 17776 22880
rect 17840 22816 17856 22880
rect 17920 22816 17936 22880
rect 18000 22816 18008 22880
rect 17688 21792 18008 22816
rect 17688 21728 17696 21792
rect 17760 21728 17776 21792
rect 17840 21728 17856 21792
rect 17920 21728 17936 21792
rect 18000 21728 18008 21792
rect 17688 20704 18008 21728
rect 17688 20640 17696 20704
rect 17760 20640 17776 20704
rect 17840 20640 17856 20704
rect 17920 20640 17936 20704
rect 18000 20640 18008 20704
rect 16987 19684 17053 19685
rect 16987 19620 16988 19684
rect 17052 19620 17053 19684
rect 16987 19619 17053 19620
rect 13502 19008 13510 19072
rect 13574 19008 13590 19072
rect 13654 19008 13670 19072
rect 13734 19008 13750 19072
rect 13814 19008 13822 19072
rect 13502 17984 13822 19008
rect 13502 17920 13510 17984
rect 13574 17920 13590 17984
rect 13654 17920 13670 17984
rect 13734 17920 13750 17984
rect 13814 17920 13822 17984
rect 13502 16896 13822 17920
rect 13502 16832 13510 16896
rect 13574 16832 13590 16896
rect 13654 16832 13670 16896
rect 13734 16832 13750 16896
rect 13814 16832 13822 16896
rect 13502 15808 13822 16832
rect 13502 15744 13510 15808
rect 13574 15744 13590 15808
rect 13654 15744 13670 15808
rect 13734 15744 13750 15808
rect 13814 15744 13822 15808
rect 12019 14788 12085 14789
rect 12019 14724 12020 14788
rect 12084 14724 12085 14788
rect 12019 14723 12085 14724
rect 9316 14112 9324 14176
rect 9388 14112 9404 14176
rect 9468 14112 9484 14176
rect 9548 14112 9564 14176
rect 9628 14112 9636 14176
rect 9316 13088 9636 14112
rect 9316 13024 9324 13088
rect 9388 13024 9404 13088
rect 9468 13024 9484 13088
rect 9548 13024 9564 13088
rect 9628 13024 9636 13088
rect 9316 12000 9636 13024
rect 9316 11936 9324 12000
rect 9388 11936 9404 12000
rect 9468 11936 9484 12000
rect 9548 11936 9564 12000
rect 9628 11936 9636 12000
rect 9316 10912 9636 11936
rect 9316 10848 9324 10912
rect 9388 10848 9404 10912
rect 9468 10848 9484 10912
rect 9548 10848 9564 10912
rect 9628 10848 9636 10912
rect 9316 9824 9636 10848
rect 9316 9760 9324 9824
rect 9388 9760 9404 9824
rect 9468 9760 9484 9824
rect 9548 9760 9564 9824
rect 9628 9760 9636 9824
rect 9316 8736 9636 9760
rect 9316 8672 9324 8736
rect 9388 8672 9404 8736
rect 9468 8672 9484 8736
rect 9548 8672 9564 8736
rect 9628 8672 9636 8736
rect 9316 7648 9636 8672
rect 9316 7584 9324 7648
rect 9388 7584 9404 7648
rect 9468 7584 9484 7648
rect 9548 7584 9564 7648
rect 9628 7584 9636 7648
rect 9316 6560 9636 7584
rect 11099 7036 11165 7037
rect 11099 6972 11100 7036
rect 11164 6972 11165 7036
rect 11099 6971 11165 6972
rect 9316 6496 9324 6560
rect 9388 6496 9404 6560
rect 9468 6496 9484 6560
rect 9548 6496 9564 6560
rect 9628 6496 9636 6560
rect 9316 5472 9636 6496
rect 9316 5408 9324 5472
rect 9388 5408 9404 5472
rect 9468 5408 9484 5472
rect 9548 5408 9564 5472
rect 9628 5408 9636 5472
rect 9075 4588 9141 4589
rect 9075 4524 9076 4588
rect 9140 4524 9141 4588
rect 9075 4523 9141 4524
rect 9316 4384 9636 5408
rect 11102 4861 11162 6971
rect 11099 4860 11165 4861
rect 11099 4796 11100 4860
rect 11164 4796 11165 4860
rect 11099 4795 11165 4796
rect 9316 4320 9324 4384
rect 9388 4320 9404 4384
rect 9468 4320 9484 4384
rect 9548 4320 9564 4384
rect 9628 4320 9636 4384
rect 8891 3636 8957 3637
rect 8891 3572 8892 3636
rect 8956 3572 8957 3636
rect 8891 3571 8957 3572
rect 8707 3364 8773 3365
rect 8707 3300 8708 3364
rect 8772 3300 8773 3364
rect 8707 3299 8773 3300
rect 5130 2688 5138 2752
rect 5202 2688 5218 2752
rect 5282 2688 5298 2752
rect 5362 2688 5378 2752
rect 5442 2688 5450 2752
rect 5130 2128 5450 2688
rect 9316 3296 9636 4320
rect 12022 3501 12082 14723
rect 13502 14720 13822 15744
rect 13502 14656 13510 14720
rect 13574 14656 13590 14720
rect 13654 14656 13670 14720
rect 13734 14656 13750 14720
rect 13814 14656 13822 14720
rect 13502 13632 13822 14656
rect 13502 13568 13510 13632
rect 13574 13568 13590 13632
rect 13654 13568 13670 13632
rect 13734 13568 13750 13632
rect 13814 13568 13822 13632
rect 13502 12544 13822 13568
rect 16803 13292 16869 13293
rect 16803 13228 16804 13292
rect 16868 13228 16869 13292
rect 16803 13227 16869 13228
rect 13502 12480 13510 12544
rect 13574 12480 13590 12544
rect 13654 12480 13670 12544
rect 13734 12480 13750 12544
rect 13814 12480 13822 12544
rect 13502 11456 13822 12480
rect 13502 11392 13510 11456
rect 13574 11392 13590 11456
rect 13654 11392 13670 11456
rect 13734 11392 13750 11456
rect 13814 11392 13822 11456
rect 13502 10368 13822 11392
rect 13502 10304 13510 10368
rect 13574 10304 13590 10368
rect 13654 10304 13670 10368
rect 13734 10304 13750 10368
rect 13814 10304 13822 10368
rect 13502 9280 13822 10304
rect 13502 9216 13510 9280
rect 13574 9216 13590 9280
rect 13654 9216 13670 9280
rect 13734 9216 13750 9280
rect 13814 9216 13822 9280
rect 13502 8192 13822 9216
rect 13502 8128 13510 8192
rect 13574 8128 13590 8192
rect 13654 8128 13670 8192
rect 13734 8128 13750 8192
rect 13814 8128 13822 8192
rect 13502 7104 13822 8128
rect 13502 7040 13510 7104
rect 13574 7040 13590 7104
rect 13654 7040 13670 7104
rect 13734 7040 13750 7104
rect 13814 7040 13822 7104
rect 13502 6016 13822 7040
rect 13502 5952 13510 6016
rect 13574 5952 13590 6016
rect 13654 5952 13670 6016
rect 13734 5952 13750 6016
rect 13814 5952 13822 6016
rect 13502 4928 13822 5952
rect 13502 4864 13510 4928
rect 13574 4864 13590 4928
rect 13654 4864 13670 4928
rect 13734 4864 13750 4928
rect 13814 4864 13822 4928
rect 13502 3840 13822 4864
rect 16806 4045 16866 13227
rect 16990 4045 17050 19619
rect 17688 19616 18008 20640
rect 17688 19552 17696 19616
rect 17760 19552 17776 19616
rect 17840 19552 17856 19616
rect 17920 19552 17936 19616
rect 18000 19552 18008 19616
rect 17688 18528 18008 19552
rect 17688 18464 17696 18528
rect 17760 18464 17776 18528
rect 17840 18464 17856 18528
rect 17920 18464 17936 18528
rect 18000 18464 18008 18528
rect 17688 17440 18008 18464
rect 17688 17376 17696 17440
rect 17760 17376 17776 17440
rect 17840 17376 17856 17440
rect 17920 17376 17936 17440
rect 18000 17376 18008 17440
rect 17688 16352 18008 17376
rect 17688 16288 17696 16352
rect 17760 16288 17776 16352
rect 17840 16288 17856 16352
rect 17920 16288 17936 16352
rect 18000 16288 18008 16352
rect 17688 15264 18008 16288
rect 17688 15200 17696 15264
rect 17760 15200 17776 15264
rect 17840 15200 17856 15264
rect 17920 15200 17936 15264
rect 18000 15200 18008 15264
rect 17688 14176 18008 15200
rect 17688 14112 17696 14176
rect 17760 14112 17776 14176
rect 17840 14112 17856 14176
rect 17920 14112 17936 14176
rect 18000 14112 18008 14176
rect 17688 13088 18008 14112
rect 17688 13024 17696 13088
rect 17760 13024 17776 13088
rect 17840 13024 17856 13088
rect 17920 13024 17936 13088
rect 18000 13024 18008 13088
rect 17688 12000 18008 13024
rect 17688 11936 17696 12000
rect 17760 11936 17776 12000
rect 17840 11936 17856 12000
rect 17920 11936 17936 12000
rect 18000 11936 18008 12000
rect 17688 10912 18008 11936
rect 17688 10848 17696 10912
rect 17760 10848 17776 10912
rect 17840 10848 17856 10912
rect 17920 10848 17936 10912
rect 18000 10848 18008 10912
rect 17688 9824 18008 10848
rect 17688 9760 17696 9824
rect 17760 9760 17776 9824
rect 17840 9760 17856 9824
rect 17920 9760 17936 9824
rect 18000 9760 18008 9824
rect 17688 8736 18008 9760
rect 17688 8672 17696 8736
rect 17760 8672 17776 8736
rect 17840 8672 17856 8736
rect 17920 8672 17936 8736
rect 18000 8672 18008 8736
rect 17688 7648 18008 8672
rect 17688 7584 17696 7648
rect 17760 7584 17776 7648
rect 17840 7584 17856 7648
rect 17920 7584 17936 7648
rect 18000 7584 18008 7648
rect 17688 6560 18008 7584
rect 17688 6496 17696 6560
rect 17760 6496 17776 6560
rect 17840 6496 17856 6560
rect 17920 6496 17936 6560
rect 18000 6496 18008 6560
rect 17688 5472 18008 6496
rect 17688 5408 17696 5472
rect 17760 5408 17776 5472
rect 17840 5408 17856 5472
rect 17920 5408 17936 5472
rect 18000 5408 18008 5472
rect 17688 4384 18008 5408
rect 17688 4320 17696 4384
rect 17760 4320 17776 4384
rect 17840 4320 17856 4384
rect 17920 4320 17936 4384
rect 18000 4320 18008 4384
rect 16803 4044 16869 4045
rect 16803 3980 16804 4044
rect 16868 3980 16869 4044
rect 16803 3979 16869 3980
rect 16987 4044 17053 4045
rect 16987 3980 16988 4044
rect 17052 3980 17053 4044
rect 16987 3979 17053 3980
rect 13502 3776 13510 3840
rect 13574 3776 13590 3840
rect 13654 3776 13670 3840
rect 13734 3776 13750 3840
rect 13814 3776 13822 3840
rect 12019 3500 12085 3501
rect 12019 3436 12020 3500
rect 12084 3436 12085 3500
rect 12019 3435 12085 3436
rect 9316 3232 9324 3296
rect 9388 3232 9404 3296
rect 9468 3232 9484 3296
rect 9548 3232 9564 3296
rect 9628 3232 9636 3296
rect 9316 2208 9636 3232
rect 9316 2144 9324 2208
rect 9388 2144 9404 2208
rect 9468 2144 9484 2208
rect 9548 2144 9564 2208
rect 9628 2144 9636 2208
rect 9316 2128 9636 2144
rect 13502 2752 13822 3776
rect 13502 2688 13510 2752
rect 13574 2688 13590 2752
rect 13654 2688 13670 2752
rect 13734 2688 13750 2752
rect 13814 2688 13822 2752
rect 13502 2128 13822 2688
rect 17688 3296 18008 4320
rect 17688 3232 17696 3296
rect 17760 3232 17776 3296
rect 17840 3232 17856 3296
rect 17920 3232 17936 3296
rect 18000 3232 18008 3296
rect 17688 2208 18008 3232
rect 17688 2144 17696 2208
rect 17760 2144 17776 2208
rect 17840 2144 17856 2208
rect 17920 2144 17936 2208
rect 18000 2144 18008 2208
rect 17688 2128 18008 2144
rect 21874 26688 22194 27248
rect 21874 26624 21882 26688
rect 21946 26624 21962 26688
rect 22026 26624 22042 26688
rect 22106 26624 22122 26688
rect 22186 26624 22194 26688
rect 21874 25600 22194 26624
rect 21874 25536 21882 25600
rect 21946 25536 21962 25600
rect 22026 25536 22042 25600
rect 22106 25536 22122 25600
rect 22186 25536 22194 25600
rect 21874 24512 22194 25536
rect 21874 24448 21882 24512
rect 21946 24448 21962 24512
rect 22026 24448 22042 24512
rect 22106 24448 22122 24512
rect 22186 24448 22194 24512
rect 21874 23424 22194 24448
rect 21874 23360 21882 23424
rect 21946 23360 21962 23424
rect 22026 23360 22042 23424
rect 22106 23360 22122 23424
rect 22186 23360 22194 23424
rect 21874 22336 22194 23360
rect 21874 22272 21882 22336
rect 21946 22272 21962 22336
rect 22026 22272 22042 22336
rect 22106 22272 22122 22336
rect 22186 22272 22194 22336
rect 21874 21248 22194 22272
rect 22507 22132 22573 22133
rect 22507 22068 22508 22132
rect 22572 22068 22573 22132
rect 22507 22067 22573 22068
rect 21874 21184 21882 21248
rect 21946 21184 21962 21248
rect 22026 21184 22042 21248
rect 22106 21184 22122 21248
rect 22186 21184 22194 21248
rect 21874 20160 22194 21184
rect 21874 20096 21882 20160
rect 21946 20096 21962 20160
rect 22026 20096 22042 20160
rect 22106 20096 22122 20160
rect 22186 20096 22194 20160
rect 21874 19072 22194 20096
rect 21874 19008 21882 19072
rect 21946 19008 21962 19072
rect 22026 19008 22042 19072
rect 22106 19008 22122 19072
rect 22186 19008 22194 19072
rect 21874 17984 22194 19008
rect 21874 17920 21882 17984
rect 21946 17920 21962 17984
rect 22026 17920 22042 17984
rect 22106 17920 22122 17984
rect 22186 17920 22194 17984
rect 21874 16896 22194 17920
rect 21874 16832 21882 16896
rect 21946 16832 21962 16896
rect 22026 16832 22042 16896
rect 22106 16832 22122 16896
rect 22186 16832 22194 16896
rect 21874 15808 22194 16832
rect 21874 15744 21882 15808
rect 21946 15744 21962 15808
rect 22026 15744 22042 15808
rect 22106 15744 22122 15808
rect 22186 15744 22194 15808
rect 21874 14720 22194 15744
rect 21874 14656 21882 14720
rect 21946 14656 21962 14720
rect 22026 14656 22042 14720
rect 22106 14656 22122 14720
rect 22186 14656 22194 14720
rect 21874 13632 22194 14656
rect 21874 13568 21882 13632
rect 21946 13568 21962 13632
rect 22026 13568 22042 13632
rect 22106 13568 22122 13632
rect 22186 13568 22194 13632
rect 21874 12544 22194 13568
rect 21874 12480 21882 12544
rect 21946 12480 21962 12544
rect 22026 12480 22042 12544
rect 22106 12480 22122 12544
rect 22186 12480 22194 12544
rect 21874 11456 22194 12480
rect 22510 12341 22570 22067
rect 22507 12340 22573 12341
rect 22507 12276 22508 12340
rect 22572 12276 22573 12340
rect 22507 12275 22573 12276
rect 21874 11392 21882 11456
rect 21946 11392 21962 11456
rect 22026 11392 22042 11456
rect 22106 11392 22122 11456
rect 22186 11392 22194 11456
rect 21874 10368 22194 11392
rect 21874 10304 21882 10368
rect 21946 10304 21962 10368
rect 22026 10304 22042 10368
rect 22106 10304 22122 10368
rect 22186 10304 22194 10368
rect 21874 9280 22194 10304
rect 21874 9216 21882 9280
rect 21946 9216 21962 9280
rect 22026 9216 22042 9280
rect 22106 9216 22122 9280
rect 22186 9216 22194 9280
rect 21874 8192 22194 9216
rect 21874 8128 21882 8192
rect 21946 8128 21962 8192
rect 22026 8128 22042 8192
rect 22106 8128 22122 8192
rect 22186 8128 22194 8192
rect 21874 7104 22194 8128
rect 21874 7040 21882 7104
rect 21946 7040 21962 7104
rect 22026 7040 22042 7104
rect 22106 7040 22122 7104
rect 22186 7040 22194 7104
rect 21874 6016 22194 7040
rect 21874 5952 21882 6016
rect 21946 5952 21962 6016
rect 22026 5952 22042 6016
rect 22106 5952 22122 6016
rect 22186 5952 22194 6016
rect 21874 4928 22194 5952
rect 21874 4864 21882 4928
rect 21946 4864 21962 4928
rect 22026 4864 22042 4928
rect 22106 4864 22122 4928
rect 22186 4864 22194 4928
rect 21874 3840 22194 4864
rect 21874 3776 21882 3840
rect 21946 3776 21962 3840
rect 22026 3776 22042 3840
rect 22106 3776 22122 3840
rect 22186 3776 22194 3840
rect 21874 2752 22194 3776
rect 21874 2688 21882 2752
rect 21946 2688 21962 2752
rect 22026 2688 22042 2752
rect 22106 2688 22122 2752
rect 22186 2688 22194 2752
rect 21874 2128 22194 2688
use sky130_fd_sc_hd__decap_12  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1640608721
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1640608721
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1640608721
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1640608721
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1640608721
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1640608721
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1640608721
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1640608721
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1640608721
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1640608721
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1640608721
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1640608721
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1640608721
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 6348 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 8372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1640608721
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1640608721
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1640608721
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1640608721
transform 1 0 8280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0695_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B
timestamp 1640608721
transform 1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1640608721
transform -1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__B
timestamp 1640608721
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_93 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_98
timestamp 1640608721
transform 1 0 10120 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1640608721
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1011_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1344_
timestamp 1640608721
transform 1 0 9384 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_1  _1013_
timestamp 1640608721
transform -1 0 11224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0665_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 11500 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1640608721
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1640608721
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1640608721
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1640608721
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1009_
timestamp 1640608721
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_122
timestamp 1640608721
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1640608721
transform 1 0 11960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1640608721
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1640608721
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1640608721
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_126
timestamp 1640608721
transform 1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1640608721
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0666_
timestamp 1640608721
transform 1 0 13156 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1346_
timestamp 1640608721
transform 1 0 13064 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1640608721
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1640608721
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_152
timestamp 1640608721
transform 1 0 15088 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1640608721
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1068_
timestamp 1640608721
transform 1 0 14628 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1640608721
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1640608721
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1640608721
transform 1 0 16928 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1640608721
transform 1 0 18032 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1640608721
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1640608721
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0999_
timestamp 1640608721
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1640608721
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1640608721
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_208
timestamp 1640608721
transform 1 0 20240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_196
timestamp 1640608721
transform 1 0 19136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_201
timestamp 1640608721
transform 1 0 19596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1640608721
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0994_
timestamp 1640608721
transform 1 0 19320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1352_
timestamp 1640608721
transform 1 0 19780 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_2  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 20792 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_0_214
timestamp 1640608721
transform 1 0 20792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1194_
timestamp 1640608721
transform -1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1640608721
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1640608721
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1640608721
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_228
timestamp 1640608721
transform 1 0 22080 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1640608721
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1640608721
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1640608721
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1640608721
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1640608721
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_234
timestamp 1640608721
transform 1 0 22632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_238
timestamp 1640608721
transform 1 0 23000 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_250
timestamp 1640608721
transform 1 0 24104 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1195_
timestamp 1640608721
transform -1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1640608721
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1640608721
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_269
timestamp 1640608721
transform 1 0 25852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_262
timestamp 1640608721
transform 1 0 25208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1640608721
transform -1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1640608721
transform -1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1640608721
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1640608721
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1640608721
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1640608721
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1640608721
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1640608721
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1640608721
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1640608721
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1640608721
transform -1 0 6440 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp 1640608721
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_58
timestamp 1640608721
transform 1 0 6440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1362_
timestamp 1640608721
transform -1 0 8280 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_2  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 8832 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A
timestamp 1640608721
transform -1 0 9844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1640608721
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_2  _0708_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 9660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1343_
timestamp 1640608721
transform 1 0 9844 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__a21bo_2  _1061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 12144 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1345_
timestamp 1640608721
transform 1 0 12144 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1640608721
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1007_
timestamp 1640608721
transform -1 0 13984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1069_
timestamp 1640608721
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _0667_
timestamp 1640608721
transform 1 0 14812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1348_
timestamp 1640608721
transform 1 0 15364 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1349_
timestamp 1640608721
transform -1 0 18492 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_2_189
timestamp 1640608721
transform 1 0 18492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp 1640608721
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1640608721
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0992_
timestamp 1640608721
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1351_
timestamp 1640608721
transform 1 0 19320 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_1  _0989_
timestamp 1640608721
transform 1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1094_
timestamp 1640608721
transform 1 0 21436 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1111_
timestamp 1640608721
transform -1 0 21436 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1353_
timestamp 1640608721
transform 1 0 22172 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_2_246
timestamp 1640608721
transform 1 0 23736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1200_
timestamp 1640608721
transform -1 0 24288 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_253
timestamp 1640608721
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_262
timestamp 1640608721
transform 1 0 25208 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1640608721
transform -1 0 26220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1640608721
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1201_
timestamp 1640608721
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B
timestamp 1640608721
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1640608721
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1640608721
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1640608721
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1640608721
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1640608721
transform 1 0 3588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_29
timestamp 1640608721
transform 1 0 3772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_41
timestamp 1640608721
transform 1 0 4876 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1022_
timestamp 1640608721
transform 1 0 3128 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_3_49
timestamp 1640608721
transform 1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1640608721
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1640608721
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _0963_
timestamp 1640608721
transform 1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 7268 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__C
timestamp 1640608721
transform -1 0 8924 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__S
timestamp 1640608721
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_67
timestamp 1640608721
transform 1 0 7268 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_76
timestamp 1640608721
transform 1 0 8096 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_82
timestamp 1640608721
transform 1 0 8648 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0845_
timestamp 1640608721
transform -1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1640608721
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1640608721
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _1010_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 9292 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1225_
timestamp 1640608721
transform 1 0 10028 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_106
timestamp 1640608721
transform 1 0 10856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1640608721
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1640608721
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0664_
timestamp 1640608721
transform 1 0 10948 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _1006_
timestamp 1640608721
transform 1 0 12420 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _1008_
timestamp 1640608721
transform -1 0 12420 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1063_
timestamp 1640608721
transform -1 0 13892 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1347_
timestamp 1640608721
transform 1 0 13892 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_3_159
timestamp 1640608721
transform 1 0 15732 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1002_
timestamp 1640608721
transform 1 0 15456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1089_
timestamp 1640608721
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_183
timestamp 1640608721
transform 1 0 17940 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1640608721
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0668_
timestamp 1640608721
transform 1 0 17388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _0998_
timestamp 1640608721
transform -1 0 17388 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1350_
timestamp 1640608721
transform 1 0 18032 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__and3b_2  _0991_
timestamp 1640608721
transform 1 0 19596 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_225
timestamp 1640608721
transform 1 0 21804 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1640608721
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _0986_
timestamp 1640608721
transform 1 0 21896 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _0988_
timestamp 1640608721
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _1112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 20332 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_3_247
timestamp 1640608721
transform 1 0 23828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1118_
timestamp 1640608721
transform 1 0 23368 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1119_
timestamp 1640608721
transform 1 0 22632 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_259
timestamp 1640608721
transform 1 0 24932 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_267
timestamp 1640608721
transform 1 0 25668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1640608721
transform -1 0 26220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_15
timestamp 1640608721
transform 1 0 2484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1640608721
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1640608721
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1640608721
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1640608721
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1640608721
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1023_
timestamp 1640608721
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1361_
timestamp 1640608721
transform 1 0 3864 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_4_47
timestamp 1640608721
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1043_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 5980 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1044_
timestamp 1640608721
transform -1 0 5980 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_2  _1046_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 6624 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A1
timestamp 1640608721
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1640608721
transform 1 0 7452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0846_
timestamp 1640608721
transform 1 0 7728 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1042_
timestamp 1640608721
transform -1 0 8648 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__C1
timestamp 1640608721
transform -1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__S
timestamp 1640608721
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__S
timestamp 1640608721
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_87
timestamp 1640608721
transform 1 0 9108 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1640608721
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1223_
timestamp 1640608721
transform 1 0 10212 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__S
timestamp 1640608721
transform 1 0 11960 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_116
timestamp 1640608721
transform 1 0 11776 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_2  _1058_
timestamp 1640608721
transform 1 0 11040 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1229_
timestamp 1640608721
transform 1 0 12144 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1640608721
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1640608721
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _1001_
timestamp 1640608721
transform 1 0 14260 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _1003_
timestamp 1640608721
transform -1 0 13984 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1004_
timestamp 1640608721
transform 1 0 12972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_159
timestamp 1640608721
transform 1 0 15732 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1076_
timestamp 1640608721
transform -1 0 15732 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1082_
timestamp 1640608721
transform 1 0 15824 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1222_
timestamp 1640608721
transform -1 0 17112 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_185
timestamp 1640608721
transform 1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0996_
timestamp 1640608721
transform 1 0 17112 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0997_
timestamp 1640608721
transform 1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__S
timestamp 1640608721
transform 1 0 19412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1640608721
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1640608721
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _0993_
timestamp 1640608721
transform 1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1282_
timestamp 1640608721
transform 1 0 19596 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_217
timestamp 1640608721
transform 1 0 21068 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_225
timestamp 1640608721
transform 1 0 21804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _0662_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 21804 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 20424 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1276_
timestamp 1640608721
transform 1 0 21896 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1354_
timestamp 1640608721
transform 1 0 22724 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_4_256
timestamp 1640608721
transform 1 0 24656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_268
timestamp 1640608721
transform 1 0 25760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1640608721
transform -1 0 26220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1640608721
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0987_
timestamp 1640608721
transform -1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1640608721
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1640608721
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1640608721
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1640608721
transform 1 0 3220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1338_
timestamp 1640608721
transform 1 0 3404 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1640608721
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0659_
timestamp 1640608721
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_2  _0962_
timestamp 1640608721
transform 1 0 6624 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0967_
timestamp 1640608721
transform -1 0 5428 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1247_
timestamp 1640608721
transform -1 0 6256 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _0661_
timestamp 1640608721
transform 1 0 8280 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _0965_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 7452 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_91
timestamp 1640608721
transform 1 0 9476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _1012_
timestamp 1640608721
transform 1 0 10028 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1045_
timestamp 1640608721
transform -1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1048_
timestamp 1640608721
transform -1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1640608721
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1640608721
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_117
timestamp 1640608721
transform 1 0 11868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1640608721
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1000_
timestamp 1640608721
transform -1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1005_
timestamp 1640608721
transform -1 0 11868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1059_
timestamp 1640608721
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1060_
timestamp 1640608721
transform -1 0 11316 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0995_
timestamp 1640608721
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1237_
timestamp 1640608721
transform 1 0 13156 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1327_
timestamp 1640608721
transform 1 0 13984 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__S
timestamp 1640608721
transform 1 0 16100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__S
timestamp 1640608721
transform 1 0 14812 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_160
timestamp 1640608721
transform 1 0 15824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1640608721
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1253_
timestamp 1640608721
transform 1 0 14996 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__S
timestamp 1640608721
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1640608721
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1083_
timestamp 1640608721
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1295_
timestamp 1640608721
transform 1 0 17572 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__S
timestamp 1640608721
transform 1 0 18860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_191
timestamp 1640608721
transform 1 0 18676 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0990_
timestamp 1640608721
transform -1 0 18676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1095_
timestamp 1640608721
transform 1 0 19872 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1301_
timestamp 1640608721
transform 1 0 19044 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__S
timestamp 1640608721
transform 1 0 22172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__S
timestamp 1640608721
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_212
timestamp 1640608721
transform 1 0 20608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1640608721
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_227
timestamp 1640608721
transform 1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1640608721
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _0669_
timestamp 1640608721
transform -1 0 21436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1124_
timestamp 1640608721
transform 1 0 23920 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1125_
timestamp 1640608721
transform 1 0 23184 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1232_
timestamp 1640608721
transform 1 0 22356 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_253
timestamp 1640608721
transform 1 0 24380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_265
timestamp 1640608721
transform 1 0 25484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_269
timestamp 1640608721
transform 1 0 25852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1640608721
transform -1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1640608721
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1640608721
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1640608721
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1640608721
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1640608721
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1640608721
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1640608721
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1640608721
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp 1640608721
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1640608721
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1640608721
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1640608721
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1041_
timestamp 1640608721
transform -1 0 6072 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0856_
timestamp 1640608721
transform 1 0 5336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp 1640608721
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A
timestamp 1640608721
transform 1 0 5152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1047_
timestamp 1640608721
transform -1 0 6808 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_2  _0966_
timestamp 1640608721
transform 1 0 6532 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0964_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 6072 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1640608721
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__S
timestamp 1640608721
transform 1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A
timestamp 1640608721
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1640608721
transform 1 0 6808 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1249_
timestamp 1640608721
transform 1 0 7360 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0849_
timestamp 1640608721
transform -1 0 7360 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1640608721
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A2
timestamp 1640608721
transform 1 0 7636 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1040_
timestamp 1640608721
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1640608721
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 1640608721
transform 1 0 8464 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__S
timestamp 1640608721
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A2
timestamp 1640608721
transform 1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A3
timestamp 1640608721
transform 1 0 7820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_79
timestamp 1640608721
transform 1 0 8372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__S
timestamp 1640608721
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_90
timestamp 1640608721
transform 1 0 9384 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_91
timestamp 1640608721
transform 1 0 9476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1640608721
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1054_
timestamp 1640608721
transform 1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1055_
timestamp 1640608721
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1056_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 10580 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1224_
timestamp 1640608721
transform 1 0 10212 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__S
timestamp 1640608721
transform 1 0 11316 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_108
timestamp 1640608721
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_113
timestamp 1640608721
transform 1 0 11500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_125
timestamp 1640608721
transform 1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_122
timestamp 1640608721
transform 1 0 12328 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1640608721
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1640608721
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1226_
timestamp 1640608721
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__S
timestamp 1640608721
transform 1 0 12972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__S
timestamp 1640608721
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_131
timestamp 1640608721
transform 1 0 13156 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_137
timestamp 1640608721
transform 1 0 13708 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1640608721
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_134
timestamp 1640608721
transform 1 0 13432 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1640608721
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1640608721
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1640608721
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_146
timestamp 1640608721
transform 1 0 14536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1640608721
transform 1 0 14996 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1640608721
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 14996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1640608721
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1640608721
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1640608721
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1640608721
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1640608721
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1151_
timestamp 1640608721
transform -1 0 18584 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1150_
timestamp 1640608721
transform -1 0 19044 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0985_
timestamp 1640608721
transform 1 0 18584 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0979_
timestamp 1640608721
transform 1 0 19228 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1640608721
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp 1640608721
transform 1 0 19044 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1640608721
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_189
timestamp 1640608721
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0980_
timestamp 1640608721
transform 1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1640608721
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_204
timestamp 1640608721
transform 1 0 19872 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_200
timestamp 1640608721
transform 1 0 19504 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1640608721
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp 1640608721
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_217
timestamp 1640608721
transform 1 0 21068 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1640608721
transform 1 0 21988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1640608721
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1640608721
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1640608721
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _0663_
timestamp 1640608721
transform 1 0 21344 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1139_
timestamp 1640608721
transform 1 0 22172 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1145_
timestamp 1640608721
transform 1 0 20608 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1640608721
transform 1 0 23092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_248
timestamp 1640608721
transform 1 0 23920 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1131_
timestamp 1640608721
transform -1 0 23920 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1138_
timestamp 1640608721
transform -1 0 23460 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1640608721
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1640608721
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp 1640608721
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_269
timestamp 1640608721
transform 1 0 25852 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_260
timestamp 1640608721
transform 1 0 25024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_268
timestamp 1640608721
transform 1 0 25760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1640608721
transform -1 0 26220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1640608721
transform -1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1640608721
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1640608721
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1640608721
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1640608721
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1640608721
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1640608721
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1640608721
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1640608721
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_53
timestamp 1640608721
transform 1 0 5980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_62
timestamp 1640608721
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1052_
timestamp 1640608721
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_68
timestamp 1640608721
transform 1 0 7360 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1640608721
transform 1 0 7912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1640608721
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1640608721
transform -1 0 8280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0861_
timestamp 1640608721
transform -1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1640608721
transform -1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_88
timestamp 1640608721
transform 1 0 9200 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1640608721
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0960_
timestamp 1640608721
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1014_
timestamp 1640608721
transform 1 0 9936 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1342_
timestamp 1640608721
transform -1 0 12236 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_1  _0744_
timestamp 1640608721
transform 1 0 12236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1640608721
transform 1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1640608721
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1640608721
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1640608721
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _0971_
timestamp 1640608721
transform -1 0 14812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1640608721
transform 1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_161
timestamp 1640608721
transform 1 0 15916 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0671_
timestamp 1640608721
transform -1 0 15916 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _1163_
timestamp 1640608721
transform 1 0 14812 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0670_
timestamp 1640608721
transform -1 0 17204 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1358_
timestamp 1640608721
transform -1 0 18768 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1640608721
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0975_
timestamp 1640608721
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1357_
timestamp 1640608721
transform 1 0 19504 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_clk
timestamp 1640608721
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_217
timestamp 1640608721
transform 1 0 21068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1356_
timestamp 1640608721
transform -1 0 23184 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1640608721
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_2  _1132_
timestamp 1640608721
transform 1 0 23184 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1640608721
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_265
timestamp 1640608721
transform 1 0 25484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_269
timestamp 1640608721
transform 1 0 25852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1640608721
transform -1 0 26220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1640608721
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_15
timestamp 1640608721
transform 1 0 2484 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1640608721
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1640608721
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_21
timestamp 1640608721
transform 1 0 3036 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_39
timestamp 1640608721
transform 1 0 4692 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1396_
timestamp 1640608721
transform 1 0 3128 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_clk
timestamp 1640608721
transform -1 0 5152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_A
timestamp 1640608721
transform -1 0 6164 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_44
timestamp 1640608721
transform 1 0 5152 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_52
timestamp 1640608721
transform 1 0 5888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1640608721
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1640608721
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1049_
timestamp 1640608721
transform 1 0 6808 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1050_
timestamp 1640608721
transform -1 0 6808 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__S
timestamp 1640608721
transform 1 0 8004 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__and3_2  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 8004 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0853_
timestamp 1640608721
transform 1 0 8556 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_clk
timestamp 1640608721
transform 1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1640608721
transform -1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_100
timestamp 1640608721
transform 1 0 10304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0672_
timestamp 1640608721
transform -1 0 10304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1640608721
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1640608721
transform -1 0 9476 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0968_
timestamp 1640608721
transform 1 0 9476 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_122
timestamp 1640608721
transform 1 0 12328 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1640608721
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0678_
timestamp 1640608721
transform -1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0701_
timestamp 1640608721
transform -1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0843_
timestamp 1640608721
transform 1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1015_
timestamp 1640608721
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1057_
timestamp 1640608721
transform 1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_134
timestamp 1640608721
transform 1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0972_
timestamp 1640608721
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1360_
timestamp 1640608721
transform 1 0 13984 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__and3b_2  _0973_
timestamp 1640608721
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0974_
timestamp 1640608721
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1640608721
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1246_
timestamp 1640608721
transform 1 0 18216 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1359_
timestamp 1640608721
transform 1 0 16652 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__and3b_2  _0978_
timestamp 1640608721
transform 1 0 19044 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1288_
timestamp 1640608721
transform 1 0 19780 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_212
timestamp 1640608721
transform 1 0 20608 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1640608721
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_2  _0981_
timestamp 1640608721
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _0983_
timestamp 1640608721
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_236
timestamp 1640608721
transform 1 0 22816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0982_
timestamp 1640608721
transform 1 0 22540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1355_
timestamp 1640608721
transform 1 0 22908 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_9_254
timestamp 1640608721
transform 1 0 24472 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_266
timestamp 1640608721
transform 1 0 25576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1640608721
transform -1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_15
timestamp 1640608721
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1640608721
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1640608721
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0865_
timestamp 1640608721
transform -1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B1
timestamp 1640608721
transform -1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1640608721
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 3956 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0864_
timestamp 1640608721
transform -1 0 5244 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_45
timestamp 1640608721
transform 1 0 5244 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0862_
timestamp 1640608721
transform -1 0 5612 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1051_
timestamp 1640608721
transform -1 0 6440 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1248_
timestamp 1640608721
transform 1 0 6440 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clk
timestamp 1640608721
transform -1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _0673_
timestamp 1640608721
transform -1 0 8832 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1640608721
transform -1 0 7544 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0957_
timestamp 1640608721
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__C
timestamp 1640608721
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_100
timestamp 1640608721
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1640608721
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _0854_
timestamp 1640608721
transform -1 0 9568 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0952_
timestamp 1640608721
transform 1 0 9568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0956_
timestamp 1640608721
transform 1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__S
timestamp 1640608721
transform 1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_112
timestamp 1640608721
transform 1 0 11408 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1228_
timestamp 1640608721
transform -1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__S
timestamp 1640608721
transform 1 0 13248 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__S
timestamp 1640608721
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_129
timestamp 1640608721
transform 1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_134
timestamp 1640608721
transform 1 0 13432 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1640608721
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1236_
timestamp 1640608721
transform 1 0 14076 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_159
timestamp 1640608721
transform 1 0 15732 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1219_
timestamp 1640608721
transform 1 0 16192 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1243_
timestamp 1640608721
transform 1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clk
timestamp 1640608721
transform -1 0 16192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _0976_
timestamp 1640608721
transform 1 0 17756 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1157_
timestamp 1640608721
transform 1 0 17020 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__S
timestamp 1640608721
transform 1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__S
timestamp 1640608721
transform 1 0 19596 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1640608721
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1640608721
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_203
timestamp 1640608721
transform 1 0 19780 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1640608721
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0977_
timestamp 1640608721
transform -1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__S
timestamp 1640608721
transform 1 0 21160 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp 1640608721
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1273_
timestamp 1640608721
transform 1 0 22172 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1279_
timestamp 1640608721
transform -1 0 22172 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_241
timestamp 1640608721
transform 1 0 23276 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 1640608721
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0984_
timestamp 1640608721
transform 1 0 23000 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1640608721
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1640608721
transform 1 0 25484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_269
timestamp 1640608721
transform 1 0 25852 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1640608721
transform -1 0 26220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1640608721
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1640608721
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1640608721
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1394_
timestamp 1640608721
transform -1 0 3036 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1395_
timestamp 1640608721
transform 1 0 3036 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1397_
timestamp 1640608721
transform 1 0 4600 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1640608721
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1640608721
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1640608721
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0955_
timestamp 1640608721
transform 1 0 6532 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0954_
timestamp 1640608721
transform 1 0 8648 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1364_
timestamp 1640608721
transform 1 0 7084 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1640608721
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_103
timestamp 1640608721
transform 1 0 10580 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_91
timestamp 1640608721
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A1
timestamp 1640608721
transform 1 0 12328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__S
timestamp 1640608721
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_109
timestamp 1640608721
transform 1 0 11132 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_124
timestamp 1640608721
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1640608721
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1227_
timestamp 1640608721
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A2
timestamp 1640608721
transform 1 0 12880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__B1
timestamp 1640608721
transform 1 0 12696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_133
timestamp 1640608721
transform 1 0 13340 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1070_
timestamp 1640608721
transform -1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1072_
timestamp 1640608721
transform -1 0 14536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1235_
timestamp 1640608721
transform -1 0 14260 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__S
timestamp 1640608721
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__S
timestamp 1640608721
transform 1 0 14720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__S
timestamp 1640608721
transform 1 0 14536 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_A
timestamp 1640608721
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_150
timestamp 1640608721
transform 1 0 14904 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_160
timestamp 1640608721
transform 1 0 15824 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1640608721
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1640608721
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1640608721
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1640608721
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__S
timestamp 1640608721
transform 1 0 19044 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1640608721
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_197
timestamp 1640608721
transform 1 0 19228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__S
timestamp 1640608721
transform 1 0 21988 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_209
timestamp 1640608721
transform 1 0 20332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1640608721
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1640608721
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_229
timestamp 1640608721
transform 1 0 22172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1640608721
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_241
timestamp 1640608721
transform 1 0 23276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_253
timestamp 1640608721
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_265
timestamp 1640608721
transform 1 0 25484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_269
timestamp 1640608721
transform 1 0 25852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1640608721
transform -1 0 26220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_11
timestamp 1640608721
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1640608721
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1640608721
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0871_
timestamp 1640608721
transform 1 0 2668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0872_
timestamp 1640608721
transform 1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_40
timestamp 1640608721
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1640608721
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0855_
timestamp 1640608721
transform -1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1640608721
transform -1 0 3680 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0869_
timestamp 1640608721
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_47
timestamp 1640608721
transform 1 0 5428 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_56
timestamp 1640608721
transform 1 0 6256 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0857_
timestamp 1640608721
transform -1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0863_
timestamp 1640608721
transform 1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A
timestamp 1640608721
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_64
timestamp 1640608721
transform 1 0 6992 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_74
timestamp 1640608721
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1640608721
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _0958_
timestamp 1640608721
transform -1 0 7728 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1640608721
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1640608721
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1640608721
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_109
timestamp 1640608721
transform 1 0 11132 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _1017_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 11408 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_2  _1191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 12236 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1640608721
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1016_
timestamp 1640608721
transform -1 0 13984 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1190_
timestamp 1640608721
transform 1 0 13064 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1326_
timestamp 1640608721
transform 1 0 14076 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__S
timestamp 1640608721
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_155
timestamp 1640608721
transform 1 0 15364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1096_
timestamp 1640608721
transform 1 0 14904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__S
timestamp 1640608721
transform 1 0 17296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_167
timestamp 1640608721
transform 1 0 16468 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_175
timestamp 1640608721
transform 1 0 17204 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1158_
timestamp 1640608721
transform 1 0 18308 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1294_
timestamp 1640608721
transform -1 0 18308 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1640608721
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1152_
timestamp 1640608721
transform 1 0 20056 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1159_
timestamp 1640608721
transform -1 0 19136 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1245_
timestamp 1640608721
transform 1 0 19228 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__S
timestamp 1640608721
transform 1 0 21620 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__S
timestamp 1640608721
transform 1 0 20884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__S
timestamp 1640608721
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1640608721
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_225
timestamp 1640608721
transform 1 0 21804 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_229
timestamp 1640608721
transform 1 0 22172 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1153_
timestamp 1640608721
transform -1 0 20884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__S
timestamp 1640608721
transform 1 0 22264 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_244
timestamp 1640608721
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1141_
timestamp 1640608721
transform -1 0 23552 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1272_
timestamp 1640608721
transform 1 0 22448 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1640608721
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_265
timestamp 1640608721
transform 1 0 25484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_269
timestamp 1640608721
transform 1 0 25852 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1640608721
transform -1 0 26220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1640608721
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_11
timestamp 1640608721
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1640608721
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1640608721
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1640608721
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1640608721
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0874_
timestamp 1640608721
transform 1 0 2392 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1393_
timestamp 1640608721
transform 1 0 1472 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_13_37
timestamp 1640608721
transform 1 0 4508 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1640608721
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1640608721
transform 1 0 4048 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1640608721
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0859_
timestamp 1640608721
transform -1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0867_
timestamp 1640608721
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0868_
timestamp 1640608721
transform 1 0 3404 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0870_
timestamp 1640608721
transform -1 0 4508 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0873_
timestamp 1640608721
transform -1 0 3588 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 1640608721
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1640608721
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1640608721
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_44
timestamp 1640608721
transform 1 0 5152 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1640608721
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0676_
timestamp 1640608721
transform -1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1459_
timestamp 1640608721
transform 1 0 5796 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1640608721
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1640608721
transform 1 0 8556 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_68
timestamp 1640608721
transform 1 0 7360 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_74
timestamp 1640608721
transform 1 0 7912 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0833_
timestamp 1640608721
transform -1 0 8832 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1405_
timestamp 1640608721
transform -1 0 10212 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__B
timestamp 1640608721
transform 1 0 10304 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_99
timestamp 1640608721
transform 1 0 10212 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1640608721
transform 1 0 10488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1640608721
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1064_
timestamp 1640608721
transform 1 0 10488 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1404_
timestamp 1640608721
transform -1 0 10488 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_13_107
timestamp 1640608721
transform 1 0 10948 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1640608721
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0702_
timestamp 1640608721
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1018_
timestamp 1640608721
transform 1 0 12420 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1403_
timestamp 1640608721
transform 1 0 10856 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1461_
timestamp 1640608721
transform 1 0 11500 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _1077_
timestamp 1640608721
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1071_
timestamp 1640608721
transform 1 0 13156 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_126
timestamp 1640608721
transform 1 0 12696 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_130
timestamp 1640608721
transform 1 0 13064 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__S
timestamp 1640608721
transform 1 0 13248 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1325_
timestamp 1640608721
transform -1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1085_
timestamp 1640608721
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1078_
timestamp 1640608721
transform 1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1640608721
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__S
timestamp 1640608721
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__S
timestamp 1640608721
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_164
timestamp 1640608721
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__and2_2  _1084_
timestamp 1640608721
transform 1 0 15640 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1220_
timestamp 1640608721
transform -1 0 16192 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1221_
timestamp 1640608721
transform -1 0 17020 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1251_
timestamp 1640608721
transform -1 0 15364 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1252_
timestamp 1640608721
transform -1 0 15640 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__S
timestamp 1640608721
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1640608721
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1217_
timestamp 1640608721
transform 1 0 17664 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1218_
timestamp 1640608721
transform 1 0 16836 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1241_
timestamp 1640608721
transform 1 0 17020 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1293_
timestamp 1640608721
transform 1 0 17848 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1299_
timestamp 1640608721
transform -1 0 19504 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1104_
timestamp 1640608721
transform -1 0 19780 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1098_
timestamp 1640608721
transform -1 0 18952 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1640608721
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__S
timestamp 1640608721
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__S
timestamp 1640608721
transform 1 0 18492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1280_
timestamp 1640608721
transform -1 0 20700 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1244_
timestamp 1640608721
transform 1 0 19596 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_203
timestamp 1640608721
transform 1 0 19780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_200
timestamp 1640608721
transform 1 0 19504 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1287_
timestamp 1640608721
transform 1 0 20424 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1281_
timestamp 1640608721
transform 1 0 20700 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1278_
timestamp 1640608721
transform 1 0 21804 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1275_
timestamp 1640608721
transform -1 0 22724 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1114_
timestamp 1640608721
transform -1 0 21804 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1640608721
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_225
timestamp 1640608721
transform 1 0 21804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1640608721
transform 1 0 21252 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__S
timestamp 1640608721
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__S
timestamp 1640608721
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__S
timestamp 1640608721
transform -1 0 24288 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1640608721
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _1126_
timestamp 1640608721
transform 1 0 23552 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1140_
timestamp 1640608721
transform 1 0 23460 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1230_
timestamp 1640608721
transform 1 0 22724 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1231_
timestamp 1640608721
transform 1 0 22632 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_261
timestamp 1640608721
transform 1 0 25116 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_269
timestamp 1640608721
transform 1 0 25852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_256
timestamp 1640608721
transform 1 0 24656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_268
timestamp 1640608721
transform 1 0 25760 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1640608721
transform -1 0 26220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1640608721
transform -1 0 26220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1640608721
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1127_
timestamp 1640608721
transform -1 0 24656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_15
timestamp 1640608721
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1640608721
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1640608721
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0875_
timestamp 1640608721
transform -1 0 3312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_24
timestamp 1640608721
transform 1 0 3312 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1640608721
transform 1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _0682_
timestamp 1640608721
transform 1 0 4600 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1640608721
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0681_
timestamp 1640608721
transform 1 0 5428 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1458_
timestamp 1640608721
transform 1 0 6348 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1339_
timestamp 1640608721
transform 1 0 7912 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__o221a_2  _0834_
timestamp 1640608721
transform 1 0 9476 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0835_
timestamp 1640608721
transform 1 0 10304 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1640608721
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1640608721
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_122
timestamp 1640608721
transform 1 0 12328 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1640608721
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0679_
timestamp 1640608721
transform 1 0 12052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1341_
timestamp 1640608721
transform 1 0 12420 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_15_140
timestamp 1640608721
transform 1 0 13984 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A
timestamp 1640608721
transform 1 0 15088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__S
timestamp 1640608721
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__S
timestamp 1640608721
transform -1 0 16192 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__S
timestamp 1640608721
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__S
timestamp 1640608721
transform -1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_161
timestamp 1640608721
transform 1 0 15916 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1090_
timestamp 1640608721
transform 1 0 15272 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__S
timestamp 1640608721
transform 1 0 18032 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_186
timestamp 1640608721
transform 1 0 18216 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1640608721
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1097_
timestamp 1640608721
transform 1 0 17480 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1242_
timestamp 1640608721
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__S
timestamp 1640608721
transform 1 0 20056 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__S
timestamp 1640608721
transform 1 0 19872 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__S
timestamp 1640608721
transform -1 0 18768 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1105_
timestamp 1640608721
transform 1 0 18768 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1274_
timestamp 1640608721
transform -1 0 21068 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1300_
timestamp 1640608721
transform -1 0 19872 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_217
timestamp 1640608721
transform 1 0 21068 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1640608721
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1640608721
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1146_
timestamp 1640608721
transform 1 0 21160 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1286_
timestamp 1640608721
transform 1 0 21804 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A
timestamp 1640608721
transform -1 0 24104 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_250
timestamp 1640608721
transform 1 0 24104 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1133_
timestamp 1640608721
transform -1 0 23920 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1271_
timestamp 1640608721
transform 1 0 22632 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_262
timestamp 1640608721
transform 1 0 25208 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1640608721
transform -1 0 26220 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1640608721
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1640608721
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1640608721
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0876_
timestamp 1640608721
transform 1 0 2300 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1640608721
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1640608721
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1640608721
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_39
timestamp 1640608721
transform 1 0 4692 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1640608721
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0687_
timestamp 1640608721
transform 1 0 3864 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0683_
timestamp 1640608721
transform 1 0 5244 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1460_
timestamp 1640608721
transform 1 0 6072 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_16_74
timestamp 1640608721
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1640608721
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0680_
timestamp 1640608721
transform -1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1640608721
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1640608721
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1259_
timestamp 1640608721
transform -1 0 9936 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1264_
timestamp 1640608721
transform -1 0 10764 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__S
timestamp 1640608721
transform -1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_107
timestamp 1640608721
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_119
timestamp 1640608721
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1640608721
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1640608721
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1640608721
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1640608721
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_A
timestamp 1640608721
transform 1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1640608721
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1640608721
transform 1 0 16100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1640608721
transform 1 0 15548 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1640608721
transform -1 0 16100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clk
timestamp 1640608721
transform -1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A
timestamp 1640608721
transform -1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_167
timestamp 1640608721
transform 1 0 16468 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1640608721
transform 1 0 17480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1640608721
transform 1 0 17204 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1164_
timestamp 1640608721
transform 1 0 16744 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1640608721
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1640608721
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1640608721
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1640608721
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _1113_
timestamp 1640608721
transform 1 0 19688 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1120_
timestamp 1640608721
transform 1 0 20240 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A
timestamp 1640608721
transform -1 0 20884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1640608721
transform -1 0 21160 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__S
timestamp 1640608721
transform 1 0 21620 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_215
timestamp 1640608721
transform 1 0 20884 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_218
timestamp 1640608721
transform 1 0 21160 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_225
timestamp 1640608721
transform 1 0 21804 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_229
timestamp 1640608721
transform 1 0 22172 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1640608721
transform 1 0 21344 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__S
timestamp 1640608721
transform 1 0 23276 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__S
timestamp 1640608721
transform 1 0 22264 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_243
timestamp 1640608721
transform 1 0 23460 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1277_
timestamp 1640608721
transform 1 0 22448 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1640608721
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1640608721
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_265
timestamp 1640608721
transform 1 0 25484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_269
timestamp 1640608721
transform 1 0 25852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1640608721
transform -1 0 26220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1640608721
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1640608721
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1640608721
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1392_
timestamp 1640608721
transform 1 0 1472 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_17_21
timestamp 1640608721
transform 1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1457_
timestamp 1640608721
transform 1 0 3772 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1640608721
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1640608721
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1640608721
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1640608721
transform 1 0 5336 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0675_
timestamp 1640608721
transform -1 0 5888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1021_
timestamp 1640608721
transform 1 0 6716 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1640608721
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_68
timestamp 1640608721
transform 1 0 7360 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_80
timestamp 1640608721
transform 1 0 8464 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__S
timestamp 1640608721
transform 1 0 9844 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_103
timestamp 1640608721
transform 1 0 10580 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0685_
timestamp 1640608721
transform -1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1019_
timestamp 1640608721
transform 1 0 10028 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1290_
timestamp 1640608721
transform 1 0 9016 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1640608721
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1640608721
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1640608721
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 1640608721
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1640608721
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1437_
timestamp 1640608721
transform 1 0 11960 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_17_139
timestamp 1640608721
transform 1 0 13892 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_clk
timestamp 1640608721
transform -1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__S
timestamp 1640608721
transform -1 0 16560 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_147
timestamp 1640608721
transform 1 0 14628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1640608721
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_2  _1087_
timestamp 1640608721
transform 1 0 14904 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1093_
timestamp 1640608721
transform 1 0 15732 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1640608721
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_185
timestamp 1640608721
transform 1 0 18124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1640608721
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1101_
timestamp 1640608721
transform -1 0 18124 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1161_
timestamp 1640608721
transform -1 0 17480 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_clk
timestamp 1640608721
transform 1 0 17480 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_197
timestamp 1640608721
transform 1 0 19228 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_205
timestamp 1640608721
transform 1 0 19964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1640608721
transform -1 0 20424 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_213
timestamp 1640608721
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1640608721
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1640608721
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1640608721
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1107_
timestamp 1640608721
transform -1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_233
timestamp 1640608721
transform 1 0 22540 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_239
timestamp 1640608721
transform 1 0 23092 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1130_
timestamp 1640608721
transform -1 0 23092 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_251
timestamp 1640608721
transform 1 0 24196 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_263
timestamp 1640608721
transform 1 0 25300 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_269
timestamp 1640608721
transform 1 0 25852 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1640608721
transform -1 0 26220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1640608721
transform 1 0 2116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1640608721
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1640608721
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0877_
timestamp 1640608721
transform 1 0 2944 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _0880_
timestamp 1640608721
transform 1 0 2208 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1640608721
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 1640608721
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1640608721
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1456_
timestamp 1640608721
transform 1 0 3864 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_A
timestamp 1640608721
transform 1 0 6440 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_50
timestamp 1640608721
transform 1 0 5704 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_60
timestamp 1640608721
transform 1 0 6624 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0686_
timestamp 1640608721
transform -1 0 5704 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0688_
timestamp 1640608721
transform -1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clk
timestamp 1640608721
transform 1 0 5796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__S
timestamp 1640608721
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__S
timestamp 1640608721
transform 1 0 8464 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_76
timestamp 1640608721
transform 1 0 8096 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0838_
timestamp 1640608721
transform -1 0 8464 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_clk
timestamp 1640608721
transform 1 0 7728 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B1
timestamp 1640608721
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__S
timestamp 1640608721
transform 1 0 10304 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1640608721
transform 1 0 10488 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1640608721
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0831_
timestamp 1640608721
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0832_
timestamp 1640608721
transform -1 0 9476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1233_
timestamp 1640608721
transform 1 0 9476 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0739_
timestamp 1640608721
transform 1 0 10856 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1436_
timestamp 1640608721
transform 1 0 11684 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_18_132
timestamp 1640608721
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1640608721
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1640608721
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__S
timestamp 1640608721
transform 1 0 14720 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_147
timestamp 1640608721
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1086_
timestamp 1640608721
transform -1 0 16192 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1207_
timestamp 1640608721
transform 1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1210_
timestamp 1640608721
transform -1 0 17020 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_178
timestamp 1640608721
transform 1 0 17480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1099_
timestamp 1640608721
transform 1 0 18308 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1100_
timestamp 1640608721
transform -1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1160_
timestamp 1640608721
transform -1 0 17480 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1640608721
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 1640608721
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_201
timestamp 1640608721
transform 1 0 19596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1640608721
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1109_
timestamp 1640608721
transform -1 0 19596 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1116_
timestamp 1640608721
transform 1 0 19964 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_217
timestamp 1640608721
transform 1 0 21068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_228
timestamp 1640608721
transform 1 0 22080 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _1115_
timestamp 1640608721
transform 1 0 20608 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1640608721
transform -1 0 22080 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1122_
timestamp 1640608721
transform 1 0 21252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__S
timestamp 1640608721
transform -1 0 22448 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_241
timestamp 1640608721
transform 1 0 23276 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1640608721
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1308_
timestamp 1640608721
transform 1 0 22448 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1640608721
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_265
timestamp 1640608721
transform 1 0 25484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_269
timestamp 1640608721
transform 1 0 25852 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1640608721
transform -1 0 26220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1640608721
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1640608721
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1640608721
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1640608721
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1640608721
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1640608721
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0690_
timestamp 1640608721
transform 1 0 2760 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _0878_
timestamp 1640608721
transform 1 0 2024 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1391_
timestamp 1640608721
transform 1 0 1472 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1640608721
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1640608721
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0689_
timestamp 1640608721
transform 1 0 3588 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0691_
timestamp 1640608721
transform -1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _0879_
timestamp 1640608721
transform -1 0 3588 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1455_
timestamp 1640608721
transform 1 0 3772 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1640608721
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_46
timestamp 1640608721
transform 1 0 5336 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1640608721
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0684_
timestamp 1640608721
transform -1 0 5888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1398_
timestamp 1640608721
transform -1 0 7912 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1400_
timestamp 1640608721
transform -1 0 8004 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_clk
timestamp 1640608721
transform -1 0 5612 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B1
timestamp 1640608721
transform 1 0 8740 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _0844_
timestamp 1640608721
transform -1 0 8832 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1269_
timestamp 1640608721
transform 1 0 7912 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__C1
timestamp 1640608721
transform 1 0 9200 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1640608721
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0738_
timestamp 1640608721
transform 1 0 10580 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0740_
timestamp 1640608721
transform 1 0 9752 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1640608721
transform -1 0 9200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0837_
timestamp 1640608721
transform 1 0 8924 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1402_
timestamp 1640608721
transform 1 0 9384 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B1
timestamp 1640608721
transform -1 0 12696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__B1
timestamp 1640608721
transform -1 0 11592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1640608721
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1640608721
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_111
timestamp 1640608721
transform 1 0 11316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_114
timestamp 1640608721
transform 1 0 11592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1640608721
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0736_
timestamp 1640608721
transform 1 0 11684 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1435_
timestamp 1640608721
transform 1 0 11592 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__S
timestamp 1640608721
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_126
timestamp 1640608721
transform 1 0 12696 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_132
timestamp 1640608721
transform 1 0 13248 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1640608721
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1640608721
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0827_
timestamp 1640608721
transform -1 0 14536 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1081_
timestamp 1640608721
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1438_
timestamp 1640608721
transform 1 0 13156 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_19_148
timestamp 1640608721
transform 1 0 14720 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_164
timestamp 1640608721
transform 1 0 16192 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0828_
timestamp 1640608721
transform 1 0 15364 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1208_
timestamp 1640608721
transform 1 0 14536 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1211_
timestamp 1640608721
transform 1 0 16284 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1406_
timestamp 1640608721
transform -1 0 16560 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_19_175
timestamp 1640608721
transform 1 0 17204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1640608721
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0733_
timestamp 1640608721
transform 1 0 17112 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1092_
timestamp 1640608721
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1204_
timestamp 1640608721
transform -1 0 18124 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1205_
timestamp 1640608721
transform 1 0 17940 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1439_
timestamp 1640608721
transform 1 0 18124 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_20_192
timestamp 1640608721
transform 1 0 18768 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1640608721
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1640608721
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0732_
timestamp 1640608721
transform -1 0 19136 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1108_
timestamp 1640608721
transform 1 0 19688 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1313_
timestamp 1640608721
transform 1 0 19320 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1319_
timestamp 1640608721
transform 1 0 20148 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__S
timestamp 1640608721
transform 1 0 20976 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_215
timestamp 1640608721
transform 1 0 20884 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1640608721
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1640608721
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0730_
timestamp 1640608721
transform -1 0 22264 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0731_
timestamp 1640608721
transform 1 0 21160 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _1106_
timestamp 1640608721
transform 1 0 20424 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1123_
timestamp 1640608721
transform 1 0 21068 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1440_
timestamp 1640608721
transform 1 0 21988 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1640608721
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0826_
timestamp 1640608721
transform 1 0 22264 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1128_
timestamp 1640608721
transform 1 0 23552 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1129_
timestamp 1640608721
transform -1 0 23736 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1407_
timestamp 1640608721
transform 1 0 23736 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_19_263
timestamp 1640608721
transform 1 0 25300 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_269
timestamp 1640608721
transform 1 0 25852 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1640608721
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_265
timestamp 1640608721
transform 1 0 25484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_269
timestamp 1640608721
transform 1 0 25852 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1640608721
transform -1 0 26220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1640608721
transform -1 0 26220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1640608721
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1640608721
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1640608721
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1390_
timestamp 1640608721
transform 1 0 1472 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1640608721
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1454_
timestamp 1640608721
transform 1 0 3404 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_21_42
timestamp 1640608721
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1640608721
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1640608721
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1640608721
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0841_
timestamp 1640608721
transform -1 0 7544 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0840_
timestamp 1640608721
transform 1 0 7544 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1234_
timestamp 1640608721
transform 1 0 8372 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__S
timestamp 1640608721
transform 1 0 9476 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1640608721
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0839_
timestamp 1640608721
transform -1 0 9476 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1640608721
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1640608721
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_116
timestamp 1640608721
transform 1 0 11776 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_124
timestamp 1640608721
transform 1 0 12512 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1640608721
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0735_
timestamp 1640608721
transform -1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_129
timestamp 1640608721
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0728_
timestamp 1640608721
transform 1 0 12696 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0836_
timestamp 1640608721
transform -1 0 13432 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1073_
timestamp 1640608721
transform -1 0 13892 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1080_
timestamp 1640608721
transform 1 0 13892 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__S
timestamp 1640608721
transform 1 0 16100 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_152
timestamp 1640608721
transform 1 0 15088 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_160
timestamp 1640608721
transform 1 0 15824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1640608721
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1079_
timestamp 1640608721
transform 1 0 14628 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__B1
timestamp 1640608721
transform -1 0 17112 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__S
timestamp 1640608721
transform 1 0 17112 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__S
timestamp 1640608721
transform 1 0 17756 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_169
timestamp 1640608721
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_176
timestamp 1640608721
transform 1 0 17296 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_180
timestamp 1640608721
transform 1 0 17664 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_183
timestamp 1640608721
transform 1 0 17940 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1640608721
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__S
timestamp 1640608721
transform 1 0 19044 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__S
timestamp 1640608721
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_191
timestamp 1640608721
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1314_
timestamp 1640608721
transform -1 0 20056 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1320_
timestamp 1640608721
transform -1 0 20884 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__S
timestamp 1640608721
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_215
timestamp 1640608721
transform 1 0 20884 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_221
timestamp 1640608721
transform 1 0 21436 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1640608721
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__or4_2  _1136_
timestamp 1640608721
transform 1 0 21804 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B1
timestamp 1640608721
transform -1 0 22632 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_243
timestamp 1640608721
transform 1 0 23460 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1307_
timestamp 1640608721
transform 1 0 22632 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_255
timestamp 1640608721
transform 1 0 24564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_267
timestamp 1640608721
transform 1 0 25668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1640608721
transform -1 0 26220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1640608721
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1640608721
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1640608721
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1640608721
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1640608721
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1453_
timestamp 1640608721
transform 1 0 3772 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1399_
timestamp 1640608721
transform -1 0 6900 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_22_63
timestamp 1640608721
transform 1 0 6900 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1401_
timestamp 1640608721
transform -1 0 8832 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1640608721
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1640608721
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1640608721
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1434_
timestamp 1640608721
transform 1 0 10396 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_22_124
timestamp 1640608721
transform 1 0 12512 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0734_
timestamp 1640608721
transform -1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0737_
timestamp 1640608721
transform -1 0 12512 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1065_
timestamp 1640608721
transform 1 0 12604 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__S
timestamp 1640608721
transform 1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1640608721
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1074_
timestamp 1640608721
transform -1 0 13984 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1214_
timestamp 1640608721
transform -1 0 14904 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_150
timestamp 1640608721
transform 1 0 14904 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_162
timestamp 1640608721
transform 1 0 16008 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_174
timestamp 1640608721
transform 1 0 17112 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_186
timestamp 1640608721
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__S
timestamp 1640608721
transform 1 0 19872 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1640608721
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 1640608721
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_203
timestamp 1640608721
transform 1 0 19780 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_206
timestamp 1640608721
transform 1 0 20056 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1640608721
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_213
timestamp 1640608721
transform 1 0 20700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_225
timestamp 1640608721
transform 1 0 21804 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0822_
timestamp 1640608721
transform 1 0 20424 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1137_
timestamp 1640608721
transform -1 0 22816 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_244
timestamp 1640608721
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1134_
timestamp 1640608721
transform -1 0 23552 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1135_
timestamp 1640608721
transform -1 0 23276 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1640608721
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_265
timestamp 1640608721
transform 1 0 25484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_269
timestamp 1640608721
transform 1 0 25852 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1640608721
transform -1 0 26220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1640608721
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1640608721
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1640608721
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1640608721
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1640608721
transform 1 0 3588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_31
timestamp 1640608721
transform 1 0 3956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0692_
timestamp 1640608721
transform -1 0 5152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0693_
timestamp 1640608721
transform -1 0 4876 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_44
timestamp 1640608721
transform 1 0 5152 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1640608721
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1640608721
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0842_
timestamp 1640608721
transform -1 0 7268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__S
timestamp 1640608721
transform 1 0 8096 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_78
timestamp 1640608721
transform 1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1267_
timestamp 1640608721
transform 1 0 7268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__B1
timestamp 1640608721
transform 1 0 9476 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_90
timestamp 1640608721
transform 1 0 9384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0743_
timestamp 1640608721
transform 1 0 9660 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0749_
timestamp 1640608721
transform -1 0 10764 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1640608721
transform 1 0 11960 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1640608721
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1640608721
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1640608721
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1640608721
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1640608721
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_2  _1066_
timestamp 1640608721
transform -1 0 12880 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 12880 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp 1640608721
transform 1 0 15548 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1640608721
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1213_
timestamp 1640608721
transform 1 0 14720 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 1640608721
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_176
timestamp 1640608721
transform 1 0 17296 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1640608721
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0724_
timestamp 1640608721
transform 1 0 16744 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0725_
timestamp 1640608721
transform 1 0 17020 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1155_
timestamp 1640608721
transform 1 0 18032 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_195
timestamp 1640608721
transform 1 0 19044 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_207
timestamp 1640608721
transform 1 0 20148 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0814_
timestamp 1640608721
transform 1 0 18768 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B1
timestamp 1640608721
transform -1 0 20884 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_225
timestamp 1640608721
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1640608721
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0729_
timestamp 1640608721
transform 1 0 20884 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1441_
timestamp 1640608721
transform 1 0 21896 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_23_246
timestamp 1640608721
transform 1 0 23736 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0727_
timestamp 1640608721
transform 1 0 23460 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_258
timestamp 1640608721
transform 1 0 24840 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1640608721
transform -1 0 26220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_15
timestamp 1640608721
transform 1 0 2484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1640608721
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1640608721
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1031_
timestamp 1640608721
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1640608721
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1640608721
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1640608721
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1640608721
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_53
timestamp 1640608721
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_61
timestamp 1640608721
transform 1 0 6716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__S
timestamp 1640608721
transform 1 0 7728 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1640608721
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1640608721
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1303_
timestamp 1640608721
transform -1 0 7728 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B1
timestamp 1640608721
transform 1 0 9752 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1640608721
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_93
timestamp 1640608721
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1640608721
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1433_
timestamp 1640608721
transform 1 0 9936 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__S
timestamp 1640608721
transform 1 0 12236 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_113
timestamp 1640608721
transform 1 0 11500 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1067_
timestamp 1640608721
transform -1 0 12696 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1640608721
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1640608721
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1640608721
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1640608721
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1075_
timestamp 1640608721
transform -1 0 13800 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1260_
timestamp 1640608721
transform -1 0 13524 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__S
timestamp 1640608721
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_151
timestamp 1640608721
transform 1 0 14996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0719_
timestamp 1640608721
transform 1 0 14536 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1446_
timestamp 1640608721
transform 1 0 15548 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1445_
timestamp 1640608721
transform 1 0 17112 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_24_200
timestamp 1640608721
transform 1 0 19504 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_208
timestamp 1640608721
transform 1 0 20240 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1640608721
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1154_
timestamp 1640608721
transform -1 0 19136 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1156_
timestamp 1640608721
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B1
timestamp 1640608721
transform 1 0 22172 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1640608721
transform 1 0 21252 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0726_
timestamp 1640608721
transform 1 0 21344 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1143_
timestamp 1640608721
transform -1 0 21252 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1640608721
transform -1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__S
timestamp 1640608721
transform 1 0 22632 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_231
timestamp 1640608721
transform 1 0 22356 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1640608721
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1322_
timestamp 1640608721
transform 1 0 22816 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1640608721
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1640608721
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1640608721
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_269
timestamp 1640608721
transform 1 0 25852 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1640608721
transform -1 0 26220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1640608721
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1640608721
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1640608721
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1640608721
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1334_
timestamp 1640608721
transform 1 0 1840 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__S
timestamp 1640608721
transform 1 0 4324 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_25
timestamp 1640608721
transform 1 0 3404 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1640608721
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1289_
timestamp 1640608721
transform -1 0 4324 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1640608721
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1640608721
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1640608721
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0790_
timestamp 1640608721
transform -1 0 7176 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1640608721
transform 1 0 8004 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B1
timestamp 1640608721
transform 1 0 8188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_79
timestamp 1640608721
transform 1 0 8372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _0791_
timestamp 1640608721
transform -1 0 8004 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0747_
timestamp 1640608721
transform 1 0 8924 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1431_
timestamp 1640608721
transform 1 0 9752 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__S
timestamp 1640608721
transform 1 0 12236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1640608721
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_116
timestamp 1640608721
transform 1 0 11776 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_120
timestamp 1640608721
transform 1 0 12144 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1640608721
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0741_
timestamp 1640608721
transform -1 0 11776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0745_
timestamp 1640608721
transform -1 0 12696 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0703_
timestamp 1640608721
transform -1 0 14628 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1255_
timestamp 1640608721
transform 1 0 13524 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1256_
timestamp 1640608721
transform -1 0 13524 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B1
timestamp 1640608721
transform 1 0 15088 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_147
timestamp 1640608721
transform 1 0 14628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_151
timestamp 1640608721
transform 1 0 14996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1640608721
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0715_
timestamp 1640608721
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0718_
timestamp 1640608721
transform 1 0 15272 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__S
timestamp 1640608721
transform 1 0 18216 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1640608721
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1444_
timestamp 1640608721
transform 1 0 16652 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_25_197
timestamp 1640608721
transform 1 0 19228 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0815_
timestamp 1640608721
transform -1 0 19780 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1142_
timestamp 1640608721
transform 1 0 19780 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1149_
timestamp 1640608721
transform 1 0 20240 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1304_
timestamp 1640608721
transform 1 0 18400 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1640608721
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1640608721
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1640608721
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1148_
timestamp 1640608721
transform -1 0 21436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1442_
timestamp 1640608721
transform 1 0 22080 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_25_245
timestamp 1640608721
transform 1 0 23644 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1408_
timestamp 1640608721
transform 1 0 24012 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_25_266
timestamp 1640608721
transform 1 0 25576 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1640608721
transform -1 0 26220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1640608721
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1640608721
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1640608721
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1640608721
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1640608721
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1333_
timestamp 1640608721
transform 1 0 2116 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1335_
timestamp 1640608721
transform 1 0 1840 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__S
timestamp 1640608721
transform 1 0 4600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_25
timestamp 1640608721
transform 1 0 3404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1640608721
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1033_
timestamp 1640608721
transform -1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1268_
timestamp 1640608721
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1292_
timestamp 1640608721
transform 1 0 3772 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1426_
timestamp 1640608721
transform 1 0 4784 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_27_46
timestamp 1640608721
transform 1 0 5336 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1640608721
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0792_
timestamp 1640608721
transform -1 0 6256 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1424_
timestamp 1640608721
transform -1 0 7912 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1425_
timestamp 1640608721
transform -1 0 7912 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__B1
timestamp 1640608721
transform -1 0 8832 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_74
timestamp 1640608721
transform 1 0 7912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_80
timestamp 1640608721
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_83
timestamp 1640608721
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0746_
timestamp 1640608721
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0788_
timestamp 1640608721
transform -1 0 8740 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B1
timestamp 1640608721
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_102
timestamp 1640608721
transform 1 0 10488 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1640608721
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0742_
timestamp 1640608721
transform -1 0 9384 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0748_
timestamp 1640608721
transform 1 0 8832 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0750_
timestamp 1640608721
transform 1 0 9660 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1432_
timestamp 1640608721
transform 1 0 9384 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__S
timestamp 1640608721
transform 1 0 12512 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_110
timestamp 1640608721
transform 1 0 11224 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_122
timestamp 1640608721
transform 1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1640608721
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1640608721
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_125
timestamp 1640608721
transform 1 0 12604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1640608721
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1640608721
transform 1 0 10948 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1020_
timestamp 1640608721
transform 1 0 11040 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1261_
timestamp 1640608721
transform 1 0 12696 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0706_
timestamp 1640608721
transform 1 0 13432 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_131
timestamp 1640608721
transform 1 0 13156 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__S
timestamp 1640608721
transform 1 0 13524 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A1
timestamp 1640608721
transform 1 0 13248 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A1
timestamp 1640608721
transform 1 0 12972 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1640608721
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1640608721
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_143
timestamp 1640608721
transform 1 0 14260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1640608721
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B1
timestamp 1640608721
transform -1 0 15548 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_153
timestamp 1640608721
transform 1 0 15180 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_155
timestamp 1640608721
transform 1 0 15364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0717_
timestamp 1640608721
transform 1 0 15548 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0721_
timestamp 1640608721
transform 1 0 15824 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0720_
timestamp 1640608721
transform 1 0 16652 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1640608721
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_175
timestamp 1640608721
transform 1 0 17204 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp 1640608721
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1640608721
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B1
timestamp 1640608721
transform 1 0 17296 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_2  _0818_
timestamp 1640608721
transform 1 0 17664 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0723_
timestamp 1640608721
transform 1 0 17480 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B1
timestamp 1640608721
transform -1 0 17664 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1305_
timestamp 1640608721
transform 1 0 18308 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1
timestamp 1640608721
transform 1 0 18492 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__S
timestamp 1640608721
transform 1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1640608721
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_205
timestamp 1640608721
transform 1 0 19964 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1640608721
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1443_
timestamp 1640608721
transform 1 0 19228 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1283_
timestamp 1640608721
transform -1 0 21804 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0722_
timestamp 1640608721
transform -1 0 20792 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1640608721
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__S
timestamp 1640608721
transform 1 0 20792 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A1
timestamp 1640608721
transform -1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1284_
timestamp 1640608721
transform 1 0 21804 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1640608721
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_220
timestamp 1640608721
transform 1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_225
timestamp 1640608721
transform 1 0 21804 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__S
timestamp 1640608721
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__S
timestamp 1640608721
transform 1 0 22448 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_231
timestamp 1640608721
transform 1 0 22356 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_234
timestamp 1640608721
transform 1 0 22632 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1640608721
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_243
timestamp 1640608721
transform 1 0 23460 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _0825_
timestamp 1640608721
transform 1 0 22816 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1323_
timestamp 1640608721
transform 1 0 22632 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1640608721
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1640608721
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_265
timestamp 1640608721
transform 1 0 25484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_269
timestamp 1640608721
transform 1 0 25852 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_255
timestamp 1640608721
transform 1 0 24564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_267
timestamp 1640608721
transform 1 0 25668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1640608721
transform -1 0 26220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1640608721
transform -1 0 26220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1640608721
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_15
timestamp 1640608721
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1640608721
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1640608721
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1030_
timestamp 1640608721
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__S
timestamp 1640608721
transform 1 0 4600 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__S
timestamp 1640608721
transform 1 0 4784 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1640608721
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1640608721
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1291_
timestamp 1640608721
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B1
timestamp 1640608721
transform -1 0 6440 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1640608721
transform 1 0 4968 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_54
timestamp 1640608721
transform 1 0 6072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_58
timestamp 1640608721
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1427_
timestamp 1640608721
transform -1 0 8280 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1640608721
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__B1
timestamp 1640608721
transform 1 0 9568 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B
timestamp 1640608721
transform 1 0 10304 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_102
timestamp 1640608721
transform 1 0 10488 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1640608721
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1640608721
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0716_
timestamp 1640608721
transform 1 0 10580 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0800_
timestamp 1640608721
transform 1 0 9752 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0829_
timestamp 1640608721
transform -1 0 9568 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_28_106
timestamp 1640608721
transform 1 0 10856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1340_
timestamp 1640608721
transform 1 0 11592 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1640608721
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0705_
timestamp 1640608721
transform 1 0 13156 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1448_
timestamp 1640608721
transform 1 0 14076 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_28_158
timestamp 1640608721
transform 1 0 15640 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_170
timestamp 1640608721
transform 1 0 16744 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_177
timestamp 1640608721
transform 1 0 17388 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1412_
timestamp 1640608721
transform -1 0 19136 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_clk
timestamp 1640608721
transform -1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__S
timestamp 1640608721
transform 1 0 19964 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1640608721
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1640608721
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1296_
timestamp 1640608721
transform 1 0 20148 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_216
timestamp 1640608721
transform 1 0 20976 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0819_
timestamp 1640608721
transform 1 0 22172 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0820_
timestamp 1640608721
transform 1 0 21068 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0823_
timestamp 1640608721
transform 1 0 21344 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_241
timestamp 1640608721
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1640608721
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0821_
timestamp 1640608721
transform 1 0 22448 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1640608721
transform -1 0 26220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1640608721
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1411_
timestamp 1640608721
transform 1 0 24380 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1640608721
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1640608721
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1640608721
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1336_
timestamp 1640608721
transform 1 0 1840 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_29_33
timestamp 1640608721
transform 1 0 4140 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_41
timestamp 1640608721
transform 1 0 4876 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_2  _1034_
timestamp 1640608721
transform 1 0 3404 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_46
timestamp 1640608721
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1640608721
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1640608721
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1640608721
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0786_
timestamp 1640608721
transform 1 0 6532 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0787_
timestamp 1640608721
transform -1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_clk
timestamp 1640608721
transform -1 0 5336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A
timestamp 1640608721
transform -1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_A
timestamp 1640608721
transform 1 0 7636 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_65
timestamp 1640608721
transform 1 0 7084 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_73
timestamp 1640608721
transform 1 0 7820 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_81
timestamp 1640608721
transform 1 0 8556 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_103
timestamp 1640608721
transform 1 0 10580 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_94
timestamp 1640608721
transform 1 0 9752 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0707_
timestamp 1640608721
transform 1 0 8832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1640608721
transform -1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0713_
timestamp 1640608721
transform -1 0 10304 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1640608721
transform 1 0 10304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_clk
timestamp 1640608721
transform 1 0 9108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1640608721
transform 1 0 11684 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1640608721
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1640608721
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1640608721
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0694_
timestamp 1640608721
transform 1 0 11868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1449_
timestamp 1640608721
transform 1 0 12144 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_29_137
timestamp 1640608721
transform 1 0 13708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_141
timestamp 1640608721
transform 1 0 14076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1447_
timestamp 1640608721
transform 1 0 14168 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1640608721
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1640608721
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1640608721
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_177
timestamp 1640608721
transform 1 0 17388 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1640608721
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0811_
timestamp 1640608721
transform 1 0 18308 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0817_
timestamp 1640608721
transform 1 0 17480 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__S
timestamp 1640608721
transform 1 0 19596 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_193
timestamp 1640608721
transform 1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0812_
timestamp 1640608721
transform -1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1297_
timestamp 1640608721
transform 1 0 19780 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_29_212
timestamp 1640608721
transform 1 0 20608 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_228
timestamp 1640608721
transform 1 0 22080 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1640608721
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1640608721
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0802_
timestamp 1640608721
transform -1 0 22080 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0804_
timestamp 1640608721
transform -1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A1
timestamp 1640608721
transform -1 0 23368 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_242
timestamp 1640608721
transform 1 0 23368 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _0824_
timestamp 1640608721
transform 1 0 22356 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_254
timestamp 1640608721
transform 1 0 24472 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_266
timestamp 1640608721
transform 1 0 25576 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1640608721
transform -1 0 26220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1640608721
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1640608721
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1332_
timestamp 1640608721
transform 1 0 2116 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1640608721
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1640608721
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1640608721
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B1
timestamp 1640608721
transform 1 0 6808 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_53
timestamp 1640608721
transform 1 0 5980 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_58
timestamp 1640608721
transform 1 0 6440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1640608721
transform -1 0 6808 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0793_
timestamp 1640608721
transform -1 0 6440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A
timestamp 1640608721
transform 1 0 8188 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B
timestamp 1640608721
transform -1 0 8188 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_64
timestamp 1640608721
transform 1 0 6992 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_74
timestamp 1640608721
transform 1 0 7912 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _0711_
timestamp 1640608721
transform 1 0 8372 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0789_
timestamp 1640608721
transform -1 0 7912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clk
timestamp 1640608721
transform -1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A2
timestamp 1640608721
transform -1 0 10120 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1640608721
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0696_
timestamp 1640608721
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _0712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 9200 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _0779_
timestamp 1640608721
transform 1 0 10120 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_106
timestamp 1640608721
transform 1 0 10856 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_116
timestamp 1640608721
transform 1 0 11776 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_2  _0704_
timestamp 1640608721
transform -1 0 13156 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1302_
timestamp 1640608721
transform -1 0 11776 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_131
timestamp 1640608721
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1640608721
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1640608721
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1416_
timestamp 1640608721
transform -1 0 15640 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__S
timestamp 1640608721
transform 1 0 16284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_164
timestamp 1640608721
transform 1 0 16192 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0803_
timestamp 1640608721
transform -1 0 15916 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0805_
timestamp 1640608721
transform -1 0 16192 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_176
timestamp 1640608721
transform 1 0 17296 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0813_
timestamp 1640608721
transform 1 0 17388 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0816_
timestamp 1640608721
transform 1 0 18216 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1317_
timestamp 1640608721
transform -1 0 17296 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1640608721
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1640608721
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1414_
timestamp 1640608721
transform 1 0 19228 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1410_
timestamp 1640608721
transform -1 0 22724 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_clk
timestamp 1640608721
transform 1 0 20792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1409_
timestamp 1640608721
transform -1 0 24288 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1640608721
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_265
timestamp 1640608721
transform 1 0 25484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_269
timestamp 1640608721
transform 1 0 25852 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1640608721
transform -1 0 26220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1640608721
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_15
timestamp 1640608721
transform 1 0 2484 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1640608721
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1640608721
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1028_
timestamp 1640608721
transform 1 0 2668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A1
timestamp 1640608721
transform 1 0 3404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__S
timestamp 1640608721
transform 1 0 4416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_38
timestamp 1640608721
transform 1 0 4600 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1238_
timestamp 1640608721
transform -1 0 4416 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1423_
timestamp 1640608721
transform 1 0 4692 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1640608721
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0795_
timestamp 1640608721
transform -1 0 7176 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A
timestamp 1640608721
transform 1 0 7912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_72
timestamp 1640608721
transform 1 0 7728 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_81
timestamp 1640608721
transform 1 0 8556 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _0780_
timestamp 1640608721
transform 1 0 8648 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0784_
timestamp 1640608721
transform -1 0 8556 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0794_
timestamp 1640608721
transform -1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0959_
timestamp 1640608721
transform -1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1640608721
transform 1 0 10672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1429_
timestamp 1640608721
transform 1 0 9108 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_31_107
timestamp 1640608721
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1640608721
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1640608721
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0697_
timestamp 1640608721
transform 1 0 12328 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0698_
timestamp 1640608721
transform 1 0 11500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0796_
timestamp 1640608721
transform -1 0 12880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_128
timestamp 1640608721
transform 1 0 12880 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_132
timestamp 1640608721
transform 1 0 13248 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_136
timestamp 1640608721
transform 1 0 13616 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0807_
timestamp 1640608721
transform 1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0810_
timestamp 1640608721
transform 1 0 13984 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A1
timestamp 1640608721
transform 1 0 15456 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_149
timestamp 1640608721
transform 1 0 14812 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_155
timestamp 1640608721
transform 1 0 15364 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_158
timestamp 1640608721
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1640608721
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__S
timestamp 1640608721
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1640608721
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_173
timestamp 1640608721
transform 1 0 17020 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1640608721
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1413_
timestamp 1640608721
transform -1 0 18952 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1415_
timestamp 1640608721
transform 1 0 18952 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__S
timestamp 1640608721
transform 1 0 22172 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_211
timestamp 1640608721
transform 1 0 20516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1640608721
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1640608721
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1640608721
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__S
timestamp 1640608721
transform 1 0 22356 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_242
timestamp 1640608721
transform 1 0 23368 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1310_
timestamp 1640608721
transform 1 0 22540 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_31_254
timestamp 1640608721
transform 1 0 24472 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_266
timestamp 1640608721
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1640608721
transform -1 0 26220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1640608721
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1640608721
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1331_
timestamp 1640608721
transform 1 0 1748 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1640608721
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_37
timestamp 1640608721
transform 1 0 4508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1640608721
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1029_
timestamp 1640608721
transform -1 0 3588 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1035_
timestamp 1640608721
transform -1 0 4508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_45
timestamp 1640608721
transform 1 0 5244 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1422_
timestamp 1640608721
transform -1 0 6900 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A
timestamp 1640608721
transform 1 0 7360 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_63
timestamp 1640608721
transform 1 0 6900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_67
timestamp 1640608721
transform 1 0 7268 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_73
timestamp 1640608721
transform 1 0 7820 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1640608721
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0775_
timestamp 1640608721
transform 1 0 7544 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0776_
timestamp 1640608721
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0782_
timestamp 1640608721
transform -1 0 8372 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__S
timestamp 1640608721
transform 1 0 9384 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_95
timestamp 1640608721
transform 1 0 9844 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1640608721
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0781_
timestamp 1640608721
transform -1 0 9384 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1640608721
transform -1 0 9844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1265_
timestamp 1640608721
transform -1 0 10764 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_105
timestamp 1640608721
transform 1 0 10764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_113
timestamp 1640608721
transform 1 0 11500 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1452_
timestamp 1640608721
transform 1 0 11776 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1640608721
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1640608721
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1640608721
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1640608721
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0809_
timestamp 1640608721
transform 1 0 14628 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1417_
timestamp 1640608721
transform 1 0 15456 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_A
timestamp 1640608721
transform 1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_182
timestamp 1640608721
transform 1 0 17848 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1316_
timestamp 1640608721
transform 1 0 17020 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clk
timestamp 1640608721
transform 1 0 18216 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_190
timestamp 1640608721
transform 1 0 18584 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1640608721
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1640608721
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1640608721
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_221
timestamp 1640608721
transform 1 0 21436 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0917_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 21712 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_32_240
timestamp 1640608721
transform 1 0 23184 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1311_
timestamp 1640608721
transform 1 0 22356 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 1640608721
transform 1 0 25208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_253
timestamp 1640608721
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_264
timestamp 1640608721
transform 1 0 25392 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1640608721
transform -1 0 26220 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1640608721
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1640608721
transform -1 0 25208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_11
timestamp 1640608721
transform 1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1640608721
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1640608721
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1640608721
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1640608721
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1036_
timestamp 1640608721
transform 1 0 2392 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1330_
timestamp 1640608721
transform 1 0 1472 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _1239_
timestamp 1640608721
transform 1 0 3128 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1216_
timestamp 1640608721
transform 1 0 3772 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1640608721
transform -1 0 3496 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1025_
timestamp 1640608721
transform 1 0 3956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1640608721
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1640608721
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_21
timestamp 1640608721
transform 1 0 3036 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1032_
timestamp 1640608721
transform 1 0 4600 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _0799_
timestamp 1640608721
transform -1 0 5428 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__S
timestamp 1640608721
transform 1 0 4232 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__B1
timestamp 1640608721
transform 1 0 4416 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1420_
timestamp 1640608721
transform -1 0 6440 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1640608721
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0797_
timestamp 1640608721
transform -1 0 7176 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0798_
timestamp 1640608721
transform 1 0 5428 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1421_
timestamp 1640608721
transform -1 0 8004 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B1
timestamp 1640608721
transform 1 0 7176 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__B1
timestamp 1640608721
transform 1 0 7360 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_70
timestamp 1640608721
transform 1 0 7544 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_2  _0783_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 8004 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1024_
timestamp 1640608721
transform -1 0 8648 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1270_
timestamp 1640608721
transform 1 0 8648 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1640608721
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1640608721
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1640608721
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_93
timestamp 1640608721
transform 1 0 9660 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A2
timestamp 1640608721
transform -1 0 9752 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B
timestamp 1640608721
transform 1 0 9476 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_2  _1170_
timestamp 1640608721
transform -1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1640608721
transform -1 0 10028 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_104
timestamp 1640608721
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__S
timestamp 1640608721
transform 1 0 10028 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A0
timestamp 1640608721
transform 1 0 10488 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1640608721
transform 1 0 10212 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1640608721
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_111
timestamp 1640608721
transform 1 0 11316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1640608721
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0699_
timestamp 1640608721
transform 1 0 11592 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1450_
timestamp 1640608721
transform 1 0 12420 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1451_
timestamp 1640608721
transform 1 0 12236 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1640608721
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1640608721
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _0700_
timestamp 1640608721
transform 1 0 13800 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1419_
timestamp 1640608721
transform 1 0 14444 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1640608721
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_162
timestamp 1640608721
transform 1 0 16008 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_2  _0806_
timestamp 1640608721
transform 1 0 14628 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _0808_
timestamp 1640608721
transform 1 0 15456 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__S
timestamp 1640608721
transform 1 0 17940 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__S
timestamp 1640608721
transform 1 0 17480 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1640608721
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1640608721
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_174
timestamp 1640608721
transform 1 0 17112 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_180
timestamp 1640608721
transform 1 0 17664 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_185
timestamp 1640608721
transform 1 0 18124 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1640608721
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0911_
timestamp 1640608721
transform 1 0 18216 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1298_
timestamp 1640608721
transform 1 0 19228 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0912_
timestamp 1640608721
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1640608721
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_197
timestamp 1640608721
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_193
timestamp 1640608721
transform 1 0 18860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__S
timestamp 1640608721
transform 1 0 19044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _1186_
timestamp 1640608721
transform -1 0 20148 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _0915_
timestamp 1640608721
transform 1 0 20056 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_33_207
timestamp 1640608721
transform 1 0 20148 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_201
timestamp 1640608721
transform 1 0 19596 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__S
timestamp 1640608721
transform 1 0 20700 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__S
timestamp 1640608721
transform 1 0 21896 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_225
timestamp 1640608721
transform 1 0 21804 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1640608721
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1285_
timestamp 1640608721
transform 1 0 20884 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1312_
timestamp 1640608721
transform 1 0 22080 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1381_
timestamp 1640608721
transform -1 0 22264 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_33_237
timestamp 1640608721
transform 1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1640608721
transform 1 0 23644 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1640608721
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _0767_
timestamp 1640608721
transform -1 0 23644 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0916_
timestamp 1640608721
transform -1 0 22540 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1380_
timestamp 1640608721
transform 1 0 22540 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1640608721
transform 1 0 24748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_269
timestamp 1640608721
transform 1 0 25852 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1640608721
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1640608721
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_269
timestamp 1640608721
transform 1 0 25852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1640608721
transform -1 0 26220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1640608721
transform -1 0 26220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1640608721
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_15
timestamp 1640608721
transform 1 0 2484 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1640608721
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1640608721
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1037_
timestamp 1640608721
transform 1 0 2576 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__S
timestamp 1640608721
transform 1 0 4600 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__S
timestamp 1640608721
transform 1 0 4784 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_27
timestamp 1640608721
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_37
timestamp 1640608721
transform 1 0 4508 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1027_
timestamp 1640608721
transform -1 0 3588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1240_
timestamp 1640608721
transform 1 0 3680 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_35_42
timestamp 1640608721
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1640608721
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1640608721
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1640608721
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_A
timestamp 1640608721
transform 1 0 7268 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_65
timestamp 1640608721
transform 1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1640608721
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0773_
timestamp 1640608721
transform -1 0 8832 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A2
timestamp 1640608721
transform 1 0 10304 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_102
timestamp 1640608721
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _0756_
timestamp 1640608721
transform 1 0 8832 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_2  _0774_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 9384 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1640608721
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1640608721
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1365_
timestamp 1640608721
transform -1 0 13064 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_35_130
timestamp 1640608721
transform 1 0 13064 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_142
timestamp 1640608721
transform 1 0 14168 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_150
timestamp 1640608721
transform 1 0 14904 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1418_
timestamp 1640608721
transform 1 0 14996 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1640608721
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0909_
timestamp 1640608721
transform 1 0 17480 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1306_
timestamp 1640608721
transform 1 0 18124 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1318_
timestamp 1640608721
transform 1 0 16652 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _0769_
timestamp 1640608721
transform -1 0 19504 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _1187_
timestamp 1640608721
transform 1 0 19504 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1188_
timestamp 1640608721
transform -1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_216
timestamp 1640608721
transform 1 0 20976 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1640608721
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0768_
timestamp 1640608721
transform -1 0 21712 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1185_
timestamp 1640608721
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_244
timestamp 1640608721
transform 1 0 23552 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0918_
timestamp 1640608721
transform 1 0 22540 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1184_
timestamp 1640608721
transform 1 0 22816 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_256
timestamp 1640608721
transform 1 0 24656 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_268
timestamp 1640608721
transform 1 0 25760 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1640608721
transform -1 0 26220 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1640608721
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1640608721
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1329_
timestamp 1640608721
transform 1 0 1932 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1640608721
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_37
timestamp 1640608721
transform 1 0 4508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1640608721
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _1038_
timestamp 1640608721
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_49
timestamp 1640608721
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_61
timestamp 1640608721
transform 1 0 6716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1428_
timestamp 1640608721
transform -1 0 8832 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clk
timestamp 1640608721
transform -1 0 7268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1640608721
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1640608721
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0753_
timestamp 1640608721
transform 1 0 9200 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1430_
timestamp 1640608721
transform 1 0 9476 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A2
timestamp 1640608721
transform -1 0 11776 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_111
timestamp 1640608721
transform 1 0 11316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0906_
timestamp 1640608721
transform 1 0 11040 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0950_
timestamp 1640608721
transform 1 0 11776 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0951_
timestamp 1640608721
transform 1 0 12420 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_36_128
timestamp 1640608721
transform 1 0 12880 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1640608721
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1640608721
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_153
timestamp 1640608721
transform 1 0 15180 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0908_
timestamp 1640608721
transform 1 0 15456 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1384_
timestamp 1640608721
transform 1 0 15732 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_1  _0771_
timestamp 1640608721
transform 1 0 17296 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1383_
timestamp 1640608721
transform 1 0 17572 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1640608721
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1382_
timestamp 1640608721
transform 1 0 19228 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__S
timestamp 1640608721
transform 1 0 22080 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_214
timestamp 1640608721
transform 1 0 20792 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_226
timestamp 1640608721
transform 1 0 21896 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_239
timestamp 1640608721
transform 1 0 23092 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_247
timestamp 1640608721
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0766_
timestamp 1640608721
transform -1 0 23828 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1324_
timestamp 1640608721
transform 1 0 22264 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1640608721
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1640608721
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_265
timestamp 1640608721
transform 1 0 25484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_269
timestamp 1640608721
transform 1 0 25852 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1640608721
transform -1 0 26220 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1640608721
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_15
timestamp 1640608721
transform 1 0 2484 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1640608721
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1640608721
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_23
timestamp 1640608721
transform 1 0 3220 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_41
timestamp 1640608721
transform 1 0 4876 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1328_
timestamp 1640608721
transform 1 0 3312 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A
timestamp 1640608721
transform 1 0 5980 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_51
timestamp 1640608721
transform 1 0 5796 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1640608721
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1640608721
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1640608721
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1640608721
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0886_
timestamp 1640608721
transform 1 0 6808 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_clk
timestamp 1640608721
transform -1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__B1
timestamp 1640608721
transform 1 0 7912 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_73
timestamp 1640608721
transform 1 0 7820 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1640608721
transform 1 0 8740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0881_
timestamp 1640608721
transform 1 0 8096 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0882_
timestamp 1640608721
transform -1 0 7544 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0884_
timestamp 1640608721
transform 1 0 7544 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A
timestamp 1640608721
transform 1 0 9936 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_101
timestamp 1640608721
transform 1 0 10396 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1640608721
transform -1 0 9936 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _0905_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform -1 0 9660 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0913_
timestamp 1640608721
transform -1 0 10396 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_109
timestamp 1640608721
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1640608721
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_125
timestamp 1640608721
transform 1 0 12604 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1640608721
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_140
timestamp 1640608721
transform 1 0 13984 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_145
timestamp 1640608721
transform 1 0 14444 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_2  _0933_
timestamp 1640608721
transform 1 0 13340 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_clk
timestamp 1640608721
transform -1 0 14444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_157
timestamp 1640608721
transform 1 0 15548 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1640608721
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0907_
timestamp 1640608721
transform -1 0 16284 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_37_181
timestamp 1640608721
transform 1 0 17756 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1640608721
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0770_
timestamp 1640608721
transform -1 0 17756 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0910_
timestamp 1640608721
transform -1 0 18584 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1189_
timestamp 1640608721
transform 1 0 16652 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_37_190
timestamp 1640608721
transform 1 0 18584 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_202
timestamp 1640608721
transform 1 0 19688 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_214
timestamp 1640608721
transform 1 0 20792 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1640608721
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1640608721
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0919_
timestamp 1640608721
transform 1 0 21804 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0920_
timestamp 1640608721
transform 1 0 22448 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1379_
timestamp 1640608721
transform 1 0 22724 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_37_252
timestamp 1640608721
transform 1 0 24288 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_264
timestamp 1640608721
transform 1 0 25392 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1640608721
transform -1 0 26220 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1640608721
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1640608721
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1640608721
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1640608721
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_29
timestamp 1640608721
transform 1 0 3772 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1640608721
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_2  _0888_
timestamp 1640608721
transform -1 0 5336 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _0889_
timestamp 1640608721
transform 1 0 3864 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_38_46
timestamp 1640608721
transform 1 0 5336 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _0904_
timestamp 1640608721
transform 1 0 5520 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1385_
timestamp 1640608721
transform 1 0 5980 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_38_81
timestamp 1640608721
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1640608721
transform 1 0 8280 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0903_
timestamp 1640608721
transform 1 0 7544 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_89
timestamp 1640608721
transform 1 0 9292 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_93
timestamp 1640608721
transform 1 0 9660 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1640608721
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1640608721
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1640608721
transform -1 0 10028 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_clk
timestamp 1640608721
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1640608721
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1640608721
transform 1 0 12236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1262_
timestamp 1640608721
transform 1 0 12604 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__S
timestamp 1640608721
transform 1 0 13432 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_136
timestamp 1640608721
transform 1 0 13616 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1640608721
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0934_
timestamp 1640608721
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1209_
timestamp 1640608721
transform 1 0 14076 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__S
timestamp 1640608721
transform 1 0 14904 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_A
timestamp 1640608721
transform -1 0 16468 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_152
timestamp 1640608721
transform 1 0 15088 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_164
timestamp 1640608721
transform 1 0 16192 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_171
timestamp 1640608721
transform 1 0 16836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_183
timestamp 1640608721
transform 1 0 17940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clk
timestamp 1640608721
transform 1 0 16468 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__S
timestamp 1640608721
transform 1 0 20056 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1640608721
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1640608721
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_208
timestamp 1640608721
transform 1 0 20240 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1640608721
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0914_
timestamp 1640608721
transform 1 0 19780 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__S
timestamp 1640608721
transform 1 0 21252 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_216
timestamp 1640608721
transform 1 0 20976 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0921_
timestamp 1640608721
transform 1 0 21436 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1309_
timestamp 1640608721
transform 1 0 22080 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_38_237
timestamp 1640608721
transform 1 0 22908 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1640608721
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _1183_
timestamp 1640608721
transform 1 0 23000 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1640608721
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_262
timestamp 1640608721
transform 1 0 25208 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1640608721
transform -1 0 26220 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1640608721
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1192_
timestamp 1640608721
transform 1 0 24932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1640608721
transform 1 0 1380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1640608721
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1640608721
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1640608721
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1640608721
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1337_
timestamp 1640608721
transform -1 0 3036 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_39_21
timestamp 1640608721
transform 1 0 3036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_29
timestamp 1640608721
transform 1 0 3772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_37
timestamp 1640608721
transform 1 0 4508 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1640608721
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1640608721
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_2  _0890_
timestamp 1640608721
transform 1 0 3864 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1386_
timestamp 1640608721
transform 1 0 4692 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1389_
timestamp 1640608721
transform 1 0 3772 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_40_46
timestamp 1640608721
transform 1 0 5336 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_55
timestamp 1640608721
transform 1 0 6164 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1640608721
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_2  _0900_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 6348 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0901_
timestamp 1640608721
transform 1 0 6348 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _0902_
timestamp 1640608721
transform 1 0 5520 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_39_64
timestamp 1640608721
transform 1 0 6992 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_79
timestamp 1640608721
transform 1 0 8372 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_73
timestamp 1640608721
transform 1 0 7820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 1640608721
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0751_
timestamp 1640608721
transform 1 0 7176 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0883_
timestamp 1640608721
transform -1 0 7544 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0887_
timestamp 1640608721
transform 1 0 7544 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0892_
timestamp 1640608721
transform -1 0 8372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_87
timestamp 1640608721
transform 1 0 9108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_85
timestamp 1640608721
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1640608721
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0942_
timestamp 1640608721
transform 1 0 9292 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0943_
timestamp 1640608721
transform 1 0 9844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0944_
timestamp 1640608721
transform 1 0 9200 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1266_
timestamp 1640608721
transform 1 0 9936 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1369_
timestamp 1640608721
transform 1 0 10120 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1640608721
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1640608721
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1640608721
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_107
timestamp 1640608721
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__S
timestamp 1640608721
transform 1 0 10764 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_2  _1169_
timestamp 1640608721
transform 1 0 11684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0940_
timestamp 1640608721
transform 1 0 11868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0939_
timestamp 1640608721
transform -1 0 13064 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0932_
timestamp 1640608721
transform 1 0 12144 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1370_
timestamp 1640608721
transform 1 0 12420 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_40_130
timestamp 1640608721
transform 1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_134
timestamp 1640608721
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1640608721
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0757_
timestamp 1640608721
transform -1 0 13984 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1172_
timestamp 1640608721
transform -1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1373_
timestamp 1640608721
transform 1 0 13984 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_39_157
timestamp 1640608721
transform 1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1640608721
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_157
timestamp 1640608721
transform 1 0 15548 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _1177_
timestamp 1640608721
transform 1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1212_
timestamp 1640608721
transform -1 0 16928 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__S
timestamp 1640608721
transform 1 0 18216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__S
timestamp 1640608721
transform 1 0 17296 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_178
timestamp 1640608721
transform 1 0 17480 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1640608721
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0762_
timestamp 1640608721
transform -1 0 18216 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _0930_
timestamp 1640608721
transform -1 0 17296 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1206_
timestamp 1640608721
transform 1 0 16928 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_clk
timestamp 1640608721
transform 1 0 18216 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1315_
timestamp 1640608721
transform 1 0 19228 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _0924_
timestamp 1640608721
transform 1 0 18492 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0923_
timestamp 1640608721
transform -1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1640608721
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_197
timestamp 1640608721
transform 1 0 19228 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_188
timestamp 1640608721
transform 1 0 18400 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_193
timestamp 1640608721
transform 1 0 18860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__S
timestamp 1640608721
transform 1 0 19044 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1321_
timestamp 1640608721
transform 1 0 20056 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0925_
timestamp 1640608721
transform 1 0 19320 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1377_
timestamp 1640608721
transform 1 0 19596 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1640608721
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_226
timestamp 1640608721
transform 1 0 21896 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1640608721
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0764_
timestamp 1640608721
transform 1 0 20884 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0922_
timestamp 1640608721
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1181_
timestamp 1640608721
transform -1 0 21896 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1378_
timestamp 1640608721
transform 1 0 22080 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_39_250
timestamp 1640608721
transform 1 0 24104 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_242
timestamp 1640608721
transform 1 0 23368 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1640608721
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _0765_
timestamp 1640608721
transform 1 0 23644 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1182_
timestamp 1640608721
transform 1 0 22632 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_262
timestamp 1640608721
transform 1 0 25208 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1640608721
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_265
timestamp 1640608721
transform 1 0 25484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_269
timestamp 1640608721
transform 1 0 25852 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1640608721
transform -1 0 26220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1640608721
transform -1 0 26220 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1640608721
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1640608721
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1640608721
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1640608721
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1640608721
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1640608721
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1640608721
transform 1 0 5796 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1640608721
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__o311a_2  _0895_
timestamp 1640608721
transform 1 0 6348 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1640608721
transform -1 0 6256 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__B1
timestamp 1640608721
transform 1 0 8096 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__S
timestamp 1640608721
transform 1 0 8740 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_78
timestamp 1640608721
transform 1 0 8280 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_82
timestamp 1640608721
transform 1 0 8648 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _0894_
timestamp 1640608721
transform -1 0 7820 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1640608721
transform 1 0 7820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_94
timestamp 1640608721
transform 1 0 9752 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1263_
timestamp 1640608721
transform 1 0 8924 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1368_
timestamp 1640608721
transform 1 0 9844 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1640608721
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1167_
timestamp 1640608721
transform 1 0 12236 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _1168_
timestamp 1640608721
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__S
timestamp 1640608721
transform 1 0 14260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_126
timestamp 1640608721
transform 1 0 12696 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_2  _0760_
timestamp 1640608721
transform 1 0 14444 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1171_
timestamp 1640608721
transform 1 0 13800 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_41_158
timestamp 1640608721
transform 1 0 15640 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0928_
timestamp 1640608721
transform -1 0 16560 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1175_
timestamp 1640608721
transform 1 0 15088 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1640608721
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0761_
timestamp 1640608721
transform 1 0 18216 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1374_
timestamp 1640608721
transform 1 0 16652 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_41_191
timestamp 1640608721
transform 1 0 18676 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__and2b_2  _0926_
timestamp 1640608721
transform 1 0 18860 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0927_
timestamp 1640608721
transform 1 0 19504 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1180_
timestamp 1640608721
transform 1 0 19780 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1640608721
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1640608721
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1640608721
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0763_
timestamp 1640608721
transform 1 0 20516 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1640608721
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1640608721
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_261
timestamp 1640608721
transform 1 0 25116 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_269
timestamp 1640608721
transform 1 0 25852 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1640608721
transform -1 0 26220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1640608721
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1640608721
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1640608721
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1640608721
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1640608721
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_41
timestamp 1640608721
transform 1 0 4876 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1640608721
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_45
timestamp 1640608721
transform 1 0 5244 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _0899_
timestamp 1640608721
transform 1 0 5336 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1388_
timestamp 1640608721
transform 1 0 5796 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__o32a_2  _0898_
timestamp 1640608721
transform 1 0 7360 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _0948_
timestamp 1640608721
transform -1 0 8832 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__S
timestamp 1640608721
transform 1 0 10672 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1640608721
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0945_
timestamp 1640608721
transform -1 0 10672 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0946_
timestamp 1640608721
transform 1 0 8924 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1254_
timestamp 1640608721
transform 1 0 9568 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_106
timestamp 1640608721
transform 1 0 10856 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_110
timestamp 1640608721
transform 1 0 11224 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_117
timestamp 1640608721
transform 1 0 11868 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_125
timestamp 1640608721
transform 1 0 12604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0759_
timestamp 1640608721
transform 1 0 11316 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1640608721
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0938_
timestamp 1640608721
transform 1 0 12880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1215_
timestamp 1640608721
transform 1 0 14076 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1257_
timestamp 1640608721
transform 1 0 13156 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__S
timestamp 1640608721
transform 1 0 15640 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_160
timestamp 1640608721
transform 1 0 15824 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0931_
timestamp 1640608721
transform 1 0 16192 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1176_
timestamp 1640608721
transform -1 0 15640 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_186
timestamp 1640608721
transform 1 0 18216 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0929_
timestamp 1640608721
transform 1 0 16468 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1178_
timestamp 1640608721
transform 1 0 16744 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1179_
timestamp 1640608721
transform 1 0 17480 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1640608721
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_197
timestamp 1640608721
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1640608721
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1376_
timestamp 1640608721
transform 1 0 19320 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_42_215
timestamp 1640608721
transform 1 0 20884 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1640608721
transform 1 0 21988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_239
timestamp 1640608721
transform 1 0 23092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1640608721
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1640608721
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_265
timestamp 1640608721
transform 1 0 25484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_269
timestamp 1640608721
transform 1 0 25852 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1640608721
transform -1 0 26220 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1640608721
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_14
timestamp 1640608721
transform 1 0 2392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_3
timestamp 1640608721
transform 1 0 1380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_9
timestamp 1640608721
transform 1 0 1932 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1640608721
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1640608721
transform 1 0 2024 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_26
timestamp 1640608721
transform 1 0 3496 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_36
timestamp 1640608721
transform 1 0 4416 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1202_
timestamp 1640608721
transform -1 0 4416 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_48
timestamp 1640608721
transform 1 0 5520 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1640608721
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1387_
timestamp 1640608721
transform 1 0 6348 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_43_74
timestamp 1640608721
transform 1 0 7912 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0949_
timestamp 1640608721
transform 1 0 8004 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1366_
timestamp 1640608721
transform 1 0 8280 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1367_
timestamp 1640608721
transform 1 0 9844 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_43_118
timestamp 1640608721
transform 1 0 11960 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1640608721
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0758_
timestamp 1640608721
transform 1 0 11500 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _0937_
timestamp 1640608721
transform 1 0 12144 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _1371_
timestamp 1640608721
transform 1 0 12788 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1372_
timestamp 1640608721
transform 1 0 14352 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1640608721
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1640608721
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_186
timestamp 1640608721
transform 1 0 18216 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1640608721
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1375_
timestamp 1640608721
transform 1 0 16652 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_43_198
timestamp 1640608721
transform 1 0 19320 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_210
timestamp 1640608721
transform 1 0 20424 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1640608721
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1640608721
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1640608721
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_237
timestamp 1640608721
transform 1 0 22908 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_245
timestamp 1640608721
transform 1 0 23644 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_249
timestamp 1640608721
transform 1 0 24012 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1196_
timestamp 1640608721
transform 1 0 23736 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_266
timestamp 1640608721
transform 1 0 25576 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1640608721
transform -1 0 26220 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1197_
timestamp 1640608721
transform 1 0 24748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1198_
timestamp 1640608721
transform 1 0 25024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1199_
timestamp 1640608721
transform 1 0 25300 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1640608721
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1640608721
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1640608721
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1640608721
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1640608721
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1640608721
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1640608721
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_53
timestamp 1640608721
transform 1 0 5980 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_61
timestamp 1640608721
transform 1 0 6716 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0891_
timestamp 1640608721
transform -1 0 7084 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_68
timestamp 1640608721
transform 1 0 7360 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1640608721
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1640608721
transform -1 0 7360 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_85
timestamp 1640608721
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1640608721
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1640608721
transform -1 0 9476 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_2  _1166_
timestamp 1640608721
transform 1 0 10304 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1258_
timestamp 1640608721
transform 1 0 9476 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__S
timestamp 1640608721
transform 1 0 11040 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_110
timestamp 1640608721
transform 1 0 11224 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_122
timestamp 1640608721
transform 1 0 12328 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_130
timestamp 1640608721
transform 1 0 13064 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1640608721
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1640608721
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_2  _0935_
timestamp 1640608721
transform 1 0 13156 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1174_
timestamp 1640608721
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_154
timestamp 1640608721
transform 1 0 15272 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_166
timestamp 1640608721
transform 1 0 16376 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1173_
timestamp 1640608721
transform -1 0 15272 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_44_178
timestamp 1640608721
transform 1 0 17480 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_190
timestamp 1640608721
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1640608721
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1640608721
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1640608721
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1640608721
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1640608721
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1640608721
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1640608721
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1640608721
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 1640608721
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_269
timestamp 1640608721
transform 1 0 25852 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1640608721
transform -1 0 26220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1640608721
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1640608721
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1640608721
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1640608721
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_27
timestamp 1640608721
transform 1 0 3588 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_29
timestamp 1640608721
transform 1 0 3772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_41
timestamp 1640608721
transform 1 0 4876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1640608721
transform 1 0 3680 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1640608721
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1640608721
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1640608721
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1640608721
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_81
timestamp 1640608721
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_85
timestamp 1640608721
transform 1 0 8924 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_93
timestamp 1640608721
transform 1 0 9660 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_97
timestamp 1640608721
transform 1 0 10028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1640608721
transform 1 0 8832 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0947_
timestamp 1640608721
transform 1 0 9752 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1640608721
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1640608721
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1640608721
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1640608721
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_137
timestamp 1640608721
transform 1 0 13708 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_144
timestamp 1640608721
transform 1 0 14352 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1640608721
transform 1 0 13984 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0936_
timestamp 1640608721
transform 1 0 14076 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_156
timestamp 1640608721
transform 1 0 15456 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1640608721
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1640608721
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1640608721
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_193
timestamp 1640608721
transform 1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_197
timestamp 1640608721
transform 1 0 19228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1640608721
transform 1 0 19136 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_209
timestamp 1640608721
transform 1 0 20332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1640608721
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1640608721
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1640608721
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1640608721
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_249
timestamp 1640608721
transform 1 0 24012 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1640608721
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_265
timestamp 1640608721
transform 1 0 25484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_269
timestamp 1640608721
transform 1 0 25852 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1640608721
transform -1 0 26220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1640608721
transform 1 0 24288 0 -1 27200
box -38 -48 130 592
<< labels >>
rlabel metal2 s 662 0 718 800 6 clk
port 0 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 data_req_i
port 1 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 reset
port 2 nsew signal input
rlabel metal3 s 0 824 800 944 6 rxd_uart
port 3 nsew signal input
rlabel metal3 s 26595 688 27395 808 6 slave_data_addr_i[0]
port 4 nsew signal input
rlabel metal3 s 26595 3408 27395 3528 6 slave_data_addr_i[1]
port 5 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 slave_data_addr_i[2]
port 6 nsew signal input
rlabel metal3 s 26595 7624 27395 7744 6 slave_data_addr_i[3]
port 7 nsew signal input
rlabel metal2 s 9218 28739 9274 29539 6 slave_data_addr_i[4]
port 8 nsew signal input
rlabel metal2 s 11242 28739 11298 29539 6 slave_data_addr_i[5]
port 9 nsew signal input
rlabel metal3 s 26595 10480 27395 10600 6 slave_data_addr_i[6]
port 10 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 slave_data_addr_i[7]
port 11 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 slave_data_addr_i[8]
port 12 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 slave_data_addr_i[9]
port 13 nsew signal input
rlabel metal3 s 26595 2048 27395 2168 6 slave_data_be_i[0]
port 14 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 slave_data_be_i[1]
port 15 nsew signal input
rlabel metal3 s 26595 4904 27395 5024 6 slave_data_be_i[2]
port 16 nsew signal input
rlabel metal2 s 7286 28739 7342 29539 6 slave_data_be_i[3]
port 17 nsew signal input
rlabel metal2 s 478 28739 534 29539 6 slave_data_gnt_o
port 18 nsew signal tristate
rlabel metal2 s 4526 0 4582 800 6 slave_data_rdata_o[0]
port 19 nsew signal tristate
rlabel metal3 s 26595 14696 27395 14816 6 slave_data_rdata_o[10]
port 20 nsew signal tristate
rlabel metal2 s 14186 28739 14242 29539 6 slave_data_rdata_o[11]
port 21 nsew signal tristate
rlabel metal2 s 15106 28739 15162 29539 6 slave_data_rdata_o[12]
port 22 nsew signal tristate
rlabel metal3 s 26595 17552 27395 17672 6 slave_data_rdata_o[13]
port 23 nsew signal tristate
rlabel metal3 s 0 13608 800 13728 6 slave_data_rdata_o[14]
port 24 nsew signal tristate
rlabel metal2 s 18050 28739 18106 29539 6 slave_data_rdata_o[15]
port 25 nsew signal tristate
rlabel metal3 s 26595 18912 27395 19032 6 slave_data_rdata_o[16]
port 26 nsew signal tristate
rlabel metal2 s 19982 28739 20038 29539 6 slave_data_rdata_o[17]
port 27 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 slave_data_rdata_o[18]
port 28 nsew signal tristate
rlabel metal2 s 18878 0 18934 800 6 slave_data_rdata_o[19]
port 29 nsew signal tristate
rlabel metal2 s 5354 28739 5410 29539 6 slave_data_rdata_o[1]
port 30 nsew signal tristate
rlabel metal2 s 22006 28739 22062 29539 6 slave_data_rdata_o[20]
port 31 nsew signal tristate
rlabel metal3 s 26595 21768 27395 21888 6 slave_data_rdata_o[21]
port 32 nsew signal tristate
rlabel metal3 s 26595 23128 27395 23248 6 slave_data_rdata_o[22]
port 33 nsew signal tristate
rlabel metal2 s 20166 0 20222 800 6 slave_data_rdata_o[23]
port 34 nsew signal tristate
rlabel metal2 s 21546 0 21602 800 6 slave_data_rdata_o[24]
port 35 nsew signal tristate
rlabel metal2 s 22834 0 22890 800 6 slave_data_rdata_o[25]
port 36 nsew signal tristate
rlabel metal2 s 23938 28739 23994 29539 6 slave_data_rdata_o[26]
port 37 nsew signal tristate
rlabel metal2 s 24950 28739 25006 29539 6 slave_data_rdata_o[27]
port 38 nsew signal tristate
rlabel metal3 s 26595 28704 27395 28824 6 slave_data_rdata_o[28]
port 39 nsew signal tristate
rlabel metal2 s 26882 28739 26938 29539 6 slave_data_rdata_o[29]
port 40 nsew signal tristate
rlabel metal2 s 7102 0 7158 800 6 slave_data_rdata_o[2]
port 41 nsew signal tristate
rlabel metal2 s 24122 0 24178 800 6 slave_data_rdata_o[30]
port 42 nsew signal tristate
rlabel metal2 s 26698 0 26754 800 6 slave_data_rdata_o[31]
port 43 nsew signal tristate
rlabel metal2 s 8298 28739 8354 29539 6 slave_data_rdata_o[3]
port 44 nsew signal tristate
rlabel metal2 s 10230 28739 10286 29539 6 slave_data_rdata_o[4]
port 45 nsew signal tristate
rlabel metal3 s 26595 9120 27395 9240 6 slave_data_rdata_o[5]
port 46 nsew signal tristate
rlabel metal3 s 0 6264 800 6384 6 slave_data_rdata_o[6]
port 47 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 slave_data_rdata_o[7]
port 48 nsew signal tristate
rlabel metal2 s 15014 0 15070 800 6 slave_data_rdata_o[8]
port 49 nsew signal tristate
rlabel metal3 s 26595 11840 27395 11960 6 slave_data_rdata_o[9]
port 50 nsew signal tristate
rlabel metal2 s 1398 28739 1454 29539 6 slave_data_rvalid_o
port 51 nsew signal tristate
rlabel metal2 s 4342 28739 4398 29539 6 slave_data_wdata_i[0]
port 52 nsew signal input
rlabel metal2 s 13174 28739 13230 29539 6 slave_data_wdata_i[10]
port 53 nsew signal input
rlabel metal3 s 26595 16056 27395 16176 6 slave_data_wdata_i[11]
port 54 nsew signal input
rlabel metal2 s 16118 28739 16174 29539 6 slave_data_wdata_i[12]
port 55 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 slave_data_wdata_i[13]
port 56 nsew signal input
rlabel metal2 s 17038 28739 17094 29539 6 slave_data_wdata_i[14]
port 57 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 slave_data_wdata_i[15]
port 58 nsew signal input
rlabel metal2 s 19062 28739 19118 29539 6 slave_data_wdata_i[16]
port 59 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 slave_data_wdata_i[17]
port 60 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 slave_data_wdata_i[18]
port 61 nsew signal input
rlabel metal2 s 20994 28739 21050 29539 6 slave_data_wdata_i[19]
port 62 nsew signal input
rlabel metal2 s 6274 28739 6330 29539 6 slave_data_wdata_i[1]
port 63 nsew signal input
rlabel metal3 s 26595 20272 27395 20392 6 slave_data_wdata_i[20]
port 64 nsew signal input
rlabel metal2 s 22926 28739 22982 29539 6 slave_data_wdata_i[21]
port 65 nsew signal input
rlabel metal3 s 26595 24488 27395 24608 6 slave_data_wdata_i[22]
port 66 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 slave_data_wdata_i[23]
port 67 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 slave_data_wdata_i[24]
port 68 nsew signal input
rlabel metal3 s 26595 25984 27395 26104 6 slave_data_wdata_i[25]
port 69 nsew signal input
rlabel metal3 s 26595 27344 27395 27464 6 slave_data_wdata_i[26]
port 70 nsew signal input
rlabel metal2 s 25870 28739 25926 29539 6 slave_data_wdata_i[27]
port 71 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 slave_data_wdata_i[28]
port 72 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 slave_data_wdata_i[29]
port 73 nsew signal input
rlabel metal3 s 26595 6264 27395 6384 6 slave_data_wdata_i[2]
port 74 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 slave_data_wdata_i[30]
port 75 nsew signal input
rlabel metal3 s 0 28432 800 28552 6 slave_data_wdata_i[31]
port 76 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 slave_data_wdata_i[3]
port 77 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 slave_data_wdata_i[4]
port 78 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 slave_data_wdata_i[5]
port 79 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 slave_data_wdata_i[6]
port 80 nsew signal input
rlabel metal2 s 12162 28739 12218 29539 6 slave_data_wdata_i[7]
port 81 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 slave_data_wdata_i[8]
port 82 nsew signal input
rlabel metal3 s 26595 13336 27395 13456 6 slave_data_wdata_i[9]
port 83 nsew signal input
rlabel metal2 s 2410 28739 2466 29539 6 slave_data_we_i
port 84 nsew signal input
rlabel metal2 s 3330 28739 3386 29539 6 txd_uart
port 85 nsew signal tristate
rlabel metal4 s 5130 2128 5450 27248 6 vccd1
port 86 nsew power input
rlabel metal4 s 13502 2128 13822 27248 6 vccd1
port 86 nsew power input
rlabel metal4 s 21874 2128 22194 27248 6 vccd1
port 86 nsew power input
rlabel metal4 s 9316 2128 9636 27248 6 vssd1
port 87 nsew ground input
rlabel metal4 s 17688 2128 18008 27248 6 vssd1
port 87 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 27395 29539
<< end >>
